

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946;

  OAI221_X1 U3532 ( .B1(n4527), .B2(keyinput56), .C1(n6171), .C2(keyinput122), 
        .A(n4383), .ZN(n4387) );
  NAND2_X1 U3533 ( .A1(n3897), .A2(n3896), .ZN(n5147) );
  NAND2_X1 U3534 ( .A1(n4748), .A2(n3827), .ZN(n4709) );
  OR2_X1 U3535 ( .A1(n3840), .A2(n4047), .ZN(n3847) );
  CLKBUF_X2 U3536 ( .A(n3366), .Z(n4217) );
  CLKBUF_X2 U3537 ( .A(n3304), .Z(n5436) );
  CLKBUF_X1 U3538 ( .A(n4127), .Z(n5440) );
  CLKBUF_X2 U3539 ( .A(n3296), .Z(n5448) );
  CLKBUF_X2 U3540 ( .A(n4243), .Z(n3088) );
  CLKBUF_X2 U3541 ( .A(n3218), .Z(n3086) );
  CLKBUF_X2 U3542 ( .A(n3297), .Z(n5447) );
  AND4_X1 U3543 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3181)
         );
  AND4_X1 U3544 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3182)
         );
  INV_X1 U3545 ( .A(n3319), .ZN(n4737) );
  AND2_X1 U3546 ( .A1(n3119), .A2(n3112), .ZN(n3296) );
  AND2_X1 U3547 ( .A1(n3112), .A2(n4788), .ZN(n4243) );
  AND2_X2 U3548 ( .A1(n3124), .A2(n4760), .ZN(n3304) );
  AOI22_X1 U3549 ( .A1(n4662), .A2(keyinput28), .B1(keyinput120), .B2(n4401), 
        .ZN(n4400) );
  AOI22_X1 U3550 ( .A1(n4527), .A2(keyinput56), .B1(keyinput122), .B2(n6171), 
        .ZN(n4383) );
  AND2_X1 U3552 ( .A1(n4760), .A2(n4788), .ZN(n3297) );
  OAI221_X1 U3553 ( .B1(n4662), .B2(keyinput28), .C1(n4401), .C2(keyinput120), 
        .A(n4400), .ZN(n4409) );
  AND4_X1 U3554 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3180)
         );
  AND2_X1 U3556 ( .A1(n4999), .A2(n4886), .ZN(n3865) );
  INV_X1 U3558 ( .A(n4289), .ZN(n3513) );
  INV_X2 U3559 ( .A(n4948), .ZN(n4699) );
  AND2_X1 U3560 ( .A1(n4710), .A2(n4711), .ZN(n3827) );
  INV_X1 U3563 ( .A(n6495), .ZN(n6483) );
  AND2_X4 U3565 ( .A1(n3124), .A2(n3112), .ZN(n3364) );
  AND2_X4 U3566 ( .A1(n3124), .A2(n3118), .ZN(n3302) );
  OAI21_X2 U3567 ( .B1(n4722), .B2(STATE2_REG_0__SCAN_IN), .A(n3377), .ZN(
        n3380) );
  AND2_X4 U3570 ( .A1(n4615), .A2(n4788), .ZN(n3397) );
  INV_X1 U3571 ( .A(n6128), .ZN(n6213) );
  OR2_X1 U3572 ( .A1(n5155), .A2(n3952), .ZN(n3953) );
  AND2_X1 U3573 ( .A1(n3291), .A2(n3344), .ZN(n4648) );
  NAND2_X2 U3574 ( .A1(n6261), .A2(n5686), .ZN(n6014) );
  CLKBUF_X2 U3575 ( .A(n3316), .Z(n3618) );
  NAND2_X1 U3576 ( .A1(n3363), .A2(n3362), .ZN(n3603) );
  NAND2_X4 U3577 ( .A1(n4737), .A2(n5184), .ZN(n3642) );
  BUF_X1 U3578 ( .A(n3320), .Z(n5303) );
  INV_X1 U3579 ( .A(n5184), .ZN(n4744) );
  AND4_X1 U3580 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3132)
         );
  BUF_X2 U3581 ( .A(n4159), .Z(n3152) );
  BUF_X2 U3582 ( .A(n3446), .Z(n5427) );
  AND2_X2 U3583 ( .A1(n3119), .A2(n3118), .ZN(n3366) );
  AOI21_X1 U3584 ( .B1(n5510), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5509), 
        .ZN(n5511) );
  NOR2_X1 U3585 ( .A1(n5714), .A2(n4282), .ZN(n5508) );
  OR2_X1 U3586 ( .A1(n3780), .A2(n5720), .ZN(n5714) );
  AND3_X1 U3587 ( .A1(n4296), .A2(n4295), .A3(n4294), .ZN(n4297) );
  AOI221_X1 U3588 ( .B1(n6002), .B2(REIP_REG_22__SCAN_IN), .C1(n5992), .C2(
        REIP_REG_22__SCAN_IN), .A(n5984), .ZN(n5985) );
  NAND2_X1 U3589 ( .A1(n5603), .A2(n4254), .ZN(n5479) );
  AND4_X1 U3590 ( .A1(n5527), .A2(n3100), .A3(n5526), .A4(n3104), .ZN(n5528)
         );
  AND2_X1 U3591 ( .A1(n3529), .A2(n3528), .ZN(n3530) );
  INV_X1 U3592 ( .A(n5052), .ZN(n3897) );
  OR2_X1 U3593 ( .A1(n3521), .A2(n3520), .ZN(n5808) );
  NAND2_X1 U3594 ( .A1(n3835), .A2(n3834), .ZN(n4754) );
  NAND2_X1 U3595 ( .A1(n3804), .A2(n4693), .ZN(n4750) );
  XNOR2_X1 U3596 ( .A(n3455), .B(n3463), .ZN(n3828) );
  AND2_X1 U3597 ( .A1(n3788), .A2(n4026), .ZN(n3804) );
  NAND2_X1 U3598 ( .A1(n3441), .A2(n3464), .ZN(n3455) );
  CLKBUF_X1 U3599 ( .A(n4719), .Z(n6583) );
  NOR2_X2 U3600 ( .A1(n5574), .A2(n5575), .ZN(n5573) );
  OR2_X1 U3601 ( .A1(n4231), .A2(n4230), .ZN(n5170) );
  OR2_X1 U3603 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  NAND2_X1 U3604 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  XNOR2_X1 U3605 ( .A(n3333), .B(n3331), .ZN(n3795) );
  AND2_X1 U3606 ( .A1(n3250), .A2(n3249), .ZN(n3331) );
  NOR2_X1 U3607 ( .A1(n5053), .A2(n5014), .ZN(n3896) );
  AND3_X1 U3608 ( .A1(n3653), .A2(n3710), .A3(n3652), .ZN(n4713) );
  OR2_X1 U3610 ( .A1(n4620), .A2(n5683), .ZN(n3632) );
  INV_X1 U3611 ( .A(n5659), .ZN(n3091) );
  INV_X1 U3612 ( .A(n5686), .ZN(n5682) );
  AND4_X1 U3613 ( .A1(n3178), .A2(n3177), .A3(n3176), .A4(n3175), .ZN(n3179)
         );
  AND4_X1 U3614 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3202)
         );
  AND4_X1 U3615 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .ZN(n3201)
         );
  AND4_X1 U3616 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3199)
         );
  AND4_X1 U3618 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3133)
         );
  INV_X2 U3619 ( .A(n3261), .ZN(n3084) );
  INV_X2 U3620 ( .A(n6696), .ZN(n3085) );
  AND2_X2 U3621 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4788) );
  AND2_X2 U3622 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U3623 ( .A1(n3319), .A2(n3628), .ZN(n3634) );
  NAND2_X1 U3624 ( .A1(n4934), .A2(n3579), .ZN(n4705) );
  OR2_X4 U3625 ( .A1(n3162), .A2(n3161), .ZN(n5686) );
  AND2_X2 U3626 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  XNOR2_X1 U3627 ( .A(n3439), .B(n6482), .ZN(n4981) );
  NOR2_X2 U3628 ( .A1(n4430), .A2(n3933), .ZN(n3994) );
  NAND2_X1 U3629 ( .A1(n3438), .A2(n3437), .ZN(n3439) );
  OR3_X4 U3630 ( .A1(n4686), .A2(n4687), .A3(n5336), .ZN(n4714) );
  AOI21_X2 U3631 ( .B1(n5545), .B2(n5495), .A(n5494), .ZN(n5496) );
  OR2_X1 U3632 ( .A1(n3626), .A2(n3634), .ZN(n4619) );
  AND2_X1 U3633 ( .A1(n3112), .A2(n3125), .ZN(n3218) );
  NAND4_X1 U3634 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3087)
         );
  NAND2_X2 U3635 ( .A1(n5157), .A2(n5156), .ZN(n5155) );
  NOR2_X4 U3636 ( .A1(n5147), .A2(n5148), .ZN(n5157) );
  OR2_X4 U3637 ( .A1(n5613), .A2(n5604), .ZN(n5606) );
  AND2_X1 U3638 ( .A1(n4615), .A2(n3125), .ZN(n3089) );
  INV_X1 U3639 ( .A(n3634), .ZN(n3090) );
  AND2_X1 U3640 ( .A1(n6147), .A2(n5183), .ZN(n3092) );
  AND2_X2 U3642 ( .A1(n6147), .A2(n5183), .ZN(n6233) );
  INV_X4 U3643 ( .A(n6233), .ZN(n6229) );
  AND2_X4 U3644 ( .A1(n4615), .A2(n3119), .ZN(n3303) );
  AND2_X4 U3645 ( .A1(n3124), .A2(n4615), .ZN(n3425) );
  AND2_X1 U3646 ( .A1(n3314), .A2(n5686), .ZN(n3227) );
  OR2_X1 U3647 ( .A1(n4699), .A2(n6809), .ZN(n3363) );
  OR2_X1 U3648 ( .A1(n5184), .A2(n6809), .ZN(n3362) );
  NAND2_X1 U3649 ( .A1(n3779), .A2(n3540), .ZN(n4283) );
  NAND2_X1 U3650 ( .A1(n3482), .A2(n3481), .ZN(n3506) );
  AND2_X1 U3651 ( .A1(n5374), .A2(n3524), .ZN(n3517) );
  OR2_X1 U3652 ( .A1(n4635), .A2(n3734), .ZN(n4641) );
  AND2_X1 U3653 ( .A1(n3628), .A2(n3579), .ZN(n3569) );
  NAND2_X1 U3654 ( .A1(n3274), .A2(n3280), .ZN(n3293) );
  NAND2_X1 U3655 ( .A1(n3795), .A2(n6809), .ZN(n3274) );
  INV_X1 U3656 ( .A(n3317), .ZN(n3318) );
  NAND2_X1 U3657 ( .A1(n3409), .A2(n3408), .ZN(n4819) );
  AND2_X1 U3658 ( .A1(n3597), .A2(n3569), .ZN(n3607) );
  INV_X1 U3659 ( .A(n3642), .ZN(n4680) );
  NAND2_X1 U3660 ( .A1(n5675), .A2(n5664), .ZN(n5666) );
  AND2_X1 U3661 ( .A1(n5795), .A2(n4269), .ZN(n3541) );
  OR2_X1 U3662 ( .A1(n5749), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4296)
         );
  OAI21_X1 U3663 ( .B1(n3513), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5753), 
        .ZN(n5749) );
  CLKBUF_X1 U3664 ( .A(n3634), .Z(n5659) );
  INV_X1 U3665 ( .A(n3292), .ZN(n3281) );
  XNOR2_X1 U3666 ( .A(n4794), .B(n5202), .ZN(n4721) );
  INV_X1 U3667 ( .A(n5259), .ZN(n6551) );
  AND2_X1 U3668 ( .A1(n6276), .A2(n5687), .ZN(n6268) );
  INV_X1 U3669 ( .A(n6276), .ZN(n6267) );
  OR2_X1 U3670 ( .A1(n6425), .A2(n4611), .ZN(n6434) );
  OR2_X1 U3671 ( .A1(n4658), .A2(n6778), .ZN(n6410) );
  INV_X1 U3672 ( .A(n6410), .ZN(n6429) );
  CLKBUF_X1 U3673 ( .A(n3446), .Z(n4105) );
  AND2_X1 U3674 ( .A1(n5784), .A2(n3096), .ZN(n3524) );
  OR2_X1 U3675 ( .A1(n3260), .A2(n3259), .ZN(n3508) );
  INV_X1 U3676 ( .A(n3615), .ZN(n3230) );
  NAND2_X1 U3677 ( .A1(n3231), .A2(n4948), .ZN(n3233) );
  NAND2_X1 U3678 ( .A1(n4939), .A2(n3319), .ZN(n3735) );
  NAND2_X1 U3679 ( .A1(n4744), .A2(n3628), .ZN(n3244) );
  NAND2_X1 U3680 ( .A1(n3994), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4033)
         );
  OR2_X1 U3681 ( .A1(n3516), .A2(n5804), .ZN(n3519) );
  AND2_X1 U3682 ( .A1(n5402), .A2(n3519), .ZN(n5806) );
  OR2_X1 U3683 ( .A1(n5401), .A2(n5400), .ZN(n5807) );
  NAND2_X1 U3684 ( .A1(n3241), .A2(n3240), .ZN(n3333) );
  NAND2_X1 U3685 ( .A1(n3327), .A2(n3102), .ZN(n3352) );
  NAND2_X1 U3686 ( .A1(n3379), .A2(n3378), .ZN(n3785) );
  OR2_X1 U3687 ( .A1(n3321), .A2(n4698), .ZN(n4620) );
  OAI21_X1 U3688 ( .B1(n3358), .B2(n5505), .A(n3357), .ZN(n3359) );
  INV_X1 U3689 ( .A(n4819), .ZN(n4820) );
  OAI21_X1 U3690 ( .B1(n6940), .B2(n4801), .A(n6797), .ZN(n4727) );
  INV_X1 U3691 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U3692 ( .A1(n4728), .A2(n5184), .ZN(n6788) );
  NAND2_X1 U3693 ( .A1(n6790), .A2(n5184), .ZN(n4587) );
  OR2_X1 U3694 ( .A1(n4658), .A2(n4587), .ZN(n4594) );
  NOR2_X2 U3695 ( .A1(n5479), .A2(n5480), .ZN(n5533) );
  NOR2_X1 U3696 ( .A1(n4190), .A2(n4189), .ZN(n4229) );
  NAND2_X1 U3697 ( .A1(n5621), .A2(n4152), .ZN(n5622) );
  AND2_X1 U3698 ( .A1(n4151), .A2(n5620), .ZN(n4152) );
  OR2_X1 U3699 ( .A1(n4066), .A2(n3995), .ZN(n4167) );
  NAND2_X1 U3700 ( .A1(n4085), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4066)
         );
  AND2_X1 U3701 ( .A1(n4083), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4085)
         );
  AND2_X1 U3702 ( .A1(n5657), .A2(n5632), .ZN(n5643) );
  NOR2_X1 U3703 ( .A1(n4144), .A2(n5791), .ZN(n4120) );
  OR2_X1 U3704 ( .A1(n5778), .A2(n5779), .ZN(n5776) );
  OR2_X1 U3705 ( .A1(n5666), .A2(n5655), .ZN(n5778) );
  AND2_X1 U3706 ( .A1(n4032), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4012)
         );
  NAND2_X1 U3707 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n4012), .ZN(n4144)
         );
  NOR2_X1 U3708 ( .A1(n4401), .A2(n4033), .ZN(n4032) );
  INV_X1 U3709 ( .A(n3898), .ZN(n3899) );
  NOR2_X1 U3710 ( .A1(n6171), .A2(n3900), .ZN(n3932) );
  NAND2_X1 U3711 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n3866), .ZN(n3898)
         );
  NOR2_X1 U3712 ( .A1(n5181), .A2(n3848), .ZN(n3866) );
  NOR2_X1 U3713 ( .A1(n3841), .A2(n5252), .ZN(n3842) );
  OAI211_X1 U3714 ( .C1(n5255), .C2(n5473), .A(n3838), .B(n3837), .ZN(n4753)
         );
  NAND2_X1 U3715 ( .A1(n3829), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3841)
         );
  INV_X1 U3716 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3813) );
  NOR2_X1 U3717 ( .A1(n3819), .A2(n3813), .ZN(n3829) );
  NOR2_X1 U3718 ( .A1(n4471), .A2(n4350), .ZN(n3820) );
  NAND2_X1 U3719 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3820), .ZN(n3819)
         );
  INV_X1 U3720 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4350) );
  INV_X1 U3721 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4471) );
  OAI221_X1 U3722 ( .B1(n4430), .B2(keyinput107), .C1(n6849), .C2(keyinput93), 
        .A(n4429), .ZN(n4431) );
  AOI22_X1 U3723 ( .A1(n4430), .A2(keyinput107), .B1(n6849), .B2(keyinput93), 
        .ZN(n4429) );
  AOI22_X1 U3724 ( .A1(n5772), .A2(n4292), .B1(n3513), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5755) );
  INV_X1 U3725 ( .A(n5658), .ZN(n5669) );
  AND2_X1 U3727 ( .A1(n5319), .A2(n5321), .ZN(n3515) );
  OR2_X1 U3728 ( .A1(n5795), .A2(n6441), .ZN(n5321) );
  OR2_X1 U3729 ( .A1(n5795), .A2(n3669), .ZN(n5319) );
  AND2_X1 U3730 ( .A1(n5795), .A2(n6441), .ZN(n5322) );
  AND3_X1 U3731 ( .A1(n3657), .A2(n3710), .A3(n3656), .ZN(n4806) );
  AND2_X1 U3732 ( .A1(n3655), .A2(n3654), .ZN(n4564) );
  AND2_X1 U3733 ( .A1(n3624), .A2(n6802), .ZN(n3761) );
  OR2_X1 U3734 ( .A1(n3794), .A2(n4948), .ZN(n6756) );
  OR2_X1 U3735 ( .A1(n4925), .A2(n4720), .ZN(n4726) );
  NAND2_X1 U3736 ( .A1(n3390), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3396) );
  INV_X1 U3737 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6759) );
  INV_X1 U3738 ( .A(n3628), .ZN(n4728) );
  INV_X2 U3739 ( .A(n3968), .ZN(n4939) );
  NAND2_X2 U3740 ( .A1(n3609), .A2(n3608), .ZN(n4635) );
  NAND2_X1 U3741 ( .A1(n5311), .A2(n5187), .ZN(n6183) );
  AND2_X1 U3742 ( .A1(n6147), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6234) );
  INV_X1 U3743 ( .A(n6216), .ZN(n6209) );
  NAND2_X1 U3744 ( .A1(n6147), .A2(n5173), .ZN(n6128) );
  INV_X1 U3745 ( .A(n6240), .ZN(n6219) );
  INV_X1 U3746 ( .A(n5663), .ZN(n6257) );
  INV_X1 U3747 ( .A(n6277), .ZN(n6272) );
  NAND2_X1 U3748 ( .A1(n4704), .A2(n6380), .ZN(n6276) );
  INV_X1 U3749 ( .A(n6279), .ZN(n6298) );
  INV_X1 U3750 ( .A(n6327), .ZN(n6330) );
  INV_X1 U3751 ( .A(n6323), .ZN(n6332) );
  OAI21_X1 U3752 ( .B1(n5551), .B2(n5562), .A(n5550), .ZN(n6025) );
  OAI21_X1 U3753 ( .B1(n5643), .B2(n5634), .A(n5633), .ZN(n5983) );
  AND2_X1 U3754 ( .A1(n5666), .A2(n5665), .ZN(n6266) );
  XNOR2_X1 U3755 ( .A(n3545), .B(n3544), .ZN(n5478) );
  OR2_X1 U3756 ( .A1(n5848), .A2(n3774), .ZN(n5833) );
  NAND2_X1 U3757 ( .A1(n5749), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4295) );
  OR2_X1 U3758 ( .A1(n4555), .A2(n3759), .ZN(n4650) );
  INV_X1 U3759 ( .A(n6485), .ZN(n6497) );
  INV_X1 U3760 ( .A(n6476), .ZN(n6503) );
  NAND2_X1 U3761 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  NAND2_X1 U3762 ( .A1(n3279), .A2(n3292), .ZN(n3284) );
  CLKBUF_X1 U3763 ( .A(n4617), .Z(n4618) );
  CLKBUF_X1 U3764 ( .A(n4718), .Z(n4960) );
  INV_X1 U3765 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6770) );
  INV_X1 U3766 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6777) );
  CLKBUF_X1 U3767 ( .A(n4721), .Z(n6553) );
  INV_X1 U3768 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3113) );
  INV_X1 U3769 ( .A(n5260), .ZN(n5299) );
  OR3_X1 U3770 ( .A1(n6652), .A2(n5259), .A3(n5258), .ZN(n6687) );
  INV_X1 U3771 ( .A(n5227), .ZN(n5243) );
  NAND2_X1 U3772 ( .A1(n4635), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6797) );
  INV_X1 U3773 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6809) );
  AND2_X1 U3774 ( .A1(n4261), .A2(n4260), .ZN(n4262) );
  NOR2_X1 U3775 ( .A1(n3626), .A2(n5184), .ZN(n3094) );
  NAND2_X1 U3777 ( .A1(n5728), .A2(n5727), .ZN(n3780) );
  NAND2_X1 U3778 ( .A1(n5795), .A2(n3690), .ZN(n3096) );
  NOR2_X1 U3779 ( .A1(n4925), .A2(n4810), .ZN(n3097) );
  NOR4_X2 U3780 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n6928)
         );
  OAI21_X2 U3781 ( .B1(n5320), .B2(n5322), .A(n3515), .ZN(n5375) );
  AND2_X4 U3782 ( .A1(n3628), .A2(n3087), .ZN(n5179) );
  AND2_X1 U3783 ( .A1(n4302), .A2(n4301), .ZN(n3098) );
  NAND2_X1 U3784 ( .A1(n6276), .A2(n4707), .ZN(n6277) );
  AND3_X1 U3785 ( .A1(n3533), .A2(n5872), .A3(n4492), .ZN(n3099) );
  OR2_X1 U3786 ( .A1(n5543), .A2(n6497), .ZN(n3100) );
  AND4_X1 U3787 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3101)
         );
  OR2_X1 U3788 ( .A1(n3326), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3102)
         );
  AND4_X1 U3789 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3103)
         );
  OR3_X1 U3790 ( .A1(n5525), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n3544), 
        .ZN(n3104) );
  AND3_X1 U3791 ( .A1(n5854), .A2(n3536), .A3(n5871), .ZN(n3105) );
  AND2_X1 U3792 ( .A1(n3333), .A2(n3332), .ZN(n3106) );
  AND2_X1 U3793 ( .A1(n3593), .A2(n3578), .ZN(n3584) );
  NOR2_X1 U3794 ( .A1(n5303), .A2(n3570), .ZN(n3593) );
  OR2_X1 U3795 ( .A1(n3558), .A2(n3574), .ZN(n3560) );
  INV_X1 U3796 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3328) );
  AND2_X1 U3797 ( .A1(n5184), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3576) );
  OR2_X1 U3798 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  AND2_X1 U3799 ( .A1(n3523), .A2(n5785), .ZN(n3529) );
  NAND2_X1 U3800 ( .A1(n3614), .A2(n4696), .ZN(n3321) );
  OR2_X1 U3801 ( .A1(n3272), .A2(n3271), .ZN(n3382) );
  AND2_X1 U3802 ( .A1(n3576), .A2(n4699), .ZN(n3597) );
  INV_X1 U3803 ( .A(n3647), .ZN(n3730) );
  INV_X1 U3804 ( .A(n5457), .ZN(n5470) );
  NAND2_X1 U3805 ( .A1(n3932), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3933)
         );
  INV_X1 U3806 ( .A(n5882), .ZN(n3700) );
  AND2_X1 U3807 ( .A1(n5806), .A2(n3518), .ZN(n5784) );
  NOR2_X1 U3808 ( .A1(n4991), .A2(n3491), .ZN(n3492) );
  AND2_X1 U3809 ( .A1(n3119), .A2(n4760), .ZN(n3365) );
  NAND2_X1 U3810 ( .A1(n4721), .A2(n6809), .ZN(n3409) );
  INV_X1 U3811 ( .A(n4806), .ZN(n3658) );
  OR2_X1 U3812 ( .A1(n4719), .A2(n4047), .ZN(n3788) );
  OR2_X1 U3813 ( .A1(n5463), .A2(n5491), .ZN(n5172) );
  NOR2_X1 U3814 ( .A1(n5170), .A2(n5169), .ZN(n5464) );
  OR2_X1 U3815 ( .A1(n4167), .A2(n5564), .ZN(n4190) );
  NOR2_X1 U3816 ( .A1(n4123), .A2(n5767), .ZN(n4083) );
  NAND2_X1 U3817 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3900)
         );
  INV_X1 U3818 ( .A(n5179), .ZN(n5520) );
  OR2_X1 U3819 ( .A1(n3522), .A2(n5808), .ZN(n5785) );
  AND2_X1 U3820 ( .A1(n3651), .A2(n3650), .ZN(n5336) );
  XNOR2_X1 U3821 ( .A(n3348), .B(n3347), .ZN(n3338) );
  XNOR2_X1 U3822 ( .A(n3786), .B(n4819), .ZN(n3818) );
  AND2_X1 U3823 ( .A1(n5709), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U3824 ( .A1(n4754), .A2(n4753), .ZN(n3839) );
  XNOR2_X1 U3825 ( .A(n5172), .B(n5171), .ZN(n5709) );
  AND2_X1 U3826 ( .A1(n5570), .A2(n5569), .ZN(n5621) );
  NAND2_X1 U3827 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4120), .ZN(n4123)
         );
  NAND2_X1 U3828 ( .A1(n5570), .A2(n5569), .ZN(n5631) );
  NAND2_X1 U3829 ( .A1(n3579), .A2(n4948), .ZN(n3626) );
  OR2_X1 U3830 ( .A1(n5862), .A2(n5853), .ZN(n5845) );
  AND2_X1 U3831 ( .A1(n5786), .A2(n5785), .ZN(n5797) );
  INV_X1 U3832 ( .A(n4726), .ZN(n4729) );
  INV_X1 U3833 ( .A(n5024), .ZN(n4905) );
  OR2_X1 U3834 ( .A1(n4839), .A2(n6551), .ZN(n5260) );
  BUF_X1 U3835 ( .A(n3818), .Z(n4925) );
  NAND2_X1 U3836 ( .A1(n3396), .A2(n3395), .ZN(n5202) );
  INV_X1 U3837 ( .A(n5473), .ZN(n5467) );
  INV_X1 U3838 ( .A(n3244), .ZN(n5310) );
  INV_X1 U3839 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6912) );
  AND2_X1 U3840 ( .A1(n5311), .A2(n5176), .ZN(n6235) );
  AND2_X1 U3841 ( .A1(n5540), .A2(n5180), .ZN(n6240) );
  NAND2_X1 U3842 ( .A1(n3642), .A2(n3634), .ZN(n5521) );
  AND2_X1 U3843 ( .A1(n5776), .A2(n5649), .ZN(n5651) );
  AND2_X1 U3844 ( .A1(n4660), .A2(n6789), .ZN(n6323) );
  INV_X1 U3845 ( .A(n6334), .ZN(n6383) );
  OR2_X1 U3846 ( .A1(n5693), .A2(n6696), .ZN(n4261) );
  AOI21_X1 U3847 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n6036) );
  NOR2_X1 U3848 ( .A1(n5631), .A2(n5630), .ZN(n5675) );
  INV_X1 U3849 ( .A(n6434), .ZN(n6387) );
  NAND2_X1 U3850 ( .A1(n3842), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3848)
         );
  NAND2_X1 U3851 ( .A1(n4635), .A2(n6802), .ZN(n4658) );
  INV_X1 U3852 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3544) );
  AND2_X1 U3853 ( .A1(n6437), .A2(n3768), .ZN(n6060) );
  AND2_X1 U3854 ( .A1(n3770), .A2(n3769), .ZN(n6061) );
  OAI21_X1 U3855 ( .B1(n3765), .B2(n5380), .A(n3754), .ZN(n6437) );
  AND2_X1 U3856 ( .A1(n3761), .A2(n3633), .ZN(n6485) );
  NAND2_X1 U3857 ( .A1(n6809), .A2(n4727), .ZN(n5024) );
  INV_X1 U3858 ( .A(n6512), .ZN(n6546) );
  INV_X1 U3859 ( .A(n6617), .ZN(n6605) );
  AND2_X1 U3860 ( .A1(n4873), .A2(n5259), .ZN(n5932) );
  AND2_X1 U3861 ( .A1(n4958), .A2(n4960), .ZN(n6635) );
  OR2_X1 U3862 ( .A1(n6652), .A2(n4960), .ZN(n4839) );
  INV_X1 U3863 ( .A(n4960), .ZN(n5258) );
  INV_X1 U3864 ( .A(n6679), .ZN(n6681) );
  NOR2_X1 U3865 ( .A1(n4826), .A2(n5259), .ZN(n5227) );
  NAND2_X1 U3866 ( .A1(n4594), .A2(n4589), .ZN(n6936) );
  INV_X1 U3867 ( .A(n6234), .ZN(n6170) );
  INV_X1 U3868 ( .A(n6235), .ZN(n6203) );
  AND2_X1 U3869 ( .A1(n5304), .A2(n6128), .ZN(n6243) );
  OR2_X1 U3870 ( .A1(n5600), .A2(n5610), .ZN(n5959) );
  OR2_X1 U3871 ( .A1(n5651), .A2(n5650), .ZN(n5999) );
  OR2_X1 U3872 ( .A1(n6323), .A2(n6932), .ZN(n6327) );
  OR2_X1 U3873 ( .A1(n5603), .A2(n5602), .ZN(n6021) );
  OR2_X1 U3874 ( .A1(n5643), .A2(n5642), .ZN(n6032) );
  AND2_X1 U3875 ( .A1(n4271), .A2(n4270), .ZN(n4272) );
  AND2_X1 U3876 ( .A1(n3767), .A2(n3766), .ZN(n6442) );
  INV_X1 U3877 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6764) );
  INV_X1 U3878 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U3879 ( .A1(n3097), .A2(n6551), .ZN(n6617) );
  INV_X1 U3880 ( .A(n5932), .ZN(n5373) );
  INV_X1 U3881 ( .A(n6635), .ZN(n6649) );
  OR2_X1 U3882 ( .A1(n4839), .A2(n5259), .ZN(n5116) );
  OR3_X1 U3883 ( .A1(n6652), .A2(n5258), .A3(n6551), .ZN(n6679) );
  OR2_X1 U3884 ( .A1(n4826), .A2(n6551), .ZN(n5120) );
  OR2_X1 U3885 ( .A1(n6694), .A2(n5259), .ZN(n6753) );
  OAI21_X1 U3886 ( .B1(n5478), .B2(n6476), .A(n3778), .ZN(U2988) );
  AND2_X2 U3887 ( .A1(n3111), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3119)
         );
  NAND2_X1 U3888 ( .A1(n3365), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3110) );
  NOR2_X4 U3889 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U3890 ( .A1(n3296), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3109) );
  INV_X1 U3891 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3798) );
  AND2_X2 U3892 ( .A1(n3798), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3118)
         );
  AND2_X2 U3893 ( .A1(n3118), .A2(n4788), .ZN(n3217) );
  NAND2_X1 U3894 ( .A1(n3217), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3108)
         );
  NAND2_X1 U3896 ( .A1(n3218), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3897 ( .A1(n3366), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3117) );
  INV_X1 U3898 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3111) );
  NOR2_X2 U3899 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3111), .ZN(n3124)
         );
  NAND2_X1 U3900 ( .A1(n3364), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3116) );
  AND2_X2 U3901 ( .A1(n3118), .A2(n3125), .ZN(n3446) );
  NAND2_X1 U3902 ( .A1(n5427), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3115) );
  NOR2_X2 U3903 ( .A1(n3113), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4615)
         );
  NAND2_X1 U3904 ( .A1(n3397), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3114)
         );
  NAND2_X1 U3905 ( .A1(n3302), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3123)
         );
  NAND2_X1 U3906 ( .A1(n3303), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U3907 ( .A1(n3304), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3121)
         );
  AND2_X2 U3908 ( .A1(n3125), .A2(n4760), .ZN(n4127) );
  NAND2_X1 U3909 ( .A1(n4127), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3120) );
  NAND2_X1 U3910 ( .A1(n3425), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3129) );
  AND2_X2 U3911 ( .A1(n4615), .A2(n3125), .ZN(n4159) );
  NAND2_X1 U3912 ( .A1(n3089), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U3913 ( .A1(n4243), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3127)
         );
  NAND2_X1 U3914 ( .A1(n3297), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3126)
         );
  NAND4_X4 U3915 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3579)
         );
  INV_X2 U3916 ( .A(n3579), .ZN(n3614) );
  AOI22_X1 U3917 ( .A1(n3365), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U3918 ( .A1(n3425), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U3919 ( .A1(n4159), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U3920 ( .A1(n3296), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3134) );
  NAND4_X1 U3921 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3143)
         );
  AOI22_X1 U3922 ( .A1(n3364), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U3923 ( .A1(n3303), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U3924 ( .A1(n3366), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3139) );
  BUF_X2 U3925 ( .A(n3446), .Z(n4238) );
  AOI22_X1 U3926 ( .A1(n4238), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3138) );
  NAND4_X1 U3927 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3142)
         );
  OR2_X2 U3928 ( .A1(n3143), .A2(n3142), .ZN(n3787) );
  NAND2_X1 U3929 ( .A1(n3614), .A2(n3787), .ZN(n4679) );
  AOI22_X1 U3930 ( .A1(n3364), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U3931 ( .A1(n3303), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U3932 ( .A1(n3366), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U3933 ( .A1(n5427), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U3934 ( .A1(n3365), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U3935 ( .A1(n3425), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U3936 ( .A1(n4159), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U3937 ( .A1(n3296), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3148) );
  AND2_X2 U3938 ( .A1(n3101), .A2(n3103), .ZN(n4948) );
  NAND2_X1 U3939 ( .A1(n4679), .A2(n4948), .ZN(n3225) );
  AOI22_X1 U3940 ( .A1(n3217), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4159), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U3941 ( .A1(n3366), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U3942 ( .A1(n3425), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U3943 ( .A1(n4238), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3153) );
  NAND4_X1 U3944 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3162)
         );
  AOI22_X1 U3945 ( .A1(n3303), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U3946 ( .A1(n3364), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U3947 ( .A1(n3365), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U3948 ( .A1(n3296), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3157) );
  NAND4_X1 U3949 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3161)
         );
  OR2_X2 U3950 ( .A1(n3225), .A2(n5682), .ZN(n3615) );
  NAND2_X1 U3951 ( .A1(n3364), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U3952 ( .A1(n3304), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3165)
         );
  NAND2_X1 U3953 ( .A1(n3366), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U3954 ( .A1(n3397), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3163)
         );
  NAND2_X1 U3955 ( .A1(n3303), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U3956 ( .A1(n3302), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3169)
         );
  NAND2_X1 U3957 ( .A1(n5427), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U3958 ( .A1(n4127), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U3959 ( .A1(n3365), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3174) );
  NAND2_X1 U3960 ( .A1(n3425), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U3961 ( .A1(n3217), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3172)
         );
  NAND2_X1 U3962 ( .A1(n3218), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U3963 ( .A1(n3089), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U3964 ( .A1(n3296), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U3965 ( .A1(n4243), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3176)
         );
  NAND2_X1 U3966 ( .A1(n3297), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3175)
         );
  NAND4_X4 U3967 ( .A1(n3182), .A2(n3181), .A3(n3180), .A4(n3179), .ZN(n3628)
         );
  NAND2_X1 U3968 ( .A1(n3425), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U3969 ( .A1(n3296), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U3970 ( .A1(n3365), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U3971 ( .A1(n3218), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U3972 ( .A1(n3364), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U3973 ( .A1(n3304), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3189)
         );
  NAND2_X1 U3974 ( .A1(n3302), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3188)
         );
  NAND2_X1 U3975 ( .A1(n3397), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3187)
         );
  NAND2_X1 U3976 ( .A1(n3303), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U3977 ( .A1(n3366), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U3978 ( .A1(n5427), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U3979 ( .A1(n4127), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3191) );
  AND4_X2 U3980 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3200)
         );
  NAND2_X1 U3981 ( .A1(n3217), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U3982 ( .A1(n3089), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U3983 ( .A1(n4243), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U3984 ( .A1(n3297), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3195)
         );
  NAND4_X4 U3985 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n5184)
         );
  AOI22_X1 U3986 ( .A1(n3365), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U3987 ( .A1(n3304), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U3988 ( .A1(n3303), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U3989 ( .A1(n4238), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3203) );
  NAND4_X1 U3990 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3212)
         );
  AOI22_X1 U3991 ( .A1(n3302), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U3992 ( .A1(n3425), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U3993 ( .A1(n3089), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U3994 ( .A1(n3366), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3207) );
  NAND4_X1 U3995 ( .A1(n3210), .A2(n3209), .A3(n3208), .A4(n3207), .ZN(n3211)
         );
  OR2_X2 U3996 ( .A1(n3212), .A2(n3211), .ZN(n3319) );
  AOI22_X1 U3997 ( .A1(n3366), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U3998 ( .A1(n3303), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U3999 ( .A1(n3364), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4000 ( .A1(n4238), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3213) );
  NAND4_X1 U4001 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3224)
         );
  AOI22_X1 U4002 ( .A1(n3365), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4003 ( .A1(n3425), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4004 ( .A1(n4159), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4005 ( .A1(n3296), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3219) );
  NAND4_X1 U4006 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3223)
         );
  OR2_X2 U4007 ( .A1(n3224), .A2(n3223), .ZN(n3968) );
  NAND2_X1 U4008 ( .A1(n3225), .A2(n3968), .ZN(n3229) );
  NAND2_X1 U4009 ( .A1(n4939), .A2(n3579), .ZN(n3340) );
  NAND2_X1 U4010 ( .A1(n3340), .A2(n4737), .ZN(n3226) );
  INV_X2 U4011 ( .A(n3787), .ZN(n4934) );
  NAND2_X1 U4012 ( .A1(n3226), .A2(n4705), .ZN(n3228) );
  NAND2_X1 U4013 ( .A1(n4948), .A2(n4934), .ZN(n3314) );
  NAND3_X1 U4014 ( .A1(n3229), .A2(n3228), .A3(n3227), .ZN(n3317) );
  NOR2_X1 U4015 ( .A1(n3628), .A2(n5184), .ZN(n3320) );
  NAND2_X1 U4016 ( .A1(n3317), .A2(n5303), .ZN(n3745) );
  OAI211_X1 U4017 ( .C1(n3230), .C2(n6788), .A(n4619), .B(n3745), .ZN(n3242)
         );
  INV_X1 U4018 ( .A(n4705), .ZN(n3231) );
  AND2_X1 U4019 ( .A1(n4679), .A2(n5686), .ZN(n3232) );
  AND2_X2 U4020 ( .A1(n3233), .A2(n3232), .ZN(n3316) );
  NAND2_X1 U4021 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6830) );
  OAI21_X1 U4022 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6830), .ZN(n3546) );
  INV_X1 U4023 ( .A(n3546), .ZN(n3234) );
  NOR2_X1 U4024 ( .A1(n3628), .A2(n3234), .ZN(n3322) );
  INV_X1 U4025 ( .A(n3735), .ZN(n3235) );
  OAI211_X1 U4026 ( .C1(n3322), .C2(n3579), .A(n3235), .B(n3244), .ZN(n3236)
         );
  INV_X1 U4027 ( .A(n3236), .ZN(n3237) );
  NAND2_X1 U4028 ( .A1(n4705), .A2(n4699), .ZN(n3243) );
  NAND3_X1 U4029 ( .A1(n3618), .A2(n3237), .A3(n3243), .ZN(n3238) );
  OAI21_X1 U4030 ( .B1(n3242), .B2(n3238), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3239) );
  INV_X1 U4031 ( .A(n3239), .ZN(n3390) );
  NAND2_X1 U4032 ( .A1(n3390), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3241) );
  AND2_X1 U4033 ( .A1(n6912), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3623) );
  NOR2_X1 U4034 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6906) );
  NAND2_X1 U4035 ( .A1(n6906), .A2(n6809), .ZN(n6933) );
  MUX2_X1 U4036 ( .A(n3623), .B(n6933), .S(n6759), .Z(n3240) );
  INV_X1 U4037 ( .A(n3242), .ZN(n3250) );
  NAND3_X1 U4038 ( .A1(n3618), .A2(n3319), .A3(n3243), .ZN(n3248) );
  NAND2_X1 U4039 ( .A1(n4934), .A2(n5686), .ZN(n3794) );
  NAND2_X1 U4040 ( .A1(n6756), .A2(n5303), .ZN(n3247) );
  NAND2_X1 U4041 ( .A1(n5310), .A2(n3626), .ZN(n3739) );
  NAND2_X1 U4042 ( .A1(n3968), .A2(n5184), .ZN(n3245) );
  NAND4_X1 U4043 ( .A1(n3739), .A2(n6906), .A3(STATE2_REG_0__SCAN_IN), .A4(
        n3245), .ZN(n3246) );
  AOI21_X1 U4044 ( .B1(n3248), .B2(n3247), .A(n3246), .ZN(n3249) );
  INV_X1 U4046 ( .A(n3365), .ZN(n3261) );
  AOI22_X1 U4047 ( .A1(n3425), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3084), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4048 ( .A1(n5436), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3253) );
  BUF_X1 U4049 ( .A(n3302), .Z(n3266) );
  AOI22_X1 U4050 ( .A1(n3266), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4052 ( .A1(n3303), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3251) );
  NAND4_X1 U4053 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3260)
         );
  AOI22_X1 U4054 ( .A1(n4217), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4055 ( .A1(n5445), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4056 ( .A1(n4159), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4057 ( .A1(n5437), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3255) );
  NAND4_X1 U4058 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3259)
         );
  INV_X1 U4059 ( .A(n3508), .ZN(n3278) );
  AOI22_X1 U4060 ( .A1(n3084), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4061 ( .A1(n3364), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4062 ( .A1(n5438), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4063 ( .A1(n3088), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3262) );
  NAND4_X1 U4064 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3272)
         );
  AOI22_X1 U4065 ( .A1(n4159), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4066 ( .A1(n4217), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4067 ( .A1(n3295), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4068 ( .A1(n3266), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3267) );
  NAND4_X1 U4069 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3271)
         );
  XNOR2_X1 U4070 ( .A(n3278), .B(n3382), .ZN(n3273) );
  INV_X1 U4071 ( .A(n3363), .ZN(n3335) );
  NAND2_X1 U4072 ( .A1(n3273), .A2(n3335), .ZN(n3280) );
  INV_X1 U4073 ( .A(n3293), .ZN(n3279) );
  NAND2_X1 U4074 ( .A1(n3597), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3277) );
  INV_X1 U4075 ( .A(n3576), .ZN(n3275) );
  OAI21_X1 U4076 ( .B1(n6809), .B2(n3382), .A(n3275), .ZN(n3276) );
  OAI211_X1 U4077 ( .C1(n3278), .C2(n4699), .A(n3277), .B(n3276), .ZN(n3292)
         );
  INV_X1 U4078 ( .A(n3280), .ZN(n3282) );
  NAND2_X2 U4079 ( .A1(n3284), .A2(n3283), .ZN(n5259) );
  NAND2_X1 U4080 ( .A1(n5259), .A2(n3569), .ZN(n3288) );
  AND2_X1 U4081 ( .A1(n4744), .A2(n3319), .ZN(n3385) );
  INV_X1 U4082 ( .A(n3385), .ZN(n3285) );
  OAI21_X1 U4083 ( .B1(n6788), .B2(n3382), .A(n3285), .ZN(n3286) );
  INV_X1 U4084 ( .A(n3286), .ZN(n3287) );
  NAND2_X1 U4085 ( .A1(n3288), .A2(n3287), .ZN(n4605) );
  NAND2_X1 U4086 ( .A1(n4605), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3289)
         );
  INV_X1 U4087 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U4088 ( .A1(n3289), .A2(n6501), .ZN(n3291) );
  AND2_X1 U4089 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4090 ( .A1(n4605), .A2(n3290), .ZN(n3344) );
  NAND2_X1 U4091 ( .A1(n3335), .A2(n3508), .ZN(n3504) );
  NAND2_X1 U4092 ( .A1(n3597), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3313) );
  INV_X1 U4093 ( .A(n3362), .ZN(n3311) );
  AOI22_X1 U4094 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3295), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4095 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n3084), .B1(n4159), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4096 ( .A1(n4217), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4097 ( .A1(n5448), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4098 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3310)
         );
  AOI22_X1 U4099 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3266), .B1(n5438), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4100 ( .A1(n5436), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4101 ( .A1(n3086), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4102 ( .A1(n4238), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3305) );
  NAND4_X1 U4103 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3309)
         );
  OR2_X1 U4104 ( .A1(n3310), .A2(n3309), .ZN(n3383) );
  NAND2_X1 U4105 ( .A1(n3311), .A2(n3383), .ZN(n3312) );
  OAI211_X1 U4106 ( .C1(n3363), .C2(n3508), .A(n3313), .B(n3312), .ZN(n3347)
         );
  NOR2_X1 U4107 ( .A1(n3314), .A2(n3735), .ZN(n3315) );
  NAND2_X1 U4108 ( .A1(n3316), .A2(n3315), .ZN(n4621) );
  INV_X2 U4109 ( .A(n4621), .ZN(n6790) );
  NAND2_X2 U4110 ( .A1(n3318), .A2(n3094), .ZN(n4571) );
  INV_X2 U4111 ( .A(n4571), .ZN(n4579) );
  NAND2_X2 U4112 ( .A1(n4579), .A2(n4728), .ZN(n4636) );
  NOR2_X1 U4113 ( .A1(n3968), .A2(n3319), .ZN(n4696) );
  INV_X1 U4114 ( .A(n3320), .ZN(n4698) );
  NAND2_X1 U4115 ( .A1(n3787), .A2(n5686), .ZN(n5683) );
  OAI211_X1 U4116 ( .C1(n4587), .C2(n3322), .A(n4636), .B(n3632), .ZN(n3323)
         );
  NAND2_X1 U4117 ( .A1(n3323), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3329) );
  INV_X1 U4118 ( .A(n3329), .ZN(n3327) );
  XNOR2_X1 U4119 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5022) );
  OR2_X1 U4120 ( .A1(n5022), .A2(n6933), .ZN(n3325) );
  INV_X1 U4121 ( .A(n3623), .ZN(n3393) );
  NAND2_X1 U4122 ( .A1(n3393), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3324) );
  AND2_X1 U4123 ( .A1(n3325), .A2(n3324), .ZN(n3330) );
  INV_X1 U4124 ( .A(n3330), .ZN(n3326) );
  INV_X1 U4125 ( .A(n3390), .ZN(n3358) );
  OAI211_X1 U4126 ( .C1(n3358), .C2(n3328), .A(n3330), .B(n3329), .ZN(n3351)
         );
  NAND2_X1 U4127 ( .A1(n3352), .A2(n3351), .ZN(n3334) );
  INV_X1 U4128 ( .A(n3331), .ZN(n3332) );
  XNOR2_X1 U4129 ( .A(n3334), .B(n3106), .ZN(n4617) );
  NAND2_X1 U4130 ( .A1(n4617), .A2(n6809), .ZN(n3337) );
  NAND2_X1 U4131 ( .A1(n3335), .A2(n3383), .ZN(n3336) );
  NAND2_X1 U4132 ( .A1(n3337), .A2(n3336), .ZN(n3346) );
  XNOR2_X1 U4133 ( .A(n3338), .B(n3346), .ZN(n4718) );
  NAND2_X1 U4134 ( .A1(n4718), .A2(n3569), .ZN(n3343) );
  INV_X1 U4135 ( .A(n3382), .ZN(n3339) );
  XNOR2_X1 U4136 ( .A(n3339), .B(n3383), .ZN(n3341) );
  INV_X1 U4137 ( .A(n6788), .ZN(n4596) );
  AOI21_X1 U4138 ( .B1(n3341), .B2(n4596), .A(n3340), .ZN(n3342) );
  NAND2_X1 U4139 ( .A1(n3343), .A2(n3342), .ZN(n4647) );
  NAND2_X1 U4140 ( .A1(n4648), .A2(n4647), .ZN(n3345) );
  OAI21_X1 U4141 ( .B1(n3348), .B2(n3347), .A(n3346), .ZN(n3350) );
  NAND2_X1 U4142 ( .A1(n3348), .A2(n3347), .ZN(n3349) );
  NAND2_X1 U4143 ( .A1(n3350), .A2(n3349), .ZN(n3381) );
  INV_X1 U4144 ( .A(n3381), .ZN(n3379) );
  NAND2_X1 U4145 ( .A1(n3106), .A2(n3351), .ZN(n3353) );
  NAND2_X1 U4146 ( .A1(n3353), .A2(n3352), .ZN(n3360) );
  INV_X1 U4147 ( .A(n6933), .ZN(n3394) );
  AND2_X1 U4148 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4149 ( .A1(n3354), .A2(n6770), .ZN(n6650) );
  INV_X1 U4150 ( .A(n3354), .ZN(n3355) );
  NAND2_X1 U4151 ( .A1(n3355), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4152 ( .A1(n6650), .A2(n3356), .ZN(n5347) );
  AOI22_X1 U4153 ( .A1(n3394), .A2(n5347), .B1(n3393), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3357) );
  BUF_X1 U4155 ( .A(n3364), .Z(n5437) );
  AOI22_X1 U4156 ( .A1(n5437), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3084), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4157 ( .A1(n4217), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4158 ( .A1(n5438), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4159 ( .A1(n3295), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3367) );
  NAND4_X1 U4160 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3376)
         );
  AOI22_X1 U4161 ( .A1(n5436), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4162 ( .A1(n5445), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4163 ( .A1(n3266), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4164 ( .A1(n3152), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4165 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3375)
         );
  OR2_X1 U4166 ( .A1(n3376), .A2(n3375), .ZN(n3384) );
  AOI22_X1 U4167 ( .A1(n3597), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3603), 
        .B2(n3384), .ZN(n3377) );
  INV_X1 U4168 ( .A(n3380), .ZN(n3378) );
  NAND2_X2 U4169 ( .A1(n3381), .A2(n3380), .ZN(n3786) );
  NAND3_X1 U4170 ( .A1(n3785), .A2(n3569), .A3(n3786), .ZN(n3388) );
  NAND2_X1 U4171 ( .A1(n3383), .A2(n3382), .ZN(n3411) );
  INV_X1 U4172 ( .A(n3384), .ZN(n3410) );
  XNOR2_X1 U4173 ( .A(n3411), .B(n3410), .ZN(n3386) );
  AOI21_X1 U4174 ( .B1(n3386), .B2(n4596), .A(n3385), .ZN(n3387) );
  NAND2_X1 U4175 ( .A1(n3388), .A2(n3387), .ZN(n6426) );
  AND2_X1 U4176 ( .A1(n6426), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3389)
         );
  OAI22_X1 U4177 ( .A1(n6427), .A2(n3389), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6426), .ZN(n6418) );
  INV_X1 U4178 ( .A(n6418), .ZN(n3417) );
  NAND3_X1 U4179 ( .A1(n6777), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5345) );
  INV_X1 U4180 ( .A(n5345), .ZN(n3391) );
  NAND2_X1 U4181 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3391), .ZN(n4957) );
  NAND2_X1 U4182 ( .A1(n6777), .A2(n4957), .ZN(n3392) );
  NAND3_X1 U4183 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6691) );
  INV_X1 U4184 ( .A(n6691), .ZN(n6702) );
  NAND2_X1 U4185 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6702), .ZN(n6688) );
  AND2_X1 U4186 ( .A1(n3392), .A2(n6688), .ZN(n5023) );
  AOI22_X1 U4187 ( .A1(n3394), .A2(n5023), .B1(n3393), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4188 ( .A1(n3364), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4189 ( .A1(n5438), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3400) );
  BUF_X8 U4190 ( .A(n3397), .Z(n5439) );
  AOI22_X1 U4191 ( .A1(n4217), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4192 ( .A1(n4238), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3398) );
  NAND4_X1 U4193 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3407)
         );
  INV_X1 U4194 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U4195 ( .A1(n3084), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4196 ( .A1(n3295), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4197 ( .A1(n3152), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4198 ( .A1(n5448), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4199 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3406)
         );
  OR2_X1 U4200 ( .A1(n3407), .A2(n3406), .ZN(n3434) );
  AOI22_X1 U4201 ( .A1(n3597), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3603), 
        .B2(n3434), .ZN(n3408) );
  NAND2_X1 U4202 ( .A1(n3818), .A2(n3569), .ZN(n3415) );
  NAND2_X1 U4203 ( .A1(n3411), .A2(n3410), .ZN(n3435) );
  INV_X1 U4204 ( .A(n3434), .ZN(n3412) );
  XNOR2_X1 U4205 ( .A(n3435), .B(n3412), .ZN(n3413) );
  NAND2_X1 U4206 ( .A1(n3413), .A2(n4596), .ZN(n3414) );
  NAND2_X1 U4207 ( .A1(n3415), .A2(n3414), .ZN(n3418) );
  XNOR2_X1 U4208 ( .A(n3418), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6419)
         );
  INV_X1 U4209 ( .A(n6419), .ZN(n3416) );
  NAND2_X1 U4210 ( .A1(n3417), .A2(n3416), .ZN(n6416) );
  NAND2_X1 U4211 ( .A1(n3418), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3419)
         );
  NAND2_X1 U4212 ( .A1(n6416), .A2(n3419), .ZN(n4982) );
  INV_X1 U4213 ( .A(n3786), .ZN(n3420) );
  NAND2_X1 U4214 ( .A1(n3420), .A2(n4819), .ZN(n3466) );
  NAND2_X1 U4215 ( .A1(n3597), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4216 ( .A1(n5437), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4217 ( .A1(n5438), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4218 ( .A1(n4217), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4219 ( .A1(n4238), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4220 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3431)
         );
  AOI22_X1 U4221 ( .A1(n3084), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4222 ( .A1(n3295), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4223 ( .A1(n3152), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4224 ( .A1(n5448), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4225 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3430)
         );
  OR2_X1 U4226 ( .A1(n3431), .A2(n3430), .ZN(n3456) );
  NAND2_X1 U4227 ( .A1(n3603), .A2(n3456), .ZN(n3432) );
  NAND2_X1 U4228 ( .A1(n3433), .A2(n3432), .ZN(n3464) );
  XNOR2_X1 U4229 ( .A(n3466), .B(n3464), .ZN(n3809) );
  NAND2_X1 U4230 ( .A1(n3809), .A2(n3569), .ZN(n3438) );
  NAND2_X1 U4231 ( .A1(n3435), .A2(n3434), .ZN(n3458) );
  XNOR2_X1 U4232 ( .A(n3458), .B(n3456), .ZN(n3436) );
  NAND2_X1 U4233 ( .A1(n3436), .A2(n4596), .ZN(n3437) );
  INV_X1 U4234 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U4235 ( .A1(n4982), .A2(n4981), .ZN(n4980) );
  NAND2_X1 U4236 ( .A1(n3439), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3440)
         );
  NAND2_X1 U4237 ( .A1(n4980), .A2(n3440), .ZN(n4561) );
  INV_X1 U4238 ( .A(n3466), .ZN(n3441) );
  NAND2_X1 U4239 ( .A1(n3597), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4240 ( .A1(n3084), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4241 ( .A1(n5437), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4242 ( .A1(n4217), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4243 ( .A1(n3295), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4244 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3452)
         );
  AOI22_X1 U4245 ( .A1(n3266), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4246 ( .A1(n4105), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4247 ( .A1(n5438), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3448) );
  INV_X1 U4248 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U4249 ( .A1(n5448), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4250 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3451)
         );
  OR2_X1 U4251 ( .A1(n3452), .A2(n3451), .ZN(n3484) );
  NAND2_X1 U4252 ( .A1(n3603), .A2(n3484), .ZN(n3453) );
  NAND2_X1 U4253 ( .A1(n3454), .A2(n3453), .ZN(n3463) );
  NAND2_X1 U4254 ( .A1(n3828), .A2(n3569), .ZN(n3461) );
  INV_X1 U4255 ( .A(n3456), .ZN(n3457) );
  OR2_X1 U4256 ( .A1(n3458), .A2(n3457), .ZN(n3483) );
  XNOR2_X1 U4257 ( .A(n3483), .B(n3484), .ZN(n3459) );
  NAND2_X1 U4258 ( .A1(n3459), .A2(n4596), .ZN(n3460) );
  NAND2_X1 U4259 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  INV_X1 U4260 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4558) );
  XNOR2_X1 U4261 ( .A(n3462), .B(n4558), .ZN(n4560) );
  NAND2_X1 U4262 ( .A1(n4561), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U4263 ( .A1(n3462), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4988)
         );
  NAND2_X1 U4264 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  NOR2_X2 U4265 ( .A1(n3466), .A2(n3465), .ZN(n3482) );
  INV_X1 U4266 ( .A(n3482), .ZN(n3480) );
  NAND2_X1 U4267 ( .A1(n3597), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4268 ( .A1(n5437), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4269 ( .A1(n5438), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4270 ( .A1(n4217), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4271 ( .A1(n4105), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3467) );
  NAND4_X1 U4272 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3476)
         );
  AOI22_X1 U4273 ( .A1(n3084), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4274 ( .A1(n3295), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4275 ( .A1(n3152), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4276 ( .A1(n5448), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3471) );
  NAND4_X1 U4277 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3475)
         );
  OR2_X1 U4278 ( .A1(n3476), .A2(n3475), .ZN(n3496) );
  NAND2_X1 U4279 ( .A1(n3603), .A2(n3496), .ZN(n3477) );
  NAND2_X1 U4280 ( .A1(n3478), .A2(n3477), .ZN(n3481) );
  INV_X1 U4281 ( .A(n3481), .ZN(n3479) );
  NAND2_X1 U4282 ( .A1(n3480), .A2(n3479), .ZN(n3836) );
  NAND3_X1 U4283 ( .A1(n3836), .A2(n3506), .A3(n3569), .ZN(n3488) );
  INV_X1 U4284 ( .A(n3483), .ZN(n3485) );
  NAND2_X1 U4285 ( .A1(n3485), .A2(n3484), .ZN(n3495) );
  XNOR2_X1 U4286 ( .A(n3495), .B(n3496), .ZN(n3486) );
  NAND2_X1 U4287 ( .A1(n3486), .A2(n4596), .ZN(n3487) );
  NAND2_X1 U4288 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  NAND2_X1 U4289 ( .A1(n3489), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3490)
         );
  AND2_X1 U4290 ( .A1(n4988), .A2(n3490), .ZN(n3493) );
  INV_X1 U4291 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6473) );
  XNOR2_X1 U4292 ( .A(n3489), .B(n6473), .ZN(n4991) );
  INV_X1 U4293 ( .A(n3490), .ZN(n3491) );
  AOI21_X2 U4294 ( .B1(n4559), .B2(n3493), .A(n3492), .ZN(n6403) );
  AOI22_X1 U4295 ( .A1(n3597), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3603), 
        .B2(n3508), .ZN(n3494) );
  XNOR2_X1 U4296 ( .A(n3506), .B(n3494), .ZN(n3840) );
  INV_X1 U4297 ( .A(n3569), .ZN(n3503) );
  OR2_X1 U4298 ( .A1(n3840), .A2(n3503), .ZN(n3500) );
  INV_X1 U4299 ( .A(n3495), .ZN(n3497) );
  NAND2_X1 U4300 ( .A1(n3497), .A2(n3496), .ZN(n3507) );
  XNOR2_X1 U4301 ( .A(n3507), .B(n3508), .ZN(n3498) );
  NAND2_X1 U4302 ( .A1(n3498), .A2(n4596), .ZN(n3499) );
  NAND2_X1 U4303 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  INV_X1 U4304 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6466) );
  XNOR2_X1 U4305 ( .A(n3501), .B(n6466), .ZN(n6402) );
  NAND2_X1 U4306 ( .A1(n6403), .A2(n6402), .ZN(n6401) );
  NAND2_X1 U4307 ( .A1(n3501), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3502)
         );
  NAND2_X1 U4308 ( .A1(n6401), .A2(n3502), .ZN(n5003) );
  NOR2_X1 U4309 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  NAND2_X2 U4310 ( .A1(n3506), .A2(n3505), .ZN(n4289) );
  INV_X1 U4311 ( .A(n3507), .ZN(n3509) );
  NAND3_X1 U4312 ( .A1(n3509), .A2(n4596), .A3(n3508), .ZN(n3510) );
  NAND2_X1 U4313 ( .A1(n4289), .A2(n3510), .ZN(n3511) );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6458) );
  XNOR2_X1 U4315 ( .A(n3511), .B(n6458), .ZN(n5002) );
  NAND2_X1 U4316 ( .A1(n5003), .A2(n5002), .ZN(n5001) );
  NAND2_X1 U4317 ( .A1(n3511), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3512)
         );
  NAND2_X1 U4318 ( .A1(n5001), .A2(n3512), .ZN(n6395) );
  INV_X4 U4319 ( .A(n3513), .ZN(n5795) );
  XNOR2_X1 U4320 ( .A(n5795), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6394)
         );
  NAND2_X1 U4321 ( .A1(n6395), .A2(n6394), .ZN(n6393) );
  INV_X1 U4322 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6449) );
  OR2_X1 U4323 ( .A1(n5795), .A2(n6449), .ZN(n3514) );
  NAND2_X1 U4324 ( .A1(n6393), .A2(n3514), .ZN(n5193) );
  INV_X1 U4325 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4326 ( .A1(n4289), .A2(n3669), .ZN(n5194) );
  NAND2_X1 U4327 ( .A1(n5193), .A2(n5194), .ZN(n5320) );
  INV_X1 U4328 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6441) );
  INV_X1 U4329 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4531) );
  NAND2_X1 U4330 ( .A1(n5795), .A2(n4531), .ZN(n5374) );
  INV_X1 U4331 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4332 ( .A1(n5795), .A2(n3755), .ZN(n5402) );
  XNOR2_X1 U4333 ( .A(n4289), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5811)
         );
  INV_X1 U4334 ( .A(n5811), .ZN(n3516) );
  INV_X1 U4335 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U4336 ( .A1(n4289), .A2(n6072), .ZN(n5804) );
  INV_X1 U4337 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U4338 ( .A1(n4289), .A2(n5903), .ZN(n3518) );
  INV_X1 U4339 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U4340 ( .A1(n5375), .A2(n3517), .ZN(n5788) );
  OR2_X1 U4341 ( .A1(n5795), .A2(n3690), .ZN(n3523) );
  INV_X1 U4342 ( .A(n3518), .ZN(n3522) );
  INV_X1 U4343 ( .A(n3519), .ZN(n3521) );
  XNOR2_X1 U4344 ( .A(n5795), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5403)
         );
  AND2_X1 U4345 ( .A1(n5403), .A2(n5811), .ZN(n3520) );
  INV_X1 U4346 ( .A(n3524), .ZN(n3527) );
  OR2_X1 U4347 ( .A1(n5795), .A2(n4531), .ZN(n5376) );
  XNOR2_X1 U4348 ( .A(n5795), .B(n3755), .ZN(n5400) );
  INV_X1 U4349 ( .A(n5400), .ZN(n3525) );
  AND2_X1 U4350 ( .A1(n5376), .A2(n3525), .ZN(n3526) );
  NAND2_X2 U4351 ( .A1(n5788), .A2(n3530), .ZN(n6042) );
  NOR2_X1 U4352 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3531) );
  NOR2_X1 U4353 ( .A1(n5795), .A2(n3531), .ZN(n5760) );
  NAND2_X1 U4354 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U4355 ( .A1(n4289), .A2(n5876), .ZN(n3532) );
  OAI21_X2 U4356 ( .B1(n6042), .B2(n5760), .A(n3532), .ZN(n4290) );
  INV_X1 U4357 ( .A(n4290), .ZN(n3534) );
  NAND2_X1 U4358 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5853) );
  INV_X1 U4359 ( .A(n5853), .ZN(n3533) );
  NAND2_X1 U4360 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4291) );
  AND2_X1 U4361 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U4362 ( .A1(n3534), .A2(n3099), .ZN(n3535) );
  NAND2_X1 U4363 ( .A1(n3535), .A2(n5795), .ZN(n3538) );
  NOR2_X1 U4365 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5854) );
  NOR2_X1 U4366 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3536) );
  NOR2_X1 U4367 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U4368 ( .A1(n5774), .A2(n3105), .ZN(n3537) );
  NAND2_X1 U4369 ( .A1(n3538), .A2(n3537), .ZN(n5728) );
  XNOR2_X1 U4370 ( .A(n5795), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5727)
         );
  INV_X1 U4371 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U4372 ( .A1(n4289), .A2(n5843), .ZN(n3539) );
  INV_X1 U4373 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4453) );
  INV_X1 U4374 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5821) );
  OAI21_X1 U4375 ( .B1(n4453), .B2(n5821), .A(n5795), .ZN(n3540) );
  INV_X1 U4376 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4269) );
  NOR2_X2 U4377 ( .A1(n4283), .A2(n3541), .ZN(n4285) );
  INV_X1 U4378 ( .A(n4285), .ZN(n5510) );
  NAND2_X1 U4379 ( .A1(n4269), .A2(n5821), .ZN(n4282) );
  NOR3_X1 U4380 ( .A1(n4282), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3542) );
  MUX2_X1 U4381 ( .A(n3542), .B(n4285), .S(n5795), .Z(n3543) );
  OAI21_X1 U4382 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5510), .A(n3543), 
        .ZN(n3545) );
  OR2_X1 U4383 ( .A1(n3546), .A2(STATE_REG_0__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U4384 ( .A1(n3628), .A2(n6824), .ZN(n3567) );
  NAND2_X1 U4385 ( .A1(n6764), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4386 ( .A1(n3328), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3547) );
  NAND2_X1 U4387 ( .A1(n3548), .A2(n3547), .ZN(n3558) );
  NAND2_X1 U4388 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6759), .ZN(n3574) );
  NAND2_X1 U4389 ( .A1(n3560), .A2(n3548), .ZN(n3557) );
  NAND2_X1 U4390 ( .A1(n6770), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4391 ( .A1(n5505), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3549) );
  AND2_X1 U4392 ( .A1(n3550), .A2(n3549), .ZN(n3555) );
  NAND2_X1 U4393 ( .A1(n3557), .A2(n3555), .ZN(n3551) );
  NAND2_X1 U4394 ( .A1(n3551), .A2(n3550), .ZN(n3562) );
  OR2_X1 U4395 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6777), .ZN(n3553)
         );
  NOR2_X1 U4396 ( .A1(n4771), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3552)
         );
  AOI21_X1 U4397 ( .B1(n3562), .B2(n3553), .A(n3552), .ZN(n3565) );
  INV_X1 U4398 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U4399 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6774), .ZN(n3554) );
  INV_X1 U4400 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3812) );
  AND2_X1 U4401 ( .A1(n3812), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3564)
         );
  AOI21_X1 U4402 ( .B1(n3565), .B2(n3554), .A(n3564), .ZN(n3606) );
  INV_X1 U4403 ( .A(n3555), .ZN(n3556) );
  XNOR2_X1 U4404 ( .A(n3557), .B(n3556), .ZN(n3571) );
  NAND2_X1 U4405 ( .A1(n3558), .A2(n3574), .ZN(n3559) );
  AND2_X1 U4406 ( .A1(n3560), .A2(n3559), .ZN(n3588) );
  XNOR2_X1 U4407 ( .A(n4771), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3561)
         );
  XNOR2_X1 U4408 ( .A(n3562), .B(n3561), .ZN(n3568) );
  AND3_X1 U4409 ( .A1(n3571), .A2(n3588), .A3(n3568), .ZN(n3563) );
  OR2_X1 U4410 ( .A1(n3606), .A2(n3563), .ZN(n3566) );
  NAND2_X1 U4411 ( .A1(n3565), .A2(n3564), .ZN(n3598) );
  AND2_X1 U4412 ( .A1(n3566), .A2(n3598), .ZN(n4578) );
  NOR2_X1 U4413 ( .A1(READY_N), .A2(n4578), .ZN(n4637) );
  NAND2_X1 U4414 ( .A1(n3567), .A2(n4637), .ZN(n3613) );
  INV_X1 U4415 ( .A(n3568), .ZN(n3596) );
  AND2_X1 U4416 ( .A1(n4728), .A2(n3579), .ZN(n3570) );
  NAND2_X1 U4417 ( .A1(n3603), .A2(n3571), .ZN(n3592) );
  AND2_X1 U4418 ( .A1(n3593), .A2(n3592), .ZN(n3573) );
  INV_X1 U4419 ( .A(n3597), .ZN(n3572) );
  OAI22_X1 U4420 ( .A1(n3573), .A2(n3596), .B1(n3572), .B2(n3571), .ZN(n3595)
         );
  OAI21_X1 U4421 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6759), .A(n3574), 
        .ZN(n3581) );
  INV_X1 U4422 ( .A(n3581), .ZN(n3575) );
  NAND2_X1 U4423 ( .A1(n3626), .A2(n3575), .ZN(n3577) );
  NAND2_X1 U4424 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  NAND2_X1 U4425 ( .A1(n3603), .A2(n3628), .ZN(n3580) );
  NAND2_X1 U4426 ( .A1(n3580), .A2(n3579), .ZN(n3589) );
  NOR2_X1 U4427 ( .A1(n3589), .A2(n3588), .ZN(n3583) );
  INV_X1 U4428 ( .A(n3603), .ZN(n3582) );
  NOR4_X1 U4429 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3587)
         );
  INV_X1 U4430 ( .A(n3584), .ZN(n3586) );
  INV_X1 U4431 ( .A(n3588), .ZN(n3585) );
  OAI22_X1 U4432 ( .A1(n3587), .A2(n3607), .B1(n3586), .B2(n3585), .ZN(n3591)
         );
  NAND3_X1 U4433 ( .A1(n3589), .A2(n3588), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3590) );
  OAI211_X1 U4434 ( .C1(n3593), .C2(n3592), .A(n3591), .B(n3590), .ZN(n3594)
         );
  AOI22_X1 U4435 ( .A1(n3596), .A2(n3607), .B1(n3595), .B2(n3594), .ZN(n3601)
         );
  NOR2_X1 U4436 ( .A1(n3597), .A2(n3598), .ZN(n3600) );
  INV_X1 U4437 ( .A(n3607), .ZN(n3599) );
  OAI22_X1 U4438 ( .A1(n3601), .A2(n3600), .B1(n3599), .B2(n3598), .ZN(n3602)
         );
  AOI21_X1 U4439 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6809), .A(n3602), 
        .ZN(n3605) );
  NAND2_X1 U4440 ( .A1(n3606), .A2(n3603), .ZN(n3604) );
  NAND2_X1 U4441 ( .A1(n3605), .A2(n3604), .ZN(n3609) );
  NAND2_X1 U4442 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  INV_X1 U4443 ( .A(n6824), .ZN(n6789) );
  OR2_X1 U4444 ( .A1(n3628), .A2(n6789), .ZN(n5186) );
  INV_X1 U4445 ( .A(READY_N), .ZN(n6827) );
  NAND2_X1 U4446 ( .A1(n5186), .A2(n6827), .ZN(n3610) );
  OAI211_X1 U4447 ( .C1(n4621), .C2(n3610), .A(n5184), .B(n5683), .ZN(n3611)
         );
  NAND2_X1 U4448 ( .A1(n4635), .A2(n3611), .ZN(n3612) );
  MUX2_X1 U4449 ( .A(n3613), .B(n3612), .S(n4939), .Z(n3622) );
  NOR2_X1 U4450 ( .A1(n6756), .A2(n3614), .ZN(n3970) );
  AND2_X1 U4451 ( .A1(n4939), .A2(n3628), .ZN(n4681) );
  NAND2_X1 U4452 ( .A1(n3970), .A2(n4681), .ZN(n3734) );
  NAND2_X1 U4453 ( .A1(n3615), .A2(n5184), .ZN(n3616) );
  MUX2_X1 U4454 ( .A(n6788), .B(n3616), .S(n4705), .Z(n3747) );
  INV_X1 U4455 ( .A(n3970), .ZN(n3617) );
  NAND2_X1 U4456 ( .A1(n3617), .A2(n4744), .ZN(n3620) );
  INV_X1 U4457 ( .A(n3618), .ZN(n3744) );
  NOR2_X1 U4458 ( .A1(n3744), .A2(n3735), .ZN(n3619) );
  AND2_X1 U4459 ( .A1(n3620), .A2(n3619), .ZN(n3625) );
  NAND2_X1 U4460 ( .A1(n3747), .A2(n3625), .ZN(n3621) );
  NAND2_X1 U4461 ( .A1(n3621), .A2(n4571), .ZN(n4632) );
  NAND3_X1 U4462 ( .A1(n3622), .A2(n4641), .A3(n4632), .ZN(n3624) );
  AND2_X1 U4463 ( .A1(n3623), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6802) );
  INV_X1 U4464 ( .A(n3625), .ZN(n3627) );
  OR2_X1 U4465 ( .A1(n3627), .A2(n3626), .ZN(n6778) );
  OR2_X1 U4466 ( .A1(n3627), .A2(n4698), .ZN(n4758) );
  AND2_X1 U4467 ( .A1(n6778), .A2(n4758), .ZN(n4576) );
  NAND2_X1 U4468 ( .A1(n6790), .A2(n5179), .ZN(n4629) );
  INV_X1 U4469 ( .A(n3632), .ZN(n3629) );
  NAND2_X1 U4470 ( .A1(n3629), .A2(n4699), .ZN(n3630) );
  NAND4_X1 U4471 ( .A1(n4576), .A2(n4629), .A3(n4636), .A4(n3630), .ZN(n3631)
         );
  NAND2_X1 U4472 ( .A1(n3761), .A2(n3631), .ZN(n6476) );
  NAND2_X1 U4473 ( .A1(n6790), .A2(n4596), .ZN(n4597) );
  OAI21_X1 U4474 ( .B1(n3632), .B2(n4699), .A(n4597), .ZN(n3633) );
  INV_X1 U4475 ( .A(n5521), .ZN(n3636) );
  INV_X1 U4476 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4318) );
  NOR2_X1 U4477 ( .A1(n5520), .A2(EBX_REG_29__SCAN_IN), .ZN(n3635) );
  AOI21_X1 U4478 ( .B1(n3636), .B2(n4318), .A(n3635), .ZN(n4275) );
  AND2_X2 U4479 ( .A1(n3090), .A2(n5179), .ZN(n3647) );
  INV_X1 U4480 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4481 ( .A1(n3647), .A2(n3637), .ZN(n3641) );
  NAND2_X1 U4482 ( .A1(n3642), .A2(n6501), .ZN(n3639) );
  NAND2_X1 U4483 ( .A1(n5179), .A2(n3637), .ZN(n3638) );
  NAND3_X1 U4484 ( .A1(n3639), .A2(n3634), .A3(n3638), .ZN(n3640) );
  NAND2_X1 U4485 ( .A1(n3642), .A2(EBX_REG_0__SCAN_IN), .ZN(n3644) );
  INV_X1 U4486 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U4487 ( .A1(n3634), .A2(n5588), .ZN(n3643) );
  NAND2_X1 U4488 ( .A1(n3644), .A2(n3643), .ZN(n4672) );
  XNOR2_X1 U4489 ( .A(n3645), .B(n4672), .ZN(n4651) );
  NAND2_X1 U4490 ( .A1(n4651), .A2(n5179), .ZN(n4652) );
  NAND2_X1 U4491 ( .A1(n4652), .A2(n3645), .ZN(n4686) );
  NAND2_X1 U4492 ( .A1(n5179), .A2(n3634), .ZN(n3728) );
  MUX2_X1 U4493 ( .A(n3728), .B(n3634), .S(EBX_REG_3__SCAN_IN), .Z(n3646) );
  OAI21_X1 U4494 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5521), .A(n3646), 
        .ZN(n4687) );
  INV_X1 U4495 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U4496 ( .A1(n3647), .A2(n6260), .ZN(n3651) );
  INV_X1 U4497 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U4498 ( .A1(n3642), .A2(n6507), .ZN(n3649) );
  NAND2_X1 U4499 ( .A1(n5179), .A2(n6260), .ZN(n3648) );
  NAND3_X1 U4500 ( .A1(n3649), .A2(n3634), .A3(n3648), .ZN(n3650) );
  MUX2_X1 U4501 ( .A(n3730), .B(n3642), .S(EBX_REG_4__SCAN_IN), .Z(n3653) );
  NAND2_X1 U4502 ( .A1(n4680), .A2(n5520), .ZN(n3710) );
  NAND2_X1 U4503 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n5520), .ZN(n3652)
         );
  NOR2_X2 U4504 ( .A1(n4714), .A2(n4713), .ZN(n4715) );
  MUX2_X1 U4505 ( .A(n3728), .B(n5659), .S(EBX_REG_5__SCAN_IN), .Z(n3655) );
  OR2_X1 U4506 ( .A1(n5521), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3654)
         );
  NAND2_X1 U4507 ( .A1(n4715), .A2(n4564), .ZN(n4563) );
  INV_X1 U4508 ( .A(n4563), .ZN(n3659) );
  MUX2_X1 U4509 ( .A(n3730), .B(n3642), .S(EBX_REG_6__SCAN_IN), .Z(n3657) );
  NAND2_X1 U4510 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5520), .ZN(n3656)
         );
  NAND2_X1 U4511 ( .A1(n3659), .A2(n3658), .ZN(n4805) );
  INV_X1 U4512 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U4513 ( .A1(n5179), .A2(n6254), .ZN(n3660) );
  OAI211_X1 U4514 ( .C1(n3091), .C2(n6466), .A(n3660), .B(n3642), .ZN(n3661)
         );
  OAI21_X1 U4515 ( .B1(n3728), .B2(EBX_REG_7__SCAN_IN), .A(n3661), .ZN(n6205)
         );
  NOR2_X2 U4516 ( .A1(n4805), .A2(n6205), .ZN(n6204) );
  INV_X1 U4517 ( .A(EBX_REG_8__SCAN_IN), .ZN(n3662) );
  NAND2_X1 U4518 ( .A1(n3647), .A2(n3662), .ZN(n3666) );
  NAND2_X1 U4519 ( .A1(n3642), .A2(n6458), .ZN(n3664) );
  NAND2_X1 U4520 ( .A1(n5179), .A2(n3662), .ZN(n3663) );
  NAND3_X1 U4521 ( .A1(n3664), .A2(n5659), .A3(n3663), .ZN(n3665) );
  NAND2_X1 U4522 ( .A1(n3666), .A2(n3665), .ZN(n4889) );
  AND2_X2 U4523 ( .A1(n6204), .A2(n4889), .ZN(n6195) );
  MUX2_X1 U4524 ( .A(n3728), .B(n5659), .S(EBX_REG_9__SCAN_IN), .Z(n3667) );
  OAI21_X1 U4525 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5521), .A(n3667), 
        .ZN(n6198) );
  INV_X1 U4526 ( .A(n6198), .ZN(n3668) );
  NAND2_X1 U4527 ( .A1(n6195), .A2(n3668), .ZN(n5017) );
  INV_X1 U4528 ( .A(EBX_REG_10__SCAN_IN), .ZN(n3670) );
  NAND2_X1 U4529 ( .A1(n3647), .A2(n3670), .ZN(n3674) );
  NAND2_X1 U4530 ( .A1(n3642), .A2(n3669), .ZN(n3672) );
  NAND2_X1 U4531 ( .A1(n5179), .A2(n3670), .ZN(n3671) );
  NAND3_X1 U4532 ( .A1(n3672), .A2(n5659), .A3(n3671), .ZN(n3673) );
  AND2_X1 U4533 ( .A1(n3674), .A2(n3673), .ZN(n5019) );
  OR2_X2 U4534 ( .A1(n5017), .A2(n5019), .ZN(n5150) );
  INV_X1 U4535 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U4536 ( .A1(n5179), .A2(n6172), .ZN(n3675) );
  OAI211_X1 U4537 ( .C1(n3091), .C2(n6441), .A(n3675), .B(n3642), .ZN(n3676)
         );
  OAI21_X1 U4538 ( .B1(n3728), .B2(EBX_REG_11__SCAN_IN), .A(n3676), .ZN(n5149)
         );
  NOR2_X4 U4539 ( .A1(n5150), .A2(n5149), .ZN(n5159) );
  INV_X1 U4540 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U4541 ( .A1(n3647), .A2(n6162), .ZN(n3680) );
  NAND2_X1 U4542 ( .A1(n3642), .A2(n4531), .ZN(n3678) );
  NAND2_X1 U4543 ( .A1(n5179), .A2(n6162), .ZN(n3677) );
  NAND3_X1 U4544 ( .A1(n3678), .A2(n5659), .A3(n3677), .ZN(n3679) );
  NAND2_X1 U4545 ( .A1(n3680), .A2(n3679), .ZN(n5158) );
  MUX2_X1 U4546 ( .A(n3730), .B(n3642), .S(EBX_REG_14__SCAN_IN), .Z(n3682) );
  NAND2_X1 U4547 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5520), .ZN(n3681) );
  AND3_X1 U4548 ( .A1(n3682), .A2(n3710), .A3(n3681), .ZN(n5395) );
  INV_X1 U4549 ( .A(n5395), .ZN(n3686) );
  INV_X1 U4550 ( .A(n3728), .ZN(n3713) );
  INV_X1 U4551 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U4552 ( .A1(n3713), .A2(n6250), .ZN(n3685) );
  NAND2_X1 U4553 ( .A1(n5179), .A2(n6250), .ZN(n3683) );
  OAI211_X1 U4554 ( .C1(n3091), .C2(n3755), .A(n3683), .B(n3642), .ZN(n3684)
         );
  AND2_X1 U4555 ( .A1(n3685), .A2(n3684), .ZN(n5382) );
  AND2_X1 U4556 ( .A1(n3686), .A2(n5382), .ZN(n3687) );
  INV_X1 U4557 ( .A(EBX_REG_15__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U4558 ( .A1(n5179), .A2(n4530), .ZN(n3688) );
  OAI211_X1 U4559 ( .C1(n3091), .C2(n5903), .A(n3688), .B(n3642), .ZN(n3689)
         );
  OAI21_X1 U4560 ( .B1(n3728), .B2(EBX_REG_15__SCAN_IN), .A(n3689), .ZN(n5575)
         );
  INV_X1 U4561 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U4562 ( .A1(n3647), .A2(n6134), .ZN(n3694) );
  NAND2_X1 U4563 ( .A1(n3642), .A2(n3690), .ZN(n3692) );
  NAND2_X1 U4564 ( .A1(n5179), .A2(n6134), .ZN(n3691) );
  NAND3_X1 U4565 ( .A1(n3692), .A2(n5659), .A3(n3691), .ZN(n3693) );
  NAND2_X1 U4566 ( .A1(n3694), .A2(n3693), .ZN(n5676) );
  NAND2_X1 U4567 ( .A1(n5573), .A2(n5676), .ZN(n5678) );
  MUX2_X1 U4568 ( .A(n3728), .B(n5659), .S(EBX_REG_17__SCAN_IN), .Z(n3695) );
  OAI21_X1 U4569 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5521), .A(n3695), 
        .ZN(n5667) );
  NOR2_X2 U4570 ( .A1(n5678), .A2(n5667), .ZN(n5658) );
  INV_X1 U4571 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U4572 ( .A1(n3647), .A2(n6017), .ZN(n3699) );
  INV_X1 U4573 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U4574 ( .A1(n3642), .A2(n5761), .ZN(n3697) );
  NAND2_X1 U4575 ( .A1(n5179), .A2(n6017), .ZN(n3696) );
  NAND3_X1 U4576 ( .A1(n3697), .A2(n5659), .A3(n3696), .ZN(n3698) );
  AND2_X1 U4577 ( .A1(n3699), .A2(n3698), .ZN(n5882) );
  NAND2_X1 U4578 ( .A1(n5658), .A2(n3700), .ZN(n5652) );
  OR2_X1 U4579 ( .A1(n5521), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3703)
         );
  INV_X1 U4580 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4581 ( .A1(n5179), .A2(n3701), .ZN(n3702) );
  NAND2_X1 U4582 ( .A1(n3703), .A2(n3702), .ZN(n5654) );
  AND2_X1 U4583 ( .A1(n5520), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3704)
         );
  AOI21_X1 U4584 ( .B1(n5521), .B2(EBX_REG_18__SCAN_IN), .A(n3704), .ZN(n5660)
         );
  MUX2_X1 U4585 ( .A(n5654), .B(n5659), .S(n5660), .Z(n3705) );
  INV_X1 U4586 ( .A(n3705), .ZN(n3707) );
  NAND2_X1 U4587 ( .A1(n3091), .A2(EBX_REG_20__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4588 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  NOR2_X2 U4589 ( .A1(n5652), .A2(n3708), .ZN(n5645) );
  NAND2_X1 U4590 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n5520), .ZN(n3709) );
  AND2_X1 U4591 ( .A1(n3710), .A2(n3709), .ZN(n3712) );
  MUX2_X1 U4592 ( .A(n3730), .B(n3642), .S(EBX_REG_21__SCAN_IN), .Z(n3711) );
  NAND2_X1 U4593 ( .A1(n3712), .A2(n3711), .ZN(n5644) );
  INV_X1 U4594 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U4595 ( .A1(n3713), .A2(n5637), .ZN(n3716) );
  INV_X1 U4596 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U4597 ( .A1(n5179), .A2(n5637), .ZN(n3714) );
  OAI211_X1 U4598 ( .C1(n3091), .C2(n5860), .A(n3714), .B(n3642), .ZN(n3715)
         );
  AND2_X1 U4599 ( .A1(n3716), .A2(n3715), .ZN(n5635) );
  NAND2_X1 U4600 ( .A1(n5647), .A2(n5635), .ZN(n5625) );
  INV_X1 U4601 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U4602 ( .A1(n3647), .A2(n4416), .ZN(n3720) );
  INV_X1 U4603 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U4604 ( .A1(n3642), .A2(n4314), .ZN(n3718) );
  NAND2_X1 U4605 ( .A1(n5179), .A2(n4416), .ZN(n3717) );
  NAND3_X1 U4606 ( .A1(n3718), .A2(n5659), .A3(n3717), .ZN(n3719) );
  AND2_X1 U4607 ( .A1(n3720), .A2(n3719), .ZN(n5628) );
  OR2_X2 U4608 ( .A1(n5625), .A2(n5628), .ZN(n5626) );
  INV_X1 U4609 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4404) );
  INV_X1 U4610 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U4611 ( .A1(n5179), .A2(n5616), .ZN(n3721) );
  OAI211_X1 U4612 ( .C1(n3091), .C2(n4404), .A(n3721), .B(n3642), .ZN(n3722)
         );
  OAI21_X1 U4613 ( .B1(n3728), .B2(EBX_REG_24__SCAN_IN), .A(n3722), .ZN(n4298)
         );
  NOR2_X2 U4614 ( .A1(n5626), .A2(n4298), .ZN(n5556) );
  NAND2_X1 U4615 ( .A1(n5521), .A2(EBX_REG_25__SCAN_IN), .ZN(n3724) );
  NAND2_X1 U4616 ( .A1(n5520), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4617 ( .A1(n3724), .A2(n3723), .ZN(n3725) );
  XNOR2_X1 U4618 ( .A(n3725), .B(n5659), .ZN(n5555) );
  NAND2_X1 U4619 ( .A1(n5556), .A2(n5555), .ZN(n5554) );
  NAND2_X1 U4620 ( .A1(n5520), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3727) );
  MUX2_X1 U4621 ( .A(n3730), .B(n3642), .S(EBX_REG_26__SCAN_IN), .Z(n3726) );
  AND2_X1 U4622 ( .A1(n3727), .A2(n3726), .ZN(n5611) );
  OR2_X2 U4623 ( .A1(n5554), .A2(n5611), .ZN(n5613) );
  MUX2_X1 U4624 ( .A(n3728), .B(n5659), .S(EBX_REG_27__SCAN_IN), .Z(n3729) );
  OAI21_X1 U4625 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5521), .A(n3729), 
        .ZN(n5604) );
  NAND2_X1 U4626 ( .A1(n5520), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3732) );
  MUX2_X1 U4627 ( .A(n3730), .B(n3642), .S(EBX_REG_28__SCAN_IN), .Z(n3731) );
  AND2_X1 U4628 ( .A1(n3732), .A2(n3731), .ZN(n4265) );
  NOR2_X4 U4629 ( .A1(n5606), .A2(n4265), .ZN(n5514) );
  MUX2_X1 U4630 ( .A(n3091), .B(n4275), .S(n5514), .Z(n3733) );
  AOI22_X1 U4631 ( .A1(n5521), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5520), .ZN(n5518) );
  XNOR2_X1 U4632 ( .A(n3733), .B(n5518), .ZN(n5489) );
  NOR2_X2 U4633 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6703) );
  NAND2_X1 U4634 ( .A1(n6703), .A2(n6912), .ZN(n6085) );
  OR2_X2 U4635 ( .A1(n6085), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6495) );
  INV_X1 U4636 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6892) );
  NOR2_X1 U4637 ( .A1(n6495), .A2(n6892), .ZN(n5474) );
  NAND2_X1 U4638 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6479) );
  NOR2_X1 U4639 ( .A1(n4558), .A2(n6479), .ZN(n6467) );
  NAND2_X1 U4640 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6467), .ZN(n5913)
         );
  NAND2_X1 U4641 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U4642 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5917) );
  NOR3_X1 U4643 ( .A1(n5913), .A2(n5916), .A3(n5917), .ZN(n3760) );
  NAND3_X1 U4644 ( .A1(n3760), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3765) );
  NOR2_X1 U4645 ( .A1(n4571), .A2(n4728), .ZN(n6755) );
  NAND2_X1 U4646 ( .A1(n3761), .A2(n6755), .ZN(n5380) );
  INV_X1 U4647 ( .A(n3734), .ZN(n3741) );
  NAND2_X1 U4648 ( .A1(n5521), .A2(n3735), .ZN(n3740) );
  OAI21_X1 U4649 ( .B1(n5683), .B2(n5184), .A(n3968), .ZN(n3738) );
  INV_X1 U4650 ( .A(n4681), .ZN(n3736) );
  OR2_X1 U4651 ( .A1(n3736), .A2(n3319), .ZN(n3737) );
  NAND4_X1 U4652 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3743)
         );
  INV_X1 U4653 ( .A(n3743), .ZN(n4642) );
  AND2_X1 U4654 ( .A1(n3741), .A2(n4642), .ZN(n4757) );
  NAND2_X1 U4655 ( .A1(n3761), .A2(n4757), .ZN(n6492) );
  INV_X1 U4656 ( .A(n6492), .ZN(n3759) );
  NAND2_X1 U4657 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U4658 ( .A1(n6507), .A2(n3742), .ZN(n6494) );
  NAND2_X1 U4659 ( .A1(n3759), .A2(n6494), .ZN(n5914) );
  AOI21_X1 U4660 ( .B1(n3091), .B2(n3744), .A(n3743), .ZN(n3746) );
  AND3_X1 U4661 ( .A1(n3747), .A2(n3746), .A3(n3745), .ZN(n4623) );
  AND3_X1 U4662 ( .A1(n4737), .A2(n4939), .A3(n4744), .ZN(n3748) );
  AND2_X1 U4663 ( .A1(n3970), .A2(n3748), .ZN(n4778) );
  OAI22_X1 U4664 ( .A1(n4620), .A2(n3794), .B1(n5184), .B2(n4619), .ZN(n3749)
         );
  NOR2_X1 U4665 ( .A1(n4778), .A2(n3749), .ZN(n3750) );
  NAND2_X1 U4666 ( .A1(n4623), .A2(n3750), .ZN(n3751) );
  NAND2_X1 U4667 ( .A1(n3761), .A2(n3751), .ZN(n4653) );
  NAND3_X1 U4668 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6493) );
  OR2_X1 U4669 ( .A1(n4653), .A2(n6493), .ZN(n3753) );
  INV_X1 U4670 ( .A(n3760), .ZN(n3752) );
  AOI21_X1 U4671 ( .B1(n5914), .B2(n3753), .A(n3752), .ZN(n6066) );
  INV_X1 U4672 ( .A(n6066), .ZN(n3754) );
  NAND2_X1 U4673 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5381) );
  NOR2_X1 U4674 ( .A1(n3755), .A2(n5381), .ZN(n6067) );
  NAND2_X1 U4675 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6067), .ZN(n5891) );
  NAND2_X1 U4676 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5892) );
  NOR2_X1 U4677 ( .A1(n5891), .A2(n5892), .ZN(n3768) );
  INV_X1 U4678 ( .A(n6060), .ZN(n3756) );
  NOR2_X1 U4679 ( .A1(n5876), .A2(n3756), .ZN(n5870) );
  INV_X1 U4680 ( .A(n4291), .ZN(n5872) );
  NAND2_X1 U4681 ( .A1(n5870), .A2(n5872), .ZN(n5862) );
  NAND2_X1 U4682 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5829) );
  INV_X1 U4683 ( .A(n5829), .ZN(n3757) );
  NAND2_X1 U4684 ( .A1(n4492), .A2(n3757), .ZN(n3758) );
  NOR2_X1 U4685 ( .A1(n5845), .A2(n3758), .ZN(n5822) );
  NAND2_X1 U4686 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4266) );
  INV_X1 U4687 ( .A(n4266), .ZN(n4279) );
  NAND3_X1 U4688 ( .A1(n5822), .A2(n4279), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U4689 ( .A1(n5380), .A2(n4653), .ZN(n4555) );
  AOI21_X1 U4690 ( .B1(n3760), .B2(n6494), .A(n6492), .ZN(n3764) );
  OR2_X1 U4691 ( .A1(n4653), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3763)
         );
  INV_X1 U4692 ( .A(n3761), .ZN(n3762) );
  NAND2_X1 U4693 ( .A1(n3762), .A2(n6495), .ZN(n4671) );
  NAND2_X1 U4694 ( .A1(n3763), .A2(n4671), .ZN(n4554) );
  NOR2_X1 U4695 ( .A1(n3764), .A2(n4554), .ZN(n3767) );
  NAND2_X1 U4696 ( .A1(n4555), .A2(n3765), .ZN(n3766) );
  NAND2_X1 U4697 ( .A1(n6442), .A2(n3768), .ZN(n3770) );
  NOR2_X1 U4698 ( .A1(n4650), .A2(n4554), .ZN(n5918) );
  INV_X1 U4699 ( .A(n5918), .ZN(n3769) );
  OAI21_X1 U4700 ( .B1(n4291), .B2(n5876), .A(n4650), .ZN(n3771) );
  INV_X1 U4701 ( .A(n3771), .ZN(n3772) );
  NOR2_X1 U4702 ( .A1(n6061), .A2(n3772), .ZN(n5869) );
  NAND2_X1 U4703 ( .A1(n4650), .A2(n5853), .ZN(n3773) );
  NAND2_X1 U4704 ( .A1(n5869), .A2(n3773), .ZN(n5848) );
  INV_X1 U4705 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4670) );
  NAND2_X1 U4706 ( .A1(n5380), .A2(n4670), .ZN(n4649) );
  NAND2_X1 U4707 ( .A1(n4555), .A2(n4649), .ZN(n6500) );
  NAND2_X1 U4708 ( .A1(n6500), .A2(n6492), .ZN(n6051) );
  INV_X1 U4709 ( .A(n4492), .ZN(n5828) );
  AND2_X1 U4710 ( .A1(n6051), .A2(n5828), .ZN(n3774) );
  AND2_X1 U4711 ( .A1(n4650), .A2(n5829), .ZN(n3775) );
  NOR2_X1 U4712 ( .A1(n5833), .A2(n3775), .ZN(n5819) );
  NAND2_X1 U4713 ( .A1(n4650), .A2(n4266), .ZN(n3776) );
  NAND2_X1 U4714 ( .A1(n5819), .A2(n3776), .ZN(n4274) );
  AOI211_X1 U4715 ( .C1(n4650), .C2(n4318), .A(n3544), .B(n4274), .ZN(n5512)
         );
  AOI21_X1 U4716 ( .B1(n3544), .B2(n5525), .A(n5512), .ZN(n3777) );
  AOI211_X1 U4717 ( .C1(n6485), .C2(n5489), .A(n5474), .B(n3777), .ZN(n3778)
         );
  AND2_X1 U4718 ( .A1(n5795), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5721)
         );
  NAND2_X1 U4719 ( .A1(n3779), .A2(n5721), .ZN(n5715) );
  INV_X1 U4720 ( .A(n5715), .ZN(n3784) );
  NOR2_X1 U4721 ( .A1(n4269), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3782)
         );
  OR2_X1 U4722 ( .A1(n5795), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5720)
         );
  NOR3_X1 U4723 ( .A1(n5715), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5821), 
        .ZN(n3781) );
  AOI211_X1 U4724 ( .C1(n3782), .C2(n5714), .A(n5508), .B(n3781), .ZN(n3783)
         );
  OAI21_X1 U4725 ( .B1(n3784), .B2(n4266), .A(n3783), .ZN(n4264) );
  NAND2_X1 U4726 ( .A1(n4264), .A2(n6429), .ZN(n4263) );
  NAND2_X1 U4727 ( .A1(n3786), .A2(n3785), .ZN(n4719) );
  INV_X2 U4728 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6937) );
  NOR2_X1 U4729 ( .A1(n3787), .A2(n6937), .ZN(n3950) );
  INV_X1 U4730 ( .A(n3950), .ZN(n4047) );
  AND2_X1 U4731 ( .A1(n6937), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5530) );
  INV_X1 U4732 ( .A(n5530), .ZN(n4026) );
  NAND2_X1 U4733 ( .A1(n4718), .A2(n3950), .ZN(n3793) );
  OR2_X1 U4734 ( .A1(n5683), .A2(n6937), .ZN(n3823) );
  OR2_X1 U4735 ( .A1(n5686), .A2(n6937), .ZN(n4171) );
  NAND2_X1 U4736 ( .A1(n5531), .A2(EAX_REG_1__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4737 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3789)
         );
  OAI211_X1 U4738 ( .C1(n3823), .C2(n3328), .A(n3790), .B(n3789), .ZN(n3791)
         );
  INV_X1 U4739 ( .A(n3791), .ZN(n3792) );
  NAND2_X1 U4740 ( .A1(n3793), .A2(n3792), .ZN(n4690) );
  OAI21_X1 U4741 ( .B1(n5259), .B2(n3794), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4607) );
  BUF_X1 U4742 ( .A(n3795), .Z(n6653) );
  INV_X2 U4743 ( .A(n4171), .ZN(n5531) );
  NAND2_X1 U4744 ( .A1(n5531), .A2(EAX_REG_0__SCAN_IN), .ZN(n3797) );
  NAND2_X1 U4745 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3796)
         );
  OAI211_X1 U4746 ( .C1(n3823), .C2(n3798), .A(n3797), .B(n3796), .ZN(n3799)
         );
  AOI21_X1 U4747 ( .B1(n6653), .B2(n3950), .A(n3799), .ZN(n4606) );
  OR2_X1 U4748 ( .A1(n4607), .A2(n4606), .ZN(n4609) );
  INV_X1 U4749 ( .A(n4606), .ZN(n3800) );
  INV_X1 U4750 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6089) );
  NAND2_X1 U4751 ( .A1(n6937), .A2(n6089), .ZN(n5473) );
  OR2_X1 U4752 ( .A1(n3800), .A2(n5473), .ZN(n3801) );
  NAND2_X1 U4753 ( .A1(n4609), .A2(n3801), .ZN(n4691) );
  NAND2_X1 U4754 ( .A1(n4690), .A2(n4691), .ZN(n4693) );
  AOI22_X1 U4755 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n4350), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4471), .ZN(n6433) );
  AOI22_X1 U4756 ( .A1(n6433), .A2(n5467), .B1(n5530), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4757 ( .A1(n5531), .A2(EAX_REG_2__SCAN_IN), .ZN(n3802) );
  OAI211_X1 U4758 ( .C1(n3823), .C2(n5505), .A(n3803), .B(n3802), .ZN(n4751)
         );
  NAND2_X1 U4759 ( .A1(n4750), .A2(n4751), .ZN(n3808) );
  INV_X1 U4760 ( .A(n4693), .ZN(n3806) );
  INV_X1 U4761 ( .A(n3804), .ZN(n3805) );
  NAND2_X1 U4762 ( .A1(n3806), .A2(n3805), .ZN(n3807) );
  NAND2_X2 U4763 ( .A1(n3808), .A2(n3807), .ZN(n4748) );
  NAND2_X1 U4764 ( .A1(n3809), .A2(n3950), .ZN(n3817) );
  NAND2_X1 U4765 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3811)
         );
  NAND2_X1 U4766 ( .A1(n5531), .A2(EAX_REG_4__SCAN_IN), .ZN(n3810) );
  OAI211_X1 U4767 ( .C1(n3823), .C2(n3812), .A(n3811), .B(n3810), .ZN(n3815)
         );
  AOI21_X1 U4768 ( .B1(n3819), .B2(n3813), .A(n3829), .ZN(n5308) );
  NOR2_X1 U4769 ( .A1(n5308), .A2(n5473), .ZN(n3814) );
  AOI21_X1 U4770 ( .B1(n3815), .B2(n5473), .A(n3814), .ZN(n3816) );
  NAND2_X1 U4771 ( .A1(n3817), .A2(n3816), .ZN(n4710) );
  NAND2_X1 U4772 ( .A1(n4925), .A2(n3950), .ZN(n3826) );
  OAI21_X1 U4773 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3820), .A(n3819), 
        .ZN(n6424) );
  AOI22_X1 U4774 ( .A1(n6424), .A2(n5467), .B1(n5530), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4775 ( .A1(n5531), .A2(EAX_REG_3__SCAN_IN), .ZN(n3821) );
  OAI211_X1 U4776 ( .C1(n3823), .C2(n4771), .A(n3822), .B(n3821), .ZN(n3824)
         );
  INV_X1 U4777 ( .A(n3824), .ZN(n3825) );
  NAND2_X1 U4778 ( .A1(n3826), .A2(n3825), .ZN(n4711) );
  NAND2_X1 U4779 ( .A1(n3828), .A2(n3950), .ZN(n3835) );
  INV_X1 U4780 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3832) );
  OAI21_X1 U4781 ( .B1(n3829), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3841), 
        .ZN(n6415) );
  NAND2_X1 U4782 ( .A1(n6415), .A2(n5467), .ZN(n3831) );
  NAND2_X1 U4783 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3830)
         );
  OAI211_X1 U4784 ( .C1(n4171), .C2(n3832), .A(n3831), .B(n3830), .ZN(n3833)
         );
  INV_X1 U4785 ( .A(n3833), .ZN(n3834) );
  XNOR2_X1 U4786 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3841), .ZN(n5255) );
  NAND2_X1 U4787 ( .A1(n3836), .A2(n3950), .ZN(n3838) );
  AOI22_X1 U4788 ( .A1(n5531), .A2(EAX_REG_6__SCAN_IN), .B1(n5530), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3837) );
  NOR2_X4 U4789 ( .A1(n4709), .A2(n3839), .ZN(n4998) );
  INV_X1 U4790 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5252) );
  OAI21_X1 U4791 ( .B1(n3842), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3848), 
        .ZN(n6408) );
  INV_X1 U4792 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3844) );
  INV_X1 U4793 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3843) );
  OAI22_X1 U4794 ( .A1(n4171), .A2(n3844), .B1(n4026), .B2(n3843), .ZN(n3845)
         );
  AOI21_X1 U4795 ( .B1(n6408), .B2(n5467), .A(n3845), .ZN(n3846) );
  NAND2_X2 U4796 ( .A1(n3847), .A2(n3846), .ZN(n4999) );
  INV_X1 U4797 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5181) );
  AOI21_X1 U4798 ( .B1(n5181), .B2(n3848), .A(n3866), .ZN(n5189) );
  OR2_X1 U4799 ( .A1(n5189), .A2(n5473), .ZN(n3864) );
  BUF_X1 U4800 ( .A(n3217), .Z(n5445) );
  AOI22_X1 U4801 ( .A1(n3084), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4802 ( .A1(n3152), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4803 ( .A1(n3266), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4804 ( .A1(n4238), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4805 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3858)
         );
  AOI22_X1 U4806 ( .A1(n4217), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5438), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4807 ( .A1(n5437), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4808 ( .A1(n3295), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4809 ( .A1(n3088), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4810 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  NOR2_X1 U4811 ( .A1(n3858), .A2(n3857), .ZN(n3861) );
  NAND2_X1 U4812 ( .A1(n5531), .A2(EAX_REG_8__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4813 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3859)
         );
  OAI211_X1 U4814 ( .C1(n4047), .C2(n3861), .A(n3860), .B(n3859), .ZN(n3862)
         );
  INV_X1 U4815 ( .A(n3862), .ZN(n3863) );
  NAND2_X1 U4816 ( .A1(n3864), .A2(n3863), .ZN(n4886) );
  NAND2_X2 U4817 ( .A1(n4998), .A2(n3865), .ZN(n5052) );
  OAI21_X1 U4818 ( .B1(PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n3866), .A(n3898), 
        .ZN(n6400) );
  AOI22_X1 U4819 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3295), .B1(n5445), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4820 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n3152), .B1(n3084), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4821 ( .A1(n5438), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4822 ( .A1(n5448), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4823 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3876)
         );
  AOI22_X1 U4824 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n4217), .B1(n5437), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4825 ( .A1(n3266), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4826 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n3086), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4827 ( .A1(n4105), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4828 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3875)
         );
  NOR2_X1 U4829 ( .A1(n3876), .A2(n3875), .ZN(n3879) );
  NAND2_X1 U4830 ( .A1(n5531), .A2(EAX_REG_9__SCAN_IN), .ZN(n3878) );
  NAND2_X1 U4831 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3877)
         );
  OAI211_X1 U4832 ( .C1(n4047), .C2(n3879), .A(n3878), .B(n3877), .ZN(n3880)
         );
  AOI21_X1 U4833 ( .B1(n6400), .B2(n5467), .A(n3880), .ZN(n5053) );
  XNOR2_X1 U4834 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3898), .ZN(n6186)
         );
  INV_X1 U4835 ( .A(n6186), .ZN(n3895) );
  AOI22_X1 U4836 ( .A1(n5437), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4837 ( .A1(n4217), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4838 ( .A1(n3295), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4839 ( .A1(n5448), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4840 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3890)
         );
  AOI22_X1 U4841 ( .A1(n5438), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4842 ( .A1(n3084), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4843 ( .A1(n3152), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4844 ( .A1(n4105), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4845 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3889)
         );
  NOR2_X1 U4846 ( .A1(n3890), .A2(n3889), .ZN(n3893) );
  NAND2_X1 U4847 ( .A1(n5531), .A2(EAX_REG_10__SCAN_IN), .ZN(n3892) );
  NAND2_X1 U4848 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3891)
         );
  OAI211_X1 U4849 ( .C1(n4047), .C2(n3893), .A(n3892), .B(n3891), .ZN(n3894)
         );
  AOI21_X1 U4850 ( .B1(n3895), .B2(n5467), .A(n3894), .ZN(n5014) );
  INV_X1 U4851 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U4852 ( .A1(n3900), .A2(n6171), .ZN(n3902) );
  INV_X1 U4853 ( .A(n3932), .ZN(n3901) );
  NAND2_X1 U4854 ( .A1(n3902), .A2(n3901), .ZN(n6174) );
  AOI22_X1 U4855 ( .A1(n4217), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4856 ( .A1(n3266), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4857 ( .A1(n5445), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4858 ( .A1(n5448), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4859 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3912)
         );
  AOI22_X1 U4860 ( .A1(n3295), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3084), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4861 ( .A1(n5437), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4862 ( .A1(n3152), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4863 ( .A1(n5438), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4864 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3911)
         );
  NOR2_X1 U4865 ( .A1(n3912), .A2(n3911), .ZN(n3915) );
  NAND2_X1 U4866 ( .A1(n5531), .A2(EAX_REG_11__SCAN_IN), .ZN(n3914) );
  NAND2_X1 U4867 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3913)
         );
  OAI211_X1 U4868 ( .C1(n4047), .C2(n3915), .A(n3914), .B(n3913), .ZN(n3916)
         );
  AOI21_X1 U4869 ( .B1(n6174), .B2(n5467), .A(n3916), .ZN(n5148) );
  XOR2_X1 U4870 ( .A(n3932), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .Z(n6388) );
  NAND2_X1 U4871 ( .A1(n6388), .A2(n5467), .ZN(n3919) );
  INV_X1 U4872 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5164) );
  OAI21_X1 U4873 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6089), .A(n6937), 
        .ZN(n3917) );
  OAI21_X1 U4874 ( .B1(n4171), .B2(n5164), .A(n3917), .ZN(n3918) );
  NAND2_X1 U4875 ( .A1(n3919), .A2(n3918), .ZN(n3931) );
  AOI22_X1 U4876 ( .A1(n3084), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4877 ( .A1(n3364), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4878 ( .A1(n3295), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4879 ( .A1(n5439), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4880 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3929)
         );
  AOI22_X1 U4881 ( .A1(n4217), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4882 ( .A1(n5438), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4883 ( .A1(n3152), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4884 ( .A1(n5448), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3924) );
  NAND4_X1 U4885 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3928)
         );
  OAI21_X1 U4886 ( .B1(n3929), .B2(n3928), .A(n3950), .ZN(n3930) );
  NAND2_X1 U4887 ( .A1(n3931), .A2(n3930), .ZN(n5156) );
  INV_X1 U4888 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U4889 ( .A1(n3933), .A2(n4430), .ZN(n3935) );
  INV_X1 U4890 ( .A(n3994), .ZN(n3934) );
  NAND2_X1 U4891 ( .A1(n3935), .A2(n3934), .ZN(n6152) );
  NAND2_X1 U4892 ( .A1(n6152), .A2(n5467), .ZN(n3938) );
  NOR2_X1 U4893 ( .A1(n4026), .A2(n4430), .ZN(n3936) );
  AOI21_X1 U4894 ( .B1(n5531), .B2(EAX_REG_13__SCAN_IN), .A(n3936), .ZN(n3937)
         );
  NAND2_X1 U4895 ( .A1(n3938), .A2(n3937), .ZN(n3951) );
  XNOR2_X2 U4896 ( .A(n5155), .B(n3951), .ZN(n5388) );
  AOI22_X1 U4897 ( .A1(n3364), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4898 ( .A1(n3303), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4899 ( .A1(n4217), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4900 ( .A1(n4105), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4901 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3948)
         );
  AOI22_X1 U4902 ( .A1(n3084), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4903 ( .A1(n3425), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4904 ( .A1(n3152), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4905 ( .A1(n5448), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4906 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3947)
         );
  OR2_X1 U4907 ( .A1(n3948), .A2(n3947), .ZN(n3949) );
  AND2_X1 U4908 ( .A1(n3950), .A2(n3949), .ZN(n5389) );
  NAND2_X1 U4909 ( .A1(n5388), .A2(n5389), .ZN(n3954) );
  INV_X1 U4910 ( .A(n3951), .ZN(n3952) );
  NAND2_X2 U4911 ( .A1(n3954), .A2(n3953), .ZN(n5570) );
  AOI22_X1 U4912 ( .A1(n5436), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4913 ( .A1(n3302), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4914 ( .A1(n3152), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4915 ( .A1(n4105), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4916 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3964)
         );
  AOI22_X1 U4917 ( .A1(n3084), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4918 ( .A1(n3303), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4919 ( .A1(n3425), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4920 ( .A1(n4217), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4921 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3963)
         );
  NOR2_X1 U4922 ( .A1(n3964), .A2(n3963), .ZN(n3967) );
  XNOR2_X1 U4923 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3994), .ZN(n6139)
         );
  AOI22_X1 U4924 ( .A1(n5467), .A2(n6139), .B1(n5530), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4925 ( .A1(n5531), .A2(EAX_REG_14__SCAN_IN), .ZN(n3965) );
  OAI211_X1 U4926 ( .C1(n4047), .C2(n3967), .A(n3966), .B(n3965), .ZN(n5569)
         );
  NOR2_X1 U4927 ( .A1(n3968), .A2(n6809), .ZN(n3969) );
  AND2_X1 U4928 ( .A1(n3970), .A2(n3969), .ZN(n5457) );
  AOI22_X1 U4929 ( .A1(n3295), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4930 ( .A1(n3084), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4931 ( .A1(n4217), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4932 ( .A1(n5438), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4933 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4934 ( .A1(n5437), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4935 ( .A1(n3086), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4936 ( .A1(n3266), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4937 ( .A1(n5448), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4938 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  NOR2_X1 U4939 ( .A1(n3980), .A2(n3979), .ZN(n4153) );
  AOI22_X1 U4940 ( .A1(n5438), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4941 ( .A1(n4217), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4942 ( .A1(n3152), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4943 ( .A1(n5427), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4944 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3990)
         );
  AOI22_X1 U4945 ( .A1(n3084), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4946 ( .A1(n5436), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4947 ( .A1(n3295), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4948 ( .A1(n5448), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3985) );
  NAND4_X1 U4949 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3989)
         );
  NOR2_X1 U4950 ( .A1(n3990), .A2(n3989), .ZN(n4154) );
  XNOR2_X1 U4951 ( .A(n4153), .B(n4154), .ZN(n3993) );
  INV_X1 U4952 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3995) );
  OAI21_X1 U4953 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3995), .A(n5473), .ZN(
        n3991) );
  AOI21_X1 U4954 ( .B1(n5531), .B2(EAX_REG_23__SCAN_IN), .A(n3991), .ZN(n3992)
         );
  OAI21_X1 U4955 ( .B1(n5470), .B2(n3993), .A(n3992), .ZN(n3998) );
  INV_X1 U4956 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4401) );
  INV_X1 U4957 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5791) );
  INV_X1 U4958 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U4959 ( .A1(n4066), .A2(n3995), .ZN(n3996) );
  NAND2_X1 U4960 ( .A1(n4167), .A2(n3996), .ZN(n5966) );
  OR2_X1 U4961 ( .A1(n5966), .A2(n5473), .ZN(n3997) );
  NAND2_X1 U4962 ( .A1(n3998), .A2(n3997), .ZN(n5624) );
  INV_X1 U4963 ( .A(n5624), .ZN(n4151) );
  AOI22_X1 U4964 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3084), .B1(n5445), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4965 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3266), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4966 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5448), .B1(n3152), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4967 ( .A1(n5438), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4968 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4008)
         );
  AOI22_X1 U4969 ( .A1(n3364), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4970 ( .A1(n5439), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4971 ( .A1(n3295), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4972 ( .A1(n3088), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4003) );
  NAND4_X1 U4973 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4007)
         );
  NOR2_X1 U4974 ( .A1(n4008), .A2(n4007), .ZN(n4009) );
  OR2_X1 U4975 ( .A1(n5470), .A2(n4009), .ZN(n4015) );
  NAND2_X1 U4976 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4010)
         );
  NAND2_X1 U4977 ( .A1(n5473), .A2(n4010), .ZN(n4011) );
  AOI21_X1 U4978 ( .B1(n5531), .B2(EAX_REG_17__SCAN_IN), .A(n4011), .ZN(n4014)
         );
  OAI21_X1 U4979 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4012), .A(n4144), 
        .ZN(n6113) );
  NOR2_X1 U4980 ( .A1(n6113), .A2(n5473), .ZN(n4013) );
  AOI21_X1 U4981 ( .B1(n4015), .B2(n4014), .A(n4013), .ZN(n5664) );
  INV_X1 U4982 ( .A(n5664), .ZN(n4051) );
  INV_X1 U4983 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U4984 ( .A(n4032), .B(n5799), .ZN(n6131) );
  OR2_X1 U4985 ( .A1(n6131), .A2(n5473), .ZN(n4031) );
  AOI22_X1 U4986 ( .A1(n3084), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4987 ( .A1(n5437), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4988 ( .A1(n5438), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4989 ( .A1(n3152), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4990 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4025)
         );
  AOI22_X1 U4991 ( .A1(n4217), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4992 ( .A1(n3295), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4993 ( .A1(n5448), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4994 ( .A1(n3266), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4995 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  OR2_X1 U4996 ( .A1(n4025), .A2(n4024), .ZN(n4029) );
  INV_X1 U4997 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4027) );
  OAI22_X1 U4998 ( .A1(n4171), .A2(n4027), .B1(n4026), .B2(n5799), .ZN(n4028)
         );
  AOI21_X1 U4999 ( .B1(n5457), .B2(n4029), .A(n4028), .ZN(n4030) );
  AND2_X1 U5000 ( .A1(n4031), .A2(n4030), .ZN(n5672) );
  AOI21_X1 U5001 ( .B1(n4401), .B2(n4033), .A(n4032), .ZN(n5576) );
  OR2_X1 U5002 ( .A1(n5576), .A2(n5473), .ZN(n4050) );
  AOI22_X1 U5003 ( .A1(n5445), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5004 ( .A1(n5438), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5005 ( .A1(n4217), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5006 ( .A1(n4105), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U5007 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4043)
         );
  AOI22_X1 U5008 ( .A1(n5437), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5009 ( .A1(n3295), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5010 ( .A1(n3084), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5011 ( .A1(n5448), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U5012 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4042)
         );
  NOR2_X1 U5013 ( .A1(n4043), .A2(n4042), .ZN(n4046) );
  NAND2_X1 U5014 ( .A1(n5531), .A2(EAX_REG_15__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U5015 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4044)
         );
  OAI211_X1 U5016 ( .C1(n4047), .C2(n4046), .A(n4045), .B(n4044), .ZN(n4048)
         );
  INV_X1 U5017 ( .A(n4048), .ZN(n4049) );
  AND2_X1 U5018 ( .A1(n4050), .A2(n4049), .ZN(n5572) );
  OR2_X1 U5019 ( .A1(n5672), .A2(n5572), .ZN(n5630) );
  OR2_X1 U5020 ( .A1(n4051), .A2(n5630), .ZN(n4150) );
  NAND2_X1 U5021 ( .A1(n5470), .A2(n5473), .ZN(n4138) );
  AOI22_X1 U5022 ( .A1(n4217), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5023 ( .A1(n3303), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4056) );
  NAND2_X1 U5024 ( .A1(n3295), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4053)
         );
  NAND2_X1 U5025 ( .A1(n4127), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4052) );
  AND3_X1 U5026 ( .A1(n4053), .A2(n5473), .A3(n4052), .ZN(n4055) );
  AOI22_X1 U5027 ( .A1(n5445), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U5028 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4063)
         );
  AOI22_X1 U5029 ( .A1(n5437), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5030 ( .A1(n3266), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3084), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5031 ( .A1(n5436), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5032 ( .A1(n5439), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5033 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4062)
         );
  OR2_X1 U5034 ( .A1(n4063), .A2(n4062), .ZN(n4064) );
  NAND2_X1 U5035 ( .A1(n4138), .A2(n4064), .ZN(n4069) );
  AOI22_X1 U5036 ( .A1(n5531), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6937), .ZN(n4068) );
  OR2_X1 U5037 ( .A1(n4085), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4065)
         );
  NAND2_X1 U5038 ( .A1(n4066), .A2(n4065), .ZN(n5977) );
  NOR2_X1 U5039 ( .A1(n5977), .A2(n5473), .ZN(n4067) );
  AOI21_X1 U5040 ( .B1(n4069), .B2(n4068), .A(n4067), .ZN(n5634) );
  AOI22_X1 U5041 ( .A1(n3295), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5042 ( .A1(n4217), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5438), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5043 ( .A1(n3152), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5044 ( .A1(n4105), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U5045 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4079)
         );
  AOI22_X1 U5046 ( .A1(n5437), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5047 ( .A1(n3266), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5048 ( .A1(n3084), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5049 ( .A1(n3088), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5050 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4078)
         );
  NOR2_X1 U5051 ( .A1(n4079), .A2(n4078), .ZN(n4082) );
  INV_X1 U5052 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5756) );
  AOI21_X1 U5053 ( .B1(n5756), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4080) );
  AOI21_X1 U5054 ( .B1(n5531), .B2(EAX_REG_21__SCAN_IN), .A(n4080), .ZN(n4081)
         );
  OAI21_X1 U5055 ( .B1(n5470), .B2(n4082), .A(n4081), .ZN(n4087) );
  NOR2_X1 U5056 ( .A1(n4083), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4084)
         );
  NOR2_X1 U5057 ( .A1(n4085), .A2(n4084), .ZN(n5987) );
  NAND2_X1 U5058 ( .A1(n5987), .A2(n5467), .ZN(n4086) );
  AND2_X1 U5059 ( .A1(n4087), .A2(n4086), .ZN(n5641) );
  INV_X1 U5060 ( .A(n5641), .ZN(n4148) );
  AOI22_X1 U5061 ( .A1(n3295), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5062 ( .A1(n5438), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5063 ( .A1(n4217), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5064 ( .A1(n5445), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5065 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4099)
         );
  AOI22_X1 U5066 ( .A1(n5437), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3084), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5067 ( .A1(n5436), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4096) );
  AOI21_X1 U5068 ( .B1(n3088), .B2(INSTQUEUE_REG_15__4__SCAN_IN), .A(n5467), 
        .ZN(n4093) );
  NAND2_X1 U5069 ( .A1(n3266), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4092)
         );
  AND2_X1 U5070 ( .A1(n4093), .A2(n4092), .ZN(n4095) );
  AOI22_X1 U5071 ( .A1(n3086), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4094) );
  NAND4_X1 U5072 ( .A1(n4097), .A2(n4096), .A3(n4095), .A4(n4094), .ZN(n4098)
         );
  OAI21_X1 U5073 ( .B1(n4099), .B2(n4098), .A(n4138), .ZN(n4102) );
  NOR2_X1 U5074 ( .A1(n5767), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4100) );
  AOI21_X1 U5075 ( .B1(n5531), .B2(EAX_REG_20__SCAN_IN), .A(n4100), .ZN(n4101)
         );
  NAND2_X1 U5076 ( .A1(n4102), .A2(n4101), .ZN(n4104) );
  XNOR2_X1 U5077 ( .A(n4123), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5997)
         );
  NAND2_X1 U5078 ( .A1(n5997), .A2(n5467), .ZN(n4103) );
  NAND2_X1 U5079 ( .A1(n4104), .A2(n4103), .ZN(n5649) );
  AOI22_X1 U5080 ( .A1(n5436), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5081 ( .A1(n5438), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5082 ( .A1(n3152), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5083 ( .A1(n5448), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5084 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4115)
         );
  AOI22_X1 U5085 ( .A1(n3084), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5086 ( .A1(n4217), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5087 ( .A1(n3295), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5088 ( .A1(n3266), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4110) );
  NAND4_X1 U5089 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4114)
         );
  NOR2_X1 U5090 ( .A1(n4115), .A2(n4114), .ZN(n4119) );
  NAND2_X1 U5091 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4116)
         );
  NAND2_X1 U5092 ( .A1(n5473), .A2(n4116), .ZN(n4117) );
  AOI21_X1 U5093 ( .B1(n5531), .B2(EAX_REG_19__SCAN_IN), .A(n4117), .ZN(n4118)
         );
  OAI21_X1 U5094 ( .B1(n5470), .B2(n4119), .A(n4118), .ZN(n4126) );
  INV_X1 U5095 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4122) );
  INV_X1 U5096 ( .A(n4120), .ZN(n4121) );
  NAND2_X1 U5097 ( .A1(n4122), .A2(n4121), .ZN(n4124) );
  AND2_X1 U5098 ( .A1(n4124), .A2(n4123), .ZN(n6008) );
  NAND2_X1 U5099 ( .A1(n6008), .A2(n5467), .ZN(n4125) );
  NAND2_X1 U5100 ( .A1(n4126), .A2(n4125), .ZN(n5779) );
  OR2_X1 U5101 ( .A1(n5649), .A2(n5779), .ZN(n4147) );
  AOI22_X1 U5102 ( .A1(n3266), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5103 ( .A1(n5438), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5104 ( .A1(n5437), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5105 ( .A1(n4217), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5106 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4140)
         );
  AOI22_X1 U5107 ( .A1(n5436), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3084), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5108 ( .A1(n5439), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5109 ( .A1(n3295), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4135) );
  NAND2_X1 U5110 ( .A1(n5427), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4133) );
  AOI21_X1 U5111 ( .B1(n5447), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n5467), 
        .ZN(n4132) );
  AND2_X1 U5112 ( .A1(n4133), .A2(n4132), .ZN(n4134) );
  NAND4_X1 U5113 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4139)
         );
  OAI21_X1 U5114 ( .B1(n4140), .B2(n4139), .A(n4138), .ZN(n4143) );
  NOR2_X1 U5115 ( .A1(n5791), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4141) );
  AOI21_X1 U5116 ( .B1(n5531), .B2(EAX_REG_18__SCAN_IN), .A(n4141), .ZN(n4142)
         );
  NAND2_X1 U5117 ( .A1(n4143), .A2(n4142), .ZN(n4146) );
  XNOR2_X1 U5118 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4144), .ZN(n6104)
         );
  NAND2_X1 U5119 ( .A1(n6104), .A2(n5467), .ZN(n4145) );
  NAND2_X1 U5120 ( .A1(n4146), .A2(n4145), .ZN(n5655) );
  OR2_X1 U5121 ( .A1(n4147), .A2(n5655), .ZN(n5640) );
  NOR2_X1 U5122 ( .A1(n4148), .A2(n5640), .ZN(n5632) );
  NAND2_X1 U5123 ( .A1(n5634), .A2(n5632), .ZN(n4149) );
  NOR2_X1 U5124 ( .A1(n4150), .A2(n4149), .ZN(n5620) );
  NOR2_X1 U5125 ( .A1(n4154), .A2(n4153), .ZN(n4185) );
  AOI22_X1 U5126 ( .A1(n5437), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5127 ( .A1(n3303), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5128 ( .A1(n4217), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5129 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n4105), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4155) );
  NAND4_X1 U5130 ( .A1(n4158), .A2(n4157), .A3(n4156), .A4(n4155), .ZN(n4165)
         );
  INV_X1 U5131 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4497) );
  AOI22_X1 U5132 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3084), .B1(n5445), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5133 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3425), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5134 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n3152), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5135 ( .A1(n5448), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4160) );
  NAND4_X1 U5136 ( .A1(n4163), .A2(n4162), .A3(n4161), .A4(n4160), .ZN(n4164)
         );
  OR2_X1 U5137 ( .A1(n4165), .A2(n4164), .ZN(n4184) );
  INV_X1 U5138 ( .A(n4184), .ZN(n4166) );
  XNOR2_X1 U5139 ( .A(n4185), .B(n4166), .ZN(n4173) );
  INV_X1 U5140 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4662) );
  NAND2_X1 U5141 ( .A1(n5530), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4170)
         );
  INV_X1 U5142 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U5143 ( .A1(n4167), .A2(n5564), .ZN(n4168) );
  NAND2_X1 U5144 ( .A1(n4190), .A2(n4168), .ZN(n5735) );
  NAND2_X1 U5145 ( .A1(n5735), .A2(n5467), .ZN(n4169) );
  OAI211_X1 U5146 ( .C1(n4171), .C2(n4662), .A(n4170), .B(n4169), .ZN(n4172)
         );
  AOI21_X1 U5147 ( .B1(n4173), .B2(n5457), .A(n4172), .ZN(n5563) );
  OR2_X2 U5148 ( .A1(n5622), .A2(n5563), .ZN(n5549) );
  AOI22_X1 U5149 ( .A1(n3303), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5150 ( .A1(n4217), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5151 ( .A1(n3084), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5152 ( .A1(n3152), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4174) );
  NAND4_X1 U5153 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4183)
         );
  AOI22_X1 U5154 ( .A1(n5445), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5155 ( .A1(n5437), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5156 ( .A1(n3425), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5157 ( .A1(n5427), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4178) );
  NAND4_X1 U5158 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4182)
         );
  NOR2_X1 U5159 ( .A1(n4183), .A2(n4182), .ZN(n4196) );
  NAND2_X1 U5160 ( .A1(n4185), .A2(n4184), .ZN(n4195) );
  XNOR2_X1 U5161 ( .A(n4196), .B(n4195), .ZN(n4188) );
  INV_X1 U5162 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4189) );
  OAI21_X1 U5163 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4189), .A(n5473), .ZN(
        n4186) );
  AOI21_X1 U5164 ( .B1(n5531), .B2(EAX_REG_25__SCAN_IN), .A(n4186), .ZN(n4187)
         );
  OAI21_X1 U5165 ( .B1(n4188), .B2(n5470), .A(n4187), .ZN(n4194) );
  INV_X1 U5166 ( .A(n4229), .ZN(n4192) );
  NAND2_X1 U5167 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  NAND2_X1 U5168 ( .A1(n4192), .A2(n4191), .ZN(n5729) );
  OR2_X1 U5169 ( .A1(n5729), .A2(n5473), .ZN(n4193) );
  NAND2_X1 U5170 ( .A1(n4194), .A2(n4193), .ZN(n5548) );
  NOR2_X4 U5171 ( .A1(n5549), .A2(n5548), .ZN(n5609) );
  NOR2_X1 U5172 ( .A1(n4196), .A2(n4195), .ZN(n4225) );
  AOI22_X1 U5173 ( .A1(n3364), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5174 ( .A1(n3303), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5175 ( .A1(n4217), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5176 ( .A1(n5427), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4197) );
  NAND4_X1 U5177 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4206)
         );
  AOI22_X1 U5178 ( .A1(n3084), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5179 ( .A1(n3295), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5180 ( .A1(n3152), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5181 ( .A1(n5448), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4201) );
  NAND4_X1 U5182 ( .A1(n4204), .A2(n4203), .A3(n4202), .A4(n4201), .ZN(n4205)
         );
  OR2_X1 U5183 ( .A1(n4206), .A2(n4205), .ZN(n4224) );
  INV_X1 U5184 ( .A(n4224), .ZN(n4207) );
  XNOR2_X1 U5185 ( .A(n4225), .B(n4207), .ZN(n4208) );
  NAND2_X1 U5186 ( .A1(n4208), .A2(n5457), .ZN(n4212) );
  INV_X1 U5187 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U5188 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5965), .A(n5473), .ZN(
        n4209) );
  AOI21_X1 U5189 ( .B1(n5531), .B2(EAX_REG_26__SCAN_IN), .A(n4209), .ZN(n4211)
         );
  XNOR2_X1 U5190 ( .A(n4229), .B(n5965), .ZN(n5956) );
  AND2_X1 U5191 ( .A1(n5956), .A2(n5467), .ZN(n4210) );
  AOI21_X1 U5192 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n5608) );
  AND2_X2 U5193 ( .A1(n5609), .A2(n5608), .ZN(n5600) );
  AOI22_X1 U5194 ( .A1(n3084), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5195 ( .A1(n3303), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5196 ( .A1(n3425), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5197 ( .A1(n3152), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U5198 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4223)
         );
  AOI22_X1 U5199 ( .A1(n4217), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5200 ( .A1(n3302), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5201 ( .A1(n5448), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5202 ( .A1(n4238), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4218) );
  NAND4_X1 U5203 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(n4222)
         );
  NOR2_X1 U5204 ( .A1(n4223), .A2(n4222), .ZN(n4237) );
  NAND2_X1 U5205 ( .A1(n4225), .A2(n4224), .ZN(n4236) );
  XNOR2_X1 U5206 ( .A(n4237), .B(n4236), .ZN(n4228) );
  INV_X1 U5207 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4230) );
  OAI21_X1 U5208 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4230), .A(n5473), .ZN(
        n4226) );
  AOI21_X1 U5209 ( .B1(n5531), .B2(EAX_REG_27__SCAN_IN), .A(n4226), .ZN(n4227)
         );
  OAI21_X1 U5210 ( .B1(n4228), .B2(n5470), .A(n4227), .ZN(n4235) );
  NAND2_X1 U5211 ( .A1(n4229), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4231)
         );
  NAND2_X1 U5212 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  NAND2_X1 U5213 ( .A1(n5170), .A2(n4232), .ZN(n5949) );
  INV_X1 U5214 ( .A(n5949), .ZN(n4233) );
  NAND2_X1 U5215 ( .A1(n4233), .A2(n5467), .ZN(n4234) );
  AND2_X1 U5216 ( .A1(n4235), .A2(n4234), .ZN(n5601) );
  AND2_X2 U5217 ( .A1(n5600), .A2(n5601), .ZN(n5603) );
  XNOR2_X1 U5218 ( .A(n5170), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5415)
         );
  INV_X1 U5219 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5169) );
  OAI21_X1 U5220 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5169), .A(n5473), .ZN(
        n4252) );
  NOR2_X1 U5221 ( .A1(n4237), .A2(n4236), .ZN(n5435) );
  AOI22_X1 U5222 ( .A1(n5437), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5223 ( .A1(n5438), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5224 ( .A1(n4217), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U5225 ( .A1(n4238), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4239) );
  NAND4_X1 U5226 ( .A1(n4242), .A2(n4241), .A3(n4240), .A4(n4239), .ZN(n4249)
         );
  INV_X1 U5227 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U5228 ( .A1(n3084), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U5229 ( .A1(n3425), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U5230 ( .A1(n3152), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4245) );
  AOI22_X1 U5231 ( .A1(n5448), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4244) );
  NAND4_X1 U5232 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(n4248)
         );
  OR2_X1 U5233 ( .A1(n4249), .A2(n4248), .ZN(n5434) );
  XNOR2_X1 U5234 ( .A(n5435), .B(n5434), .ZN(n4250) );
  NOR2_X1 U5235 ( .A1(n4250), .A2(n5470), .ZN(n4251) );
  AOI211_X1 U5236 ( .C1(n5531), .C2(EAX_REG_28__SCAN_IN), .A(n4252), .B(n4251), 
        .ZN(n4253) );
  AOI21_X1 U5237 ( .B1(n5467), .B2(n5415), .A(n4253), .ZN(n4254) );
  OAI21_X1 U5238 ( .B1(n5603), .B2(n4254), .A(n5479), .ZN(n5693) );
  AND2_X1 U5239 ( .A1(n6809), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5165) );
  NAND3_X1 U5240 ( .A1(n5165), .A2(n6703), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n6696) );
  INV_X1 U5241 ( .A(n6703), .ZN(n6934) );
  NAND2_X1 U5242 ( .A1(n6934), .A2(n6933), .ZN(n4255) );
  NAND2_X1 U5243 ( .A1(n4255), .A2(n6809), .ZN(n4256) );
  AND2_X2 U5244 ( .A1(n6410), .A2(n4256), .ZN(n6425) );
  NAND2_X1 U5245 ( .A1(n6809), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U5246 ( .A1(n6089), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4257) );
  AND2_X1 U5247 ( .A1(n4258), .A2(n4257), .ZN(n4611) );
  INV_X1 U5248 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6886) );
  NOR2_X1 U5249 ( .A1(n6495), .A2(n6886), .ZN(n4268) );
  INV_X1 U5250 ( .A(n6425), .ZN(n5800) );
  NOR2_X1 U5251 ( .A1(n5800), .A2(n5169), .ZN(n4259) );
  AOI211_X1 U5252 ( .C1(n6387), .C2(n5415), .A(n4268), .B(n4259), .ZN(n4260)
         );
  NAND2_X1 U5253 ( .A1(n4263), .A2(n4262), .ZN(U2958) );
  NAND2_X1 U5254 ( .A1(n4264), .A2(n6503), .ZN(n4273) );
  AOI21_X1 U5255 ( .B1(n4265), .B2(n5606), .A(n5514), .ZN(n5417) );
  AND3_X1 U5256 ( .A1(n5822), .A2(n4282), .A3(n4266), .ZN(n4267) );
  AOI211_X1 U5257 ( .C1(n5417), .C2(n6485), .A(n4268), .B(n4267), .ZN(n4271)
         );
  OR2_X1 U5258 ( .A1(n5819), .A2(n4269), .ZN(n4270) );
  NAND2_X1 U5259 ( .A1(n4273), .A2(n4272), .ZN(U2990) );
  INV_X1 U5260 ( .A(n4274), .ZN(n4288) );
  OR2_X1 U5261 ( .A1(n4275), .A2(n3091), .ZN(n4276) );
  INV_X1 U5262 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5596) );
  OR2_X1 U5263 ( .A1(n5659), .A2(n5596), .ZN(n5516) );
  AND2_X1 U5264 ( .A1(n4276), .A2(n5516), .ZN(n4277) );
  NAND2_X1 U5265 ( .A1(n5514), .A2(n4277), .ZN(n5519) );
  OR2_X1 U5266 ( .A1(n5514), .A2(n4277), .ZN(n4278) );
  NAND2_X1 U5267 ( .A1(n5519), .A2(n4278), .ZN(n5947) );
  INV_X1 U5268 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6888) );
  OR2_X1 U5269 ( .A1(n6495), .A2(n6888), .ZN(n5482) );
  NAND3_X1 U5270 ( .A1(n5822), .A2(n4279), .A3(n4318), .ZN(n4280) );
  OAI211_X1 U5271 ( .C1(n5947), .C2(n6497), .A(n5482), .B(n4280), .ZN(n4281)
         );
  INV_X1 U5272 ( .A(n4281), .ZN(n4287) );
  NOR2_X1 U5273 ( .A1(n5720), .A2(n4282), .ZN(n4284) );
  AOI22_X1 U5274 ( .A1(n4285), .A2(n5795), .B1(n4284), .B2(n4283), .ZN(n4286)
         );
  XNOR2_X1 U5275 ( .A(n4286), .B(n4318), .ZN(n5485) );
  OAI211_X1 U5276 ( .C1(n4318), .C2(n4288), .A(n4287), .B(n3095), .ZN(U2989)
         );
  XNOR2_X1 U5277 ( .A(n5795), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5773)
         );
  NAND2_X1 U5278 ( .A1(n4290), .A2(n5773), .ZN(n5772) );
  NAND2_X1 U5279 ( .A1(n4289), .A2(n4291), .ZN(n4292) );
  XNOR2_X1 U5280 ( .A(n5795), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5754)
         );
  NAND2_X1 U5281 ( .A1(n5755), .A2(n5754), .ZN(n5753) );
  MUX2_X1 U5282 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .B(n4314), .S(n5795), 
        .Z(n4293) );
  INV_X1 U5283 ( .A(n4293), .ZN(n4294) );
  XNOR2_X1 U5284 ( .A(n4297), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5739)
         );
  INV_X1 U5285 ( .A(n4298), .ZN(n4299) );
  XNOR2_X1 U5286 ( .A(n5626), .B(n4299), .ZN(n5618) );
  INV_X1 U5287 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U5288 ( .A1(n6495), .A2(n6873), .ZN(n5733) );
  AOI21_X1 U5289 ( .B1(n5618), .B2(n6485), .A(n5733), .ZN(n4302) );
  NOR2_X1 U5290 ( .A1(n5845), .A2(n4314), .ZN(n4300) );
  OAI21_X1 U5291 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4300), .A(n5833), 
        .ZN(n4301) );
  OAI21_X1 U5292 ( .B1(n5739), .B2(n6476), .A(n3098), .ZN(n4553) );
  INV_X1 U5293 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5305) );
  AOI22_X1 U5294 ( .A1(n5305), .A2(keyinput58), .B1(keyinput114), .B2(n5756), 
        .ZN(n4303) );
  OAI221_X1 U5295 ( .B1(n5305), .B2(keyinput58), .C1(n5756), .C2(keyinput114), 
        .A(n4303), .ZN(n4312) );
  INV_X1 U5296 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4306) );
  INV_X1 U5297 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U5298 ( .A1(n4306), .A2(keyinput92), .B1(n4305), .B2(keyinput42), 
        .ZN(n4304) );
  OAI221_X1 U5299 ( .B1(n4306), .B2(keyinput92), .C1(n4305), .C2(keyinput42), 
        .A(n4304), .ZN(n4311) );
  INV_X1 U5300 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6285) );
  INV_X1 U5301 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6326) );
  AOI22_X1 U5302 ( .A1(n6285), .A2(keyinput10), .B1(keyinput103), .B2(n6326), 
        .ZN(n4307) );
  OAI221_X1 U5303 ( .B1(n6285), .B2(keyinput10), .C1(n6326), .C2(keyinput103), 
        .A(n4307), .ZN(n4310) );
  INV_X1 U5304 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6843) );
  INV_X1 U5305 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6854) );
  AOI22_X1 U5306 ( .A1(n6843), .A2(keyinput105), .B1(keyinput22), .B2(n6854), 
        .ZN(n4308) );
  OAI221_X1 U5307 ( .B1(n6843), .B2(keyinput105), .C1(n6854), .C2(keyinput22), 
        .A(n4308), .ZN(n4309) );
  NOR4_X1 U5308 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4324)
         );
  INV_X1 U5309 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6816) );
  AOI22_X1 U5310 ( .A1(n4314), .A2(keyinput81), .B1(keyinput8), .B2(n6816), 
        .ZN(n4313) );
  OAI221_X1 U5311 ( .B1(n4314), .B2(keyinput81), .C1(n6816), .C2(keyinput8), 
        .A(n4313), .ZN(n4322) );
  INV_X1 U5312 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U5313 ( .A1(n6867), .A2(keyinput17), .B1(n3701), .B2(keyinput45), 
        .ZN(n4315) );
  OAI221_X1 U5314 ( .B1(n6867), .B2(keyinput17), .C1(n3701), .C2(keyinput45), 
        .A(n4315), .ZN(n4321) );
  OAI221_X1 U5315 ( .B1(n6162), .B2(keyinput11), .C1(n5181), .C2(keyinput78), 
        .A(n4316), .ZN(n4320) );
  AOI22_X1 U5316 ( .A1(n6473), .A2(keyinput64), .B1(keyinput116), .B2(n4318), 
        .ZN(n4317) );
  OAI221_X1 U5317 ( .B1(n6473), .B2(keyinput64), .C1(n4318), .C2(keyinput116), 
        .A(n4317), .ZN(n4319) );
  NOR4_X1 U5318 ( .A1(n4322), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(n4323)
         );
  NAND2_X1 U5319 ( .A1(n4324), .A2(n4323), .ZN(n4491) );
  INV_X1 U5320 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n4326) );
  INV_X1 U5321 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U5322 ( .A1(n4326), .A2(keyinput43), .B1(keyinput48), .B2(n6895), 
        .ZN(n4325) );
  OAI221_X1 U5323 ( .B1(n4326), .B2(keyinput43), .C1(n6895), .C2(keyinput48), 
        .A(n4325), .ZN(n4336) );
  INV_X1 U5324 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4328) );
  INV_X1 U5325 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6310) );
  AOI22_X1 U5326 ( .A1(n4328), .A2(keyinput80), .B1(keyinput111), .B2(n6310), 
        .ZN(n4327) );
  OAI221_X1 U5327 ( .B1(n4328), .B2(keyinput80), .C1(n6310), .C2(keyinput111), 
        .A(n4327), .ZN(n4335) );
  INV_X1 U5328 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6305) );
  INV_X1 U5329 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U5330 ( .A1(n6305), .A2(keyinput112), .B1(n4330), .B2(keyinput50), 
        .ZN(n4329) );
  OAI221_X1 U5331 ( .B1(n6305), .B2(keyinput112), .C1(n4330), .C2(keyinput50), 
        .A(n4329), .ZN(n4334) );
  INV_X1 U5332 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4496) );
  INV_X1 U5333 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U5334 ( .A1(n4496), .A2(keyinput35), .B1(n4332), .B2(keyinput18), 
        .ZN(n4331) );
  OAI221_X1 U5335 ( .B1(n4496), .B2(keyinput35), .C1(n4332), .C2(keyinput18), 
        .A(n4331), .ZN(n4333) );
  NOR4_X1 U5336 ( .A1(n4336), .A2(n4335), .A3(n4334), .A4(n4333), .ZN(n4371)
         );
  INV_X1 U5337 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4804) );
  INV_X1 U5338 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6880) );
  AOI22_X1 U5339 ( .A1(n4804), .A2(keyinput51), .B1(keyinput49), .B2(n6880), 
        .ZN(n4337) );
  OAI221_X1 U5340 ( .B1(n4804), .B2(keyinput51), .C1(n6880), .C2(keyinput49), 
        .A(n4337), .ZN(n4347) );
  INV_X1 U5341 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6885) );
  AOI22_X1 U5342 ( .A1(n6885), .A2(keyinput1), .B1(n5588), .B2(keyinput74), 
        .ZN(n4338) );
  OAI221_X1 U5343 ( .B1(n6885), .B2(keyinput1), .C1(n5588), .C2(keyinput74), 
        .A(n4338), .ZN(n4346) );
  INV_X1 U5344 ( .A(DATAI_29_), .ZN(n4340) );
  INV_X1 U5345 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U5346 ( .A1(n4340), .A2(keyinput123), .B1(keyinput37), .B2(n6814), 
        .ZN(n4339) );
  OAI221_X1 U5347 ( .B1(n4340), .B2(keyinput123), .C1(n6814), .C2(keyinput37), 
        .A(n4339), .ZN(n4345) );
  INV_X1 U5348 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4343) );
  INV_X1 U5349 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U5350 ( .A1(n4343), .A2(keyinput73), .B1(n4342), .B2(keyinput67), 
        .ZN(n4341) );
  OAI221_X1 U5351 ( .B1(n4343), .B2(keyinput73), .C1(n4342), .C2(keyinput67), 
        .A(n4341), .ZN(n4344) );
  NOR4_X1 U5352 ( .A1(n4347), .A2(n4346), .A3(n4345), .A4(n4344), .ZN(n4370)
         );
  INV_X1 U5353 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6281) );
  INV_X1 U5354 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6313) );
  AOI22_X1 U5355 ( .A1(n6281), .A2(keyinput27), .B1(n6313), .B2(keyinput84), 
        .ZN(n4348) );
  OAI221_X1 U5356 ( .B1(n6281), .B2(keyinput27), .C1(n6313), .C2(keyinput84), 
        .A(n4348), .ZN(n4358) );
  INV_X1 U5357 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U5358 ( .A1(n4350), .A2(keyinput113), .B1(n6840), .B2(keyinput72), 
        .ZN(n4349) );
  OAI221_X1 U5359 ( .B1(n4350), .B2(keyinput113), .C1(n6840), .C2(keyinput72), 
        .A(n4349), .ZN(n4357) );
  INV_X1 U5360 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4352) );
  AOI22_X1 U5361 ( .A1(n3995), .A2(keyinput65), .B1(n4352), .B2(keyinput60), 
        .ZN(n4351) );
  OAI221_X1 U5362 ( .B1(n3995), .B2(keyinput65), .C1(n4352), .C2(keyinput60), 
        .A(n4351), .ZN(n4356) );
  INV_X1 U5363 ( .A(DATAI_14_), .ZN(n6381) );
  INV_X1 U5364 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U5365 ( .A1(n6381), .A2(keyinput89), .B1(n4354), .B2(keyinput13), 
        .ZN(n4353) );
  OAI221_X1 U5366 ( .B1(n6381), .B2(keyinput89), .C1(n4354), .C2(keyinput13), 
        .A(n4353), .ZN(n4355) );
  NOR4_X1 U5367 ( .A1(n4358), .A2(n4357), .A3(n4356), .A4(n4355), .ZN(n4369)
         );
  INV_X1 U5368 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5615) );
  AOI22_X1 U5369 ( .A1(n4530), .A2(keyinput21), .B1(keyinput121), .B2(n5615), 
        .ZN(n4359) );
  OAI221_X1 U5370 ( .B1(n4530), .B2(keyinput21), .C1(n5615), .C2(keyinput121), 
        .A(n4359), .ZN(n4367) );
  INV_X1 U5371 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6295) );
  INV_X1 U5372 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6080) );
  AOI22_X1 U5373 ( .A1(n6295), .A2(keyinput94), .B1(n6080), .B2(keyinput6), 
        .ZN(n4360) );
  OAI221_X1 U5374 ( .B1(n6295), .B2(keyinput94), .C1(n6080), .C2(keyinput6), 
        .A(n4360), .ZN(n4366) );
  INV_X1 U5375 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U5376 ( .A1(n4362), .A2(keyinput55), .B1(keyinput52), .B2(n6892), 
        .ZN(n4361) );
  OAI221_X1 U5377 ( .B1(n4362), .B2(keyinput55), .C1(n6892), .C2(keyinput52), 
        .A(n4361), .ZN(n4365) );
  INV_X1 U5378 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6817) );
  AOI22_X1 U5379 ( .A1(n5843), .A2(keyinput125), .B1(n6817), .B2(keyinput82), 
        .ZN(n4363) );
  OAI221_X1 U5380 ( .B1(n5843), .B2(keyinput125), .C1(n6817), .C2(keyinput82), 
        .A(n4363), .ZN(n4364) );
  NOR4_X1 U5381 ( .A1(n4367), .A2(n4366), .A3(n4365), .A4(n4364), .ZN(n4368)
         );
  NAND4_X1 U5382 ( .A1(n4371), .A2(n4370), .A3(n4369), .A4(n4368), .ZN(n4490)
         );
  INV_X1 U5383 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6114) );
  INV_X1 U5384 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6818) );
  AOI22_X1 U5385 ( .A1(n6114), .A2(keyinput87), .B1(n6818), .B2(keyinput98), 
        .ZN(n4372) );
  OAI221_X1 U5386 ( .B1(n6114), .B2(keyinput87), .C1(n6818), .C2(keyinput98), 
        .A(n4372), .ZN(n4380) );
  INV_X1 U5387 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6312) );
  AOI22_X1 U5388 ( .A1(n6312), .A2(keyinput99), .B1(n6873), .B2(keyinput23), 
        .ZN(n4373) );
  OAI221_X1 U5389 ( .B1(n6312), .B2(keyinput99), .C1(n6873), .C2(keyinput23), 
        .A(n4373), .ZN(n4379) );
  INV_X1 U5390 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U5391 ( .A1(n4375), .A2(keyinput39), .B1(keyinput24), .B2(n6260), 
        .ZN(n4374) );
  OAI221_X1 U5392 ( .B1(n4375), .B2(keyinput39), .C1(n6260), .C2(keyinput24), 
        .A(n4374), .ZN(n4378) );
  INV_X1 U5393 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4601) );
  INV_X1 U5394 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U5395 ( .A1(n4601), .A2(keyinput77), .B1(keyinput76), .B2(n6320), 
        .ZN(n4376) );
  OAI221_X1 U5396 ( .B1(n4601), .B2(keyinput77), .C1(n6320), .C2(keyinput76), 
        .A(n4376), .ZN(n4377) );
  NOR4_X1 U5397 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), .ZN(n4413)
         );
  INV_X1 U5398 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U5399 ( .A1(n6881), .A2(keyinput75), .B1(n5235), .B2(keyinput119), 
        .ZN(n4381) );
  OAI221_X1 U5400 ( .B1(n6881), .B2(keyinput75), .C1(n5235), .C2(keyinput119), 
        .A(n4381), .ZN(n4389) );
  INV_X1 U5401 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4498) );
  AOI22_X1 U5402 ( .A1(n6827), .A2(keyinput31), .B1(keyinput12), .B2(n4498), 
        .ZN(n4382) );
  OAI221_X1 U5403 ( .B1(n6827), .B2(keyinput31), .C1(n4498), .C2(keyinput12), 
        .A(n4382), .ZN(n4388) );
  INV_X1 U5404 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4385) );
  INV_X1 U5405 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6308) );
  AOI22_X1 U5406 ( .A1(n4385), .A2(keyinput68), .B1(keyinput46), .B2(n6308), 
        .ZN(n4384) );
  OAI221_X1 U5407 ( .B1(n4385), .B2(keyinput68), .C1(n6308), .C2(keyinput46), 
        .A(n4384), .ZN(n4386) );
  NOR4_X1 U5408 ( .A1(n4389), .A2(n4388), .A3(n4387), .A4(n4386), .ZN(n4412)
         );
  INV_X1 U5409 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6848) );
  INV_X1 U5410 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U5411 ( .A1(n6848), .A2(keyinput115), .B1(n4391), .B2(keyinput34), 
        .ZN(n4390) );
  OAI221_X1 U5412 ( .B1(n6848), .B2(keyinput115), .C1(n4391), .C2(keyinput34), 
        .A(n4390), .ZN(n4399) );
  INV_X1 U5413 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5414 ( .A1(n4493), .A2(keyinput104), .B1(n4495), .B2(keyinput53), 
        .ZN(n4392) );
  OAI221_X1 U5415 ( .B1(n4493), .B2(keyinput104), .C1(n4495), .C2(keyinput53), 
        .A(n4392), .ZN(n4398) );
  INV_X1 U5416 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6289) );
  INV_X1 U5417 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U5418 ( .A1(n6289), .A2(keyinput3), .B1(n4494), .B2(keyinput108), 
        .ZN(n4393) );
  OAI221_X1 U5419 ( .B1(n6289), .B2(keyinput3), .C1(n4494), .C2(keyinput108), 
        .A(n4393), .ZN(n4397) );
  INV_X1 U5420 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4395) );
  INV_X1 U5421 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6874) );
  AOI22_X1 U5422 ( .A1(n4395), .A2(keyinput15), .B1(keyinput38), .B2(n6874), 
        .ZN(n4394) );
  OAI221_X1 U5423 ( .B1(n4395), .B2(keyinput15), .C1(n6874), .C2(keyinput38), 
        .A(n4394), .ZN(n4396) );
  NOR4_X1 U5424 ( .A1(n4399), .A2(n4398), .A3(n4397), .A4(n4396), .ZN(n4411)
         );
  INV_X1 U5425 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6287) );
  INV_X1 U5426 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5427 ( .A1(n6287), .A2(keyinput110), .B1(keyinput30), .B2(n4616), 
        .ZN(n4402) );
  OAI221_X1 U5428 ( .B1(n6287), .B2(keyinput110), .C1(n4616), .C2(keyinput30), 
        .A(n4402), .ZN(n4408) );
  INV_X1 U5429 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6869) );
  AOI22_X1 U5430 ( .A1(n6869), .A2(keyinput5), .B1(n4404), .B2(keyinput62), 
        .ZN(n4403) );
  OAI221_X1 U5431 ( .B1(n6869), .B2(keyinput5), .C1(n4404), .C2(keyinput62), 
        .A(n4403), .ZN(n4407) );
  INV_X1 U5432 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6845) );
  INV_X1 U5433 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6297) );
  AOI22_X1 U5434 ( .A1(n6845), .A2(keyinput124), .B1(n6297), .B2(keyinput29), 
        .ZN(n4405) );
  OAI221_X1 U5435 ( .B1(n6845), .B2(keyinput124), .C1(n6297), .C2(keyinput29), 
        .A(n4405), .ZN(n4406) );
  NOR4_X1 U5436 ( .A1(n4409), .A2(n4408), .A3(n4407), .A4(n4406), .ZN(n4410)
         );
  NAND4_X1 U5437 ( .A1(n4413), .A2(n4412), .A3(n4411), .A4(n4410), .ZN(n4489)
         );
  INV_X1 U5438 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6549) );
  AOI22_X1 U5439 ( .A1(n6912), .A2(keyinput88), .B1(keyinput91), .B2(n6549), 
        .ZN(n4414) );
  OAI221_X1 U5440 ( .B1(n6912), .B2(keyinput88), .C1(n6549), .C2(keyinput91), 
        .A(n4414), .ZN(n4422) );
  INV_X1 U5441 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U5442 ( .A1(n4416), .A2(keyinput20), .B1(keyinput71), .B2(n6859), 
        .ZN(n4415) );
  OAI221_X1 U5443 ( .B1(n4416), .B2(keyinput20), .C1(n6859), .C2(keyinput71), 
        .A(n4415), .ZN(n4421) );
  INV_X1 U5444 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5491) );
  INV_X1 U5445 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6868) );
  AOI22_X1 U5446 ( .A1(n5491), .A2(keyinput44), .B1(n6868), .B2(keyinput69), 
        .ZN(n4417) );
  OAI221_X1 U5447 ( .B1(n5491), .B2(keyinput44), .C1(n6868), .C2(keyinput69), 
        .A(n4417), .ZN(n4420) );
  INV_X1 U5448 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6293) );
  INV_X1 U5449 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6081) );
  AOI22_X1 U5450 ( .A1(n6293), .A2(keyinput118), .B1(n6081), .B2(keyinput127), 
        .ZN(n4418) );
  OAI221_X1 U5451 ( .B1(n6293), .B2(keyinput118), .C1(n6081), .C2(keyinput127), 
        .A(n4418), .ZN(n4419) );
  NOR4_X1 U5452 ( .A1(n4422), .A2(n4421), .A3(n4420), .A4(n4419), .ZN(n4487)
         );
  INV_X1 U5453 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U5454 ( .A1(n4425), .A2(keyinput4), .B1(n4424), .B2(keyinput117), 
        .ZN(n4423) );
  OAI221_X1 U5455 ( .B1(n4425), .B2(keyinput4), .C1(n4424), .C2(keyinput117), 
        .A(n4423), .ZN(n4434) );
  INV_X1 U5456 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4427) );
  INV_X1 U5457 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5614) );
  AOI22_X1 U5458 ( .A1(n4427), .A2(keyinput32), .B1(keyinput102), .B2(n5614), 
        .ZN(n4426) );
  OAI221_X1 U5459 ( .B1(n4427), .B2(keyinput32), .C1(n5614), .C2(keyinput102), 
        .A(n4426), .ZN(n4433) );
  INV_X1 U5460 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5446) );
  AOI22_X1 U5461 ( .A1(n5860), .A2(keyinput54), .B1(n5446), .B2(keyinput96), 
        .ZN(n4428) );
  OAI221_X1 U5462 ( .B1(n5860), .B2(keyinput54), .C1(n5446), .C2(keyinput96), 
        .A(n4428), .ZN(n4432) );
  INV_X1 U5463 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6849) );
  NOR4_X1 U5464 ( .A1(n4434), .A2(n4433), .A3(n4432), .A4(n4431), .ZN(n4486)
         );
  INV_X1 U5465 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4529) );
  INV_X1 U5466 ( .A(BS16_N), .ZN(n4436) );
  AOI22_X1 U5467 ( .A1(n4529), .A2(keyinput25), .B1(keyinput97), .B2(n4436), 
        .ZN(n4435) );
  OAI221_X1 U5468 ( .B1(n4529), .B2(keyinput25), .C1(n4436), .C2(keyinput97), 
        .A(n4435), .ZN(n4444) );
  INV_X1 U5469 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5868) );
  INV_X1 U5470 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U5471 ( .A1(n5868), .A2(keyinput36), .B1(n4438), .B2(keyinput19), 
        .ZN(n4437) );
  OAI221_X1 U5472 ( .B1(n5868), .B2(keyinput36), .C1(n4438), .C2(keyinput19), 
        .A(n4437), .ZN(n4443) );
  INV_X1 U5473 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U5474 ( .A1(n6921), .A2(keyinput47), .B1(n6501), .B2(keyinput59), 
        .ZN(n4439) );
  OAI221_X1 U5475 ( .B1(n6921), .B2(keyinput47), .C1(n6501), .C2(keyinput59), 
        .A(n4439), .ZN(n4442) );
  INV_X1 U5476 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5978) );
  AOI22_X1 U5477 ( .A1(n4531), .A2(keyinput79), .B1(keyinput16), .B2(n5978), 
        .ZN(n4440) );
  OAI221_X1 U5478 ( .B1(n4531), .B2(keyinput79), .C1(n5978), .C2(keyinput16), 
        .A(n4440), .ZN(n4441) );
  NOR4_X1 U5479 ( .A1(n4444), .A2(n4443), .A3(n4442), .A4(n4441), .ZN(n4485)
         );
  INV_X1 U5480 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6858) );
  INV_X1 U5481 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5482 ( .A1(n6858), .A2(keyinput14), .B1(n4528), .B2(keyinput83), 
        .ZN(n4445) );
  OAI221_X1 U5483 ( .B1(n6858), .B2(keyinput14), .C1(n4528), .C2(keyinput83), 
        .A(n4445), .ZN(n4450) );
  INV_X1 U5484 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6283) );
  INV_X1 U5485 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U5486 ( .A1(n6283), .A2(keyinput106), .B1(n4447), .B2(keyinput41), 
        .ZN(n4446) );
  OAI221_X1 U5487 ( .B1(n6283), .B2(keyinput106), .C1(n4447), .C2(keyinput41), 
        .A(n4446), .ZN(n4449) );
  INV_X1 U5488 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6893) );
  XNOR2_X1 U5489 ( .A(n6893), .B(keyinput40), .ZN(n4448) );
  NOR3_X1 U5490 ( .A1(n4450), .A2(n4449), .A3(n4448), .ZN(n4483) );
  INV_X1 U5491 ( .A(DATAI_25_), .ZN(n4452) );
  AOI22_X1 U5492 ( .A1(n4453), .A2(keyinput95), .B1(keyinput86), .B2(n4452), 
        .ZN(n4451) );
  OAI221_X1 U5493 ( .B1(n4453), .B2(keyinput95), .C1(n4452), .C2(keyinput86), 
        .A(n4451), .ZN(n4456) );
  INV_X1 U5494 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6621) );
  INV_X1 U5495 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n6300) );
  AOI22_X1 U5496 ( .A1(n6621), .A2(keyinput63), .B1(keyinput85), .B2(n6300), 
        .ZN(n4454) );
  OAI221_X1 U5497 ( .B1(n6621), .B2(keyinput63), .C1(n6300), .C2(keyinput85), 
        .A(n4454), .ZN(n4455) );
  NOR2_X1 U5498 ( .A1(n4456), .A2(n4455), .ZN(n4482) );
  INV_X1 U5499 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6815) );
  INV_X1 U5500 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U5501 ( .A1(n6815), .A2(keyinput33), .B1(n4458), .B2(keyinput70), 
        .ZN(n4457) );
  OAI221_X1 U5502 ( .B1(n6815), .B2(keyinput33), .C1(n4458), .C2(keyinput70), 
        .A(n4457), .ZN(n4461) );
  INV_X1 U5503 ( .A(DATAI_18_), .ZN(n4519) );
  INV_X1 U5504 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4669) );
  AOI22_X1 U5505 ( .A1(n4519), .A2(keyinput126), .B1(keyinput61), .B2(n4669), 
        .ZN(n4459) );
  OAI221_X1 U5506 ( .B1(n4519), .B2(keyinput126), .C1(n4669), .C2(keyinput61), 
        .A(n4459), .ZN(n4460) );
  NOR2_X1 U5507 ( .A1(n4461), .A2(n4460), .ZN(n4469) );
  AOI22_X1 U5508 ( .A1(n4497), .A2(keyinput109), .B1(keyinput57), .B2(n6888), 
        .ZN(n4462) );
  OAI221_X1 U5509 ( .B1(n4497), .B2(keyinput109), .C1(n6888), .C2(keyinput57), 
        .A(n4462), .ZN(n4467) );
  XNOR2_X1 U5510 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .B(keyinput7), .ZN(n4465)
         );
  XNOR2_X1 U5511 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .B(keyinput26), .ZN(n4464)
         );
  XNOR2_X1 U5512 ( .A(keyinput2), .B(UWORD_REG_7__SCAN_IN), .ZN(n4463) );
  NAND3_X1 U5513 ( .A1(n4465), .A2(n4464), .A3(n4463), .ZN(n4466) );
  NOR2_X1 U5514 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  AND2_X1 U5515 ( .A1(n4469), .A2(n4468), .ZN(n4481) );
  INV_X1 U5516 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5517 ( .A1(n4472), .A2(keyinput0), .B1(keyinput100), .B2(n4471), 
        .ZN(n4470) );
  OAI221_X1 U5518 ( .B1(n4472), .B2(keyinput0), .C1(n4471), .C2(keyinput100), 
        .A(n4470), .ZN(n4479) );
  INV_X1 U5519 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4474) );
  INV_X1 U5520 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4536) );
  AOI22_X1 U5521 ( .A1(n4474), .A2(keyinput9), .B1(keyinput101), .B2(n4536), 
        .ZN(n4473) );
  OAI221_X1 U5522 ( .B1(n4474), .B2(keyinput9), .C1(n4536), .C2(keyinput101), 
        .A(n4473), .ZN(n4478) );
  XNOR2_X1 U5523 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .B(keyinput90), .ZN(n4476)
         );
  XNOR2_X1 U5524 ( .A(keyinput66), .B(REIP_REG_10__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U5525 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  NOR3_X1 U5526 ( .A1(n4479), .A2(n4478), .A3(n4477), .ZN(n4480) );
  AND4_X1 U5527 ( .A1(n4483), .A2(n4482), .A3(n4481), .A4(n4480), .ZN(n4484)
         );
  NAND4_X1 U5528 ( .A1(n4487), .A2(n4486), .A3(n4485), .A4(n4484), .ZN(n4488)
         );
  NOR4_X1 U5529 ( .A1(n4491), .A2(n4490), .A3(n4489), .A4(n4488), .ZN(n4551)
         );
  NOR2_X1 U5530 ( .A1(n6892), .A2(n6888), .ZN(n5537) );
  NOR2_X1 U5531 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6093) );
  NAND4_X1 U5532 ( .A1(n4492), .A2(n5537), .A3(n6093), .A4(n5854), .ZN(n4507)
         );
  NAND4_X1 U5533 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(
        INSTQUEUE_REG_2__5__SCAN_IN), .A3(INSTQUEUE_REG_15__5__SCAN_IN), .A4(
        n4493), .ZN(n4506) );
  NAND4_X1 U5534 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(
        INSTQUEUE_REG_11__2__SCAN_IN), .A3(INSTQUEUE_REG_7__5__SCAN_IN), .A4(
        n4494), .ZN(n4505) );
  NOR4_X1 U5535 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(READY_N), .A3(n4495), 
        .A4(n6080), .ZN(n4503) );
  NOR4_X1 U5536 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(
        INSTQUEUE_REG_10__4__SCAN_IN), .A3(INSTQUEUE_REG_9__0__SCAN_IN), .A4(
        n4496), .ZN(n4502) );
  NOR4_X1 U5537 ( .A1(STATE2_REG_1__SCAN_IN), .A2(REIP_REG_24__SCAN_IN), .A3(
        INSTQUEUE_REG_3__1__SCAN_IN), .A4(n4497), .ZN(n4499) );
  NAND3_X1 U5538 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4499), .A3(
        INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4500) );
  NOR3_X1 U5539 ( .A1(n4500), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .A3(
        INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4501) );
  NAND3_X1 U5540 ( .A1(n4503), .A2(n4502), .A3(n4501), .ZN(n4504) );
  NOR4_X1 U5541 ( .A1(n4507), .A2(n4506), .A3(n4505), .A4(n4504), .ZN(n4518)
         );
  NOR4_X1 U5542 ( .A1(ADDRESS_REG_3__SCAN_IN), .A2(UWORD_REG_10__SCAN_IN), 
        .A3(DATAO_REG_1__SCAN_IN), .A4(BS16_N), .ZN(n4517) );
  NOR4_X1 U5543 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(ADDRESS_REG_14__SCAN_IN), 
        .A3(ADDRESS_REG_8__SCAN_IN), .A4(ADDRESS_REG_5__SCAN_IN), .ZN(n4516)
         );
  NOR4_X1 U5544 ( .A1(DATAI_25_), .A2(REIP_REG_21__SCAN_IN), .A3(
        PHYADDRPOINTER_REG_15__SCAN_IN), .A4(n6854), .ZN(n4508) );
  NAND3_X1 U5545 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(n4508), .A3(n6880), .ZN(
        n4514) );
  NOR4_X1 U5546 ( .A1(UWORD_REG_2__SCAN_IN), .A2(EBX_REG_26__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .A4(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4512)
         );
  NOR4_X1 U5547 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .A3(UWORD_REG_11__SCAN_IN), .A4(
        UWORD_REG_7__SCAN_IN), .ZN(n4511) );
  NOR4_X1 U5548 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .A3(PHYADDRPOINTER_REG_23__SCAN_IN), 
        .A4(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4510) );
  NOR4_X1 U5549 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(INSTADDRPOINTER_REG_31__SCAN_IN), .A4(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n4509) );
  NAND4_X1 U5550 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n4513)
         );
  NOR4_X1 U5551 ( .A1(EAX_REG_21__SCAN_IN), .A2(EAX_REG_24__SCAN_IN), .A3(
        n4514), .A4(n4513), .ZN(n4515) );
  NAND4_X1 U5552 ( .A1(n4518), .A2(n4517), .A3(n4516), .A4(n4515), .ZN(n4549)
         );
  NOR4_X1 U5553 ( .A1(DATAO_REG_13__SCAN_IN), .A2(BE_N_REG_1__SCAN_IN), .A3(
        BE_N_REG_0__SCAN_IN), .A4(ADDRESS_REG_27__SCAN_IN), .ZN(n4526) );
  NAND4_X1 U5554 ( .A1(DATAO_REG_30__SCAN_IN), .A2(DATAWIDTH_REG_30__SCAN_IN), 
        .A3(BYTEENABLE_REG_2__SCAN_IN), .A4(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4523) );
  NAND4_X1 U5555 ( .A1(DATAO_REG_16__SCAN_IN), .A2(DATAO_REG_12__SCAN_IN), 
        .A3(DATAO_REG_29__SCAN_IN), .A4(DATAO_REG_28__SCAN_IN), .ZN(n4522) );
  NAND4_X1 U5556 ( .A1(LWORD_REG_0__SCAN_IN), .A2(UWORD_REG_4__SCAN_IN), .A3(
        UWORD_REG_8__SCAN_IN), .A4(LWORD_REG_4__SCAN_IN), .ZN(n4521) );
  NAND4_X1 U5557 ( .A1(EAX_REG_4__SCAN_IN), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .A3(UWORD_REG_6__SCAN_IN), .A4(LWORD_REG_9__SCAN_IN), .ZN(n4520) );
  NOR4_X1 U5558 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4524)
         );
  NAND3_X1 U5559 ( .A1(n4526), .A2(n4525), .A3(n4524), .ZN(n4548) );
  NOR4_X1 U5560 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4528), .A3(n4527), 
        .A4(n6473), .ZN(n4535) );
  NOR4_X1 U5561 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(
        INSTQUEUE_REG_8__7__SCAN_IN), .A3(INSTQUEUE_REG_12__3__SCAN_IN), .A4(
        n4529), .ZN(n4534) );
  NOR4_X1 U5562 ( .A1(EBX_REG_12__SCAN_IN), .A2(EBX_REG_4__SCAN_IN), .A3(
        EBX_REG_2__SCAN_IN), .A4(n5588), .ZN(n4533) );
  NOR4_X1 U5563 ( .A1(EBX_REG_23__SCAN_IN), .A2(n4531), .A3(n6501), .A4(n4530), 
        .ZN(n4532) );
  NAND4_X1 U5564 ( .A1(n4535), .A2(n4534), .A3(n4533), .A4(n4532), .ZN(n4546)
         );
  NAND4_X1 U5565 ( .A1(DATAI_14_), .A2(DATAI_29_), .A3(ADDRESS_REG_20__SCAN_IN), .A4(DATAO_REG_2__SCAN_IN), .ZN(n4545) );
  NAND4_X1 U5566 ( .A1(ADS_N_REG_SCAN_IN), .A2(ADDRESS_REG_23__SCAN_IN), .A3(
        DATAO_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U5567 ( .A1(n4343), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4537) );
  NOR4_X1 U5568 ( .A1(n4538), .A2(n4537), .A3(n4536), .A4(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4542) );
  INV_X1 U5569 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4540) );
  NAND4_X1 U5570 ( .A1(EBX_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(REIP_REG_1__SCAN_IN), .A4(
        PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4539) );
  NOR3_X1 U5571 ( .A1(n4540), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .A3(n4539), 
        .ZN(n4541) );
  NAND4_X1 U5572 ( .A1(n4542), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .A3(n4541), 
        .A4(n4375), .ZN(n4544) );
  NAND4_X1 U5573 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        EBX_REG_25__SCAN_IN), .A3(REIP_REG_22__SCAN_IN), .A4(
        REIP_REG_15__SCAN_IN), .ZN(n4543) );
  OR4_X1 U5574 ( .A1(n4546), .A2(n4545), .A3(n4544), .A4(n4543), .ZN(n4547) );
  NOR3_X1 U5575 ( .A1(n4549), .A2(n4548), .A3(n4547), .ZN(n4550) );
  XNOR2_X1 U5576 ( .A(n4551), .B(n4550), .ZN(n4552) );
  XNOR2_X1 U5577 ( .A(n4553), .B(n4552), .ZN(U2994) );
  INV_X1 U5578 ( .A(n4650), .ZN(n5921) );
  NAND2_X1 U5579 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5915) );
  AOI21_X1 U5580 ( .B1(n4555), .B2(n5915), .A(n4554), .ZN(n6508) );
  OAI21_X1 U5581 ( .B1(n6492), .B2(n6494), .A(n6508), .ZN(n4556) );
  INV_X1 U5582 ( .A(n4556), .ZN(n6491) );
  OAI21_X1 U5583 ( .B1(n5921), .B2(n6467), .A(n6491), .ZN(n4557) );
  INV_X1 U5584 ( .A(n4557), .ZN(n6472) );
  AOI221_X1 U5585 ( .B1(n6479), .B2(n4558), .C1(n5914), .C2(n4558), .A(n6472), 
        .ZN(n4570) );
  CLKBUF_X1 U5586 ( .A(n4559), .Z(n4989) );
  OR2_X1 U5587 ( .A1(n4561), .A2(n4560), .ZN(n4562) );
  NAND2_X1 U5588 ( .A1(n4989), .A2(n4562), .ZN(n6411) );
  NOR2_X1 U5589 ( .A1(n6411), .A2(n6476), .ZN(n4569) );
  NOR4_X1 U5590 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6500), .A3(n6479), 
        .A4(n5915), .ZN(n4568) );
  OR2_X1 U5591 ( .A1(n4715), .A2(n4564), .ZN(n4565) );
  NAND2_X1 U5592 ( .A1(n4563), .A2(n4565), .ZN(n6218) );
  INV_X1 U5593 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4566) );
  OAI22_X1 U5594 ( .A1(n6497), .A2(n6218), .B1(n6495), .B2(n4566), .ZN(n4567)
         );
  OR4_X1 U5595 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(U3013) );
  OR2_X1 U5596 ( .A1(n4635), .A2(n5303), .ZN(n4574) );
  NOR2_X1 U5597 ( .A1(n4571), .A2(n4578), .ZN(n4586) );
  INV_X1 U5598 ( .A(n4586), .ZN(n4572) );
  NAND2_X1 U5599 ( .A1(n4572), .A2(n4587), .ZN(n4573) );
  AND2_X1 U5600 ( .A1(n4574), .A2(n4573), .ZN(n6082) );
  OR2_X1 U5601 ( .A1(n5310), .A2(n4596), .ZN(n4593) );
  NAND2_X1 U5602 ( .A1(n4593), .A2(n6824), .ZN(n4575) );
  NAND2_X1 U5603 ( .A1(n4575), .A2(n6827), .ZN(n6939) );
  NAND2_X1 U5604 ( .A1(n6082), .A2(n6939), .ZN(n6781) );
  AND2_X1 U5605 ( .A1(n6781), .A2(n6802), .ZN(n6091) );
  INV_X1 U5606 ( .A(MORE_REG_SCAN_IN), .ZN(n4585) );
  AND2_X1 U5607 ( .A1(n4576), .A2(n4587), .ZN(n4577) );
  OR2_X1 U5608 ( .A1(n4635), .A2(n4577), .ZN(n4582) );
  NAND2_X1 U5609 ( .A1(n4635), .A2(n4757), .ZN(n4581) );
  NAND2_X1 U5610 ( .A1(n4579), .A2(n4578), .ZN(n4580) );
  AND3_X1 U5611 ( .A1(n4582), .A2(n4581), .A3(n4580), .ZN(n6779) );
  INV_X1 U5612 ( .A(n6779), .ZN(n4583) );
  NAND2_X1 U5613 ( .A1(n6091), .A2(n4583), .ZN(n4584) );
  OAI21_X1 U5614 ( .B1(n6091), .B2(n4585), .A(n4584), .ZN(U3471) );
  NAND2_X1 U5615 ( .A1(n4586), .A2(n6802), .ZN(n4589) );
  NAND2_X1 U5616 ( .A1(n4594), .A2(n6085), .ZN(n4591) );
  AOI21_X1 U5617 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n4589), .A(n4591), .ZN(
        n4588) );
  INV_X1 U5618 ( .A(n4588), .ZN(U2788) );
  INV_X1 U5619 ( .A(n4589), .ZN(n4590) );
  NOR3_X1 U5620 ( .A1(n4591), .A2(n4590), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n4592) );
  AOI21_X1 U5621 ( .B1(n6936), .B2(n4593), .A(n4592), .ZN(U3474) );
  INV_X1 U5622 ( .A(n4594), .ZN(n4595) );
  OAI21_X1 U5623 ( .B1(n4596), .B2(n6827), .A(n4595), .ZN(n6375) );
  INV_X1 U5624 ( .A(n6375), .ZN(n6334) );
  OR2_X1 U5625 ( .A1(n4658), .A2(n4597), .ZN(n6385) );
  INV_X2 U5626 ( .A(n6385), .ZN(n6378) );
  OR3_X2 U5627 ( .A1(n4658), .A2(READY_N), .A3(n4629), .ZN(n6380) );
  INV_X1 U5628 ( .A(DATAI_9_), .ZN(n5056) );
  NOR2_X1 U5629 ( .A1(n6380), .A2(n5056), .ZN(n6343) );
  AOI21_X1 U5630 ( .B1(n6378), .B2(EAX_REG_9__SCAN_IN), .A(n6343), .ZN(n4598)
         );
  OAI21_X1 U5631 ( .B1(n6334), .B2(n6312), .A(n4598), .ZN(U2948) );
  INV_X1 U5632 ( .A(DATAI_8_), .ZN(n4599) );
  NOR2_X1 U5633 ( .A1(n6380), .A2(n4599), .ZN(n6365) );
  AOI21_X1 U5634 ( .B1(n6378), .B2(EAX_REG_24__SCAN_IN), .A(n6365), .ZN(n4600)
         );
  OAI21_X1 U5635 ( .B1(n6334), .B2(n4601), .A(n4600), .ZN(U2932) );
  INV_X1 U5636 ( .A(DATAI_10_), .ZN(n4602) );
  NOR2_X1 U5637 ( .A1(n6380), .A2(n4602), .ZN(n6368) );
  AOI21_X1 U5638 ( .B1(n6378), .B2(EAX_REG_26__SCAN_IN), .A(n6368), .ZN(n4603)
         );
  OAI21_X1 U5639 ( .B1(n6334), .B2(n6289), .A(n4603), .ZN(U2934) );
  INV_X1 U5640 ( .A(DATAI_11_), .ZN(n5153) );
  INV_X1 U5641 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4604) );
  OAI222_X1 U5642 ( .A1(n5153), .A2(n6380), .B1(n6334), .B2(n6287), .C1(n4604), 
        .C2(n6385), .ZN(U2935) );
  XOR2_X1 U5643 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .B(n4605), .Z(n4676) );
  NAND2_X1 U5644 ( .A1(n4607), .A2(n4606), .ZN(n4608) );
  NAND2_X1 U5645 ( .A1(n4609), .A2(n4608), .ZN(n6278) );
  NAND2_X1 U5646 ( .A1(n6483), .A2(REIP_REG_0__SCAN_IN), .ZN(n4673) );
  OAI21_X1 U5647 ( .B1(n6278), .B2(n6696), .A(n4673), .ZN(n4613) );
  INV_X1 U5648 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4610) );
  AOI21_X1 U5649 ( .B1(n5800), .B2(n4611), .A(n4610), .ZN(n4612) );
  AOI211_X1 U5650 ( .C1(n6429), .C2(n4676), .A(n4613), .B(n4612), .ZN(n4614)
         );
  INV_X1 U5651 ( .A(n4614), .ZN(U2986) );
  INV_X1 U5652 ( .A(n4615), .ZN(n4628) );
  NAND2_X1 U5653 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5500) );
  AOI22_X1 U5654 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4616), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6501), .ZN(n5499) );
  INV_X1 U5655 ( .A(n5499), .ZN(n4627) );
  INV_X1 U5656 ( .A(n6906), .ZN(n6918) );
  INV_X1 U5657 ( .A(n4618), .ZN(n4898) );
  AND4_X1 U5658 ( .A1(n4636), .A2(n4621), .A3(n4620), .A4(n4619), .ZN(n4622)
         );
  AND2_X1 U5659 ( .A1(n4623), .A2(n4622), .ZN(n6757) );
  NOR3_X1 U5660 ( .A1(n6756), .A2(n3112), .A3(n4760), .ZN(n4624) );
  AOI21_X1 U5661 ( .B1(n6755), .B2(n3328), .A(n4624), .ZN(n4625) );
  OAI21_X1 U5662 ( .B1(n4898), .B2(n6757), .A(n4625), .ZN(n6761) );
  INV_X1 U5663 ( .A(n6761), .ZN(n4626) );
  OAI222_X1 U5664 ( .A1(n6797), .A2(n4628), .B1(n5500), .B2(n4627), .C1(n6918), 
        .C2(n4626), .ZN(n4645) );
  INV_X1 U5665 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6904) );
  AOI21_X1 U5666 ( .B1(n4629), .B2(n6824), .A(READY_N), .ZN(n4630) );
  OAI211_X1 U5667 ( .C1(n6790), .C2(n6755), .A(n4635), .B(n4630), .ZN(n4633)
         );
  NAND2_X1 U5668 ( .A1(n5310), .A2(n4939), .ZN(n4631) );
  NAND3_X1 U5669 ( .A1(n4633), .A2(n4632), .A3(n4631), .ZN(n4640) );
  INV_X1 U5670 ( .A(n4758), .ZN(n4634) );
  NAND2_X1 U5671 ( .A1(n4635), .A2(n4634), .ZN(n4639) );
  INV_X1 U5672 ( .A(n4636), .ZN(n6076) );
  NAND2_X1 U5673 ( .A1(n6076), .A2(n4637), .ZN(n4638) );
  NAND2_X1 U5674 ( .A1(n4639), .A2(n4638), .ZN(n4703) );
  NOR2_X1 U5675 ( .A1(n4640), .A2(n4703), .ZN(n4644) );
  INV_X1 U5676 ( .A(n4641), .ZN(n4643) );
  NAND2_X1 U5677 ( .A1(n4643), .A2(n4642), .ZN(n4684) );
  NAND2_X1 U5678 ( .A1(n4644), .A2(n4684), .ZN(n6762) );
  NOR2_X1 U5679 ( .A1(n6912), .A2(n6937), .ZN(n4801) );
  NAND2_X1 U5680 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4801), .ZN(n6902) );
  INV_X1 U5681 ( .A(n6902), .ZN(n6795) );
  AOI22_X1 U5682 ( .A1(n6762), .A2(n6802), .B1(FLUSH_REG_SCAN_IN), .B2(n6795), 
        .ZN(n6074) );
  OAI21_X1 U5683 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6904), .A(n6074), .ZN(
        n6916) );
  OAI21_X1 U5684 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6797), .A(n6916), 
        .ZN(n6914) );
  AOI22_X1 U5685 ( .A1(n4645), .A2(n6916), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n6914), .ZN(n4646) );
  INV_X1 U5686 ( .A(n4646), .ZN(U3460) );
  XNOR2_X1 U5687 ( .A(n4647), .B(n4648), .ZN(n4977) );
  NAND3_X1 U5688 ( .A1(n4650), .A2(n4649), .A3(n6501), .ZN(n4656) );
  OAI21_X1 U5689 ( .B1(n4651), .B2(n5179), .A(n4652), .ZN(n4694) );
  NOR2_X1 U5690 ( .A1(n6495), .A2(n6921), .ZN(n4972) );
  NAND2_X1 U5691 ( .A1(n6492), .A2(n4653), .ZN(n5378) );
  NAND2_X1 U5692 ( .A1(n5378), .A2(n4670), .ZN(n4677) );
  AOI21_X1 U5693 ( .B1(n4671), .B2(n4677), .A(n6501), .ZN(n4654) );
  AOI211_X1 U5694 ( .C1(n6485), .C2(n4694), .A(n4972), .B(n4654), .ZN(n4655)
         );
  OAI211_X1 U5695 ( .C1(n4977), .C2(n6476), .A(n4656), .B(n4655), .ZN(U3017)
         );
  INV_X1 U5696 ( .A(n6755), .ZN(n4657) );
  OR2_X1 U5697 ( .A1(n4658), .A2(n4657), .ZN(n4659) );
  NAND2_X1 U5698 ( .A1(n6385), .A2(n4659), .ZN(n4660) );
  NAND2_X1 U5699 ( .A1(n6323), .A2(n5184), .ZN(n6279) );
  NAND2_X1 U5700 ( .A1(n6809), .A2(n4801), .ZN(n6328) );
  INV_X1 U5701 ( .A(n6328), .ZN(n6932) );
  AOI22_X1 U5702 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6932), .B1(n6330), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4661) );
  OAI21_X1 U5703 ( .B1(n4662), .B2(n6279), .A(n4661), .ZN(U2899) );
  INV_X1 U5704 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5705 ( .A1(n6932), .A2(UWORD_REG_3__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4663) );
  OAI21_X1 U5706 ( .B1(n4664), .B2(n6279), .A(n4663), .ZN(U2904) );
  INV_X1 U5707 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6345) );
  AOI22_X1 U5708 ( .A1(n6932), .A2(UWORD_REG_9__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4665) );
  OAI21_X1 U5709 ( .B1(n6345), .B2(n6279), .A(n4665), .ZN(U2898) );
  INV_X1 U5710 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4667) );
  AOI22_X1 U5711 ( .A1(n6932), .A2(UWORD_REG_1__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4666) );
  OAI21_X1 U5712 ( .B1(n4667), .B2(n6279), .A(n4666), .ZN(U2906) );
  AOI22_X1 U5713 ( .A1(n6932), .A2(UWORD_REG_5__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4668) );
  OAI21_X1 U5714 ( .B1(n4669), .B2(n6279), .A(n4668), .ZN(U2902) );
  AOI21_X1 U5715 ( .B1(n4671), .B2(n5380), .A(n4670), .ZN(n4675) );
  OAI21_X1 U5716 ( .B1(n5521), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4672), 
        .ZN(n5593) );
  OAI21_X1 U5717 ( .B1(n6497), .B2(n5593), .A(n4673), .ZN(n4674) );
  AOI211_X1 U5718 ( .C1(n6503), .C2(n4676), .A(n4675), .B(n4674), .ZN(n4678)
         );
  NAND2_X1 U5719 ( .A1(n4678), .A2(n4677), .ZN(U3018) );
  OR2_X1 U5720 ( .A1(n4679), .A2(n5686), .ZN(n4700) );
  INV_X1 U5721 ( .A(n4700), .ZN(n4682) );
  NAND4_X1 U5722 ( .A1(n4682), .A2(n4948), .A3(n4681), .A4(n4680), .ZN(n4683)
         );
  NAND2_X1 U5723 ( .A1(n4684), .A2(n4683), .ZN(n4685) );
  AND2_X2 U5724 ( .A1(n4685), .A2(n6802), .ZN(n6261) );
  NAND2_X1 U5725 ( .A1(n6261), .A2(n5682), .ZN(n5663) );
  OAI222_X1 U5726 ( .A1(n6278), .A2(n6014), .B1(n5588), .B2(n6261), .C1(n5593), 
        .C2(n5663), .ZN(U2859) );
  XNOR2_X1 U5727 ( .A(n4748), .B(n4711), .ZN(n6420) );
  OAI21_X1 U5728 ( .B1(n4686), .B2(n5336), .A(n4687), .ZN(n4688) );
  AND2_X1 U5729 ( .A1(n4688), .A2(n4714), .ZN(n6484) );
  INV_X1 U5730 ( .A(n6261), .ZN(n5680) );
  AOI22_X1 U5731 ( .A1(n6257), .A2(n6484), .B1(EBX_REG_3__SCAN_IN), .B2(n5680), 
        .ZN(n4689) );
  OAI21_X1 U5732 ( .B1(n6420), .B2(n6014), .A(n4689), .ZN(U2856) );
  OR2_X1 U5733 ( .A1(n4691), .A2(n4690), .ZN(n4692) );
  NAND2_X1 U5734 ( .A1(n4693), .A2(n4692), .ZN(n5587) );
  AOI22_X1 U5735 ( .A1(n6257), .A2(n4694), .B1(EBX_REG_1__SCAN_IN), .B2(n5680), 
        .ZN(n4695) );
  OAI21_X1 U5736 ( .B1(n6014), .B2(n5587), .A(n4695), .ZN(U2858) );
  INV_X1 U5737 ( .A(n4696), .ZN(n4697) );
  OR2_X1 U5738 ( .A1(n4698), .A2(n4697), .ZN(n4701) );
  NOR3_X1 U5739 ( .A1(n4701), .A2(n4700), .A3(n4699), .ZN(n4702) );
  OAI21_X1 U5740 ( .B1(n4703), .B2(n4702), .A(n6802), .ZN(n4704) );
  NAND2_X1 U5741 ( .A1(n4705), .A2(n5686), .ZN(n4707) );
  INV_X1 U5742 ( .A(n4754), .ZN(n4706) );
  XNOR2_X1 U5743 ( .A(n4709), .B(n4706), .ZN(n6409) );
  INV_X1 U5744 ( .A(n4707), .ZN(n4708) );
  NAND2_X1 U5745 ( .A1(n6276), .A2(n4708), .ZN(n6275) );
  INV_X1 U5746 ( .A(DATAI_5_), .ZN(n6360) );
  OAI222_X1 U5747 ( .A1(n6277), .A2(n6409), .B1(n6275), .B2(n6360), .C1(n6276), 
        .C2(n3832), .ZN(U2886) );
  INV_X1 U5748 ( .A(n4709), .ZN(n4755) );
  AOI21_X1 U5749 ( .B1(n4748), .B2(n4711), .A(n4710), .ZN(n4712) );
  NOR2_X1 U5750 ( .A1(n4755), .A2(n4712), .ZN(n4986) );
  INV_X1 U5751 ( .A(n4986), .ZN(n5318) );
  AND2_X1 U5752 ( .A1(n4714), .A2(n4713), .ZN(n4716) );
  OR2_X1 U5753 ( .A1(n4716), .A2(n4715), .ZN(n6477) );
  OAI222_X1 U5754 ( .A1(n5318), .A2(n6014), .B1(n6261), .B2(n5305), .C1(n6477), 
        .C2(n5663), .ZN(U2855) );
  INV_X1 U5755 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4717) );
  OAI222_X1 U5756 ( .A1(n6218), .A2(n5663), .B1(n6014), .B2(n6409), .C1(n4717), 
        .C2(n6261), .ZN(U2854) );
  NAND2_X1 U5757 ( .A1(n5258), .A2(n6583), .ZN(n4720) );
  AOI21_X1 U5758 ( .B1(n4729), .B2(STATEBS16_REG_SCAN_IN), .A(n6934), .ZN(
        n4731) );
  INV_X1 U5759 ( .A(n6553), .ZN(n4723) );
  AND2_X1 U5760 ( .A1(n4722), .A2(n4898), .ZN(n6511) );
  NAND3_X1 U5761 ( .A1(n4723), .A2(n6653), .A3(n6511), .ZN(n4724) );
  NAND3_X1 U5762 ( .A1(n6777), .A2(n6770), .A3(n6764), .ZN(n6510) );
  OR2_X1 U5763 ( .A1(n6759), .A2(n6510), .ZN(n5132) );
  NAND2_X1 U5764 ( .A1(n4724), .A2(n5132), .ZN(n4733) );
  INV_X1 U5765 ( .A(n6510), .ZN(n4725) );
  AOI22_X1 U5766 ( .A1(n4731), .A2(n4733), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4725), .ZN(n5138) );
  INV_X1 U5767 ( .A(DATAI_1_), .ZN(n6352) );
  NAND2_X1 U5768 ( .A1(n6912), .A2(n6937), .ZN(n6810) );
  INV_X1 U5769 ( .A(n6810), .ZN(n6940) );
  NOR2_X2 U5770 ( .A1(n6352), .A2(n5024), .ZN(n6708) );
  INV_X1 U5771 ( .A(n6708), .ZN(n5274) );
  AND2_X1 U5772 ( .A1(n3085), .A2(DATAI_17_), .ZN(n6710) );
  NOR2_X2 U5773 ( .A1(n4726), .A2(n6551), .ZN(n6577) );
  NAND3_X1 U5774 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6809), .A3(n4727), .ZN(
        n4949) );
  NOR2_X2 U5775 ( .A1(n4949), .A2(n4728), .ZN(n6709) );
  INV_X1 U5776 ( .A(n6709), .ZN(n4915) );
  AND2_X1 U5777 ( .A1(n3085), .A2(DATAI_25_), .ZN(n6622) );
  INV_X1 U5778 ( .A(n6622), .ZN(n6713) );
  NAND2_X1 U5779 ( .A1(n4729), .A2(n6551), .ZN(n6512) );
  OAI22_X1 U5780 ( .A1(n4915), .A2(n5132), .B1(n6713), .B2(n6512), .ZN(n4730)
         );
  AOI21_X1 U5781 ( .B1(n6710), .B2(n6577), .A(n4730), .ZN(n4736) );
  INV_X1 U5782 ( .A(n4731), .ZN(n4734) );
  OAI21_X1 U5783 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6904), .A(n4905), 
        .ZN(n6655) );
  AOI21_X1 U5784 ( .B1(n6934), .B2(n6510), .A(n6655), .ZN(n4732) );
  OAI21_X1 U5785 ( .B1(n4734), .B2(n4733), .A(n4732), .ZN(n5135) );
  NAND2_X1 U5786 ( .A1(n5135), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4735) );
  OAI211_X1 U5787 ( .C1(n5138), .C2(n5274), .A(n4736), .B(n4735), .ZN(U3029)
         );
  INV_X1 U5788 ( .A(DATAI_3_), .ZN(n6356) );
  NOR2_X2 U5789 ( .A1(n6356), .A2(n5024), .ZN(n6720) );
  INV_X1 U5790 ( .A(n6720), .ZN(n5294) );
  AND2_X1 U5791 ( .A1(n3085), .A2(DATAI_19_), .ZN(n6722) );
  NOR2_X2 U5792 ( .A1(n4949), .A2(n4737), .ZN(n6721) );
  INV_X1 U5793 ( .A(n6721), .ZN(n4911) );
  NAND2_X1 U5794 ( .A1(n3085), .A2(DATAI_27_), .ZN(n6725) );
  OAI22_X1 U5795 ( .A1(n4911), .A2(n5132), .B1(n6725), .B2(n6512), .ZN(n4738)
         );
  AOI21_X1 U5796 ( .B1(n6722), .B2(n6577), .A(n4738), .ZN(n4740) );
  NAND2_X1 U5797 ( .A1(n5135), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4739) );
  OAI211_X1 U5798 ( .C1(n5138), .C2(n5294), .A(n4740), .B(n4739), .ZN(U3031)
         );
  INV_X1 U5799 ( .A(DATAI_7_), .ZN(n6364) );
  NOR2_X2 U5800 ( .A1(n6364), .A2(n5024), .ZN(n6745) );
  INV_X1 U5801 ( .A(n6745), .ZN(n5278) );
  AND2_X1 U5802 ( .A1(n3085), .A2(DATAI_23_), .ZN(n6749) );
  NOR2_X2 U5803 ( .A1(n4949), .A2(n5682), .ZN(n6747) );
  INV_X1 U5804 ( .A(n6747), .ZN(n4919) );
  NAND2_X1 U5805 ( .A1(n3085), .A2(DATAI_31_), .ZN(n6754) );
  OAI22_X1 U5806 ( .A1(n4919), .A2(n5132), .B1(n6754), .B2(n6512), .ZN(n4741)
         );
  AOI21_X1 U5807 ( .B1(n6749), .B2(n6577), .A(n4741), .ZN(n4743) );
  NAND2_X1 U5808 ( .A1(n5135), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4742) );
  OAI211_X1 U5809 ( .C1(n5138), .C2(n5278), .A(n4743), .B(n4742), .ZN(U3035)
         );
  INV_X1 U5810 ( .A(DATAI_0_), .ZN(n6350) );
  NOR2_X2 U5811 ( .A1(n6350), .A2(n5024), .ZN(n6693) );
  INV_X1 U5812 ( .A(n6693), .ZN(n5270) );
  AND2_X1 U5813 ( .A1(n3085), .A2(DATAI_16_), .ZN(n6704) );
  NOR2_X2 U5814 ( .A1(n4949), .A2(n4744), .ZN(n6692) );
  INV_X1 U5815 ( .A(n6692), .ZN(n4901) );
  NAND2_X1 U5816 ( .A1(n3085), .A2(DATAI_24_), .ZN(n6707) );
  OAI22_X1 U5817 ( .A1(n4901), .A2(n5132), .B1(n6707), .B2(n6512), .ZN(n4745)
         );
  AOI21_X1 U5818 ( .B1(n6704), .B2(n6577), .A(n4745), .ZN(n4747) );
  NAND2_X1 U5819 ( .A1(n5135), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4746) );
  OAI211_X1 U5820 ( .C1(n5138), .C2(n5270), .A(n4747), .B(n4746), .ZN(U3028)
         );
  INV_X1 U5821 ( .A(n4748), .ZN(n4749) );
  OAI21_X1 U5822 ( .B1(n4751), .B2(n4750), .A(n4749), .ZN(n6255) );
  INV_X1 U5823 ( .A(n6275), .ZN(n6271) );
  AOI22_X1 U5824 ( .A1(n6271), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n6267), .ZN(n4752) );
  OAI21_X1 U5825 ( .B1(n6255), .B2(n6277), .A(n4752), .ZN(U2889) );
  AOI21_X1 U5826 ( .B1(n4755), .B2(n4754), .A(n4753), .ZN(n4756) );
  OR2_X1 U5827 ( .A1(n4756), .A2(n4998), .ZN(n5257) );
  INV_X1 U5828 ( .A(DATAI_6_), .ZN(n6362) );
  INV_X1 U5829 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6317) );
  OAI222_X1 U5830 ( .A1(n5257), .A2(n6277), .B1(n6275), .B2(n6362), .C1(n6276), 
        .C2(n6317), .ZN(U2885) );
  OR2_X1 U5831 ( .A1(n6762), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4769)
         );
  OR2_X1 U5832 ( .A1(n4722), .A2(n6757), .ZN(n4767) );
  INV_X1 U5833 ( .A(n4757), .ZN(n4759) );
  NAND2_X1 U5834 ( .A1(n4759), .A2(n4758), .ZN(n4774) );
  INV_X1 U5835 ( .A(n4760), .ZN(n5498) );
  NAND2_X1 U5836 ( .A1(n5498), .A2(n5505), .ZN(n4772) );
  NAND2_X1 U5837 ( .A1(n4760), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U5838 ( .A1(n4772), .A2(n4776), .ZN(n4761) );
  NAND2_X1 U5839 ( .A1(n4774), .A2(n4761), .ZN(n4765) );
  XNOR2_X1 U5840 ( .A(n5505), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4763)
         );
  INV_X1 U5841 ( .A(n4761), .ZN(n4762) );
  AOI22_X1 U5842 ( .A1(n6755), .A2(n4763), .B1(n4778), .B2(n4762), .ZN(n4764)
         );
  AND2_X1 U5843 ( .A1(n4765), .A2(n4764), .ZN(n4766) );
  AND2_X1 U5844 ( .A1(n4767), .A2(n4766), .ZN(n5501) );
  NAND2_X1 U5845 ( .A1(n6762), .A2(n5501), .ZN(n4768) );
  NAND2_X1 U5846 ( .A1(n4769), .A2(n4768), .ZN(n6768) );
  INV_X1 U5847 ( .A(n6768), .ZN(n4786) );
  OR2_X1 U5848 ( .A1(n6762), .A2(n4771), .ZN(n4785) );
  INV_X1 U5849 ( .A(n6757), .ZN(n4770) );
  NAND2_X1 U5850 ( .A1(n6553), .A2(n4770), .ZN(n4783) );
  XNOR2_X1 U5851 ( .A(n4772), .B(n4771), .ZN(n4773) );
  NAND2_X1 U5852 ( .A1(n4774), .A2(n4773), .ZN(n4781) );
  NAND2_X1 U5853 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4775) );
  XNOR2_X1 U5854 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4775), .ZN(n4779)
         );
  NAND2_X1 U5855 ( .A1(n4776), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U5856 ( .A1(n3261), .A2(n4777), .ZN(n6907) );
  AOI22_X1 U5857 ( .A1(n6755), .A2(n4779), .B1(n4778), .B2(n6907), .ZN(n4780)
         );
  AND2_X1 U5858 ( .A1(n4781), .A2(n4780), .ZN(n4782) );
  NAND2_X1 U5859 ( .A1(n4783), .A2(n4782), .ZN(n6905) );
  NAND2_X1 U5860 ( .A1(n6762), .A2(n6905), .ZN(n4784) );
  NAND2_X1 U5861 ( .A1(n4785), .A2(n4784), .ZN(n6776) );
  NAND3_X1 U5862 ( .A1(n4786), .A2(n6912), .A3(n6776), .ZN(n4790) );
  INV_X1 U5863 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6090) );
  NAND2_X1 U5864 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6090), .ZN(n4791) );
  INV_X1 U5865 ( .A(n4791), .ZN(n4787) );
  NAND2_X1 U5866 ( .A1(n4788), .A2(n4787), .ZN(n4789) );
  AND2_X1 U5867 ( .A1(n4790), .A2(n4789), .ZN(n6785) );
  INV_X1 U5868 ( .A(n6785), .ZN(n4799) );
  INV_X1 U5869 ( .A(n3112), .ZN(n4798) );
  OAI21_X1 U5870 ( .B1(n6762), .B2(STATE2_REG_1__SCAN_IN), .A(n4791), .ZN(
        n4792) );
  NAND2_X1 U5871 ( .A1(n4792), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4797) );
  INV_X1 U5872 ( .A(n5202), .ZN(n4793) );
  OR2_X1 U5873 ( .A1(n4794), .A2(n4793), .ZN(n4795) );
  XNOR2_X1 U5874 ( .A(n4795), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6075)
         );
  NAND3_X1 U5875 ( .A1(n6075), .A2(n6076), .A3(n6912), .ZN(n4796) );
  NAND2_X1 U5876 ( .A1(n4797), .A2(n4796), .ZN(n6783) );
  AOI21_X1 U5877 ( .B1(n4799), .B2(n4798), .A(n6783), .ZN(n6796) );
  AND2_X1 U5878 ( .A1(n6796), .A2(n6090), .ZN(n4800) );
  OAI21_X1 U5879 ( .B1(n4800), .B2(n6902), .A(n5024), .ZN(n6509) );
  INV_X1 U5880 ( .A(n6509), .ZN(n4923) );
  OR2_X1 U5881 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6912), .ZN(n4943) );
  AOI222_X1 U5882 ( .A1(n6796), .A2(n4801), .B1(n6653), .B2(n4943), .C1(n5259), 
        .C2(n6703), .ZN(n4803) );
  NAND2_X1 U5883 ( .A1(n4923), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4802) );
  OAI21_X1 U5884 ( .B1(n4923), .B2(n4803), .A(n4802), .ZN(U3465) );
  INV_X1 U5885 ( .A(DATAI_4_), .ZN(n6358) );
  OAI222_X1 U5886 ( .A1(n5318), .A2(n6277), .B1(n6275), .B2(n6358), .C1(n6276), 
        .C2(n4804), .ZN(U2887) );
  INV_X1 U5887 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6325) );
  OAI222_X1 U5888 ( .A1(n5587), .A2(n6277), .B1(n6275), .B2(n6352), .C1(n6276), 
        .C2(n6325), .ZN(U2890) );
  INV_X1 U5889 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6322) );
  OAI222_X1 U5890 ( .A1(n6420), .A2(n6277), .B1(n6275), .B2(n6356), .C1(n6276), 
        .C2(n6322), .ZN(U2888) );
  NAND2_X1 U5891 ( .A1(n4563), .A2(n4806), .ZN(n4807) );
  NAND2_X1 U5892 ( .A1(n4805), .A2(n4807), .ZN(n6469) );
  INV_X1 U5893 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4808) );
  OAI222_X1 U5894 ( .A1(n6469), .A2(n5663), .B1(n6261), .B2(n4808), .C1(n5257), 
        .C2(n6014), .ZN(U2853) );
  NAND3_X1 U5895 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6777), .A3(n6764), .ZN(n4869) );
  NOR2_X1 U5896 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4869), .ZN(n5095)
         );
  INV_X1 U5897 ( .A(n5095), .ZN(n4809) );
  NOR2_X1 U5898 ( .A1(n5347), .A2(n6937), .ZN(n6555) );
  INV_X1 U5899 ( .A(n5022), .ZN(n6554) );
  NOR2_X1 U5900 ( .A1(n6554), .A2(n5023), .ZN(n6518) );
  OAI21_X1 U5901 ( .B1(n6518), .B2(n6937), .A(n4905), .ZN(n6516) );
  AOI211_X1 U5902 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4809), .A(n6555), .B(
        n6516), .ZN(n4813) );
  NAND2_X1 U5903 ( .A1(n6583), .A2(n4960), .ZN(n4810) );
  NAND2_X1 U5904 ( .A1(n3097), .A2(n5259), .ZN(n6608) );
  OR2_X1 U5905 ( .A1(n6583), .A2(n4819), .ZN(n4959) );
  NOR2_X1 U5906 ( .A1(n4959), .A2(n4960), .ZN(n4873) );
  NAND2_X1 U5907 ( .A1(n4873), .A2(n6551), .ZN(n5143) );
  AOI21_X1 U5908 ( .B1(n6608), .B2(n5143), .A(n6089), .ZN(n4811) );
  OR2_X1 U5909 ( .A1(n4722), .A2(n4618), .ZN(n4821) );
  NOR2_X1 U5910 ( .A1(n4821), .A2(n5202), .ZN(n4862) );
  OR3_X1 U5911 ( .A1(n4811), .A2(n4862), .A3(n6934), .ZN(n4812) );
  NAND2_X1 U5912 ( .A1(n4813), .A2(n4812), .ZN(n5099) );
  INV_X1 U5913 ( .A(n5099), .ZN(n5088) );
  INV_X1 U5914 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4818) );
  OR2_X1 U5915 ( .A1(n6553), .A2(n6934), .ZN(n6521) );
  AND2_X1 U5916 ( .A1(n5347), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U5917 ( .A1(n6518), .A2(n6517), .ZN(n4814) );
  OAI21_X1 U5918 ( .B1(n6521), .B2(n4821), .A(n4814), .ZN(n5094) );
  INV_X1 U5919 ( .A(n5143), .ZN(n5084) );
  AOI22_X1 U5920 ( .A1(n6692), .A2(n5095), .B1(n5084), .B2(n6704), .ZN(n4815)
         );
  OAI21_X1 U5921 ( .B1(n6707), .B2(n6608), .A(n4815), .ZN(n4816) );
  AOI21_X1 U5922 ( .B1(n6693), .B2(n5094), .A(n4816), .ZN(n4817) );
  OAI21_X1 U5923 ( .B1(n5088), .B2(n4818), .A(n4817), .ZN(U3052) );
  INV_X1 U5924 ( .A(n6749), .ZN(n6582) );
  NOR2_X1 U5925 ( .A1(n6583), .A2(n4820), .ZN(n4900) );
  NAND2_X1 U5926 ( .A1(n4900), .A2(n5258), .ZN(n4826) );
  AND2_X1 U5927 ( .A1(n6553), .A2(n6653), .ZN(n6690) );
  INV_X1 U5928 ( .A(n4821), .ZN(n5207) );
  NAND3_X1 U5929 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6764), .ZN(n5203) );
  NOR2_X1 U5930 ( .A1(n6759), .A2(n5203), .ZN(n4950) );
  AOI21_X1 U5931 ( .B1(n6690), .B2(n5207), .A(n4950), .ZN(n4825) );
  INV_X1 U5932 ( .A(n4825), .ZN(n4823) );
  OR2_X1 U5933 ( .A1(n4826), .A2(n6089), .ZN(n4927) );
  NAND2_X1 U5934 ( .A1(n6703), .A2(n4927), .ZN(n4824) );
  AOI21_X1 U5935 ( .B1(n6934), .B2(n5203), .A(n6655), .ZN(n4822) );
  OAI21_X1 U5936 ( .B1(n4823), .B2(n4824), .A(n4822), .ZN(n4947) );
  OAI22_X1 U5937 ( .A1(n4825), .A2(n4824), .B1(n6937), .B2(n5203), .ZN(n4946)
         );
  AOI22_X1 U5938 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4947), .B1(n6745), 
        .B2(n4946), .ZN(n4828) );
  INV_X1 U5939 ( .A(n6754), .ZN(n6578) );
  AOI22_X1 U5940 ( .A1(n6747), .A2(n4950), .B1(n5227), .B2(n6578), .ZN(n4827)
         );
  OAI211_X1 U5941 ( .C1(n6582), .C2(n5120), .A(n4828), .B(n4827), .ZN(U3131)
         );
  INV_X1 U5942 ( .A(n6722), .ZN(n6634) );
  AOI22_X1 U5943 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4947), .B1(n6720), 
        .B2(n4946), .ZN(n4830) );
  INV_X1 U5944 ( .A(n6725), .ZN(n6630) );
  AOI22_X1 U5945 ( .A1(n6721), .A2(n4950), .B1(n5227), .B2(n6630), .ZN(n4829)
         );
  OAI211_X1 U5946 ( .C1(n6634), .C2(n5120), .A(n4830), .B(n4829), .ZN(U3127)
         );
  INV_X1 U5947 ( .A(n6704), .ZN(n6562) );
  AOI22_X1 U5948 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4947), .B1(n6693), 
        .B2(n4946), .ZN(n4832) );
  INV_X1 U5949 ( .A(n6707), .ZN(n6618) );
  AOI22_X1 U5950 ( .A1(n6692), .A2(n4950), .B1(n5227), .B2(n6618), .ZN(n4831)
         );
  OAI211_X1 U5951 ( .C1(n6562), .C2(n5120), .A(n4832), .B(n4831), .ZN(U3124)
         );
  INV_X1 U5952 ( .A(n6710), .ZN(n6597) );
  AOI22_X1 U5953 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4947), .B1(n6708), 
        .B2(n4946), .ZN(n4834) );
  AOI22_X1 U5954 ( .A1(n6709), .A2(n4950), .B1(n5227), .B2(n6622), .ZN(n4833)
         );
  OAI211_X1 U5955 ( .C1(n6597), .C2(n5120), .A(n4834), .B(n4833), .ZN(U3125)
         );
  NAND2_X1 U5956 ( .A1(n4925), .A2(n6583), .ZN(n6652) );
  NAND3_X1 U5957 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6770), .A3(n6764), .ZN(n5021) );
  NOR2_X1 U5958 ( .A1(n6759), .A2(n5021), .ZN(n5011) );
  AOI21_X1 U5959 ( .B1(n6690), .B2(n6511), .A(n5011), .ZN(n4838) );
  INV_X1 U5960 ( .A(n4838), .ZN(n4836) );
  OAI21_X1 U5961 ( .B1(n4839), .B2(n6089), .A(n6703), .ZN(n4837) );
  AOI21_X1 U5962 ( .B1(n6934), .B2(n5021), .A(n6655), .ZN(n4835) );
  OAI21_X1 U5963 ( .B1(n4836), .B2(n4837), .A(n4835), .ZN(n5010) );
  OAI22_X1 U5964 ( .A1(n4838), .A2(n4837), .B1(n6937), .B2(n5021), .ZN(n5009)
         );
  AOI22_X1 U5965 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5010), .B1(n6708), 
        .B2(n5009), .ZN(n4841) );
  AOI22_X1 U5966 ( .A1(n5299), .A2(n6710), .B1(n6709), .B2(n5011), .ZN(n4840)
         );
  OAI211_X1 U5967 ( .C1(n5116), .C2(n6713), .A(n4841), .B(n4840), .ZN(U3093)
         );
  AOI22_X1 U5968 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5010), .B1(n6693), 
        .B2(n5009), .ZN(n4843) );
  AOI22_X1 U5969 ( .A1(n5299), .A2(n6704), .B1(n6692), .B2(n5011), .ZN(n4842)
         );
  OAI211_X1 U5970 ( .C1(n5116), .C2(n6707), .A(n4843), .B(n4842), .ZN(U3092)
         );
  AOI22_X1 U5971 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5010), .B1(n6720), 
        .B2(n5009), .ZN(n4845) );
  AOI22_X1 U5972 ( .A1(n5299), .A2(n6722), .B1(n6721), .B2(n5011), .ZN(n4844)
         );
  OAI211_X1 U5973 ( .C1(n5116), .C2(n6725), .A(n4845), .B(n4844), .ZN(U3095)
         );
  AOI22_X1 U5974 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5010), .B1(n6745), 
        .B2(n5009), .ZN(n4847) );
  AOI22_X1 U5975 ( .A1(n5299), .A2(n6749), .B1(n6747), .B2(n5011), .ZN(n4846)
         );
  OAI211_X1 U5976 ( .C1(n5116), .C2(n6754), .A(n4847), .B(n4846), .ZN(U3099)
         );
  AOI22_X1 U5977 ( .A1(n6721), .A2(n5095), .B1(n6720), .B2(n5094), .ZN(n4849)
         );
  INV_X1 U5978 ( .A(n6608), .ZN(n6612) );
  NAND2_X1 U5979 ( .A1(n6612), .A2(n6630), .ZN(n4848) );
  OAI211_X1 U5980 ( .C1(n5143), .C2(n6634), .A(n4849), .B(n4848), .ZN(n4850)
         );
  AOI21_X1 U5981 ( .B1(n5099), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n4850), 
        .ZN(n4851) );
  INV_X1 U5982 ( .A(n4851), .ZN(U3055) );
  AOI22_X1 U5983 ( .A1(n6709), .A2(n5095), .B1(n6708), .B2(n5094), .ZN(n4853)
         );
  NAND2_X1 U5984 ( .A1(n6612), .A2(n6622), .ZN(n4852) );
  OAI211_X1 U5985 ( .C1(n5143), .C2(n6597), .A(n4853), .B(n4852), .ZN(n4854)
         );
  AOI21_X1 U5986 ( .B1(n5099), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n4854), 
        .ZN(n4855) );
  INV_X1 U5987 ( .A(n4855), .ZN(U3053) );
  AOI22_X1 U5988 ( .A1(n6747), .A2(n5095), .B1(n6745), .B2(n5094), .ZN(n4857)
         );
  NAND2_X1 U5989 ( .A1(n6612), .A2(n6578), .ZN(n4856) );
  OAI211_X1 U5990 ( .C1(n5143), .C2(n6582), .A(n4857), .B(n4856), .ZN(n4858)
         );
  AOI21_X1 U5991 ( .B1(n5099), .B2(INSTQUEUE_REG_4__7__SCAN_IN), .A(n4858), 
        .ZN(n4859) );
  INV_X1 U5992 ( .A(n4859), .ZN(U3059) );
  INV_X1 U5993 ( .A(n6655), .ZN(n6700) );
  INV_X1 U5994 ( .A(n4873), .ZN(n4860) );
  NAND2_X1 U5995 ( .A1(n4860), .A2(n6703), .ZN(n4861) );
  NAND2_X1 U5996 ( .A1(n6703), .A2(n6089), .ZN(n6695) );
  NAND2_X1 U5997 ( .A1(n4861), .A2(n6695), .ZN(n4868) );
  NAND2_X1 U5998 ( .A1(n4862), .A2(n6653), .ZN(n4864) );
  NOR2_X1 U5999 ( .A1(n6759), .A2(n4869), .ZN(n5139) );
  INV_X1 U6000 ( .A(n5139), .ZN(n4863) );
  NAND2_X1 U6001 ( .A1(n4864), .A2(n4863), .ZN(n4867) );
  INV_X1 U6002 ( .A(n4867), .ZN(n4865) );
  AOI22_X1 U6003 ( .A1(n4868), .A2(n4865), .B1(n4869), .B2(n6934), .ZN(n4866)
         );
  NAND2_X1 U6004 ( .A1(n6700), .A2(n4866), .ZN(n5145) );
  INV_X1 U6005 ( .A(n5145), .ZN(n5093) );
  INV_X1 U6006 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U6007 ( .A1(n4868), .A2(n4867), .ZN(n4872) );
  INV_X1 U6008 ( .A(n4869), .ZN(n4870) );
  NAND2_X1 U6009 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4870), .ZN(n4871) );
  NAND2_X1 U6010 ( .A1(n4872), .A2(n4871), .ZN(n5140) );
  AOI22_X1 U6011 ( .A1(n6692), .A2(n5139), .B1(n5932), .B2(n6704), .ZN(n4874)
         );
  OAI21_X1 U6012 ( .B1(n6707), .B2(n5143), .A(n4874), .ZN(n4875) );
  AOI21_X1 U6013 ( .B1(n6693), .B2(n5140), .A(n4875), .ZN(n4876) );
  OAI21_X1 U6014 ( .B1(n5093), .B2(n4877), .A(n4876), .ZN(U3060) );
  AOI22_X1 U6015 ( .A1(n6747), .A2(n5139), .B1(n5932), .B2(n6749), .ZN(n4879)
         );
  NAND2_X1 U6016 ( .A1(n5140), .A2(n6745), .ZN(n4878) );
  OAI211_X1 U6017 ( .C1(n5143), .C2(n6754), .A(n4879), .B(n4878), .ZN(n4880)
         );
  AOI21_X1 U6018 ( .B1(n5145), .B2(INSTQUEUE_REG_5__7__SCAN_IN), .A(n4880), 
        .ZN(n4881) );
  INV_X1 U6019 ( .A(n4881), .ZN(U3067) );
  AOI22_X1 U6020 ( .A1(n6709), .A2(n5139), .B1(n5932), .B2(n6710), .ZN(n4883)
         );
  NAND2_X1 U6021 ( .A1(n5140), .A2(n6708), .ZN(n4882) );
  OAI211_X1 U6022 ( .C1(n5143), .C2(n6713), .A(n4883), .B(n4882), .ZN(n4884)
         );
  AOI21_X1 U6023 ( .B1(n5145), .B2(INSTQUEUE_REG_5__1__SCAN_IN), .A(n4884), 
        .ZN(n4885) );
  INV_X1 U6024 ( .A(n4885), .ZN(U3061) );
  INV_X1 U6025 ( .A(n5052), .ZN(n4888) );
  AOI21_X1 U6026 ( .B1(n4998), .B2(n4999), .A(n4886), .ZN(n4887) );
  NOR2_X1 U6027 ( .A1(n4888), .A2(n4887), .ZN(n5007) );
  INV_X1 U6028 ( .A(n5007), .ZN(n5192) );
  NOR2_X1 U6029 ( .A1(n6204), .A2(n4889), .ZN(n4890) );
  OR2_X1 U6030 ( .A1(n6195), .A2(n4890), .ZN(n6452) );
  INV_X1 U6031 ( .A(n6452), .ZN(n4891) );
  AOI22_X1 U6032 ( .A1(n6257), .A2(n4891), .B1(EBX_REG_8__SCAN_IN), .B2(n5680), 
        .ZN(n4892) );
  OAI21_X1 U6033 ( .B1(n5192), .B2(n6014), .A(n4892), .ZN(U2851) );
  AOI22_X1 U6034 ( .A1(n6271), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6267), .ZN(n4893) );
  OAI21_X1 U6035 ( .B1(n5192), .B2(n6277), .A(n4893), .ZN(U2883) );
  AOI22_X1 U6036 ( .A1(n6721), .A2(n5139), .B1(n5932), .B2(n6722), .ZN(n4895)
         );
  NAND2_X1 U6037 ( .A1(n5140), .A2(n6720), .ZN(n4894) );
  OAI211_X1 U6038 ( .C1(n5143), .C2(n6725), .A(n4895), .B(n4894), .ZN(n4896)
         );
  AOI21_X1 U6039 ( .B1(n5145), .B2(INSTQUEUE_REG_5__3__SCAN_IN), .A(n4896), 
        .ZN(n4897) );
  INV_X1 U6040 ( .A(n4897), .ZN(U3063) );
  NOR2_X1 U6041 ( .A1(n4722), .A2(n4898), .ZN(n6689) );
  INV_X1 U6042 ( .A(n6689), .ZN(n5349) );
  NOR2_X1 U6043 ( .A1(n5349), .A2(n6934), .ZN(n4899) );
  NOR2_X1 U6044 ( .A1(n5022), .A2(n6777), .ZN(n5263) );
  AOI22_X1 U6045 ( .A1(n4899), .A2(n6553), .B1(n6517), .B2(n5263), .ZN(n5127)
         );
  NAND2_X1 U6046 ( .A1(n4900), .A2(n4960), .ZN(n6694) );
  INV_X1 U6047 ( .A(n6753), .ZN(n5123) );
  NOR2_X1 U6048 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6691), .ZN(n4908)
         );
  INV_X1 U6049 ( .A(n4908), .ZN(n5121) );
  OAI22_X1 U6050 ( .A1(n4901), .A2(n5121), .B1(n6707), .B2(n5120), .ZN(n4902)
         );
  AOI21_X1 U6051 ( .B1(n6704), .B2(n5123), .A(n4902), .ZN(n4910) );
  INV_X1 U6052 ( .A(n5120), .ZN(n4903) );
  OAI21_X1 U6053 ( .B1(n5123), .B2(n4903), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4904) );
  NAND3_X1 U6054 ( .A1(n5349), .A2(n6703), .A3(n4904), .ZN(n4907) );
  OAI21_X1 U6055 ( .B1(n6554), .B2(n6937), .A(n4905), .ZN(n5351) );
  NOR3_X1 U6056 ( .A1(n5351), .A2(n6777), .A3(n6555), .ZN(n4906) );
  OAI211_X1 U6057 ( .C1(n4908), .C2(n6904), .A(n4907), .B(n4906), .ZN(n5124)
         );
  NAND2_X1 U6058 ( .A1(n5124), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4909)
         );
  OAI211_X1 U6059 ( .C1(n5127), .C2(n5270), .A(n4910), .B(n4909), .ZN(U3132)
         );
  OAI22_X1 U6060 ( .A1(n6634), .A2(n6753), .B1(n5120), .B2(n6725), .ZN(n4913)
         );
  OAI22_X1 U6061 ( .A1(n4911), .A2(n5121), .B1(n5127), .B2(n5294), .ZN(n4912)
         );
  AOI211_X1 U6062 ( .C1(n5124), .C2(INSTQUEUE_REG_14__3__SCAN_IN), .A(n4913), 
        .B(n4912), .ZN(n4914) );
  INV_X1 U6063 ( .A(n4914), .ZN(U3135) );
  OAI22_X1 U6064 ( .A1(n6597), .A2(n6753), .B1(n5120), .B2(n6713), .ZN(n4917)
         );
  OAI22_X1 U6065 ( .A1(n4915), .A2(n5121), .B1(n5127), .B2(n5274), .ZN(n4916)
         );
  AOI211_X1 U6066 ( .C1(n5124), .C2(INSTQUEUE_REG_14__1__SCAN_IN), .A(n4917), 
        .B(n4916), .ZN(n4918) );
  INV_X1 U6067 ( .A(n4918), .ZN(U3133) );
  OAI22_X1 U6068 ( .A1(n6582), .A2(n6753), .B1(n5120), .B2(n6754), .ZN(n4921)
         );
  OAI22_X1 U6069 ( .A1(n4919), .A2(n5121), .B1(n5127), .B2(n5278), .ZN(n4920)
         );
  AOI211_X1 U6070 ( .C1(n5124), .C2(INSTQUEUE_REG_14__7__SCAN_IN), .A(n4921), 
        .B(n4920), .ZN(n4922) );
  INV_X1 U6071 ( .A(n4922), .ZN(U3139) );
  NOR2_X1 U6072 ( .A1(n4923), .A2(n6934), .ZN(n4942) );
  INV_X1 U6073 ( .A(n4959), .ZN(n4924) );
  NAND2_X1 U6074 ( .A1(n4960), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6651) );
  INV_X1 U6075 ( .A(n6651), .ZN(n6584) );
  NAND2_X1 U6076 ( .A1(n4924), .A2(n6584), .ZN(n4953) );
  NAND2_X1 U6077 ( .A1(n4925), .A2(n6089), .ZN(n4926) );
  NAND4_X1 U6078 ( .A1(n4927), .A2(n6652), .A3(n4953), .A4(n4926), .ZN(n4928)
         );
  NAND2_X1 U6079 ( .A1(n4942), .A2(n4928), .ZN(n4930) );
  NAND3_X1 U6080 ( .A1(n6509), .A2(n6553), .A3(n4943), .ZN(n4929) );
  OAI211_X1 U6081 ( .C1(n6509), .C2(n6777), .A(n4930), .B(n4929), .ZN(U3462)
         );
  XOR2_X1 U6082 ( .A(n6583), .B(n6651), .Z(n4931) );
  NAND2_X1 U6083 ( .A1(n4942), .A2(n4931), .ZN(n4933) );
  INV_X1 U6084 ( .A(n4722), .ZN(n5337) );
  NAND3_X1 U6085 ( .A1(n6509), .A2(n5337), .A3(n4943), .ZN(n4932) );
  OAI211_X1 U6086 ( .C1(n6509), .C2(n6770), .A(n4933), .B(n4932), .ZN(U3463)
         );
  AND2_X1 U6087 ( .A1(n3085), .A2(DATAI_22_), .ZN(n6740) );
  INV_X1 U6088 ( .A(n6740), .ZN(n6680) );
  NOR2_X2 U6089 ( .A1(n6362), .A2(n5024), .ZN(n6738) );
  AOI22_X1 U6090 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4947), .B1(n6738), 
        .B2(n4946), .ZN(n4936) );
  NOR2_X2 U6091 ( .A1(n4949), .A2(n4934), .ZN(n6739) );
  NAND2_X1 U6092 ( .A1(n3085), .A2(DATAI_30_), .ZN(n6743) );
  INV_X1 U6093 ( .A(n6743), .ZN(n6675) );
  AOI22_X1 U6094 ( .A1(n6739), .A2(n4950), .B1(n5227), .B2(n6675), .ZN(n4935)
         );
  OAI211_X1 U6095 ( .C1(n6680), .C2(n5120), .A(n4936), .B(n4935), .ZN(U3130)
         );
  AND2_X1 U6096 ( .A1(n3085), .A2(DATAI_21_), .ZN(n6734) );
  INV_X1 U6097 ( .A(n6734), .ZN(n6640) );
  NOR2_X2 U6098 ( .A1(n6360), .A2(n5024), .ZN(n6732) );
  AOI22_X1 U6099 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4947), .B1(n6732), 
        .B2(n4946), .ZN(n4938) );
  NOR2_X2 U6100 ( .A1(n4949), .A2(n3614), .ZN(n6733) );
  NAND2_X1 U6101 ( .A1(n3085), .A2(DATAI_29_), .ZN(n6737) );
  INV_X1 U6102 ( .A(n6737), .ZN(n6636) );
  AOI22_X1 U6103 ( .A1(n6733), .A2(n4950), .B1(n5227), .B2(n6636), .ZN(n4937)
         );
  OAI211_X1 U6104 ( .C1(n6640), .C2(n5120), .A(n4938), .B(n4937), .ZN(U3129)
         );
  AND2_X1 U6105 ( .A1(n3085), .A2(DATAI_18_), .ZN(n6716) );
  INV_X1 U6106 ( .A(n6716), .ZN(n6600) );
  INV_X1 U6107 ( .A(DATAI_2_), .ZN(n6354) );
  NOR2_X2 U6108 ( .A1(n6354), .A2(n5024), .ZN(n6715) );
  AOI22_X1 U6109 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4947), .B1(n6715), 
        .B2(n4946), .ZN(n4941) );
  NOR2_X2 U6110 ( .A1(n4949), .A2(n4939), .ZN(n6714) );
  AND2_X1 U6111 ( .A1(n3085), .A2(DATAI_26_), .ZN(n6626) );
  AOI22_X1 U6112 ( .A1(n6714), .A2(n4950), .B1(n5227), .B2(n6626), .ZN(n4940)
         );
  OAI211_X1 U6113 ( .C1(n6600), .C2(n5120), .A(n4941), .B(n4940), .ZN(U3126)
         );
  OAI211_X1 U6114 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4960), .A(n4942), .B(
        n6651), .ZN(n4945) );
  NAND3_X1 U6115 ( .A1(n6509), .A2(n4618), .A3(n4943), .ZN(n4944) );
  OAI211_X1 U6116 ( .C1(n6509), .C2(n6764), .A(n4945), .B(n4944), .ZN(U3464)
         );
  AND2_X1 U6117 ( .A1(n3085), .A2(DATAI_20_), .ZN(n6728) );
  INV_X1 U6118 ( .A(n6728), .ZN(n6672) );
  NOR2_X2 U6119 ( .A1(n6358), .A2(n5024), .ZN(n6726) );
  AOI22_X1 U6120 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4947), .B1(n6726), 
        .B2(n4946), .ZN(n4952) );
  NOR2_X2 U6121 ( .A1(n4949), .A2(n4948), .ZN(n6727) );
  NAND2_X1 U6122 ( .A1(n3085), .A2(DATAI_28_), .ZN(n6731) );
  INV_X1 U6123 ( .A(n6731), .ZN(n6669) );
  AOI22_X1 U6124 ( .A1(n6727), .A2(n4950), .B1(n5227), .B2(n6669), .ZN(n4951)
         );
  OAI211_X1 U6125 ( .C1(n6672), .C2(n5120), .A(n4952), .B(n4951), .ZN(U3128)
         );
  INV_X1 U6126 ( .A(n4953), .ZN(n4955) );
  NOR2_X1 U6127 ( .A1(n5349), .A2(n5202), .ZN(n5350) );
  INV_X1 U6128 ( .A(n5350), .ZN(n4954) );
  INV_X1 U6129 ( .A(n6653), .ZN(n6758) );
  OAI21_X1 U6130 ( .B1(n4954), .B2(n6758), .A(n4957), .ZN(n4963) );
  NOR3_X1 U6131 ( .A1(n4955), .A2(n6934), .A3(n4963), .ZN(n4956) );
  AOI211_X1 U6132 ( .C1(n5345), .C2(n6934), .A(n6655), .B(n4956), .ZN(n6631)
         );
  INV_X1 U6133 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4967) );
  INV_X1 U6134 ( .A(n4957), .ZN(n6644) );
  NOR2_X1 U6135 ( .A1(n4959), .A2(n5259), .ZN(n4958) );
  NOR2_X1 U6136 ( .A1(n4959), .A2(n6551), .ZN(n4961) );
  NAND2_X1 U6137 ( .A1(n4961), .A2(n4960), .ZN(n6639) );
  OAI22_X1 U6138 ( .A1(n6649), .A2(n6731), .B1(n6672), .B2(n6639), .ZN(n4962)
         );
  AOI21_X1 U6139 ( .B1(n6644), .B2(n6727), .A(n4962), .ZN(n4966) );
  NAND2_X1 U6140 ( .A1(n4963), .A2(n6703), .ZN(n4964) );
  OAI21_X1 U6141 ( .B1(n5345), .B2(n6937), .A(n4964), .ZN(n6645) );
  NAND2_X1 U6142 ( .A1(n6645), .A2(n6726), .ZN(n4965) );
  OAI211_X1 U6143 ( .C1(n6631), .C2(n4967), .A(n4966), .B(n4965), .ZN(U3080)
         );
  AOI22_X1 U6144 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5010), .B1(n6738), 
        .B2(n5009), .ZN(n4969) );
  AOI22_X1 U6145 ( .A1(n5299), .A2(n6740), .B1(n6739), .B2(n5011), .ZN(n4968)
         );
  OAI211_X1 U6146 ( .C1(n5116), .C2(n6743), .A(n4969), .B(n4968), .ZN(U3098)
         );
  AOI22_X1 U6147 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5010), .B1(n6732), 
        .B2(n5009), .ZN(n4971) );
  AOI22_X1 U6148 ( .A1(n5299), .A2(n6734), .B1(n6733), .B2(n5011), .ZN(n4970)
         );
  OAI211_X1 U6149 ( .C1(n5116), .C2(n6737), .A(n4971), .B(n4970), .ZN(U3097)
         );
  INV_X1 U6150 ( .A(n5587), .ZN(n4975) );
  AOI21_X1 U6151 ( .B1(n6425), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4972), 
        .ZN(n4973) );
  OAI21_X1 U6152 ( .B1(n6434), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4973), 
        .ZN(n4974) );
  AOI21_X1 U6153 ( .B1(n3085), .B2(n4975), .A(n4974), .ZN(n4976) );
  OAI21_X1 U6154 ( .B1(n4977), .B2(n6410), .A(n4976), .ZN(U2985) );
  INV_X1 U6155 ( .A(n6626), .ZN(n6719) );
  AOI22_X1 U6156 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5010), .B1(n6715), 
        .B2(n5009), .ZN(n4979) );
  AOI22_X1 U6157 ( .A1(n5299), .A2(n6716), .B1(n6714), .B2(n5011), .ZN(n4978)
         );
  OAI211_X1 U6158 ( .C1(n5116), .C2(n6719), .A(n4979), .B(n4978), .ZN(U3094)
         );
  OAI21_X1 U6159 ( .B1(n4982), .B2(n4981), .A(n4980), .ZN(n6475) );
  INV_X1 U6160 ( .A(n5308), .ZN(n4984) );
  AOI22_X1 U6161 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6483), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4983) );
  OAI21_X1 U6162 ( .B1(n6434), .B2(n4984), .A(n4983), .ZN(n4985) );
  AOI21_X1 U6163 ( .B1(n4986), .B2(n3085), .A(n4985), .ZN(n4987) );
  OAI21_X1 U6164 ( .B1(n6410), .B2(n6475), .A(n4987), .ZN(U2982) );
  NAND2_X1 U6165 ( .A1(n4989), .A2(n4988), .ZN(n4992) );
  NAND2_X1 U6166 ( .A1(n4992), .A2(n4991), .ZN(n4990) );
  OAI21_X1 U6167 ( .B1(n4992), .B2(n4991), .A(n4990), .ZN(n6468) );
  INV_X1 U6168 ( .A(n5257), .ZN(n4996) );
  INV_X1 U6169 ( .A(n5255), .ZN(n4994) );
  AOI22_X1 U6170 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6483), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4993) );
  OAI21_X1 U6171 ( .B1(n6434), .B2(n4994), .A(n4993), .ZN(n4995) );
  AOI21_X1 U6172 ( .B1(n4996), .B2(n3085), .A(n4995), .ZN(n4997) );
  OAI21_X1 U6173 ( .B1(n6468), .B2(n6410), .A(n4997), .ZN(U2980) );
  XOR2_X1 U6174 ( .A(n4999), .B(n4998), .Z(n6405) );
  INV_X1 U6175 ( .A(n6405), .ZN(n5000) );
  OAI222_X1 U6176 ( .A1(n6277), .A2(n5000), .B1(n6275), .B2(n6364), .C1(n6276), 
        .C2(n3844), .ZN(U2884) );
  OAI21_X1 U6177 ( .B1(n5003), .B2(n5002), .A(n5001), .ZN(n6451) );
  INV_X1 U6178 ( .A(n5189), .ZN(n5005) );
  AOI22_X1 U6179 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6483), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5004) );
  OAI21_X1 U6180 ( .B1(n6434), .B2(n5005), .A(n5004), .ZN(n5006) );
  AOI21_X1 U6181 ( .B1(n5007), .B2(n3085), .A(n5006), .ZN(n5008) );
  OAI21_X1 U6182 ( .B1(n6451), .B2(n6410), .A(n5008), .ZN(U2978) );
  AOI22_X1 U6183 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5010), .B1(n6726), 
        .B2(n5009), .ZN(n5013) );
  AOI22_X1 U6184 ( .A1(n5299), .A2(n6728), .B1(n6727), .B2(n5011), .ZN(n5012)
         );
  OAI211_X1 U6185 ( .C1(n5116), .C2(n6731), .A(n5013), .B(n5012), .ZN(U3096)
         );
  OAI21_X1 U6186 ( .B1(n5052), .B2(n5053), .A(n5014), .ZN(n5015) );
  NAND2_X1 U6187 ( .A1(n5015), .A2(n5147), .ZN(n6185) );
  AOI22_X1 U6188 ( .A1(n6271), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6267), .ZN(n5016) );
  OAI21_X1 U6189 ( .B1(n6185), .B2(n6277), .A(n5016), .ZN(U2881) );
  INV_X1 U6190 ( .A(n5150), .ZN(n5018) );
  AOI21_X1 U6191 ( .B1(n5019), .B2(n5017), .A(n5018), .ZN(n6181) );
  AOI22_X1 U6192 ( .A1(n6257), .A2(n6181), .B1(EBX_REG_10__SCAN_IN), .B2(n5680), .ZN(n5020) );
  OAI21_X1 U6193 ( .B1(n6185), .B2(n6014), .A(n5020), .ZN(U2849) );
  AOI21_X1 U6194 ( .B1(n5116), .B2(n6639), .A(n6089), .ZN(n5029) );
  NAND2_X1 U6195 ( .A1(n6511), .A2(n6553), .ZN(n5030) );
  NAND2_X1 U6196 ( .A1(n5030), .A2(n6703), .ZN(n5028) );
  NOR2_X1 U6197 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5021), .ZN(n5113)
         );
  INV_X1 U6198 ( .A(n5113), .ZN(n5026) );
  NAND2_X1 U6199 ( .A1(n5023), .A2(n5022), .ZN(n5210) );
  AOI21_X1 U6200 ( .B1(n5210), .B2(STATE2_REG_2__SCAN_IN), .A(n5024), .ZN(
        n5025) );
  INV_X1 U6201 ( .A(n5025), .ZN(n5204) );
  AOI211_X1 U6202 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5026), .A(n6517), .B(
        n5204), .ZN(n5027) );
  OAI21_X1 U6203 ( .B1(n5029), .B2(n5028), .A(n5027), .ZN(n5118) );
  OR2_X1 U6204 ( .A1(n5030), .A2(n6934), .ZN(n5033) );
  INV_X1 U6205 ( .A(n5210), .ZN(n5031) );
  NAND2_X1 U6206 ( .A1(n6555), .A2(n5031), .ZN(n5032) );
  AND2_X1 U6207 ( .A1(n5033), .A2(n5032), .ZN(n5072) );
  INV_X1 U6208 ( .A(n5072), .ZN(n5112) );
  NAND2_X1 U6209 ( .A1(n6693), .A2(n5112), .ZN(n5035) );
  INV_X1 U6210 ( .A(n6639), .ZN(n6643) );
  AOI22_X1 U6211 ( .A1(n6692), .A2(n5113), .B1(n6643), .B2(n6618), .ZN(n5034)
         );
  OAI211_X1 U6212 ( .C1(n6562), .C2(n5116), .A(n5035), .B(n5034), .ZN(n5036)
         );
  AOI21_X1 U6213 ( .B1(n5118), .B2(INSTQUEUE_REG_8__0__SCAN_IN), .A(n5036), 
        .ZN(n5037) );
  INV_X1 U6214 ( .A(n5037), .ZN(U3084) );
  AOI22_X1 U6215 ( .A1(n6733), .A2(n5095), .B1(n6732), .B2(n5094), .ZN(n5039)
         );
  NAND2_X1 U6216 ( .A1(n6612), .A2(n6636), .ZN(n5038) );
  OAI211_X1 U6217 ( .C1(n5143), .C2(n6640), .A(n5039), .B(n5038), .ZN(n5040)
         );
  AOI21_X1 U6218 ( .B1(n5099), .B2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n5040), 
        .ZN(n5041) );
  INV_X1 U6219 ( .A(n5041), .ZN(U3057) );
  AOI22_X1 U6220 ( .A1(n6739), .A2(n5095), .B1(n6738), .B2(n5094), .ZN(n5043)
         );
  NAND2_X1 U6221 ( .A1(n6612), .A2(n6675), .ZN(n5042) );
  OAI211_X1 U6222 ( .C1(n5143), .C2(n6680), .A(n5043), .B(n5042), .ZN(n5044)
         );
  AOI21_X1 U6223 ( .B1(n5099), .B2(INSTQUEUE_REG_4__6__SCAN_IN), .A(n5044), 
        .ZN(n5045) );
  INV_X1 U6224 ( .A(n5045), .ZN(U3058) );
  OAI22_X1 U6225 ( .A1(n6640), .A2(n6753), .B1(n5120), .B2(n6737), .ZN(n5047)
         );
  INV_X1 U6226 ( .A(n6733), .ZN(n5076) );
  INV_X1 U6227 ( .A(n6732), .ZN(n5290) );
  OAI22_X1 U6228 ( .A1(n5076), .A2(n5121), .B1(n5127), .B2(n5290), .ZN(n5046)
         );
  AOI211_X1 U6229 ( .C1(n5124), .C2(INSTQUEUE_REG_14__5__SCAN_IN), .A(n5047), 
        .B(n5046), .ZN(n5048) );
  INV_X1 U6230 ( .A(n5048), .ZN(U3137) );
  OAI22_X1 U6231 ( .A1(n6680), .A2(n6753), .B1(n5120), .B2(n6743), .ZN(n5050)
         );
  INV_X1 U6232 ( .A(n6739), .ZN(n5080) );
  INV_X1 U6233 ( .A(n6738), .ZN(n5282) );
  OAI22_X1 U6234 ( .A1(n5080), .A2(n5121), .B1(n5127), .B2(n5282), .ZN(n5049)
         );
  AOI211_X1 U6235 ( .C1(n5124), .C2(INSTQUEUE_REG_14__6__SCAN_IN), .A(n5050), 
        .B(n5049), .ZN(n5051) );
  INV_X1 U6236 ( .A(n5051), .ZN(U3138) );
  XOR2_X1 U6237 ( .A(n5053), .B(n5052), .Z(n6397) );
  INV_X1 U6238 ( .A(n6397), .ZN(n5055) );
  INV_X1 U6239 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5054) );
  OAI222_X1 U6240 ( .A1(n5056), .A2(n6275), .B1(n6277), .B2(n5055), .C1(n5054), 
        .C2(n6276), .ZN(U2882) );
  NAND2_X1 U6241 ( .A1(n5118), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5059) );
  OAI22_X1 U6242 ( .A1(n6639), .A2(n6737), .B1(n5072), .B2(n5290), .ZN(n5057)
         );
  AOI21_X1 U6243 ( .B1(n6733), .B2(n5113), .A(n5057), .ZN(n5058) );
  OAI211_X1 U6244 ( .C1(n6640), .C2(n5116), .A(n5059), .B(n5058), .ZN(U3089)
         );
  NAND2_X1 U6245 ( .A1(n5118), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5062) );
  OAI22_X1 U6246 ( .A1(n6639), .A2(n6725), .B1(n5072), .B2(n5294), .ZN(n5060)
         );
  AOI21_X1 U6247 ( .B1(n6721), .B2(n5113), .A(n5060), .ZN(n5061) );
  OAI211_X1 U6248 ( .C1(n6634), .C2(n5116), .A(n5062), .B(n5061), .ZN(U3087)
         );
  NAND2_X1 U6249 ( .A1(n5118), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5065) );
  OAI22_X1 U6250 ( .A1(n6639), .A2(n6713), .B1(n5072), .B2(n5274), .ZN(n5063)
         );
  AOI21_X1 U6251 ( .B1(n6709), .B2(n5113), .A(n5063), .ZN(n5064) );
  OAI211_X1 U6252 ( .C1(n6597), .C2(n5116), .A(n5065), .B(n5064), .ZN(U3085)
         );
  NAND2_X1 U6253 ( .A1(n5118), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5068) );
  OAI22_X1 U6254 ( .A1(n6639), .A2(n6743), .B1(n5072), .B2(n5282), .ZN(n5066)
         );
  AOI21_X1 U6255 ( .B1(n6739), .B2(n5113), .A(n5066), .ZN(n5067) );
  OAI211_X1 U6256 ( .C1(n6680), .C2(n5116), .A(n5068), .B(n5067), .ZN(U3090)
         );
  NAND2_X1 U6257 ( .A1(n5118), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5071) );
  OAI22_X1 U6258 ( .A1(n6639), .A2(n6754), .B1(n5072), .B2(n5278), .ZN(n5069)
         );
  AOI21_X1 U6259 ( .B1(n6747), .B2(n5113), .A(n5069), .ZN(n5070) );
  OAI211_X1 U6260 ( .C1(n6582), .C2(n5116), .A(n5071), .B(n5070), .ZN(U3091)
         );
  NAND2_X1 U6261 ( .A1(n5118), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5075) );
  INV_X1 U6262 ( .A(n6726), .ZN(n5286) );
  OAI22_X1 U6263 ( .A1(n6639), .A2(n6731), .B1(n5072), .B2(n5286), .ZN(n5073)
         );
  AOI21_X1 U6264 ( .B1(n6727), .B2(n5113), .A(n5073), .ZN(n5074) );
  OAI211_X1 U6265 ( .C1(n6672), .C2(n5116), .A(n5075), .B(n5074), .ZN(U3088)
         );
  OAI22_X1 U6266 ( .A1(n5076), .A2(n5132), .B1(n6737), .B2(n6512), .ZN(n5077)
         );
  AOI21_X1 U6267 ( .B1(n6734), .B2(n6577), .A(n5077), .ZN(n5079) );
  NAND2_X1 U6268 ( .A1(n5135), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5078) );
  OAI211_X1 U6269 ( .C1(n5138), .C2(n5290), .A(n5079), .B(n5078), .ZN(U3033)
         );
  OAI22_X1 U6270 ( .A1(n5080), .A2(n5132), .B1(n6743), .B2(n6512), .ZN(n5081)
         );
  AOI21_X1 U6271 ( .B1(n6740), .B2(n6577), .A(n5081), .ZN(n5083) );
  NAND2_X1 U6272 ( .A1(n5135), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5082) );
  OAI211_X1 U6273 ( .C1(n5138), .C2(n5282), .A(n5083), .B(n5082), .ZN(U3034)
         );
  AOI22_X1 U6274 ( .A1(n6714), .A2(n5095), .B1(n5084), .B2(n6716), .ZN(n5085)
         );
  OAI21_X1 U6275 ( .B1(n6719), .B2(n6608), .A(n5085), .ZN(n5086) );
  AOI21_X1 U6276 ( .B1(n6715), .B2(n5094), .A(n5086), .ZN(n5087) );
  OAI21_X1 U6277 ( .B1(n5088), .B2(n4494), .A(n5087), .ZN(U3054) );
  INV_X1 U6278 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5092) );
  AOI22_X1 U6279 ( .A1(n6714), .A2(n5139), .B1(n5932), .B2(n6716), .ZN(n5089)
         );
  OAI21_X1 U6280 ( .B1(n6719), .B2(n5143), .A(n5089), .ZN(n5090) );
  AOI21_X1 U6281 ( .B1(n6715), .B2(n5140), .A(n5090), .ZN(n5091) );
  OAI21_X1 U6282 ( .B1(n5093), .B2(n5092), .A(n5091), .ZN(U3062) );
  AOI22_X1 U6283 ( .A1(n6727), .A2(n5095), .B1(n6726), .B2(n5094), .ZN(n5097)
         );
  NAND2_X1 U6284 ( .A1(n6612), .A2(n6669), .ZN(n5096) );
  OAI211_X1 U6285 ( .C1(n5143), .C2(n6672), .A(n5097), .B(n5096), .ZN(n5098)
         );
  AOI21_X1 U6286 ( .B1(n5099), .B2(INSTQUEUE_REG_4__4__SCAN_IN), .A(n5098), 
        .ZN(n5100) );
  INV_X1 U6287 ( .A(n5100), .ZN(U3056) );
  AOI22_X1 U6288 ( .A1(n6733), .A2(n5139), .B1(n5932), .B2(n6734), .ZN(n5102)
         );
  NAND2_X1 U6289 ( .A1(n5140), .A2(n6732), .ZN(n5101) );
  OAI211_X1 U6290 ( .C1(n5143), .C2(n6737), .A(n5102), .B(n5101), .ZN(n5103)
         );
  AOI21_X1 U6291 ( .B1(n5145), .B2(INSTQUEUE_REG_5__5__SCAN_IN), .A(n5103), 
        .ZN(n5104) );
  INV_X1 U6292 ( .A(n5104), .ZN(U3065) );
  AOI22_X1 U6293 ( .A1(n6739), .A2(n5139), .B1(n5932), .B2(n6740), .ZN(n5106)
         );
  NAND2_X1 U6294 ( .A1(n5140), .A2(n6738), .ZN(n5105) );
  OAI211_X1 U6295 ( .C1(n5143), .C2(n6743), .A(n5106), .B(n5105), .ZN(n5107)
         );
  AOI21_X1 U6296 ( .B1(n5145), .B2(INSTQUEUE_REG_5__6__SCAN_IN), .A(n5107), 
        .ZN(n5108) );
  INV_X1 U6297 ( .A(n5108), .ZN(U3066) );
  OAI22_X1 U6298 ( .A1(n6672), .A2(n6753), .B1(n5120), .B2(n6731), .ZN(n5110)
         );
  INV_X1 U6299 ( .A(n6727), .ZN(n5133) );
  OAI22_X1 U6300 ( .A1(n5133), .A2(n5121), .B1(n5127), .B2(n5286), .ZN(n5109)
         );
  AOI211_X1 U6301 ( .C1(n5124), .C2(INSTQUEUE_REG_14__4__SCAN_IN), .A(n5110), 
        .B(n5109), .ZN(n5111) );
  INV_X1 U6302 ( .A(n5111), .ZN(U3136) );
  NAND2_X1 U6303 ( .A1(n6715), .A2(n5112), .ZN(n5115) );
  AOI22_X1 U6304 ( .A1(n6714), .A2(n5113), .B1(n6643), .B2(n6626), .ZN(n5114)
         );
  OAI211_X1 U6305 ( .C1(n6600), .C2(n5116), .A(n5115), .B(n5114), .ZN(n5117)
         );
  AOI21_X1 U6306 ( .B1(n5118), .B2(INSTQUEUE_REG_8__2__SCAN_IN), .A(n5117), 
        .ZN(n5119) );
  INV_X1 U6307 ( .A(n5119), .ZN(U3086) );
  INV_X1 U6308 ( .A(n6715), .ZN(n5301) );
  INV_X1 U6309 ( .A(n6714), .ZN(n5128) );
  OAI22_X1 U6310 ( .A1(n5128), .A2(n5121), .B1(n6719), .B2(n5120), .ZN(n5122)
         );
  AOI21_X1 U6311 ( .B1(n6716), .B2(n5123), .A(n5122), .ZN(n5126) );
  NAND2_X1 U6312 ( .A1(n5124), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5125)
         );
  OAI211_X1 U6313 ( .C1(n5127), .C2(n5301), .A(n5126), .B(n5125), .ZN(U3134)
         );
  OAI22_X1 U6314 ( .A1(n5128), .A2(n5132), .B1(n6719), .B2(n6512), .ZN(n5129)
         );
  AOI21_X1 U6315 ( .B1(n6716), .B2(n6577), .A(n5129), .ZN(n5131) );
  NAND2_X1 U6316 ( .A1(n5135), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5130) );
  OAI211_X1 U6317 ( .C1(n5138), .C2(n5301), .A(n5131), .B(n5130), .ZN(U3030)
         );
  OAI22_X1 U6318 ( .A1(n5133), .A2(n5132), .B1(n6731), .B2(n6512), .ZN(n5134)
         );
  AOI21_X1 U6319 ( .B1(n6728), .B2(n6577), .A(n5134), .ZN(n5137) );
  NAND2_X1 U6320 ( .A1(n5135), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5136) );
  OAI211_X1 U6321 ( .C1(n5138), .C2(n5286), .A(n5137), .B(n5136), .ZN(U3032)
         );
  AOI22_X1 U6322 ( .A1(n6727), .A2(n5139), .B1(n5932), .B2(n6728), .ZN(n5142)
         );
  NAND2_X1 U6323 ( .A1(n5140), .A2(n6726), .ZN(n5141) );
  OAI211_X1 U6324 ( .C1(n5143), .C2(n6731), .A(n5142), .B(n5141), .ZN(n5144)
         );
  AOI21_X1 U6325 ( .B1(n5145), .B2(INSTQUEUE_REG_5__4__SCAN_IN), .A(n5144), 
        .ZN(n5146) );
  INV_X1 U6326 ( .A(n5146), .ZN(U3064) );
  AOI21_X1 U6327 ( .B1(n5148), .B2(n5147), .A(n5157), .ZN(n6176) );
  INV_X1 U6328 ( .A(n6176), .ZN(n5330) );
  AND2_X1 U6329 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  NOR2_X1 U6330 ( .A1(n5159), .A2(n5151), .ZN(n6436) );
  AOI22_X1 U6331 ( .A1(n6257), .A2(n6436), .B1(EBX_REG_11__SCAN_IN), .B2(n5680), .ZN(n5152) );
  OAI21_X1 U6332 ( .B1(n5330), .B2(n6014), .A(n5152), .ZN(U2848) );
  INV_X1 U6333 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5154) );
  OAI222_X1 U6334 ( .A1(n5330), .A2(n6277), .B1(n6276), .B2(n5154), .C1(n6275), 
        .C2(n5153), .ZN(U2880) );
  OAI21_X1 U6335 ( .B1(n5157), .B2(n5156), .A(n5155), .ZN(n6166) );
  NOR2_X1 U6336 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  OR2_X1 U6337 ( .A1(n5383), .A2(n5160), .ZN(n6157) );
  INV_X1 U6338 ( .A(n6157), .ZN(n5161) );
  AOI22_X1 U6339 ( .A1(n6257), .A2(n5161), .B1(EBX_REG_12__SCAN_IN), .B2(n5680), .ZN(n5162) );
  OAI21_X1 U6340 ( .B1(n6166), .B2(n6014), .A(n5162), .ZN(U2847) );
  INV_X1 U6341 ( .A(DATAI_12_), .ZN(n5163) );
  OAI222_X1 U6342 ( .A1(n6166), .A2(n6277), .B1(n6276), .B2(n5164), .C1(n6275), 
        .C2(n5163), .ZN(U2879) );
  NOR3_X1 U6343 ( .A1(n6809), .A2(n6904), .A3(n6810), .ZN(n6794) );
  AND2_X1 U6344 ( .A1(n5467), .A2(n5165), .ZN(n6803) );
  INV_X1 U6345 ( .A(n6803), .ZN(n5166) );
  NAND2_X1 U6346 ( .A1(n5166), .A2(n6495), .ZN(n5167) );
  OR2_X1 U6347 ( .A1(n6794), .A2(n5167), .ZN(n5168) );
  OR2_X2 U6348 ( .A1(n6936), .A2(n5168), .ZN(n6147) );
  NAND2_X1 U6349 ( .A1(n5464), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5463)
         );
  INV_X1 U6350 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5171) );
  NOR2_X1 U6351 ( .A1(n5709), .A2(n6912), .ZN(n5173) );
  NOR2_X1 U6353 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5185) );
  INV_X1 U6354 ( .A(n5185), .ZN(n5178) );
  NOR2_X1 U6355 ( .A1(n6824), .A2(n5178), .ZN(n5174) );
  NOR2_X1 U6356 ( .A1(n6788), .A2(n5174), .ZN(n5539) );
  INV_X1 U6357 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5529) );
  AND3_X1 U6358 ( .A1(n5184), .A2(n5529), .A3(n5178), .ZN(n5175) );
  OR2_X1 U6359 ( .A1(n5539), .A2(n5175), .ZN(n5176) );
  INV_X1 U6360 ( .A(n6085), .ZN(n5177) );
  NAND2_X1 U6361 ( .A1(n6147), .A2(n5177), .ZN(n6216) );
  AND2_X1 U6362 ( .A1(n5311), .A2(EBX_REG_31__SCAN_IN), .ZN(n5540) );
  AND2_X1 U6363 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  OAI22_X1 U6364 ( .A1(n5181), .A2(n6170), .B1(n6219), .B2(n6452), .ZN(n5182)
         );
  AOI211_X1 U6365 ( .C1(n6235), .C2(EBX_REG_8__SCAN_IN), .A(n6209), .B(n5182), 
        .ZN(n5191) );
  INV_X1 U6366 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6846) );
  INV_X1 U6367 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6844) );
  NOR3_X1 U6368 ( .A1(n6848), .A2(n6846), .A3(n6844), .ZN(n5409) );
  INV_X1 U6369 ( .A(n6147), .ZN(n6161) );
  INV_X1 U6370 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6841) );
  NAND3_X1 U6371 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5309) );
  NOR2_X1 U6372 ( .A1(n6841), .A2(n5309), .ZN(n6223) );
  NAND2_X1 U6373 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6223), .ZN(n5411) );
  NOR2_X1 U6374 ( .A1(n6161), .A2(n5411), .ZN(n5249) );
  AND3_X1 U6375 ( .A1(n5186), .A2(n5185), .A3(n5184), .ZN(n5187) );
  NAND2_X1 U6376 ( .A1(n6183), .A2(n6147), .ZN(n6159) );
  INV_X1 U6377 ( .A(n6159), .ZN(n6007) );
  AOI21_X1 U6378 ( .B1(n5409), .B2(n5249), .A(n6007), .ZN(n6194) );
  NOR2_X1 U6379 ( .A1(n6183), .A2(n5411), .ZN(n5248) );
  NAND2_X1 U6380 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5248), .ZN(n6207) );
  OAI21_X1 U6381 ( .B1(n6846), .B2(n6207), .A(n6848), .ZN(n5188) );
  AOI22_X1 U6382 ( .A1(n5189), .A2(n3092), .B1(n6194), .B2(n5188), .ZN(n5190)
         );
  OAI211_X1 U6383 ( .C1(n6128), .C2(n5192), .A(n5191), .B(n5190), .ZN(U2819)
         );
  INV_X1 U6384 ( .A(n5320), .ZN(n5196) );
  AOI21_X1 U6385 ( .B1(n5194), .B2(n5319), .A(n5193), .ZN(n5195) );
  AOI21_X1 U6386 ( .B1(n5196), .B2(n5319), .A(n5195), .ZN(n5912) );
  NAND2_X1 U6387 ( .A1(n5912), .A2(n6429), .ZN(n5200) );
  INV_X1 U6388 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5197) );
  OAI22_X1 U6389 ( .A1(n5800), .A2(n5197), .B1(n6495), .B2(n6852), .ZN(n5198)
         );
  AOI21_X1 U6390 ( .B1(n6387), .B2(n6186), .A(n5198), .ZN(n5199) );
  OAI211_X1 U6391 ( .C1(n6696), .C2(n6185), .A(n5200), .B(n5199), .ZN(U2976)
         );
  AOI21_X1 U6392 ( .B1(n5243), .B2(n6679), .A(n6089), .ZN(n5201) );
  AOI211_X1 U6393 ( .C1(n5207), .C2(n5202), .A(n6934), .B(n5201), .ZN(n5206)
         );
  NOR2_X1 U6394 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5203), .ZN(n5241)
         );
  NOR2_X1 U6395 ( .A1(n5241), .A2(n6904), .ZN(n5205) );
  NOR4_X2 U6396 ( .A1(n5206), .A2(n6555), .A3(n5205), .A4(n5204), .ZN(n5247)
         );
  INV_X1 U6397 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5214) );
  INV_X1 U6398 ( .A(n6517), .ZN(n5209) );
  NAND3_X1 U6399 ( .A1(n5207), .A2(n6703), .A3(n6553), .ZN(n5208) );
  OAI21_X1 U6400 ( .B1(n5210), .B2(n5209), .A(n5208), .ZN(n5240) );
  AOI22_X1 U6401 ( .A1(n6709), .A2(n5241), .B1(n6708), .B2(n5240), .ZN(n5211)
         );
  OAI21_X1 U6402 ( .B1(n6597), .B2(n5243), .A(n5211), .ZN(n5212) );
  AOI21_X1 U6403 ( .B1(n6622), .B2(n6681), .A(n5212), .ZN(n5213) );
  OAI21_X1 U6404 ( .B1(n5247), .B2(n5214), .A(n5213), .ZN(U3117) );
  INV_X1 U6405 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5218) );
  AOI22_X1 U6406 ( .A1(n6727), .A2(n5241), .B1(n6726), .B2(n5240), .ZN(n5215)
         );
  OAI21_X1 U6407 ( .B1(n6672), .B2(n5243), .A(n5215), .ZN(n5216) );
  AOI21_X1 U6408 ( .B1(n6669), .B2(n6681), .A(n5216), .ZN(n5217) );
  OAI21_X1 U6409 ( .B1(n5247), .B2(n5218), .A(n5217), .ZN(U3120) );
  INV_X1 U6410 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5222) );
  AOI22_X1 U6411 ( .A1(n6692), .A2(n5241), .B1(n5227), .B2(n6704), .ZN(n5219)
         );
  OAI21_X1 U6412 ( .B1(n6707), .B2(n6679), .A(n5219), .ZN(n5220) );
  AOI21_X1 U6413 ( .B1(n6693), .B2(n5240), .A(n5220), .ZN(n5221) );
  OAI21_X1 U6414 ( .B1(n5247), .B2(n5222), .A(n5221), .ZN(U3116) );
  INV_X1 U6415 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5226) );
  AOI22_X1 U6416 ( .A1(n6733), .A2(n5241), .B1(n6732), .B2(n5240), .ZN(n5223)
         );
  OAI21_X1 U6417 ( .B1(n6640), .B2(n5243), .A(n5223), .ZN(n5224) );
  AOI21_X1 U6418 ( .B1(n6636), .B2(n6681), .A(n5224), .ZN(n5225) );
  OAI21_X1 U6419 ( .B1(n5247), .B2(n5226), .A(n5225), .ZN(U3121) );
  INV_X1 U6420 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5231) );
  AOI22_X1 U6421 ( .A1(n6714), .A2(n5241), .B1(n5227), .B2(n6716), .ZN(n5228)
         );
  OAI21_X1 U6422 ( .B1(n6719), .B2(n6679), .A(n5228), .ZN(n5229) );
  AOI21_X1 U6423 ( .B1(n6715), .B2(n5240), .A(n5229), .ZN(n5230) );
  OAI21_X1 U6424 ( .B1(n5247), .B2(n5231), .A(n5230), .ZN(U3118) );
  INV_X1 U6425 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5235) );
  AOI22_X1 U6426 ( .A1(n6721), .A2(n5241), .B1(n6720), .B2(n5240), .ZN(n5232)
         );
  OAI21_X1 U6427 ( .B1(n6634), .B2(n5243), .A(n5232), .ZN(n5233) );
  AOI21_X1 U6428 ( .B1(n6630), .B2(n6681), .A(n5233), .ZN(n5234) );
  OAI21_X1 U6429 ( .B1(n5247), .B2(n5235), .A(n5234), .ZN(U3119) );
  INV_X1 U6430 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5239) );
  AOI22_X1 U6431 ( .A1(n6747), .A2(n5241), .B1(n6745), .B2(n5240), .ZN(n5236)
         );
  OAI21_X1 U6432 ( .B1(n6582), .B2(n5243), .A(n5236), .ZN(n5237) );
  AOI21_X1 U6433 ( .B1(n6578), .B2(n6681), .A(n5237), .ZN(n5238) );
  OAI21_X1 U6434 ( .B1(n5247), .B2(n5239), .A(n5238), .ZN(U3123) );
  INV_X1 U6435 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U6436 ( .A1(n6739), .A2(n5241), .B1(n6738), .B2(n5240), .ZN(n5242)
         );
  OAI21_X1 U6437 ( .B1(n6680), .B2(n5243), .A(n5242), .ZN(n5244) );
  AOI21_X1 U6438 ( .B1(n6675), .B2(n6681), .A(n5244), .ZN(n5245) );
  OAI21_X1 U6439 ( .B1(n5247), .B2(n5246), .A(n5245), .ZN(U3122) );
  NAND2_X1 U6440 ( .A1(n5248), .A2(n6844), .ZN(n6211) );
  OAI21_X1 U6441 ( .B1(n6469), .B2(n6219), .A(n6211), .ZN(n5254) );
  INV_X1 U6442 ( .A(n5249), .ZN(n5250) );
  AND2_X1 U6443 ( .A1(n6159), .A2(n5250), .ZN(n6210) );
  AOI22_X1 U6444 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6235), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6210), .ZN(n5251) );
  OAI211_X1 U6445 ( .C1(n6170), .C2(n5252), .A(n5251), .B(n6216), .ZN(n5253)
         );
  AOI211_X1 U6446 ( .C1(n5255), .C2(n3092), .A(n5254), .B(n5253), .ZN(n5256)
         );
  OAI21_X1 U6447 ( .B1(n6128), .B2(n5257), .A(n5256), .ZN(U2821) );
  NAND3_X1 U6448 ( .A1(n5260), .A2(n6703), .A3(n6687), .ZN(n5261) );
  NAND2_X1 U6449 ( .A1(n5261), .A2(n6695), .ZN(n5265) );
  NAND2_X1 U6450 ( .A1(n4722), .A2(n4618), .ZN(n6552) );
  INV_X1 U6451 ( .A(n6552), .ZN(n5262) );
  AND2_X1 U6452 ( .A1(n5262), .A2(n6553), .ZN(n6654) );
  AOI22_X1 U6453 ( .A1(n5265), .A2(n6654), .B1(n5263), .B2(n6555), .ZN(n5302)
         );
  NAND3_X1 U6454 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6770), .ZN(n6658) );
  NOR2_X1 U6455 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6658), .ZN(n5296)
         );
  NOR2_X1 U6456 ( .A1(n6517), .A2(n5351), .ZN(n6558) );
  INV_X1 U6457 ( .A(n6654), .ZN(n5264) );
  NOR2_X1 U6458 ( .A1(n6937), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5346)
         );
  AOI21_X1 U6459 ( .B1(n5265), .B2(n5264), .A(n5346), .ZN(n5266) );
  OAI211_X1 U6460 ( .C1(n5296), .C2(n6904), .A(n6558), .B(n5266), .ZN(n5295)
         );
  AOI22_X1 U6461 ( .A1(n6692), .A2(n5296), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5295), .ZN(n5267) );
  OAI21_X1 U6462 ( .B1(n6562), .B2(n6687), .A(n5267), .ZN(n5268) );
  AOI21_X1 U6463 ( .B1(n6618), .B2(n5299), .A(n5268), .ZN(n5269) );
  OAI21_X1 U6464 ( .B1(n5302), .B2(n5270), .A(n5269), .ZN(U3100) );
  AOI22_X1 U6465 ( .A1(n6709), .A2(n5296), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5295), .ZN(n5271) );
  OAI21_X1 U6466 ( .B1(n6597), .B2(n6687), .A(n5271), .ZN(n5272) );
  AOI21_X1 U6467 ( .B1(n5299), .B2(n6622), .A(n5272), .ZN(n5273) );
  OAI21_X1 U6468 ( .B1(n5302), .B2(n5274), .A(n5273), .ZN(U3101) );
  AOI22_X1 U6469 ( .A1(n6747), .A2(n5296), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5295), .ZN(n5275) );
  OAI21_X1 U6470 ( .B1(n6582), .B2(n6687), .A(n5275), .ZN(n5276) );
  AOI21_X1 U6471 ( .B1(n5299), .B2(n6578), .A(n5276), .ZN(n5277) );
  OAI21_X1 U6472 ( .B1(n5302), .B2(n5278), .A(n5277), .ZN(U3107) );
  AOI22_X1 U6473 ( .A1(n6739), .A2(n5296), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5295), .ZN(n5279) );
  OAI21_X1 U6474 ( .B1(n6680), .B2(n6687), .A(n5279), .ZN(n5280) );
  AOI21_X1 U6475 ( .B1(n5299), .B2(n6675), .A(n5280), .ZN(n5281) );
  OAI21_X1 U6476 ( .B1(n5302), .B2(n5282), .A(n5281), .ZN(U3106) );
  AOI22_X1 U6477 ( .A1(n6727), .A2(n5296), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5295), .ZN(n5283) );
  OAI21_X1 U6478 ( .B1(n6672), .B2(n6687), .A(n5283), .ZN(n5284) );
  AOI21_X1 U6479 ( .B1(n5299), .B2(n6669), .A(n5284), .ZN(n5285) );
  OAI21_X1 U6480 ( .B1(n5302), .B2(n5286), .A(n5285), .ZN(U3104) );
  AOI22_X1 U6481 ( .A1(n6733), .A2(n5296), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5295), .ZN(n5287) );
  OAI21_X1 U6482 ( .B1(n6640), .B2(n6687), .A(n5287), .ZN(n5288) );
  AOI21_X1 U6483 ( .B1(n5299), .B2(n6636), .A(n5288), .ZN(n5289) );
  OAI21_X1 U6484 ( .B1(n5302), .B2(n5290), .A(n5289), .ZN(U3105) );
  AOI22_X1 U6485 ( .A1(n6721), .A2(n5296), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5295), .ZN(n5291) );
  OAI21_X1 U6486 ( .B1(n6634), .B2(n6687), .A(n5291), .ZN(n5292) );
  AOI21_X1 U6487 ( .B1(n5299), .B2(n6630), .A(n5292), .ZN(n5293) );
  OAI21_X1 U6488 ( .B1(n5302), .B2(n5294), .A(n5293), .ZN(U3103) );
  AOI22_X1 U6489 ( .A1(n6714), .A2(n5296), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5295), .ZN(n5297) );
  OAI21_X1 U6490 ( .B1(n6600), .B2(n6687), .A(n5297), .ZN(n5298) );
  AOI21_X1 U6491 ( .B1(n5299), .B2(n6626), .A(n5298), .ZN(n5300) );
  OAI21_X1 U6492 ( .B1(n5302), .B2(n5301), .A(n5300), .ZN(U3102) );
  NAND2_X1 U6493 ( .A1(n5311), .A2(n5303), .ZN(n5304) );
  OAI21_X1 U6494 ( .B1(n6161), .B2(n5309), .A(n6159), .ZN(n6247) );
  OR2_X1 U6495 ( .A1(n6247), .A2(n6841), .ZN(n5316) );
  OAI22_X1 U6496 ( .A1(n5305), .A2(n6203), .B1(n6219), .B2(n6477), .ZN(n5306)
         );
  INV_X1 U6497 ( .A(n5306), .ZN(n5307) );
  AND2_X1 U6498 ( .A1(n6216), .A2(n5307), .ZN(n5315) );
  AOI22_X1 U6499 ( .A1(n5308), .A2(n3092), .B1(n6234), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5314) );
  NOR2_X1 U6500 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5309), .ZN(n5312) );
  AND2_X1 U6501 ( .A1(n5311), .A2(n5310), .ZN(n6236) );
  AOI22_X1 U6502 ( .A1(n6946), .A2(n5312), .B1(n6236), .B2(n6075), .ZN(n5313)
         );
  AND4_X1 U6503 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n5317)
         );
  OAI21_X1 U6504 ( .B1(n6243), .B2(n5318), .A(n5317), .ZN(U2823) );
  AND2_X1 U6505 ( .A1(n5320), .A2(n5319), .ZN(n5325) );
  INV_X1 U6506 ( .A(n5321), .ZN(n5323) );
  NOR2_X1 U6507 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  XNOR2_X1 U6508 ( .A(n5325), .B(n5324), .ZN(n6438) );
  NAND2_X1 U6509 ( .A1(n6438), .A2(n6429), .ZN(n5329) );
  INV_X1 U6510 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5326) );
  NOR2_X1 U6511 ( .A1(n6495), .A2(n5326), .ZN(n6435) );
  NOR2_X1 U6512 ( .A1(n6434), .A2(n6174), .ZN(n5327) );
  AOI211_X1 U6513 ( .C1(n6425), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6435), 
        .B(n5327), .ZN(n5328) );
  OAI211_X1 U6514 ( .C1(n6696), .C2(n5330), .A(n5329), .B(n5328), .ZN(U2975)
         );
  XNOR2_X1 U6515 ( .A(n5795), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5331)
         );
  XNOR2_X1 U6516 ( .A(n5375), .B(n5331), .ZN(n6392) );
  OAI211_X1 U6517 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A(n6437), .B(n5381), .ZN(n5335) );
  INV_X1 U6518 ( .A(n6442), .ZN(n5333) );
  INV_X1 U6519 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6855) );
  OAI22_X1 U6520 ( .A1(n6497), .A2(n6157), .B1(n6855), .B2(n6495), .ZN(n5332)
         );
  AOI21_X1 U6521 ( .B1(n5333), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5332), 
        .ZN(n5334) );
  OAI211_X1 U6522 ( .C1(n6392), .C2(n6476), .A(n5335), .B(n5334), .ZN(U3006)
         );
  OAI21_X1 U6523 ( .B1(n6183), .B2(REIP_REG_1__SCAN_IN), .A(n6147), .ZN(n6231)
         );
  XNOR2_X1 U6524 ( .A(n4686), .B(n5336), .ZN(n6496) );
  INV_X1 U6525 ( .A(n6496), .ZN(n6256) );
  NAND2_X1 U6526 ( .A1(n6240), .A2(n6256), .ZN(n5342) );
  AOI22_X1 U6527 ( .A1(n6235), .A2(EBX_REG_2__SCAN_IN), .B1(n6236), .B2(n5337), 
        .ZN(n5341) );
  INV_X1 U6528 ( .A(n6433), .ZN(n5338) );
  AOI22_X1 U6529 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6234), .B1(n3092), 
        .B2(n5338), .ZN(n5340) );
  INV_X1 U6530 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6230) );
  NAND3_X1 U6531 ( .A1(n6946), .A2(REIP_REG_1__SCAN_IN), .A3(n6230), .ZN(n5339) );
  NAND4_X1 U6532 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n5343)
         );
  AOI21_X1 U6533 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6231), .A(n5343), .ZN(n5344)
         );
  OAI21_X1 U6534 ( .B1(n6243), .B2(n6255), .A(n5344), .ZN(U2825) );
  NOR2_X1 U6535 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5345), .ZN(n5933)
         );
  NAND3_X1 U6536 ( .A1(n5347), .A2(n6554), .A3(n5346), .ZN(n5348) );
  OAI21_X1 U6537 ( .B1(n5349), .B2(n6521), .A(n5348), .ZN(n5930) );
  NOR2_X1 U6538 ( .A1(n5350), .A2(n6934), .ZN(n5353) );
  OAI21_X1 U6539 ( .B1(n5932), .B2(n6635), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5352) );
  AOI211_X1 U6540 ( .C1(n5353), .C2(n5352), .A(n6555), .B(n5351), .ZN(n5354)
         );
  OAI211_X1 U6541 ( .C1(n5933), .C2(n6904), .A(n5354), .B(n6777), .ZN(n5931)
         );
  AOI22_X1 U6542 ( .A1(n5930), .A2(n6720), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n5931), .ZN(n5355) );
  OAI21_X1 U6543 ( .B1(n6649), .B2(n6634), .A(n5355), .ZN(n5356) );
  AOI21_X1 U6544 ( .B1(n6721), .B2(n5933), .A(n5356), .ZN(n5357) );
  OAI21_X1 U6545 ( .B1(n6725), .B2(n5373), .A(n5357), .ZN(U3071) );
  AOI22_X1 U6546 ( .A1(n5930), .A2(n6732), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n5931), .ZN(n5358) );
  OAI21_X1 U6547 ( .B1(n6649), .B2(n6640), .A(n5358), .ZN(n5359) );
  AOI21_X1 U6548 ( .B1(n6733), .B2(n5933), .A(n5359), .ZN(n5360) );
  OAI21_X1 U6549 ( .B1(n6737), .B2(n5373), .A(n5360), .ZN(U3073) );
  AOI22_X1 U6550 ( .A1(n5930), .A2(n6726), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n5931), .ZN(n5361) );
  OAI21_X1 U6551 ( .B1(n6649), .B2(n6672), .A(n5361), .ZN(n5362) );
  AOI21_X1 U6552 ( .B1(n6727), .B2(n5933), .A(n5362), .ZN(n5363) );
  OAI21_X1 U6553 ( .B1(n6731), .B2(n5373), .A(n5363), .ZN(U3072) );
  AOI22_X1 U6554 ( .A1(n5930), .A2(n6745), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n5931), .ZN(n5364) );
  OAI21_X1 U6555 ( .B1(n6649), .B2(n6582), .A(n5364), .ZN(n5365) );
  AOI21_X1 U6556 ( .B1(n6747), .B2(n5933), .A(n5365), .ZN(n5366) );
  OAI21_X1 U6557 ( .B1(n6754), .B2(n5373), .A(n5366), .ZN(U3075) );
  AOI22_X1 U6558 ( .A1(n5930), .A2(n6708), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n5931), .ZN(n5367) );
  OAI21_X1 U6559 ( .B1(n6649), .B2(n6597), .A(n5367), .ZN(n5368) );
  AOI21_X1 U6560 ( .B1(n6709), .B2(n5933), .A(n5368), .ZN(n5369) );
  OAI21_X1 U6561 ( .B1(n6713), .B2(n5373), .A(n5369), .ZN(U3069) );
  AOI22_X1 U6562 ( .A1(n5930), .A2(n6738), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n5931), .ZN(n5370) );
  OAI21_X1 U6563 ( .B1(n6649), .B2(n6680), .A(n5370), .ZN(n5371) );
  AOI21_X1 U6564 ( .B1(n6739), .B2(n5933), .A(n5371), .ZN(n5372) );
  OAI21_X1 U6565 ( .B1(n6743), .B2(n5373), .A(n5372), .ZN(U3074) );
  NAND2_X1 U6566 ( .A1(n5375), .A2(n5374), .ZN(n5377) );
  NAND2_X1 U6567 ( .A1(n5377), .A2(n5376), .ZN(n5401) );
  XOR2_X1 U6568 ( .A(n5400), .B(n5401), .Z(n5394) );
  NAND2_X1 U6569 ( .A1(n5381), .A2(n5378), .ZN(n5379) );
  OAI211_X1 U6570 ( .C1(n6067), .C2(n5380), .A(n6442), .B(n5379), .ZN(n6064)
         );
  NOR2_X1 U6571 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5381), .ZN(n6065)
         );
  AOI22_X1 U6572 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6064), .B1(n6065), .B2(n6437), .ZN(n5387) );
  NAND2_X1 U6573 ( .A1(n5383), .A2(n5382), .ZN(n5396) );
  OAI21_X1 U6574 ( .B1(n5383), .B2(n5382), .A(n5396), .ZN(n5384) );
  INV_X1 U6575 ( .A(n5384), .ZN(n6248) );
  INV_X1 U6576 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5385) );
  NOR2_X1 U6577 ( .A1(n6495), .A2(n5385), .ZN(n5390) );
  AOI21_X1 U6578 ( .B1(n6248), .B2(n6485), .A(n5390), .ZN(n5386) );
  OAI211_X1 U6579 ( .C1(n5394), .C2(n6476), .A(n5387), .B(n5386), .ZN(U3005)
         );
  XOR2_X1 U6580 ( .A(n5389), .B(n5388), .Z(n6273) );
  AOI21_X1 U6581 ( .B1(n6425), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5390), 
        .ZN(n5391) );
  OAI21_X1 U6582 ( .B1(n6434), .B2(n6152), .A(n5391), .ZN(n5392) );
  AOI21_X1 U6583 ( .B1(n6273), .B2(n3085), .A(n5392), .ZN(n5393) );
  OAI21_X1 U6584 ( .B1(n5394), .B2(n6410), .A(n5393), .ZN(U2973) );
  XOR2_X1 U6585 ( .A(n5569), .B(n5570), .Z(n6141) );
  INV_X1 U6586 ( .A(n6141), .ZN(n5399) );
  INV_X1 U6587 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6588 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6589 ( .A1(n5574), .A2(n5397), .ZN(n6136) );
  OAI222_X1 U6590 ( .A1(n5399), .A2(n6014), .B1(n5398), .B2(n6261), .C1(n5663), 
        .C2(n6136), .ZN(U2845) );
  INV_X1 U6591 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6303) );
  OAI222_X1 U6592 ( .A1(n5399), .A2(n6277), .B1(n6275), .B2(n6381), .C1(n6276), 
        .C2(n6303), .ZN(U2877) );
  NAND2_X1 U6593 ( .A1(n5807), .A2(n5402), .ZN(n5404) );
  NAND2_X1 U6594 ( .A1(n5404), .A2(n5403), .ZN(n5805) );
  OAI21_X1 U6595 ( .B1(n5404), .B2(n5403), .A(n5805), .ZN(n5405) );
  INV_X1 U6596 ( .A(n5405), .ZN(n6068) );
  AOI22_X1 U6597 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6483), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5406) );
  OAI21_X1 U6598 ( .B1(n6434), .B2(n6139), .A(n5406), .ZN(n5407) );
  AOI21_X1 U6599 ( .B1(n6141), .B2(n3085), .A(n5407), .ZN(n5408) );
  OAI21_X1 U6600 ( .B1(n6068), .B2(n6410), .A(n5408), .ZN(U2972) );
  INV_X1 U6601 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6872) );
  INV_X1 U6602 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6862) );
  INV_X1 U6603 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6852) );
  INV_X1 U6604 ( .A(n5409), .ZN(n5410) );
  NOR2_X1 U6605 ( .A1(n5411), .A2(n5410), .ZN(n6188) );
  NAND2_X1 U6606 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6188), .ZN(n6182) );
  NOR2_X1 U6607 ( .A1(n6852), .A2(n6182), .ZN(n6169) );
  NAND2_X1 U6608 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6169), .ZN(n6160) );
  NOR2_X1 U6609 ( .A1(n6855), .A2(n6160), .ZN(n5420) );
  NAND4_X1 U6610 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n5420), .A4(n6147), .ZN(n5577) );
  NAND2_X1 U6611 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n6122) );
  NOR3_X1 U6612 ( .A1(n6862), .A2(n5577), .A3(n6122), .ZN(n6006) );
  NAND4_X1 U6613 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6006), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5975) );
  NOR4_X1 U6614 ( .A1(n6867), .A2(n6869), .A3(n6872), .A4(n5975), .ZN(n5552)
         );
  INV_X1 U6615 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6875) );
  NOR3_X1 U6616 ( .A1(n6873), .A2(n6880), .A3(n6875), .ZN(n5412) );
  AOI21_X1 U6617 ( .B1(n5552), .B2(n5412), .A(n6007), .ZN(n5962) );
  AND2_X1 U6618 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5413) );
  NOR2_X1 U6619 ( .A1(n6183), .A2(n5413), .ZN(n5414) );
  OR2_X1 U6620 ( .A1(n5962), .A2(n5414), .ZN(n5941) );
  INV_X1 U6621 ( .A(n5941), .ZN(n5488) );
  AOI22_X1 U6622 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6234), .B1(n5415), 
        .B2(n6233), .ZN(n5416) );
  OAI21_X1 U6623 ( .B1(n5488), .B2(n6886), .A(n5416), .ZN(n5419) );
  INV_X1 U6624 ( .A(n5417), .ZN(n5598) );
  OAI22_X1 U6625 ( .A1(n5693), .A2(n6128), .B1(n5598), .B2(n6219), .ZN(n5418)
         );
  AOI211_X1 U6626 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6235), .A(n5419), .B(n5418), 
        .ZN(n5422) );
  NAND2_X1 U6627 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n6005) );
  NAND2_X1 U6628 ( .A1(n6946), .A2(n5420), .ZN(n6150) );
  NOR2_X1 U6629 ( .A1(n5385), .A2(n6150), .ZN(n6135) );
  NAND2_X1 U6630 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6135), .ZN(n6124) );
  NOR2_X1 U6631 ( .A1(n6122), .A2(n6124), .ZN(n6118) );
  NAND2_X1 U6632 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6118), .ZN(n6112) );
  NOR2_X1 U6633 ( .A1(n6005), .A2(n6112), .ZN(n6001) );
  NAND2_X1 U6634 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6001), .ZN(n5976) );
  NOR2_X1 U6635 ( .A1(n6869), .A2(n5976), .ZN(n5980) );
  NAND2_X1 U6636 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5980), .ZN(n5973) );
  NOR2_X1 U6637 ( .A1(n6872), .A2(n5973), .ZN(n5553) );
  NAND4_X1 U6638 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .A4(n5553), .ZN(n5955) );
  INV_X1 U6639 ( .A(n5955), .ZN(n5487) );
  NAND3_X1 U6640 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6886), .A3(n5487), .ZN(
        n5421) );
  NAND2_X1 U6641 ( .A1(n5422), .A2(n5421), .ZN(U2799) );
  AOI22_X1 U6642 ( .A1(n5436), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5448), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5426) );
  AOI22_X1 U6643 ( .A1(n3084), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5425) );
  AOI22_X1 U6644 ( .A1(n3303), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5424) );
  AOI22_X1 U6645 ( .A1(n3152), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5423) );
  NAND4_X1 U6646 ( .A1(n5426), .A2(n5425), .A3(n5424), .A4(n5423), .ZN(n5433)
         );
  AOI22_X1 U6647 ( .A1(n5437), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5431) );
  AOI22_X1 U6648 ( .A1(n4217), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5430) );
  AOI22_X1 U6649 ( .A1(n3302), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5429) );
  AOI22_X1 U6650 ( .A1(n3425), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5428) );
  NAND4_X1 U6651 ( .A1(n5431), .A2(n5430), .A3(n5429), .A4(n5428), .ZN(n5432)
         );
  NOR2_X1 U6652 ( .A1(n5433), .A2(n5432), .ZN(n5466) );
  NAND2_X1 U6653 ( .A1(n5435), .A2(n5434), .ZN(n5465) );
  NOR2_X1 U6654 ( .A1(n5466), .A2(n5465), .ZN(n5456) );
  AOI22_X1 U6655 ( .A1(n5437), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5444) );
  AOI22_X1 U6656 ( .A1(n5438), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5443) );
  AOI22_X1 U6657 ( .A1(n4217), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5439), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5442) );
  AOI22_X1 U6658 ( .A1(n4105), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5440), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5441) );
  NAND4_X1 U6659 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n5454)
         );
  AOI22_X1 U6660 ( .A1(n3084), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5445), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5452) );
  AOI22_X1 U6661 ( .A1(n3425), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5451) );
  AOI22_X1 U6662 ( .A1(n3152), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3088), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5450) );
  AOI22_X1 U6663 ( .A1(n5448), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5447), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5449) );
  NAND4_X1 U6664 ( .A1(n5452), .A2(n5451), .A3(n5450), .A4(n5449), .ZN(n5453)
         );
  NOR2_X1 U6665 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  XNOR2_X1 U6666 ( .A(n5456), .B(n5455), .ZN(n5458) );
  NAND2_X1 U6667 ( .A1(n5458), .A2(n5457), .ZN(n5462) );
  OAI21_X1 U6668 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5491), .A(n5473), .ZN(
        n5459) );
  AOI21_X1 U6669 ( .B1(n5531), .B2(EAX_REG_30__SCAN_IN), .A(n5459), .ZN(n5461)
         );
  XNOR2_X1 U6670 ( .A(n5463), .B(n5491), .ZN(n5490) );
  NOR2_X1 U6671 ( .A1(n5490), .A2(n5473), .ZN(n5460) );
  AOI21_X1 U6672 ( .B1(n5462), .B2(n5461), .A(n5460), .ZN(n5532) );
  OAI21_X1 U6673 ( .B1(n5464), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5463), 
        .ZN(n5938) );
  XNOR2_X1 U6674 ( .A(n5466), .B(n5465), .ZN(n5471) );
  AOI21_X1 U6675 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6937), .A(n5467), 
        .ZN(n5469) );
  NAND2_X1 U6676 ( .A1(n5531), .A2(EAX_REG_29__SCAN_IN), .ZN(n5468) );
  OAI211_X1 U6677 ( .C1(n5471), .C2(n5470), .A(n5469), .B(n5468), .ZN(n5472)
         );
  OAI21_X1 U6678 ( .B1(n5473), .B2(n5938), .A(n5472), .ZN(n5480) );
  XOR2_X1 U6679 ( .A(n5532), .B(n5533), .Z(n5486) );
  AOI21_X1 U6680 ( .B1(n6425), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5474), 
        .ZN(n5475) );
  OAI21_X1 U6681 ( .B1(n6434), .B2(n5490), .A(n5475), .ZN(n5476) );
  AOI21_X1 U6682 ( .B1(n5486), .B2(n3085), .A(n5476), .ZN(n5477) );
  OAI21_X1 U6683 ( .B1(n5478), .B2(n6410), .A(n5477), .ZN(U2956) );
  AOI21_X1 U6684 ( .B1(n5480), .B2(n5479), .A(n5533), .ZN(n6018) );
  NAND2_X1 U6685 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5481)
         );
  OAI211_X1 U6686 ( .C1(n6434), .C2(n5938), .A(n5482), .B(n5481), .ZN(n5483)
         );
  AOI21_X1 U6687 ( .B1(n6018), .B2(n3085), .A(n5483), .ZN(n5484) );
  OAI21_X1 U6688 ( .B1(n5485), .B2(n6410), .A(n5484), .ZN(U2957) );
  INV_X1 U6689 ( .A(n5486), .ZN(n5690) );
  NAND3_X1 U6690 ( .A1(n5487), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5944) );
  OAI21_X1 U6691 ( .B1(n5944), .B2(n5537), .A(n5488), .ZN(n5545) );
  OAI21_X1 U6692 ( .B1(n6888), .B2(n5944), .A(n6892), .ZN(n5495) );
  INV_X1 U6693 ( .A(n5489), .ZN(n5594) );
  OAI22_X1 U6694 ( .A1(n5491), .A2(n6170), .B1(n5490), .B2(n6229), .ZN(n5492)
         );
  AOI21_X1 U6695 ( .B1(n6235), .B2(EBX_REG_30__SCAN_IN), .A(n5492), .ZN(n5493)
         );
  OAI21_X1 U6696 ( .B1(n5594), .B2(n6219), .A(n5493), .ZN(n5494) );
  OAI21_X1 U6697 ( .B1(n5690), .B2(n6128), .A(n5496), .ZN(U2797) );
  INV_X1 U6698 ( .A(n6797), .ZN(n6908) );
  INV_X1 U6699 ( .A(n6916), .ZN(n5497) );
  AOI21_X1 U6700 ( .B1(n6908), .B2(n5498), .A(n5497), .ZN(n5506) );
  NOR3_X1 U6701 ( .A1(n6797), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5498), 
        .ZN(n5503) );
  OAI22_X1 U6702 ( .A1(n5501), .A2(n6918), .B1(n5500), .B2(n5499), .ZN(n5502)
         );
  OAI21_X1 U6703 ( .B1(n5503), .B2(n5502), .A(n6916), .ZN(n5504) );
  OAI21_X1 U6704 ( .B1(n5506), .B2(n5505), .A(n5504), .ZN(U3459) );
  OAI21_X1 U6705 ( .B1(n3513), .B2(n3544), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n5507) );
  OAI21_X1 U6706 ( .B1(n5508), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5507), 
        .ZN(n5509) );
  XNOR2_X1 U6707 ( .A(n5511), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5713)
         );
  INV_X1 U6708 ( .A(n5833), .ZN(n5844) );
  AOI211_X1 U6709 ( .C1(n5844), .C2(n5921), .A(n4616), .B(n5512), .ZN(n5513)
         );
  INV_X1 U6710 ( .A(n5513), .ZN(n5527) );
  INV_X1 U6711 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U6712 ( .A1(n5515), .A2(n3091), .ZN(n5517) );
  OAI211_X1 U6713 ( .C1(n5519), .C2(n5518), .A(n5517), .B(n5516), .ZN(n5524)
         );
  AOI22_X1 U6714 ( .A1(n5521), .A2(EBX_REG_31__SCAN_IN), .B1(n5520), .B2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5522) );
  INV_X1 U6715 ( .A(n5522), .ZN(n5523) );
  XNOR2_X1 U6716 ( .A(n5524), .B(n5523), .ZN(n5543) );
  INV_X1 U6717 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5536) );
  NOR2_X1 U6718 ( .A1(n6495), .A2(n5536), .ZN(n5707) );
  INV_X1 U6719 ( .A(n5707), .ZN(n5526) );
  OAI21_X1 U6720 ( .B1(n5713), .B2(n6476), .A(n5528), .ZN(U2987) );
  OAI22_X1 U6721 ( .A1(n5543), .A2(n5663), .B1(n6261), .B2(n5529), .ZN(U2828)
         );
  AOI22_X1 U6722 ( .A1(n5531), .A2(EAX_REG_31__SCAN_IN), .B1(n5530), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6723 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  XOR2_X1 U6724 ( .A(n5535), .B(n5534), .Z(n5711) );
  INV_X1 U6725 ( .A(n5711), .ZN(n5547) );
  INV_X1 U6726 ( .A(n5944), .ZN(n5538) );
  NAND3_X1 U6727 ( .A1(n5538), .A2(n5537), .A3(n5536), .ZN(n5542) );
  AOI22_X1 U6728 ( .A1(n5540), .A2(n5539), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n6234), .ZN(n5541) );
  OAI211_X1 U6729 ( .C1(n5543), .C2(n6219), .A(n5542), .B(n5541), .ZN(n5544)
         );
  AOI21_X1 U6730 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5545), .A(n5544), .ZN(n5546) );
  OAI21_X1 U6731 ( .B1(n5547), .B2(n6128), .A(n5546), .ZN(U2796) );
  INV_X1 U6732 ( .A(n5548), .ZN(n5551) );
  INV_X1 U6733 ( .A(n5549), .ZN(n5562) );
  INV_X1 U6734 ( .A(n5609), .ZN(n5550) );
  NAND2_X1 U6735 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5553), .ZN(n5957) );
  OAI22_X1 U6736 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5957), .B1(n5729), .B2(
        n6229), .ZN(n5560) );
  OR2_X1 U6737 ( .A1(n6007), .A2(n5552), .ZN(n5974) );
  NAND2_X1 U6738 ( .A1(n6873), .A2(n5553), .ZN(n5568) );
  AOI21_X1 U6739 ( .B1(n5974), .B2(n5568), .A(n6875), .ZN(n5559) );
  OAI21_X1 U6740 ( .B1(n5556), .B2(n5555), .A(n5554), .ZN(n5837) );
  AOI22_X1 U6741 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6235), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6234), .ZN(n5557) );
  OAI21_X1 U6742 ( .B1(n5837), .B2(n6219), .A(n5557), .ZN(n5558) );
  NOR3_X1 U6743 ( .A1(n5560), .A2(n5559), .A3(n5558), .ZN(n5561) );
  OAI21_X1 U6744 ( .B1(n6025), .B2(n6128), .A(n5561), .ZN(U2802) );
  AOI21_X1 U6745 ( .B1(n5563), .B2(n5622), .A(n5562), .ZN(n5737) );
  INV_X1 U6746 ( .A(n5737), .ZN(n5698) );
  OAI22_X1 U6747 ( .A1(n5616), .A2(n6203), .B1(n5564), .B2(n6170), .ZN(n5566)
         );
  OAI22_X1 U6748 ( .A1(n6873), .A2(n5974), .B1(n5735), .B2(n6229), .ZN(n5565)
         );
  AOI211_X1 U6749 ( .C1(n6240), .C2(n5618), .A(n5566), .B(n5565), .ZN(n5567)
         );
  OAI211_X1 U6750 ( .C1(n5698), .C2(n6128), .A(n5568), .B(n5567), .ZN(U2803)
         );
  OR2_X1 U6751 ( .A1(n5631), .A2(n5572), .ZN(n5673) );
  INV_X1 U6752 ( .A(n5673), .ZN(n5571) );
  AOI21_X1 U6753 ( .B1(n5572), .B2(n5631), .A(n5571), .ZN(n5817) );
  INV_X1 U6754 ( .A(n5817), .ZN(n5706) );
  AOI21_X1 U6755 ( .B1(n5575), .B2(n5574), .A(n5573), .ZN(n5901) );
  INV_X1 U6756 ( .A(n5576), .ZN(n5815) );
  OAI22_X1 U6757 ( .A1(n6203), .A2(n4530), .B1(n5815), .B2(n6229), .ZN(n5580)
         );
  NAND2_X1 U6758 ( .A1(n6159), .A2(n5577), .ZN(n6144) );
  AOI21_X1 U6759 ( .B1(n6234), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6209), 
        .ZN(n5578) );
  OAI221_X1 U6760 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6124), .C1(n6858), .C2(
        n6144), .A(n5578), .ZN(n5579) );
  AOI211_X1 U6761 ( .C1(n5901), .C2(n6240), .A(n5580), .B(n5579), .ZN(n5581)
         );
  OAI21_X1 U6762 ( .B1(n5706), .B2(n6128), .A(n5581), .ZN(U2812) );
  NAND2_X1 U6763 ( .A1(n6235), .A2(EBX_REG_1__SCAN_IN), .ZN(n5583) );
  AOI22_X1 U6764 ( .A1(n6234), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6161), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5582) );
  OAI211_X1 U6765 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6229), .A(n5583), 
        .B(n5582), .ZN(n5584) );
  AOI21_X1 U6766 ( .B1(n6240), .B2(n4651), .A(n5584), .ZN(n5586) );
  AOI22_X1 U6767 ( .A1(n6946), .A2(n6921), .B1(n6236), .B2(n4618), .ZN(n5585)
         );
  OAI211_X1 U6768 ( .C1(n6243), .C2(n5587), .A(n5586), .B(n5585), .ZN(U2826)
         );
  OAI22_X1 U6769 ( .A1(n6203), .A2(n5588), .B1(n6243), .B2(n6278), .ZN(n5589)
         );
  AOI21_X1 U6770 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6159), .A(n5589), .ZN(n5592)
         );
  NAND2_X1 U6771 ( .A1(n6170), .A2(n6229), .ZN(n5590) );
  AOI22_X1 U6772 ( .A1(n5590), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6236), 
        .B2(n6653), .ZN(n5591) );
  OAI211_X1 U6773 ( .C1(n6219), .C2(n5593), .A(n5592), .B(n5591), .ZN(U2827)
         );
  INV_X1 U6774 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5595) );
  OAI222_X1 U6775 ( .A1(n6014), .A2(n5690), .B1(n5595), .B2(n6261), .C1(n5663), 
        .C2(n5594), .ZN(U2829) );
  INV_X1 U6776 ( .A(n6018), .ZN(n5597) );
  OAI222_X1 U6777 ( .A1(n6014), .A2(n5597), .B1(n5596), .B2(n6261), .C1(n5947), 
        .C2(n5663), .ZN(U2830) );
  INV_X1 U6778 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5599) );
  OAI222_X1 U6779 ( .A1(n6014), .A2(n5693), .B1(n6261), .B2(n5599), .C1(n5598), 
        .C2(n5663), .ZN(U2831) );
  NOR2_X1 U6780 ( .A1(n5600), .A2(n5601), .ZN(n5602) );
  INV_X1 U6781 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U6782 ( .A1(n5613), .A2(n5604), .ZN(n5605) );
  NAND2_X1 U6783 ( .A1(n5606), .A2(n5605), .ZN(n5951) );
  OAI222_X1 U6784 ( .A1(n6014), .A2(n6021), .B1(n5607), .B2(n6261), .C1(n5951), 
        .C2(n5663), .ZN(U2832) );
  NOR2_X1 U6785 ( .A1(n5609), .A2(n5608), .ZN(n5610) );
  NAND2_X1 U6786 ( .A1(n5554), .A2(n5611), .ZN(n5612) );
  NAND2_X1 U6787 ( .A1(n5613), .A2(n5612), .ZN(n5958) );
  OAI222_X1 U6788 ( .A1(n6014), .A2(n5959), .B1(n6261), .B2(n5614), .C1(n5958), 
        .C2(n5663), .ZN(U2833) );
  OAI222_X1 U6789 ( .A1(n5663), .A2(n5837), .B1(n5615), .B2(n6261), .C1(n6014), 
        .C2(n6025), .ZN(U2834) );
  NOR2_X1 U6790 ( .A1(n6261), .A2(n5616), .ZN(n5617) );
  AOI21_X1 U6791 ( .B1(n5618), .B2(n6257), .A(n5617), .ZN(n5619) );
  OAI21_X1 U6792 ( .B1(n5698), .B2(n6014), .A(n5619), .ZN(U2835) );
  NAND2_X1 U6793 ( .A1(n5621), .A2(n5620), .ZN(n5633) );
  INV_X1 U6794 ( .A(n5622), .ZN(n5623) );
  AOI21_X1 U6795 ( .B1(n5624), .B2(n5633), .A(n5623), .ZN(n6029) );
  INV_X1 U6796 ( .A(n6029), .ZN(n5969) );
  INV_X1 U6797 ( .A(n5626), .ZN(n5627) );
  AOI21_X1 U6798 ( .B1(n5628), .B2(n5625), .A(n5627), .ZN(n5967) );
  AOI22_X1 U6799 ( .A1(n5967), .A2(n6257), .B1(EBX_REG_23__SCAN_IN), .B2(n5680), .ZN(n5629) );
  OAI21_X1 U6800 ( .B1(n5969), .B2(n6014), .A(n5629), .ZN(U2836) );
  INV_X1 U6801 ( .A(n5666), .ZN(n5657) );
  OR2_X1 U6802 ( .A1(n5647), .A2(n5635), .ZN(n5636) );
  NAND2_X1 U6803 ( .A1(n5625), .A2(n5636), .ZN(n5986) );
  OAI22_X1 U6804 ( .A1(n5986), .A2(n5663), .B1(n5637), .B2(n6261), .ZN(n5638)
         );
  INV_X1 U6805 ( .A(n5638), .ZN(n5639) );
  OAI21_X1 U6806 ( .B1(n5983), .B2(n6014), .A(n5639), .ZN(U2837) );
  NOR2_X1 U6807 ( .A1(n5666), .A2(n5640), .ZN(n5650) );
  NOR2_X1 U6808 ( .A1(n5650), .A2(n5641), .ZN(n5642) );
  INV_X1 U6809 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5648) );
  NOR2_X1 U6810 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  OR2_X1 U6811 ( .A1(n5647), .A2(n5646), .ZN(n5996) );
  OAI222_X1 U6812 ( .A1(n6014), .A2(n6032), .B1(n5648), .B2(n6261), .C1(n5996), 
        .C2(n5663), .ZN(U2838) );
  MUX2_X1 U6813 ( .A(n5660), .B(n5659), .S(n5652), .Z(n5653) );
  XOR2_X1 U6814 ( .A(n5654), .B(n5653), .Z(n5875) );
  INV_X1 U6815 ( .A(n5875), .ZN(n5998) );
  OAI222_X1 U6816 ( .A1(n5999), .A2(n6014), .B1(n6261), .B2(n3701), .C1(n5663), 
        .C2(n5998), .ZN(U2839) );
  INV_X1 U6817 ( .A(n5655), .ZN(n5656) );
  OAI21_X1 U6818 ( .B1(n5657), .B2(n5656), .A(n5778), .ZN(n6108) );
  INV_X1 U6819 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6106) );
  XNOR2_X1 U6820 ( .A(n5660), .B(n5659), .ZN(n5661) );
  NOR2_X1 U6821 ( .A1(n5669), .A2(n5661), .ZN(n5883) );
  AND2_X1 U6822 ( .A1(n5669), .A2(n5661), .ZN(n5662) );
  OR2_X1 U6823 ( .A1(n5883), .A2(n5662), .ZN(n6049) );
  OAI222_X1 U6824 ( .A1(n6108), .A2(n6014), .B1(n6106), .B2(n6261), .C1(n6049), 
        .C2(n5663), .ZN(U2841) );
  OR2_X1 U6825 ( .A1(n5675), .A2(n5664), .ZN(n5665) );
  INV_X1 U6826 ( .A(n6266), .ZN(n5671) );
  NAND2_X1 U6827 ( .A1(n5678), .A2(n5667), .ZN(n5668) );
  AND2_X1 U6828 ( .A1(n5669), .A2(n5668), .ZN(n6116) );
  AOI22_X1 U6829 ( .A1(n6116), .A2(n6257), .B1(EBX_REG_17__SCAN_IN), .B2(n5680), .ZN(n5670) );
  OAI21_X1 U6830 ( .B1(n5671), .B2(n6014), .A(n5670), .ZN(U2842) );
  AND2_X1 U6831 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  OR2_X1 U6832 ( .A1(n5675), .A2(n5674), .ZN(n6129) );
  OR2_X1 U6833 ( .A1(n5573), .A2(n5676), .ZN(n5677) );
  AND2_X1 U6834 ( .A1(n5678), .A2(n5677), .ZN(n6126) );
  AOI22_X1 U6835 ( .A1(n6126), .A2(n6257), .B1(EBX_REG_16__SCAN_IN), .B2(n5680), .ZN(n5679) );
  OAI21_X1 U6836 ( .B1(n6129), .B2(n6014), .A(n5679), .ZN(U2843) );
  AOI22_X1 U6837 ( .A1(n5901), .A2(n6257), .B1(EBX_REG_15__SCAN_IN), .B2(n5680), .ZN(n5681) );
  OAI21_X1 U6838 ( .B1(n5706), .B2(n6014), .A(n5681), .ZN(U2844) );
  NAND3_X1 U6839 ( .A1(n5711), .A2(n5682), .A3(n6276), .ZN(n5685) );
  NOR2_X2 U6840 ( .A1(n6267), .A2(n5683), .ZN(n6265) );
  AOI22_X1 U6841 ( .A1(n6265), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6267), .ZN(n5684) );
  NAND2_X1 U6842 ( .A1(n5685), .A2(n5684), .ZN(U2860) );
  AOI22_X1 U6843 ( .A1(n6265), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6267), .ZN(n5689) );
  AND2_X1 U6844 ( .A1(n3614), .A2(n5686), .ZN(n5687) );
  NAND2_X1 U6845 ( .A1(n6268), .A2(DATAI_14_), .ZN(n5688) );
  OAI211_X1 U6846 ( .C1(n5690), .C2(n6277), .A(n5689), .B(n5688), .ZN(U2861)
         );
  AOI22_X1 U6847 ( .A1(n6268), .A2(DATAI_12_), .B1(n6267), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6848 ( .A1(n6265), .A2(DATAI_28_), .ZN(n5691) );
  OAI211_X1 U6849 ( .C1(n5693), .C2(n6277), .A(n5692), .B(n5691), .ZN(U2863)
         );
  AOI22_X1 U6850 ( .A1(n6268), .A2(DATAI_10_), .B1(n6267), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U6851 ( .A1(n6265), .A2(DATAI_26_), .ZN(n5694) );
  OAI211_X1 U6852 ( .C1(n5959), .C2(n6277), .A(n5695), .B(n5694), .ZN(U2865)
         );
  AOI22_X1 U6853 ( .A1(n6265), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6267), .ZN(n5697) );
  NAND2_X1 U6854 ( .A1(n6268), .A2(DATAI_8_), .ZN(n5696) );
  OAI211_X1 U6855 ( .C1(n5698), .C2(n6277), .A(n5697), .B(n5696), .ZN(U2867)
         );
  AOI22_X1 U6856 ( .A1(n6268), .A2(DATAI_6_), .B1(n6267), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U6857 ( .A1(n6265), .A2(DATAI_22_), .ZN(n5699) );
  OAI211_X1 U6858 ( .C1(n5983), .C2(n6277), .A(n5700), .B(n5699), .ZN(U2869)
         );
  AOI22_X1 U6859 ( .A1(n6268), .A2(DATAI_4_), .B1(n6267), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6860 ( .A1(n6265), .A2(DATAI_20_), .ZN(n5701) );
  OAI211_X1 U6861 ( .C1(n5999), .C2(n6277), .A(n5702), .B(n5701), .ZN(U2871)
         );
  AOI22_X1 U6862 ( .A1(n6265), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6267), .ZN(n5704) );
  NAND2_X1 U6863 ( .A1(n6268), .A2(DATAI_0_), .ZN(n5703) );
  OAI211_X1 U6864 ( .C1(n6129), .C2(n6277), .A(n5704), .B(n5703), .ZN(U2875)
         );
  AOI22_X1 U6865 ( .A1(n6271), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6267), .ZN(n5705) );
  OAI21_X1 U6866 ( .B1(n5706), .B2(n6277), .A(n5705), .ZN(U2876) );
  AOI21_X1 U6867 ( .B1(n6425), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5707), 
        .ZN(n5708) );
  OAI21_X1 U6868 ( .B1(n5709), .B2(n6434), .A(n5708), .ZN(n5710) );
  AOI21_X1 U6869 ( .B1(n5711), .B2(n3085), .A(n5710), .ZN(n5712) );
  OAI21_X1 U6870 ( .B1(n5713), .B2(n6410), .A(n5712), .ZN(U2955) );
  NAND2_X1 U6871 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  XNOR2_X1 U6872 ( .A(n5716), .B(n5821), .ZN(n5826) );
  NAND2_X1 U6873 ( .A1(n5826), .A2(n6429), .ZN(n5719) );
  INV_X1 U6874 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6882) );
  NOR2_X1 U6875 ( .A1(n6495), .A2(n6882), .ZN(n5820) );
  NOR2_X1 U6876 ( .A1(n6434), .A2(n5949), .ZN(n5717) );
  AOI211_X1 U6877 ( .C1(n6425), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5820), 
        .B(n5717), .ZN(n5718) );
  OAI211_X1 U6878 ( .C1(n6696), .C2(n6021), .A(n5719), .B(n5718), .ZN(U2959)
         );
  INV_X1 U6879 ( .A(n5720), .ZN(n5722) );
  NOR2_X1 U6880 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  XOR2_X1 U6881 ( .A(n5723), .B(n3779), .Z(n5835) );
  OR2_X1 U6882 ( .A1(n6495), .A2(n6880), .ZN(n5831) );
  OAI21_X1 U6883 ( .B1(n5800), .B2(n5965), .A(n5831), .ZN(n5725) );
  NOR2_X1 U6884 ( .A1(n5959), .A2(n6696), .ZN(n5724) );
  AOI211_X1 U6885 ( .C1(n6387), .C2(n5956), .A(n5725), .B(n5724), .ZN(n5726)
         );
  OAI21_X1 U6886 ( .B1(n5835), .B2(n6410), .A(n5726), .ZN(U2960) );
  OAI21_X1 U6887 ( .B1(n5728), .B2(n5727), .A(n3780), .ZN(n5836) );
  NAND2_X1 U6888 ( .A1(n5836), .A2(n6429), .ZN(n5732) );
  NOR2_X1 U6889 ( .A1(n6495), .A2(n6875), .ZN(n5839) );
  NOR2_X1 U6890 ( .A1(n6434), .A2(n5729), .ZN(n5730) );
  AOI211_X1 U6891 ( .C1(n6425), .C2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5839), 
        .B(n5730), .ZN(n5731) );
  OAI211_X1 U6892 ( .C1(n6696), .C2(n6025), .A(n5732), .B(n5731), .ZN(U2961)
         );
  AOI21_X1 U6893 ( .B1(n6425), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5733), 
        .ZN(n5734) );
  OAI21_X1 U6894 ( .B1(n6434), .B2(n5735), .A(n5734), .ZN(n5736) );
  AOI21_X1 U6895 ( .B1(n5737), .B2(n3085), .A(n5736), .ZN(n5738) );
  OAI21_X1 U6896 ( .B1(n5739), .B2(n6410), .A(n5738), .ZN(U2962) );
  OR2_X1 U6897 ( .A1(n5795), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5746)
         );
  NOR2_X1 U6898 ( .A1(n3513), .A2(n5860), .ZN(n5745) );
  NAND4_X1 U6899 ( .A1(n5772), .A2(n5872), .A3(INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n5745), .ZN(n5740) );
  OAI21_X1 U6900 ( .B1(n5753), .B2(n5746), .A(n5740), .ZN(n5741) );
  XNOR2_X1 U6901 ( .A(n5741), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5851)
         );
  NOR2_X1 U6902 ( .A1(n6495), .A2(n6872), .ZN(n5847) );
  AOI21_X1 U6903 ( .B1(n6425), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5847), 
        .ZN(n5742) );
  OAI21_X1 U6904 ( .B1(n6434), .B2(n5966), .A(n5742), .ZN(n5743) );
  AOI21_X1 U6905 ( .B1(n6029), .B2(n3085), .A(n5743), .ZN(n5744) );
  OAI21_X1 U6906 ( .B1(n5851), .B2(n6410), .A(n5744), .ZN(U2963) );
  INV_X1 U6907 ( .A(n5745), .ZN(n5747) );
  NAND2_X1 U6908 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  XNOR2_X1 U6909 ( .A(n5749), .B(n5748), .ZN(n5852) );
  NAND2_X1 U6910 ( .A1(n5852), .A2(n6429), .ZN(n5752) );
  NOR2_X1 U6911 ( .A1(n6495), .A2(n6867), .ZN(n5856) );
  NOR2_X1 U6912 ( .A1(n6434), .A2(n5977), .ZN(n5750) );
  AOI211_X1 U6913 ( .C1(n6425), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5856), 
        .B(n5750), .ZN(n5751) );
  OAI211_X1 U6914 ( .C1(n6696), .C2(n5983), .A(n5752), .B(n5751), .ZN(U2964)
         );
  OAI21_X1 U6915 ( .B1(n5755), .B2(n5754), .A(n5753), .ZN(n5861) );
  NAND2_X1 U6916 ( .A1(n5861), .A2(n6429), .ZN(n5759) );
  NOR2_X1 U6917 ( .A1(n6495), .A2(n6869), .ZN(n5864) );
  NOR2_X1 U6918 ( .A1(n5800), .A2(n5756), .ZN(n5757) );
  AOI211_X1 U6919 ( .C1(n6387), .C2(n5987), .A(n5864), .B(n5757), .ZN(n5758)
         );
  OAI211_X1 U6920 ( .C1(n6696), .C2(n6032), .A(n5759), .B(n5758), .ZN(U2965)
         );
  NAND2_X1 U6921 ( .A1(n4289), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5764) );
  OR2_X1 U6922 ( .A1(n6042), .A2(n5760), .ZN(n5763) );
  NAND2_X1 U6923 ( .A1(n3513), .A2(n5761), .ZN(n5762) );
  OAI22_X1 U6924 ( .A1(n5774), .A2(n5764), .B1(n5763), .B2(n5762), .ZN(n5765)
         );
  XNOR2_X1 U6925 ( .A(n5765), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5881)
         );
  INV_X1 U6926 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5766) );
  NOR2_X1 U6927 ( .A1(n6495), .A2(n5766), .ZN(n5874) );
  NOR2_X1 U6928 ( .A1(n5800), .A2(n5767), .ZN(n5768) );
  AOI211_X1 U6929 ( .C1(n6387), .C2(n5997), .A(n5874), .B(n5768), .ZN(n5771)
         );
  INV_X1 U6930 ( .A(n5999), .ZN(n5769) );
  NAND2_X1 U6931 ( .A1(n5769), .A2(n3085), .ZN(n5770) );
  OAI211_X1 U6932 ( .C1(n5881), .C2(n6410), .A(n5771), .B(n5770), .ZN(U2966)
         );
  OAI21_X1 U6933 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5775) );
  INV_X1 U6934 ( .A(n5775), .ZN(n5890) );
  INV_X1 U6935 ( .A(n5776), .ZN(n5777) );
  INV_X1 U6936 ( .A(n6008), .ZN(n5781) );
  AOI22_X1 U6937 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6483), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5780) );
  OAI21_X1 U6938 ( .B1(n6434), .B2(n5781), .A(n5780), .ZN(n5782) );
  AOI21_X1 U6939 ( .B1(n6036), .B2(n3085), .A(n5782), .ZN(n5783) );
  OAI21_X1 U6940 ( .B1(n5890), .B2(n6410), .A(n5783), .ZN(U2967) );
  NAND2_X1 U6941 ( .A1(n5807), .A2(n5784), .ZN(n5786) );
  INV_X1 U6942 ( .A(n5797), .ZN(n5787) );
  NAND2_X1 U6943 ( .A1(n3513), .A2(n6059), .ZN(n6041) );
  NOR3_X1 U6944 ( .A1(n5787), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6041), 
        .ZN(n6043) );
  NAND2_X1 U6945 ( .A1(n4289), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6039) );
  NOR2_X1 U6946 ( .A1(n5788), .A2(n6039), .ZN(n6046) );
  NOR2_X1 U6947 ( .A1(n6043), .A2(n6046), .ZN(n5789) );
  XNOR2_X1 U6948 ( .A(n5789), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6050)
         );
  NAND2_X1 U6949 ( .A1(n6050), .A2(n6429), .ZN(n5794) );
  INV_X1 U6950 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5790) );
  OAI22_X1 U6951 ( .A1(n5800), .A2(n5791), .B1(n6495), .B2(n5790), .ZN(n5792)
         );
  AOI21_X1 U6952 ( .B1(n6387), .B2(n6104), .A(n5792), .ZN(n5793) );
  OAI211_X1 U6953 ( .C1(n6696), .C2(n6108), .A(n5794), .B(n5793), .ZN(U2968)
         );
  XNOR2_X1 U6954 ( .A(n5795), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5796)
         );
  XNOR2_X1 U6955 ( .A(n5797), .B(n5796), .ZN(n5899) );
  NAND2_X1 U6956 ( .A1(n5899), .A2(n6429), .ZN(n5803) );
  INV_X1 U6957 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5798) );
  NOR2_X1 U6958 ( .A1(n6495), .A2(n5798), .ZN(n5893) );
  NOR2_X1 U6959 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  AOI211_X1 U6960 ( .C1(n6387), .C2(n6131), .A(n5893), .B(n5801), .ZN(n5802)
         );
  OAI211_X1 U6961 ( .C1(n6696), .C2(n6129), .A(n5803), .B(n5802), .ZN(U2970)
         );
  NAND2_X1 U6962 ( .A1(n5805), .A2(n5804), .ZN(n5812) );
  NAND2_X1 U6963 ( .A1(n5807), .A2(n5806), .ZN(n5809) );
  NAND2_X1 U6964 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  OAI21_X1 U6965 ( .B1(n5812), .B2(n5811), .A(n5810), .ZN(n5813) );
  INV_X1 U6966 ( .A(n5813), .ZN(n5911) );
  NAND2_X1 U6967 ( .A1(n6483), .A2(REIP_REG_15__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U6968 ( .A1(n6425), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5814)
         );
  OAI211_X1 U6969 ( .C1(n6434), .C2(n5815), .A(n5905), .B(n5814), .ZN(n5816)
         );
  AOI21_X1 U6970 ( .B1(n5817), .B2(n3085), .A(n5816), .ZN(n5818) );
  OAI21_X1 U6971 ( .B1(n5911), .B2(n6410), .A(n5818), .ZN(U2971) );
  NOR2_X1 U6972 ( .A1(n5819), .A2(n5821), .ZN(n5825) );
  AOI21_X1 U6973 ( .B1(n5822), .B2(n5821), .A(n5820), .ZN(n5823) );
  OAI21_X1 U6974 ( .B1(n5951), .B2(n6497), .A(n5823), .ZN(n5824) );
  AOI211_X1 U6975 ( .C1(n5826), .C2(n6503), .A(n5825), .B(n5824), .ZN(n5827)
         );
  INV_X1 U6976 ( .A(n5827), .ZN(U2991) );
  NOR2_X1 U6977 ( .A1(n5845), .A2(n5828), .ZN(n5840) );
  OAI211_X1 U6978 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5840), .B(n5829), .ZN(n5830) );
  OAI211_X1 U6979 ( .C1(n5958), .C2(n6497), .A(n5831), .B(n5830), .ZN(n5832)
         );
  AOI21_X1 U6980 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5833), .A(n5832), 
        .ZN(n5834) );
  OAI21_X1 U6981 ( .B1(n5835), .B2(n6476), .A(n5834), .ZN(U2992) );
  NAND2_X1 U6982 ( .A1(n5836), .A2(n6503), .ZN(n5842) );
  NOR2_X1 U6983 ( .A1(n5837), .A2(n6497), .ZN(n5838) );
  AOI211_X1 U6984 ( .C1(n5840), .C2(n5843), .A(n5839), .B(n5838), .ZN(n5841)
         );
  OAI211_X1 U6985 ( .C1(n5844), .C2(n5843), .A(n5842), .B(n5841), .ZN(U2993)
         );
  NOR2_X1 U6986 ( .A1(n5845), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5846)
         );
  AOI211_X1 U6987 ( .C1(n5967), .C2(n6485), .A(n5847), .B(n5846), .ZN(n5850)
         );
  NAND2_X1 U6988 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5849) );
  OAI211_X1 U6989 ( .C1(n5851), .C2(n6476), .A(n5850), .B(n5849), .ZN(U2995)
         );
  NAND2_X1 U6990 ( .A1(n5852), .A2(n6503), .ZN(n5859) );
  INV_X1 U6991 ( .A(n5986), .ZN(n5857) );
  NOR3_X1 U6992 ( .A1(n5862), .A2(n3533), .A3(n5854), .ZN(n5855) );
  AOI211_X1 U6993 ( .C1(n5857), .C2(n6485), .A(n5856), .B(n5855), .ZN(n5858)
         );
  OAI211_X1 U6994 ( .C1(n5869), .C2(n5860), .A(n5859), .B(n5858), .ZN(U2996)
         );
  NAND2_X1 U6995 ( .A1(n5861), .A2(n6503), .ZN(n5867) );
  INV_X1 U6996 ( .A(n5996), .ZN(n5865) );
  NOR2_X1 U6997 ( .A1(n5862), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5863)
         );
  AOI211_X1 U6998 ( .C1(n5865), .C2(n6485), .A(n5864), .B(n5863), .ZN(n5866)
         );
  OAI211_X1 U6999 ( .C1(n5869), .C2(n5868), .A(n5867), .B(n5866), .ZN(U2997)
         );
  INV_X1 U7000 ( .A(n5870), .ZN(n5886) );
  NOR3_X1 U7001 ( .A1(n5886), .A2(n5872), .A3(n5871), .ZN(n5873) );
  AOI211_X1 U7002 ( .C1(n5875), .C2(n6485), .A(n5874), .B(n5873), .ZN(n5880)
         );
  INV_X1 U7003 ( .A(n5876), .ZN(n5878) );
  INV_X1 U7004 ( .A(n6061), .ZN(n5877) );
  OAI21_X1 U7005 ( .B1(n5878), .B2(n5921), .A(n5877), .ZN(n5888) );
  NAND2_X1 U7006 ( .A1(n5888), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5879) );
  OAI211_X1 U7007 ( .C1(n5881), .C2(n6476), .A(n5880), .B(n5879), .ZN(U2998)
         );
  XNOR2_X1 U7008 ( .A(n5883), .B(n5882), .ZN(n6015) );
  NAND2_X1 U7009 ( .A1(n6015), .A2(n6485), .ZN(n5885) );
  NAND2_X1 U7010 ( .A1(n6483), .A2(REIP_REG_19__SCAN_IN), .ZN(n5884) );
  OAI211_X1 U7011 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5886), .A(n5885), .B(n5884), .ZN(n5887) );
  AOI21_X1 U7012 ( .B1(n5888), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5887), 
        .ZN(n5889) );
  OAI21_X1 U7013 ( .B1(n5890), .B2(n6476), .A(n5889), .ZN(U2999) );
  INV_X1 U7014 ( .A(n5891), .ZN(n5902) );
  OAI211_X1 U7015 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6437), .B(n5902), .ZN(n5897) );
  INV_X1 U7016 ( .A(n5892), .ZN(n5896) );
  OAI21_X1 U7017 ( .B1(n5921), .B2(n5902), .A(n6442), .ZN(n5909) );
  NAND2_X1 U7018 ( .A1(n5909), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5895) );
  AOI21_X1 U7019 ( .B1(n6126), .B2(n6485), .A(n5893), .ZN(n5894) );
  OAI211_X1 U7020 ( .C1(n5897), .C2(n5896), .A(n5895), .B(n5894), .ZN(n5898)
         );
  AOI21_X1 U7021 ( .B1(n5899), .B2(n6503), .A(n5898), .ZN(n5900) );
  INV_X1 U7022 ( .A(n5900), .ZN(U3002) );
  INV_X1 U7023 ( .A(n5901), .ZN(n5907) );
  AND2_X1 U7024 ( .A1(n6437), .A2(n5902), .ZN(n5904) );
  NAND2_X1 U7025 ( .A1(n5904), .A2(n5903), .ZN(n5906) );
  OAI211_X1 U7026 ( .C1(n6497), .C2(n5907), .A(n5906), .B(n5905), .ZN(n5908)
         );
  AOI21_X1 U7027 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5909), .A(n5908), 
        .ZN(n5910) );
  OAI21_X1 U7028 ( .B1(n5911), .B2(n6476), .A(n5910), .ZN(U3003) );
  NAND2_X1 U7029 ( .A1(n5912), .A2(n6503), .ZN(n5925) );
  INV_X1 U7030 ( .A(n5913), .ZN(n5919) );
  OAI21_X1 U7031 ( .B1(n5915), .B2(n6500), .A(n5914), .ZN(n6487) );
  NAND2_X1 U7032 ( .A1(n5919), .A2(n6487), .ZN(n6460) );
  NOR2_X1 U7033 ( .A1(n5917), .A2(n6460), .ZN(n6445) );
  OAI211_X1 U7034 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6445), .B(n5916), .ZN(n5924) );
  AOI22_X1 U7035 ( .A1(n6485), .A2(n6181), .B1(n6483), .B2(
        REIP_REG_10__SCAN_IN), .ZN(n5923) );
  INV_X1 U7036 ( .A(n5917), .ZN(n6453) );
  AOI21_X1 U7037 ( .B1(n5919), .B2(n6491), .A(n5918), .ZN(n5920) );
  INV_X1 U7038 ( .A(n5920), .ZN(n6465) );
  OAI21_X1 U7039 ( .B1(n5921), .B2(n6453), .A(n6465), .ZN(n6443) );
  NAND2_X1 U7040 ( .A1(n6443), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5922) );
  NAND4_X1 U7041 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(U3008)
         );
  NAND2_X1 U7042 ( .A1(n6693), .A2(n5930), .ZN(n5929) );
  AOI22_X1 U7043 ( .A1(n6635), .A2(n6704), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n5931), .ZN(n5928) );
  NAND2_X1 U7044 ( .A1(n5932), .A2(n6618), .ZN(n5927) );
  NAND2_X1 U7045 ( .A1(n6692), .A2(n5933), .ZN(n5926) );
  NAND4_X1 U7046 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(U3068)
         );
  NAND2_X1 U7047 ( .A1(n6715), .A2(n5930), .ZN(n5937) );
  AOI22_X1 U7048 ( .A1(n6635), .A2(n6716), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n5931), .ZN(n5936) );
  NAND2_X1 U7049 ( .A1(n5932), .A2(n6626), .ZN(n5935) );
  NAND2_X1 U7050 ( .A1(n6714), .A2(n5933), .ZN(n5934) );
  NAND4_X1 U7051 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(U3070)
         );
  AND2_X1 U7052 ( .A1(n6330), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7053 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5939) );
  OAI22_X1 U7054 ( .A1(n5939), .A2(n6170), .B1(n5938), .B2(n6229), .ZN(n5940)
         );
  AOI21_X1 U7055 ( .B1(EBX_REG_29__SCAN_IN), .B2(n6235), .A(n5940), .ZN(n5943)
         );
  NAND2_X1 U7056 ( .A1(n5941), .A2(REIP_REG_29__SCAN_IN), .ZN(n5942) );
  OAI211_X1 U7057 ( .C1(n5944), .C2(REIP_REG_29__SCAN_IN), .A(n5943), .B(n5942), .ZN(n5945) );
  AOI21_X1 U7058 ( .B1(n6018), .B2(n6213), .A(n5945), .ZN(n5946) );
  OAI21_X1 U7059 ( .B1(n5947), .B2(n6219), .A(n5946), .ZN(U2798) );
  AOI22_X1 U7060 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6235), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6234), .ZN(n5948) );
  OAI21_X1 U7061 ( .B1(n5949), .B2(n6229), .A(n5948), .ZN(n5950) );
  AOI21_X1 U7062 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5962), .A(n5950), .ZN(n5954) );
  OAI22_X1 U7063 ( .A1(n6021), .A2(n6128), .B1(n5951), .B2(n6219), .ZN(n5952)
         );
  INV_X1 U7064 ( .A(n5952), .ZN(n5953) );
  OAI211_X1 U7065 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5955), .A(n5954), .B(n5953), .ZN(U2800) );
  AOI22_X1 U7066 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6235), .B1(n5956), .B2(n3092), .ZN(n5964) );
  OAI21_X1 U7067 ( .B1(n6875), .B2(n5957), .A(n6880), .ZN(n5961) );
  OAI22_X1 U7068 ( .A1(n5959), .A2(n6128), .B1(n5958), .B2(n6219), .ZN(n5960)
         );
  AOI21_X1 U7069 ( .B1(n5962), .B2(n5961), .A(n5960), .ZN(n5963) );
  OAI211_X1 U7070 ( .C1(n5965), .C2(n6170), .A(n5964), .B(n5963), .ZN(U2801)
         );
  OAI22_X1 U7071 ( .A1(n3995), .A2(n6170), .B1(n5966), .B2(n6229), .ZN(n5971)
         );
  INV_X1 U7072 ( .A(n5967), .ZN(n5968) );
  OAI22_X1 U7073 ( .A1(n5969), .A2(n6128), .B1(n5968), .B2(n6219), .ZN(n5970)
         );
  AOI211_X1 U7074 ( .C1(EBX_REG_23__SCAN_IN), .C2(n6235), .A(n5971), .B(n5970), 
        .ZN(n5972) );
  OAI221_X1 U7075 ( .B1(n5974), .B2(n6872), .C1(n5974), .C2(n5973), .A(n5972), 
        .ZN(U2804) );
  AND2_X1 U7076 ( .A1(n6159), .A2(n5975), .ZN(n6002) );
  NOR2_X1 U7077 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5976), .ZN(n5992) );
  OAI22_X1 U7078 ( .A1(n5978), .A2(n6170), .B1(n6229), .B2(n5977), .ZN(n5979)
         );
  AOI21_X1 U7079 ( .B1(n6235), .B2(EBX_REG_22__SCAN_IN), .A(n5979), .ZN(n5982)
         );
  NAND2_X1 U7080 ( .A1(n5980), .A2(n6867), .ZN(n5981) );
  OAI211_X1 U7081 ( .C1(n5983), .C2(n6128), .A(n5982), .B(n5981), .ZN(n5984)
         );
  OAI21_X1 U7082 ( .B1(n5986), .B2(n6219), .A(n5985), .ZN(U2805) );
  NAND2_X1 U7083 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6002), .ZN(n5990) );
  AOI22_X1 U7084 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6235), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6234), .ZN(n5989) );
  NAND2_X1 U7085 ( .A1(n6233), .A2(n5987), .ZN(n5988) );
  NAND3_X1 U7086 ( .A1(n5990), .A2(n5989), .A3(n5988), .ZN(n5991) );
  NOR2_X1 U7087 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  OAI21_X1 U7088 ( .B1(n6032), .B2(n6128), .A(n5993), .ZN(n5994) );
  INV_X1 U7089 ( .A(n5994), .ZN(n5995) );
  OAI21_X1 U7090 ( .B1(n5996), .B2(n6219), .A(n5995), .ZN(U2806) );
  AOI22_X1 U7091 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6234), .B1(n5997), 
        .B2(n6233), .ZN(n6004) );
  OAI22_X1 U7092 ( .A1(n5999), .A2(n6128), .B1(n5998), .B2(n6219), .ZN(n6000)
         );
  AOI221_X1 U7093 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6002), .C1(n6001), .C2(
        n6002), .A(n6000), .ZN(n6003) );
  OAI211_X1 U7094 ( .C1(n3701), .C2(n6203), .A(n6004), .B(n6003), .ZN(U2807)
         );
  OAI21_X1 U7095 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n6005), .ZN(n6013) );
  NOR2_X1 U7096 ( .A1(n6007), .A2(n6006), .ZN(n6117) );
  AOI22_X1 U7097 ( .A1(n6008), .A2(n3092), .B1(REIP_REG_19__SCAN_IN), .B2(
        n6117), .ZN(n6009) );
  OAI21_X1 U7098 ( .B1(n6017), .B2(n6203), .A(n6009), .ZN(n6010) );
  AOI211_X1 U7099 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6209), 
        .B(n6010), .ZN(n6012) );
  AOI22_X1 U7100 ( .A1(n6036), .A2(n6213), .B1(n6240), .B2(n6015), .ZN(n6011)
         );
  OAI211_X1 U7101 ( .C1(n6112), .C2(n6013), .A(n6012), .B(n6011), .ZN(U2808)
         );
  INV_X1 U7102 ( .A(n6014), .ZN(n6258) );
  AOI22_X1 U7103 ( .A1(n6036), .A2(n6258), .B1(n6257), .B2(n6015), .ZN(n6016)
         );
  OAI21_X1 U7104 ( .B1(n6261), .B2(n6017), .A(n6016), .ZN(U2840) );
  AOI22_X1 U7105 ( .A1(n6018), .A2(n6272), .B1(n6265), .B2(DATAI_29_), .ZN(
        n6020) );
  AOI22_X1 U7106 ( .A1(n6268), .A2(DATAI_13_), .B1(n6267), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7107 ( .A1(n6020), .A2(n6019), .ZN(U2862) );
  INV_X1 U7108 ( .A(n6021), .ZN(n6022) );
  AOI22_X1 U7109 ( .A1(n6022), .A2(n6272), .B1(n6265), .B2(DATAI_27_), .ZN(
        n6024) );
  AOI22_X1 U7110 ( .A1(n6268), .A2(DATAI_11_), .B1(n6267), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7111 ( .A1(n6024), .A2(n6023), .ZN(U2864) );
  INV_X1 U7112 ( .A(n6025), .ZN(n6026) );
  AOI22_X1 U7113 ( .A1(n6026), .A2(n6272), .B1(n6265), .B2(DATAI_25_), .ZN(
        n6028) );
  AOI22_X1 U7114 ( .A1(n6268), .A2(DATAI_9_), .B1(n6267), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7115 ( .A1(n6028), .A2(n6027), .ZN(U2866) );
  AOI22_X1 U7116 ( .A1(n6029), .A2(n6272), .B1(n6265), .B2(DATAI_23_), .ZN(
        n6031) );
  AOI22_X1 U7117 ( .A1(n6268), .A2(DATAI_7_), .B1(n6267), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7118 ( .A1(n6031), .A2(n6030), .ZN(U2868) );
  INV_X1 U7119 ( .A(n6032), .ZN(n6033) );
  AOI22_X1 U7120 ( .A1(n6033), .A2(n6272), .B1(n6265), .B2(DATAI_21_), .ZN(
        n6035) );
  AOI22_X1 U7121 ( .A1(n6268), .A2(DATAI_5_), .B1(n6267), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7122 ( .A1(n6035), .A2(n6034), .ZN(U2870) );
  AOI22_X1 U7123 ( .A1(n6036), .A2(n6272), .B1(n6265), .B2(DATAI_19_), .ZN(
        n6038) );
  AOI22_X1 U7124 ( .A1(n6268), .A2(DATAI_3_), .B1(n6267), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7125 ( .A1(n6038), .A2(n6037), .ZN(U2872) );
  AOI22_X1 U7126 ( .A1(n6483), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6425), .ZN(n6048) );
  INV_X1 U7127 ( .A(n6039), .ZN(n6040) );
  AOI21_X1 U7128 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6045) );
  INV_X1 U7129 ( .A(n6043), .ZN(n6044) );
  OAI21_X1 U7130 ( .B1(n6046), .B2(n6045), .A(n6044), .ZN(n6057) );
  AOI22_X1 U7131 ( .A1(n6057), .A2(n6429), .B1(n3085), .B2(n6266), .ZN(n6047)
         );
  OAI211_X1 U7132 ( .C1(n6434), .C2(n6113), .A(n6048), .B(n6047), .ZN(U2969)
         );
  INV_X1 U7133 ( .A(n6049), .ZN(n6109) );
  AOI22_X1 U7134 ( .A1(n6050), .A2(n6503), .B1(n6485), .B2(n6109), .ZN(n6056)
         );
  NAND2_X1 U7135 ( .A1(n6483), .A2(REIP_REG_18__SCAN_IN), .ZN(n6055) );
  INV_X1 U7136 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6059) );
  OAI221_X1 U7137 ( .B1(n6061), .B2(n6051), .C1(n6061), .C2(n6059), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6054) );
  INV_X1 U7138 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6052) );
  NAND3_X1 U7139 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6060), .A3(n6052), .ZN(n6053) );
  NAND4_X1 U7140 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(U3000)
         );
  AOI22_X1 U7141 ( .A1(n6057), .A2(n6503), .B1(n6485), .B2(n6116), .ZN(n6063)
         );
  NOR2_X1 U7142 ( .A1(n6495), .A2(n6862), .ZN(n6058) );
  AOI221_X1 U7143 ( .B1(n6061), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n6060), .C2(n6059), .A(n6058), .ZN(n6062) );
  NAND2_X1 U7144 ( .A1(n6063), .A2(n6062), .ZN(U3001) );
  AOI21_X1 U7145 ( .B1(n6066), .B2(n6065), .A(n6064), .ZN(n6073) );
  AND3_X1 U7146 ( .A1(n6072), .A2(n6437), .A3(n6067), .ZN(n6070) );
  OAI22_X1 U7147 ( .A1(n6068), .A2(n6476), .B1(n6497), .B2(n6136), .ZN(n6069)
         );
  AOI211_X1 U7148 ( .C1(REIP_REG_14__SCAN_IN), .C2(n6483), .A(n6070), .B(n6069), .ZN(n6071) );
  OAI21_X1 U7149 ( .B1(n6073), .B2(n6072), .A(n6071), .ZN(U3004) );
  INV_X1 U7150 ( .A(n6074), .ZN(n6077) );
  NAND4_X1 U7151 ( .A1(n6077), .A2(n6906), .A3(n6076), .A4(n6075), .ZN(n6078)
         );
  OAI21_X1 U7152 ( .B1(n6916), .B2(n3812), .A(n6078), .ZN(U3455) );
  INV_X1 U7153 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6079) );
  AOI21_X1 U7154 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6079), .A(n6080), .ZN(n6087) );
  NAND2_X1 U7155 ( .A1(n6080), .A2(STATE_REG_1__SCAN_IN), .ZN(n6931) );
  INV_X1 U7156 ( .A(n6931), .ZN(n6945) );
  AOI21_X1 U7157 ( .B1(n6087), .B2(n6081), .A(n6945), .ZN(U2789) );
  INV_X1 U7158 ( .A(n6082), .ZN(n6083) );
  INV_X1 U7159 ( .A(n6802), .ZN(n6800) );
  OAI21_X1 U7160 ( .B1(n6083), .B2(n6800), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6084) );
  OAI21_X1 U7161 ( .B1(n6085), .B2(n6809), .A(n6084), .ZN(U2790) );
  NOR2_X1 U7162 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6088) );
  OAI21_X1 U7163 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6088), .A(n6931), .ZN(n6086)
         );
  OAI21_X1 U7164 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6931), .A(n6086), .ZN(
        U2791) );
  NOR2_X1 U7165 ( .A1(n6945), .A2(n6087), .ZN(n6901) );
  OAI21_X1 U7166 ( .B1(BS16_N), .B2(n6088), .A(n6901), .ZN(n6899) );
  OAI21_X1 U7167 ( .B1(n6901), .B2(n6089), .A(n6899), .ZN(U2792) );
  OAI21_X1 U7168 ( .B1(n6091), .B2(n6090), .A(n6410), .ZN(U2793) );
  AOI211_X1 U7169 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_27__SCAN_IN), .B(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6092) );
  NAND4_X1 U7170 ( .A1(n6093), .A2(n6092), .A3(n6814), .A4(n6818), .ZN(n6101)
         );
  OR4_X1 U7171 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), 
        .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(
        n6100) );
  OR4_X1 U7172 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6099) );
  NOR4_X1 U7173 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6097) );
  NOR4_X1 U7174 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6096) );
  NOR4_X1 U7175 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n6095) );
  NOR4_X1 U7176 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6094) );
  NAND4_X1 U7177 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n6098)
         );
  INV_X1 U7178 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6894) );
  INV_X1 U7179 ( .A(n6928), .ZN(n6923) );
  NOR2_X1 U7180 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6923), .ZN(n6920) );
  INV_X1 U7181 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6925) );
  INV_X1 U7182 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6900) );
  NAND3_X1 U7183 ( .A1(n6920), .A2(n6925), .A3(n6900), .ZN(n6102) );
  OAI221_X1 U7184 ( .B1(n6928), .B2(n6894), .C1(n6923), .C2(n6921), .A(n6102), 
        .ZN(U2794) );
  INV_X1 U7185 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6103) );
  NAND3_X1 U7186 ( .A1(n6928), .A2(n6921), .A3(n6900), .ZN(n6926) );
  OAI211_X1 U7187 ( .C1(n6928), .C2(n6103), .A(n6102), .B(n6926), .ZN(U2795)
         );
  AOI22_X1 U7188 ( .A1(n6104), .A2(n3092), .B1(REIP_REG_18__SCAN_IN), .B2(
        n6117), .ZN(n6105) );
  OAI21_X1 U7189 ( .B1(n6106), .B2(n6203), .A(n6105), .ZN(n6107) );
  AOI211_X1 U7190 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6209), 
        .B(n6107), .ZN(n6111) );
  INV_X1 U7191 ( .A(n6108), .ZN(n6262) );
  AOI22_X1 U7192 ( .A1(n6262), .A2(n6213), .B1(n6240), .B2(n6109), .ZN(n6110)
         );
  OAI211_X1 U7193 ( .C1(REIP_REG_18__SCAN_IN), .C2(n6112), .A(n6111), .B(n6110), .ZN(U2809) );
  OAI22_X1 U7194 ( .A1(n6114), .A2(n6170), .B1(n6113), .B2(n6229), .ZN(n6115)
         );
  AOI211_X1 U7195 ( .C1(n6235), .C2(EBX_REG_17__SCAN_IN), .A(n6209), .B(n6115), 
        .ZN(n6121) );
  AOI22_X1 U7196 ( .A1(n6266), .A2(n6213), .B1(n6240), .B2(n6116), .ZN(n6120)
         );
  OAI21_X1 U7197 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6118), .A(n6117), .ZN(n6119) );
  NAND3_X1 U7198 ( .A1(n6121), .A2(n6120), .A3(n6119), .ZN(U2810) );
  OAI21_X1 U7199 ( .B1(REIP_REG_15__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .A(
        n6122), .ZN(n6123) );
  OAI22_X1 U7200 ( .A1(n5798), .A2(n6144), .B1(n6124), .B2(n6123), .ZN(n6125)
         );
  AOI211_X1 U7201 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6209), 
        .B(n6125), .ZN(n6133) );
  INV_X1 U7202 ( .A(n6126), .ZN(n6127) );
  OAI22_X1 U7203 ( .A1(n6129), .A2(n6128), .B1(n6219), .B2(n6127), .ZN(n6130)
         );
  AOI21_X1 U7204 ( .B1(n6131), .B2(n3092), .A(n6130), .ZN(n6132) );
  OAI211_X1 U7205 ( .C1(n6134), .C2(n6203), .A(n6133), .B(n6132), .ZN(U2811)
         );
  NOR2_X1 U7206 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6135), .ZN(n6145) );
  INV_X1 U7207 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6137) );
  OAI22_X1 U7208 ( .A1(n6137), .A2(n6170), .B1(n6219), .B2(n6136), .ZN(n6138)
         );
  AOI211_X1 U7209 ( .C1(n6235), .C2(EBX_REG_14__SCAN_IN), .A(n6209), .B(n6138), 
        .ZN(n6143) );
  INV_X1 U7210 ( .A(n6139), .ZN(n6140) );
  AOI22_X1 U7211 ( .A1(n6141), .A2(n6213), .B1(n6140), .B2(n3092), .ZN(n6142)
         );
  OAI211_X1 U7212 ( .C1(n6145), .C2(n6144), .A(n6143), .B(n6142), .ZN(U2813)
         );
  INV_X1 U7213 ( .A(n6160), .ZN(n6146) );
  NAND3_X1 U7214 ( .A1(n6147), .A2(REIP_REG_12__SCAN_IN), .A3(n6146), .ZN(
        n6148) );
  NAND2_X1 U7215 ( .A1(n6159), .A2(n6148), .ZN(n6156) );
  AOI22_X1 U7216 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6235), .B1(n6240), .B2(n6248), .ZN(n6149) );
  OAI21_X1 U7217 ( .B1(REIP_REG_13__SCAN_IN), .B2(n6150), .A(n6149), .ZN(n6151) );
  AOI211_X1 U7218 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6209), 
        .B(n6151), .ZN(n6155) );
  INV_X1 U7219 ( .A(n6152), .ZN(n6153) );
  AOI22_X1 U7220 ( .A1(n6273), .A2(n6213), .B1(n6153), .B2(n3092), .ZN(n6154)
         );
  OAI211_X1 U7221 ( .C1(n6156), .C2(n5385), .A(n6155), .B(n6154), .ZN(U2814)
         );
  NOR3_X1 U7222 ( .A1(n6183), .A2(n6160), .A3(REIP_REG_12__SCAN_IN), .ZN(n6165) );
  INV_X1 U7223 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6158) );
  OAI22_X1 U7224 ( .A1(n6158), .A2(n6170), .B1(n6219), .B2(n6157), .ZN(n6164)
         );
  OAI21_X1 U7225 ( .B1(n6161), .B2(n6160), .A(n6159), .ZN(n6179) );
  OAI22_X1 U7226 ( .A1(n6162), .A2(n6203), .B1(n6855), .B2(n6179), .ZN(n6163)
         );
  NOR4_X1 U7227 ( .A1(n6209), .A2(n6165), .A3(n6164), .A4(n6163), .ZN(n6168)
         );
  INV_X1 U7228 ( .A(n6166), .ZN(n6389) );
  AOI22_X1 U7229 ( .A1(n6389), .A2(n6213), .B1(n6388), .B2(n6233), .ZN(n6167)
         );
  NAND2_X1 U7230 ( .A1(n6168), .A2(n6167), .ZN(U2815) );
  AOI21_X1 U7231 ( .B1(n6946), .B2(n6169), .A(REIP_REG_11__SCAN_IN), .ZN(n6180) );
  OAI22_X1 U7232 ( .A1(n6172), .A2(n6203), .B1(n6171), .B2(n6170), .ZN(n6173)
         );
  AOI211_X1 U7233 ( .C1(n6240), .C2(n6436), .A(n6209), .B(n6173), .ZN(n6178)
         );
  INV_X1 U7234 ( .A(n6174), .ZN(n6175) );
  AOI22_X1 U7235 ( .A1(n6176), .A2(n6213), .B1(n6175), .B2(n6233), .ZN(n6177)
         );
  OAI211_X1 U7236 ( .C1(n6180), .C2(n6179), .A(n6178), .B(n6177), .ZN(U2816)
         );
  AOI22_X1 U7237 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6235), .B1(n6240), .B2(n6181), .ZN(n6192) );
  NOR3_X1 U7238 ( .A1(n6183), .A2(REIP_REG_10__SCAN_IN), .A3(n6182), .ZN(n6184) );
  AOI211_X1 U7239 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6209), 
        .B(n6184), .ZN(n6191) );
  INV_X1 U7240 ( .A(n6185), .ZN(n6187) );
  AOI22_X1 U7241 ( .A1(n6187), .A2(n6213), .B1(n3092), .B2(n6186), .ZN(n6190)
         );
  INV_X1 U7242 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6850) );
  AND3_X1 U7243 ( .A1(n6946), .A2(n6850), .A3(n6188), .ZN(n6193) );
  OAI21_X1 U7244 ( .B1(n6194), .B2(n6193), .A(REIP_REG_10__SCAN_IN), .ZN(n6189) );
  NAND4_X1 U7245 ( .A1(n6192), .A2(n6191), .A3(n6190), .A4(n6189), .ZN(U2817)
         );
  INV_X1 U7246 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6252) );
  AOI21_X1 U7247 ( .B1(n6194), .B2(REIP_REG_9__SCAN_IN), .A(n6193), .ZN(n6202)
         );
  INV_X1 U7248 ( .A(n6195), .ZN(n6197) );
  INV_X1 U7249 ( .A(n5017), .ZN(n6196) );
  AOI21_X1 U7250 ( .B1(n6198), .B2(n6197), .A(n6196), .ZN(n6444) );
  AOI22_X1 U7251 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6234), .B1(n6240), 
        .B2(n6444), .ZN(n6199) );
  OAI211_X1 U7252 ( .C1(n6229), .C2(n6400), .A(n6199), .B(n6216), .ZN(n6200)
         );
  AOI21_X1 U7253 ( .B1(n6213), .B2(n6397), .A(n6200), .ZN(n6201) );
  OAI211_X1 U7254 ( .C1(n6252), .C2(n6203), .A(n6202), .B(n6201), .ZN(U2818)
         );
  AOI21_X1 U7255 ( .B1(n4805), .B2(n6205), .A(n6204), .ZN(n6459) );
  AOI22_X1 U7256 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6235), .B1(n6240), .B2(n6459), 
        .ZN(n6206) );
  OAI21_X1 U7257 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6207), .A(n6206), .ZN(n6208)
         );
  AOI211_X1 U7258 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6209), 
        .B(n6208), .ZN(n6215) );
  INV_X1 U7259 ( .A(n6210), .ZN(n6226) );
  NAND2_X1 U7260 ( .A1(n6226), .A2(n6211), .ZN(n6212) );
  AOI22_X1 U7261 ( .A1(n6405), .A2(n6213), .B1(REIP_REG_7__SCAN_IN), .B2(n6212), .ZN(n6214) );
  OAI211_X1 U7262 ( .C1(n6408), .C2(n6229), .A(n6215), .B(n6214), .ZN(U2820)
         );
  INV_X1 U7263 ( .A(n6409), .ZN(n6222) );
  INV_X1 U7264 ( .A(n6243), .ZN(n6221) );
  AOI22_X1 U7265 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6235), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6234), .ZN(n6217) );
  OAI211_X1 U7266 ( .C1(n6219), .C2(n6218), .A(n6217), .B(n6216), .ZN(n6220)
         );
  AOI21_X1 U7267 ( .B1(n6222), .B2(n6221), .A(n6220), .ZN(n6228) );
  AOI21_X1 U7268 ( .B1(n6946), .B2(n6223), .A(REIP_REG_5__SCAN_IN), .ZN(n6225)
         );
  OR2_X1 U7269 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  OAI211_X1 U7270 ( .C1(n6229), .C2(n6415), .A(n6228), .B(n6227), .ZN(U2822)
         );
  INV_X1 U7271 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6839) );
  OR2_X1 U7272 ( .A1(n6231), .A2(n6230), .ZN(n6246) );
  INV_X1 U7273 ( .A(n6424), .ZN(n6232) );
  AOI22_X1 U7274 ( .A1(n6234), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n3092), 
        .B2(n6232), .ZN(n6239) );
  NAND2_X1 U7275 ( .A1(n6235), .A2(EBX_REG_3__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7276 ( .A1(n6236), .A2(n6553), .ZN(n6237) );
  AND3_X1 U7277 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n6242) );
  NAND2_X1 U7278 ( .A1(n6240), .A2(n6484), .ZN(n6241) );
  OAI211_X1 U7279 ( .C1(n6243), .C2(n6420), .A(n6242), .B(n6241), .ZN(n6244)
         );
  INV_X1 U7280 ( .A(n6244), .ZN(n6245) );
  OAI221_X1 U7281 ( .B1(n6247), .B2(n6839), .C1(n6247), .C2(n6246), .A(n6245), 
        .ZN(U2824) );
  AOI22_X1 U7282 ( .A1(n6273), .A2(n6258), .B1(n6257), .B2(n6248), .ZN(n6249)
         );
  OAI21_X1 U7283 ( .B1(n6261), .B2(n6250), .A(n6249), .ZN(U2846) );
  AOI22_X1 U7284 ( .A1(n6397), .A2(n6258), .B1(n6257), .B2(n6444), .ZN(n6251)
         );
  OAI21_X1 U7285 ( .B1(n6261), .B2(n6252), .A(n6251), .ZN(U2850) );
  AOI22_X1 U7286 ( .A1(n6405), .A2(n6258), .B1(n6257), .B2(n6459), .ZN(n6253)
         );
  OAI21_X1 U7287 ( .B1(n6261), .B2(n6254), .A(n6253), .ZN(U2852) );
  INV_X1 U7288 ( .A(n6255), .ZN(n6430) );
  AOI22_X1 U7289 ( .A1(n6430), .A2(n6258), .B1(n6257), .B2(n6256), .ZN(n6259)
         );
  OAI21_X1 U7290 ( .B1(n6261), .B2(n6260), .A(n6259), .ZN(U2857) );
  AOI22_X1 U7291 ( .A1(n6262), .A2(n6272), .B1(n6265), .B2(DATAI_18_), .ZN(
        n6264) );
  AOI22_X1 U7292 ( .A1(n6268), .A2(DATAI_2_), .B1(n6267), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7293 ( .A1(n6264), .A2(n6263), .ZN(U2873) );
  AOI22_X1 U7294 ( .A1(n6266), .A2(n6272), .B1(n6265), .B2(DATAI_17_), .ZN(
        n6270) );
  AOI22_X1 U7295 ( .A1(n6268), .A2(DATAI_1_), .B1(n6267), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7296 ( .A1(n6270), .A2(n6269), .ZN(U2874) );
  INV_X1 U7297 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6304) );
  AOI22_X1 U7298 ( .A1(n6273), .A2(n6272), .B1(n6271), .B2(DATAI_13_), .ZN(
        n6274) );
  OAI21_X1 U7299 ( .B1(n6304), .B2(n6276), .A(n6274), .ZN(U2878) );
  INV_X1 U7300 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6333) );
  OAI222_X1 U7301 ( .A1(n6278), .A2(n6277), .B1(n6276), .B2(n6333), .C1(n6275), 
        .C2(n6350), .ZN(U2891) );
  AOI22_X1 U7302 ( .A1(n6298), .A2(EAX_REG_30__SCAN_IN), .B1(n6932), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6280) );
  OAI21_X1 U7303 ( .B1(n6281), .B2(n6327), .A(n6280), .ZN(U2893) );
  AOI22_X1 U7304 ( .A1(n6298), .A2(EAX_REG_29__SCAN_IN), .B1(n6932), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7305 ( .B1(n6283), .B2(n6327), .A(n6282), .ZN(U2894) );
  AOI22_X1 U7306 ( .A1(n6298), .A2(EAX_REG_28__SCAN_IN), .B1(n6932), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7307 ( .B1(n6285), .B2(n6327), .A(n6284), .ZN(U2895) );
  AOI22_X1 U7308 ( .A1(n6330), .A2(DATAO_REG_27__SCAN_IN), .B1(n6298), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7309 ( .B1(n6287), .B2(n6328), .A(n6286), .ZN(U2896) );
  AOI22_X1 U7310 ( .A1(n6330), .A2(DATAO_REG_26__SCAN_IN), .B1(n6298), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6288) );
  OAI21_X1 U7311 ( .B1(n6289), .B2(n6328), .A(n6288), .ZN(U2897) );
  INV_X1 U7312 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6291) );
  AOI22_X1 U7313 ( .A1(n6330), .A2(DATAO_REG_23__SCAN_IN), .B1(n6298), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6290) );
  OAI21_X1 U7314 ( .B1(n6291), .B2(n6328), .A(n6290), .ZN(U2900) );
  AOI22_X1 U7315 ( .A1(n6330), .A2(DATAO_REG_22__SCAN_IN), .B1(n6298), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6292) );
  OAI21_X1 U7316 ( .B1(n6293), .B2(n6328), .A(n6292), .ZN(U2901) );
  AOI22_X1 U7317 ( .A1(n6330), .A2(DATAO_REG_20__SCAN_IN), .B1(n6298), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6294) );
  OAI21_X1 U7318 ( .B1(n6295), .B2(n6328), .A(n6294), .ZN(U2903) );
  AOI22_X1 U7319 ( .A1(n6330), .A2(DATAO_REG_18__SCAN_IN), .B1(n6298), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U7320 ( .B1(n6297), .B2(n6328), .A(n6296), .ZN(U2905) );
  AOI22_X1 U7321 ( .A1(n6298), .A2(EAX_REG_16__SCAN_IN), .B1(n6932), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n6299) );
  OAI21_X1 U7322 ( .B1(n6300), .B2(n6327), .A(n6299), .ZN(U2907) );
  INV_X1 U7323 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6386) );
  AOI22_X1 U7324 ( .A1(n6932), .A2(LWORD_REG_15__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U7325 ( .B1(n6386), .B2(n6332), .A(n6301), .ZN(U2908) );
  AOI22_X1 U7326 ( .A1(n6932), .A2(LWORD_REG_14__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6302) );
  OAI21_X1 U7327 ( .B1(n6303), .B2(n6332), .A(n6302), .ZN(U2909) );
  INV_X1 U7328 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6306) );
  OAI222_X1 U7329 ( .A1(n6306), .A2(n6328), .B1(n6327), .B2(n6305), .C1(n6304), 
        .C2(n6332), .ZN(U2910) );
  AOI22_X1 U7330 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6323), .B1(n6932), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6307) );
  OAI21_X1 U7331 ( .B1(n6308), .B2(n6327), .A(n6307), .ZN(U2911) );
  AOI22_X1 U7332 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6323), .B1(n6932), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6309) );
  OAI21_X1 U7333 ( .B1(n6310), .B2(n6327), .A(n6309), .ZN(U2912) );
  INV_X1 U7334 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6370) );
  AOI22_X1 U7335 ( .A1(n6932), .A2(LWORD_REG_10__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6311) );
  OAI21_X1 U7336 ( .B1(n6370), .B2(n6332), .A(n6311), .ZN(U2913) );
  OAI222_X1 U7337 ( .A1(n6332), .A2(n5054), .B1(n6327), .B2(n6313), .C1(n6328), 
        .C2(n6312), .ZN(U2914) );
  INV_X1 U7338 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6367) );
  AOI22_X1 U7339 ( .A1(n6932), .A2(LWORD_REG_8__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U7340 ( .B1(n6367), .B2(n6332), .A(n6314), .ZN(U2915) );
  AOI22_X1 U7341 ( .A1(n6932), .A2(LWORD_REG_7__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6315) );
  OAI21_X1 U7342 ( .B1(n3844), .B2(n6332), .A(n6315), .ZN(U2916) );
  AOI22_X1 U7343 ( .A1(n6932), .A2(LWORD_REG_6__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6316) );
  OAI21_X1 U7344 ( .B1(n6317), .B2(n6332), .A(n6316), .ZN(U2917) );
  AOI22_X1 U7345 ( .A1(n6932), .A2(LWORD_REG_5__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U7346 ( .B1(n3832), .B2(n6332), .A(n6318), .ZN(U2918) );
  AOI22_X1 U7347 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6323), .B1(n6330), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7348 ( .B1(n6320), .B2(n6328), .A(n6319), .ZN(U2919) );
  AOI22_X1 U7349 ( .A1(n6932), .A2(LWORD_REG_3__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6321) );
  OAI21_X1 U7350 ( .B1(n6322), .B2(n6332), .A(n6321), .ZN(U2920) );
  AOI222_X1 U7351 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6932), .B1(n6330), .B2(
        DATAO_REG_2__SCAN_IN), .C1(EAX_REG_2__SCAN_IN), .C2(n6323), .ZN(n6324)
         );
  INV_X1 U7352 ( .A(n6324), .ZN(U2921) );
  INV_X1 U7353 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6329) );
  OAI222_X1 U7354 ( .A1(n6329), .A2(n6328), .B1(n6327), .B2(n6326), .C1(n6325), 
        .C2(n6332), .ZN(U2922) );
  AOI22_X1 U7355 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6932), .B1(n6330), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6331) );
  OAI21_X1 U7356 ( .B1(n6333), .B2(n6332), .A(n6331), .ZN(U2923) );
  AOI22_X1 U7357 ( .A1(n6383), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6378), .ZN(n6335) );
  OAI21_X1 U7358 ( .B1(n6380), .B2(n6350), .A(n6335), .ZN(U2924) );
  AOI22_X1 U7359 ( .A1(n6383), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6378), .ZN(n6336) );
  OAI21_X1 U7360 ( .B1(n6380), .B2(n6352), .A(n6336), .ZN(U2925) );
  AOI22_X1 U7361 ( .A1(n6375), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6378), .ZN(n6337) );
  OAI21_X1 U7362 ( .B1(n6380), .B2(n6354), .A(n6337), .ZN(U2926) );
  AOI22_X1 U7363 ( .A1(n6375), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6378), .ZN(n6338) );
  OAI21_X1 U7364 ( .B1(n6380), .B2(n6356), .A(n6338), .ZN(U2927) );
  AOI22_X1 U7365 ( .A1(n6375), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6378), .ZN(n6339) );
  OAI21_X1 U7366 ( .B1(n6380), .B2(n6358), .A(n6339), .ZN(U2928) );
  AOI22_X1 U7367 ( .A1(n6375), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6378), .ZN(n6340) );
  OAI21_X1 U7368 ( .B1(n6380), .B2(n6360), .A(n6340), .ZN(U2929) );
  AOI22_X1 U7369 ( .A1(n6375), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6378), .ZN(n6341) );
  OAI21_X1 U7370 ( .B1(n6380), .B2(n6362), .A(n6341), .ZN(U2930) );
  AOI22_X1 U7371 ( .A1(n6383), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6378), .ZN(n6342) );
  OAI21_X1 U7372 ( .B1(n6380), .B2(n6364), .A(n6342), .ZN(U2931) );
  AOI21_X1 U7373 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6383), .A(n6343), .ZN(n6344) );
  OAI21_X1 U7374 ( .B1(n6345), .B2(n6385), .A(n6344), .ZN(U2933) );
  AOI22_X1 U7375 ( .A1(n6383), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6378), .ZN(n6346) );
  INV_X1 U7376 ( .A(n6380), .ZN(n6382) );
  NAND2_X1 U7377 ( .A1(n6382), .A2(DATAI_12_), .ZN(n6373) );
  NAND2_X1 U7378 ( .A1(n6346), .A2(n6373), .ZN(U2936) );
  AOI22_X1 U7379 ( .A1(n6383), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6378), .ZN(n6347) );
  NAND2_X1 U7380 ( .A1(n6382), .A2(DATAI_13_), .ZN(n6376) );
  NAND2_X1 U7381 ( .A1(n6347), .A2(n6376), .ZN(U2937) );
  AOI22_X1 U7382 ( .A1(n6383), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6378), .ZN(n6348) );
  OAI21_X1 U7383 ( .B1(n6381), .B2(n6380), .A(n6348), .ZN(U2938) );
  AOI22_X1 U7384 ( .A1(n6383), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6378), .ZN(n6349) );
  OAI21_X1 U7385 ( .B1(n6380), .B2(n6350), .A(n6349), .ZN(U2939) );
  AOI22_X1 U7386 ( .A1(n6383), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6378), .ZN(n6351) );
  OAI21_X1 U7387 ( .B1(n6380), .B2(n6352), .A(n6351), .ZN(U2940) );
  AOI22_X1 U7388 ( .A1(n6383), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6378), .ZN(n6353) );
  OAI21_X1 U7389 ( .B1(n6380), .B2(n6354), .A(n6353), .ZN(U2941) );
  AOI22_X1 U7390 ( .A1(n6383), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6378), .ZN(n6355) );
  OAI21_X1 U7391 ( .B1(n6380), .B2(n6356), .A(n6355), .ZN(U2942) );
  AOI22_X1 U7392 ( .A1(n6383), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6378), .ZN(n6357) );
  OAI21_X1 U7393 ( .B1(n6380), .B2(n6358), .A(n6357), .ZN(U2943) );
  AOI22_X1 U7394 ( .A1(n6383), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6378), .ZN(n6359) );
  OAI21_X1 U7395 ( .B1(n6380), .B2(n6360), .A(n6359), .ZN(U2944) );
  AOI22_X1 U7396 ( .A1(n6383), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6378), .ZN(n6361) );
  OAI21_X1 U7397 ( .B1(n6380), .B2(n6362), .A(n6361), .ZN(U2945) );
  AOI22_X1 U7398 ( .A1(n6383), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6378), .ZN(n6363) );
  OAI21_X1 U7399 ( .B1(n6380), .B2(n6364), .A(n6363), .ZN(U2946) );
  AOI21_X1 U7400 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6383), .A(n6365), .ZN(n6366) );
  OAI21_X1 U7401 ( .B1(n6367), .B2(n6385), .A(n6366), .ZN(U2947) );
  AOI21_X1 U7402 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6383), .A(n6368), .ZN(
        n6369) );
  OAI21_X1 U7403 ( .B1(n6370), .B2(n6385), .A(n6369), .ZN(U2949) );
  AOI22_X1 U7404 ( .A1(n6383), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6378), .ZN(n6372) );
  NAND2_X1 U7405 ( .A1(n6382), .A2(DATAI_11_), .ZN(n6371) );
  NAND2_X1 U7406 ( .A1(n6372), .A2(n6371), .ZN(U2950) );
  AOI22_X1 U7407 ( .A1(n6383), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6378), .ZN(n6374) );
  NAND2_X1 U7408 ( .A1(n6374), .A2(n6373), .ZN(U2951) );
  AOI22_X1 U7409 ( .A1(n6375), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6378), .ZN(n6377) );
  NAND2_X1 U7410 ( .A1(n6377), .A2(n6376), .ZN(U2952) );
  AOI22_X1 U7411 ( .A1(n6383), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6378), .ZN(n6379) );
  OAI21_X1 U7412 ( .B1(n6381), .B2(n6380), .A(n6379), .ZN(U2953) );
  AOI22_X1 U7413 ( .A1(n6383), .A2(LWORD_REG_15__SCAN_IN), .B1(n6382), .B2(
        DATAI_15_), .ZN(n6384) );
  OAI21_X1 U7414 ( .B1(n6386), .B2(n6385), .A(n6384), .ZN(U2954) );
  AOI22_X1 U7415 ( .A1(n6483), .A2(REIP_REG_12__SCAN_IN), .B1(n6425), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6391) );
  AOI22_X1 U7416 ( .A1(n6389), .A2(n3085), .B1(n6388), .B2(n6387), .ZN(n6390)
         );
  OAI211_X1 U7417 ( .C1(n6392), .C2(n6410), .A(n6391), .B(n6390), .ZN(U2974)
         );
  AOI22_X1 U7418 ( .A1(n6483), .A2(REIP_REG_9__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n6425), .ZN(n6399) );
  OAI21_X1 U7419 ( .B1(n6395), .B2(n6394), .A(n6393), .ZN(n6396) );
  INV_X1 U7420 ( .A(n6396), .ZN(n6446) );
  AOI22_X1 U7421 ( .A1(n6446), .A2(n6429), .B1(n3085), .B2(n6397), .ZN(n6398)
         );
  OAI211_X1 U7422 ( .C1(n6434), .C2(n6400), .A(n6399), .B(n6398), .ZN(U2977)
         );
  AOI22_X1 U7423 ( .A1(n6483), .A2(REIP_REG_7__SCAN_IN), .B1(n6425), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U7424 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(n6404) );
  INV_X1 U7425 ( .A(n6404), .ZN(n6462) );
  AOI22_X1 U7426 ( .A1(n6462), .A2(n6429), .B1(n3085), .B2(n6405), .ZN(n6406)
         );
  OAI211_X1 U7427 ( .C1(n6434), .C2(n6408), .A(n6407), .B(n6406), .ZN(U2979)
         );
  AOI22_X1 U7428 ( .A1(n6483), .A2(REIP_REG_5__SCAN_IN), .B1(n6425), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6414) );
  OAI22_X1 U7429 ( .A1(n6411), .A2(n6410), .B1(n6409), .B2(n6696), .ZN(n6412)
         );
  INV_X1 U7430 ( .A(n6412), .ZN(n6413) );
  OAI211_X1 U7431 ( .C1(n6434), .C2(n6415), .A(n6414), .B(n6413), .ZN(U2981)
         );
  AOI22_X1 U7432 ( .A1(n6483), .A2(REIP_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6425), .ZN(n6423) );
  INV_X1 U7433 ( .A(n6416), .ZN(n6417) );
  AOI21_X1 U7434 ( .B1(n6419), .B2(n6418), .A(n6417), .ZN(n6486) );
  INV_X1 U7435 ( .A(n6420), .ZN(n6421) );
  AOI22_X1 U7436 ( .A1(n6486), .A2(n6429), .B1(n3085), .B2(n6421), .ZN(n6422)
         );
  OAI211_X1 U7437 ( .C1(n6434), .C2(n6424), .A(n6423), .B(n6422), .ZN(U2983)
         );
  AOI22_X1 U7438 ( .A1(n6483), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6425), .ZN(n6432) );
  XNOR2_X1 U7439 ( .A(n6426), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6428)
         );
  XNOR2_X1 U7440 ( .A(n6428), .B(n6427), .ZN(n6504) );
  AOI22_X1 U7441 ( .A1(n6430), .A2(n3085), .B1(n6429), .B2(n6504), .ZN(n6431)
         );
  OAI211_X1 U7442 ( .C1(n6434), .C2(n6433), .A(n6432), .B(n6431), .ZN(U2984)
         );
  AOI21_X1 U7443 ( .B1(n6485), .B2(n6436), .A(n6435), .ZN(n6440) );
  AOI22_X1 U7444 ( .A1(n6438), .A2(n6503), .B1(n6441), .B2(n6437), .ZN(n6439)
         );
  OAI211_X1 U7445 ( .C1(n6442), .C2(n6441), .A(n6440), .B(n6439), .ZN(U3007)
         );
  INV_X1 U7446 ( .A(n6443), .ZN(n6450) );
  AOI22_X1 U7447 ( .A1(n6485), .A2(n6444), .B1(n6483), .B2(REIP_REG_9__SCAN_IN), .ZN(n6448) );
  AOI22_X1 U7448 ( .A1(n6446), .A2(n6503), .B1(n6445), .B2(n6449), .ZN(n6447)
         );
  OAI211_X1 U7449 ( .C1(n6450), .C2(n6449), .A(n6448), .B(n6447), .ZN(U3009)
         );
  INV_X1 U7450 ( .A(n6451), .ZN(n6456) );
  OAI22_X1 U7451 ( .A1(n6497), .A2(n6452), .B1(n6848), .B2(n6495), .ZN(n6455)
         );
  AOI211_X1 U7452 ( .C1(n6458), .C2(n6466), .A(n6453), .B(n6460), .ZN(n6454)
         );
  AOI211_X1 U7453 ( .C1(n6456), .C2(n6503), .A(n6455), .B(n6454), .ZN(n6457)
         );
  OAI21_X1 U7454 ( .B1(n6458), .B2(n6465), .A(n6457), .ZN(U3010) );
  AOI22_X1 U7455 ( .A1(n6485), .A2(n6459), .B1(n6483), .B2(REIP_REG_7__SCAN_IN), .ZN(n6464) );
  INV_X1 U7456 ( .A(n6460), .ZN(n6461) );
  AOI22_X1 U7457 ( .A1(n6462), .A2(n6503), .B1(n6461), .B2(n6466), .ZN(n6463)
         );
  OAI211_X1 U7458 ( .C1(n6466), .C2(n6465), .A(n6464), .B(n6463), .ZN(U3011)
         );
  NAND2_X1 U7459 ( .A1(n6467), .A2(n6487), .ZN(n6474) );
  OAI222_X1 U7460 ( .A1(n6469), .A2(n6497), .B1(n6495), .B2(n6844), .C1(n6476), 
        .C2(n6468), .ZN(n6470) );
  INV_X1 U7461 ( .A(n6470), .ZN(n6471) );
  OAI221_X1 U7462 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6474), .C1(n6473), .C2(n6472), .A(n6471), .ZN(U3012) );
  OAI222_X1 U7463 ( .A1(n6477), .A2(n6497), .B1(n6495), .B2(n6841), .C1(n6476), 
        .C2(n6475), .ZN(n6478) );
  INV_X1 U7464 ( .A(n6478), .ZN(n6481) );
  OAI211_X1 U7465 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6487), .B(n6479), .ZN(n6480) );
  OAI211_X1 U7466 ( .C1(n6491), .C2(n6482), .A(n6481), .B(n6480), .ZN(U3014)
         );
  INV_X1 U7467 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6490) );
  AOI22_X1 U7468 ( .A1(n6485), .A2(n6484), .B1(n6483), .B2(REIP_REG_3__SCAN_IN), .ZN(n6489) );
  AOI22_X1 U7469 ( .A1(n6487), .A2(n6490), .B1(n6503), .B2(n6486), .ZN(n6488)
         );
  OAI211_X1 U7470 ( .C1(n6491), .C2(n6490), .A(n6489), .B(n6488), .ZN(U3015)
         );
  AOI21_X1 U7471 ( .B1(n6494), .B2(n6493), .A(n6492), .ZN(n6499) );
  OAI22_X1 U7472 ( .A1(n6497), .A2(n6496), .B1(n6230), .B2(n6495), .ZN(n6498)
         );
  NOR2_X1 U7473 ( .A1(n6499), .A2(n6498), .ZN(n6506) );
  NOR3_X1 U7474 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6501), .A3(n6500), 
        .ZN(n6502) );
  AOI21_X1 U7475 ( .B1(n6504), .B2(n6503), .A(n6502), .ZN(n6505) );
  OAI211_X1 U7476 ( .C1(n6508), .C2(n6507), .A(n6506), .B(n6505), .ZN(U3016)
         );
  NOR2_X1 U7477 ( .A1(n6774), .A2(n6509), .ZN(U3019) );
  NOR2_X1 U7478 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6510), .ZN(n6545)
         );
  INV_X1 U7479 ( .A(n6511), .ZN(n6522) );
  NOR2_X2 U7480 ( .A1(n6694), .A2(n6551), .ZN(n6748) );
  OAI21_X1 U7481 ( .B1(n6748), .B2(n6546), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6513) );
  OAI211_X1 U7482 ( .C1(n6553), .C2(n6522), .A(n6513), .B(n6703), .ZN(n6514)
         );
  OAI21_X1 U7483 ( .B1(n6545), .B2(n6904), .A(n6514), .ZN(n6515) );
  NOR3_X2 U7484 ( .A1(n6517), .A2(n6516), .A3(n6515), .ZN(n6550) );
  INV_X1 U7485 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6525) );
  INV_X1 U7486 ( .A(n6555), .ZN(n6520) );
  INV_X1 U7487 ( .A(n6518), .ZN(n6519) );
  OAI22_X1 U7488 ( .A1(n6522), .A2(n6521), .B1(n6520), .B2(n6519), .ZN(n6544)
         );
  AOI22_X1 U7489 ( .A1(n6693), .A2(n6544), .B1(n6692), .B2(n6545), .ZN(n6524)
         );
  AOI22_X1 U7490 ( .A1(n6618), .A2(n6748), .B1(n6546), .B2(n6704), .ZN(n6523)
         );
  OAI211_X1 U7491 ( .C1(n6550), .C2(n6525), .A(n6524), .B(n6523), .ZN(U3020)
         );
  INV_X1 U7492 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7493 ( .A1(n6709), .A2(n6545), .B1(n6708), .B2(n6544), .ZN(n6527)
         );
  AOI22_X1 U7494 ( .A1(n6622), .A2(n6748), .B1(n6546), .B2(n6710), .ZN(n6526)
         );
  OAI211_X1 U7495 ( .C1(n6550), .C2(n6528), .A(n6527), .B(n6526), .ZN(U3021)
         );
  INV_X1 U7496 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7497 ( .A1(n6715), .A2(n6544), .B1(n6714), .B2(n6545), .ZN(n6530)
         );
  AOI22_X1 U7498 ( .A1(n6626), .A2(n6748), .B1(n6546), .B2(n6716), .ZN(n6529)
         );
  OAI211_X1 U7499 ( .C1(n6550), .C2(n6531), .A(n6530), .B(n6529), .ZN(U3022)
         );
  INV_X1 U7500 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6534) );
  AOI22_X1 U7501 ( .A1(n6721), .A2(n6545), .B1(n6720), .B2(n6544), .ZN(n6533)
         );
  AOI22_X1 U7502 ( .A1(n6630), .A2(n6748), .B1(n6546), .B2(n6722), .ZN(n6532)
         );
  OAI211_X1 U7503 ( .C1(n6550), .C2(n6534), .A(n6533), .B(n6532), .ZN(U3023)
         );
  INV_X1 U7504 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6537) );
  AOI22_X1 U7505 ( .A1(n6727), .A2(n6545), .B1(n6726), .B2(n6544), .ZN(n6536)
         );
  AOI22_X1 U7506 ( .A1(n6669), .A2(n6748), .B1(n6546), .B2(n6728), .ZN(n6535)
         );
  OAI211_X1 U7507 ( .C1(n6550), .C2(n6537), .A(n6536), .B(n6535), .ZN(U3024)
         );
  INV_X1 U7508 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6540) );
  AOI22_X1 U7509 ( .A1(n6733), .A2(n6545), .B1(n6732), .B2(n6544), .ZN(n6539)
         );
  AOI22_X1 U7510 ( .A1(n6636), .A2(n6748), .B1(n6546), .B2(n6734), .ZN(n6538)
         );
  OAI211_X1 U7511 ( .C1(n6550), .C2(n6540), .A(n6539), .B(n6538), .ZN(U3025)
         );
  INV_X1 U7512 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6543) );
  AOI22_X1 U7513 ( .A1(n6739), .A2(n6545), .B1(n6738), .B2(n6544), .ZN(n6542)
         );
  AOI22_X1 U7514 ( .A1(n6675), .A2(n6748), .B1(n6546), .B2(n6740), .ZN(n6541)
         );
  OAI211_X1 U7515 ( .C1(n6550), .C2(n6543), .A(n6542), .B(n6541), .ZN(U3026)
         );
  AOI22_X1 U7516 ( .A1(n6747), .A2(n6545), .B1(n6745), .B2(n6544), .ZN(n6548)
         );
  AOI22_X1 U7517 ( .A1(n6578), .A2(n6748), .B1(n6546), .B2(n6749), .ZN(n6547)
         );
  OAI211_X1 U7518 ( .C1(n6550), .C2(n6549), .A(n6548), .B(n6547), .ZN(U3027)
         );
  OR2_X1 U7519 ( .A1(n6553), .A2(n6552), .ZN(n6586) );
  NAND3_X1 U7520 ( .A1(n6555), .A2(n6554), .A3(n6777), .ZN(n6556) );
  OAI21_X1 U7521 ( .B1(n6586), .B2(n6934), .A(n6556), .ZN(n6575) );
  NAND3_X1 U7522 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6777), .A3(n6770), .ZN(n6590) );
  NOR2_X1 U7523 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6590), .ZN(n6576)
         );
  AOI22_X1 U7524 ( .A1(n6693), .A2(n6575), .B1(n6692), .B2(n6576), .ZN(n6561)
         );
  OAI21_X1 U7525 ( .B1(n6605), .B2(n6577), .A(n6695), .ZN(n6557) );
  AOI21_X1 U7526 ( .B1(n6557), .B2(n6586), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6559) );
  OAI21_X1 U7527 ( .B1(n6559), .B2(n6576), .A(n6558), .ZN(n6579) );
  AOI22_X1 U7528 ( .A1(n6579), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6618), 
        .B2(n6577), .ZN(n6560) );
  OAI211_X1 U7529 ( .C1(n6562), .C2(n6617), .A(n6561), .B(n6560), .ZN(U3036)
         );
  AOI22_X1 U7530 ( .A1(n6709), .A2(n6576), .B1(n6708), .B2(n6575), .ZN(n6564)
         );
  AOI22_X1 U7531 ( .A1(n6579), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6622), 
        .B2(n6577), .ZN(n6563) );
  OAI211_X1 U7532 ( .C1(n6617), .C2(n6597), .A(n6564), .B(n6563), .ZN(U3037)
         );
  AOI22_X1 U7533 ( .A1(n6715), .A2(n6575), .B1(n6714), .B2(n6576), .ZN(n6566)
         );
  AOI22_X1 U7534 ( .A1(n6579), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6626), 
        .B2(n6577), .ZN(n6565) );
  OAI211_X1 U7535 ( .C1(n6617), .C2(n6600), .A(n6566), .B(n6565), .ZN(U3038)
         );
  AOI22_X1 U7536 ( .A1(n6721), .A2(n6576), .B1(n6720), .B2(n6575), .ZN(n6568)
         );
  AOI22_X1 U7537 ( .A1(n6579), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6630), 
        .B2(n6577), .ZN(n6567) );
  OAI211_X1 U7538 ( .C1(n6617), .C2(n6634), .A(n6568), .B(n6567), .ZN(U3039)
         );
  AOI22_X1 U7539 ( .A1(n6727), .A2(n6576), .B1(n6726), .B2(n6575), .ZN(n6570)
         );
  AOI22_X1 U7540 ( .A1(n6579), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6669), 
        .B2(n6577), .ZN(n6569) );
  OAI211_X1 U7541 ( .C1(n6617), .C2(n6672), .A(n6570), .B(n6569), .ZN(U3040)
         );
  AOI22_X1 U7542 ( .A1(n6733), .A2(n6576), .B1(n6732), .B2(n6575), .ZN(n6572)
         );
  AOI22_X1 U7543 ( .A1(n6579), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6636), 
        .B2(n6577), .ZN(n6571) );
  OAI211_X1 U7544 ( .C1(n6617), .C2(n6640), .A(n6572), .B(n6571), .ZN(U3041)
         );
  AOI22_X1 U7545 ( .A1(n6739), .A2(n6576), .B1(n6738), .B2(n6575), .ZN(n6574)
         );
  AOI22_X1 U7546 ( .A1(n6579), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6675), 
        .B2(n6577), .ZN(n6573) );
  OAI211_X1 U7547 ( .C1(n6617), .C2(n6680), .A(n6574), .B(n6573), .ZN(U3042)
         );
  AOI22_X1 U7548 ( .A1(n6747), .A2(n6576), .B1(n6745), .B2(n6575), .ZN(n6581)
         );
  AOI22_X1 U7549 ( .A1(n6579), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6578), 
        .B2(n6577), .ZN(n6580) );
  OAI211_X1 U7550 ( .C1(n6617), .C2(n6582), .A(n6581), .B(n6580), .ZN(U3043)
         );
  NOR2_X1 U7551 ( .A1(n6650), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6611)
         );
  AOI22_X1 U7552 ( .A1(n6704), .A2(n6612), .B1(n6692), .B2(n6611), .ZN(n6594)
         );
  NAND3_X1 U7553 ( .A1(n6652), .A2(n6584), .A3(n6583), .ZN(n6585) );
  NAND2_X1 U7554 ( .A1(n6585), .A2(n6703), .ZN(n6592) );
  INV_X1 U7555 ( .A(n6586), .ZN(n6587) );
  AOI21_X1 U7556 ( .B1(n6587), .B2(n6653), .A(n6611), .ZN(n6591) );
  INV_X1 U7557 ( .A(n6591), .ZN(n6589) );
  AOI21_X1 U7558 ( .B1(n6934), .B2(n6590), .A(n6655), .ZN(n6588) );
  OAI21_X1 U7559 ( .B1(n6592), .B2(n6589), .A(n6588), .ZN(n6614) );
  OAI22_X1 U7560 ( .A1(n6592), .A2(n6591), .B1(n6590), .B2(n6937), .ZN(n6613)
         );
  AOI22_X1 U7561 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6614), .B1(n6693), 
        .B2(n6613), .ZN(n6593) );
  OAI211_X1 U7562 ( .C1(n6707), .C2(n6617), .A(n6594), .B(n6593), .ZN(U3044)
         );
  AOI22_X1 U7563 ( .A1(n6622), .A2(n6605), .B1(n6709), .B2(n6611), .ZN(n6596)
         );
  AOI22_X1 U7564 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6614), .B1(n6708), 
        .B2(n6613), .ZN(n6595) );
  OAI211_X1 U7565 ( .C1(n6597), .C2(n6608), .A(n6596), .B(n6595), .ZN(U3045)
         );
  AOI22_X1 U7566 ( .A1(n6626), .A2(n6605), .B1(n6714), .B2(n6611), .ZN(n6599)
         );
  AOI22_X1 U7567 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6614), .B1(n6715), 
        .B2(n6613), .ZN(n6598) );
  OAI211_X1 U7568 ( .C1(n6600), .C2(n6608), .A(n6599), .B(n6598), .ZN(U3046)
         );
  AOI22_X1 U7569 ( .A1(n6630), .A2(n6605), .B1(n6721), .B2(n6611), .ZN(n6602)
         );
  AOI22_X1 U7570 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6614), .B1(n6720), 
        .B2(n6613), .ZN(n6601) );
  OAI211_X1 U7571 ( .C1(n6634), .C2(n6608), .A(n6602), .B(n6601), .ZN(U3047)
         );
  AOI22_X1 U7572 ( .A1(n6669), .A2(n6605), .B1(n6727), .B2(n6611), .ZN(n6604)
         );
  AOI22_X1 U7573 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6614), .B1(n6726), 
        .B2(n6613), .ZN(n6603) );
  OAI211_X1 U7574 ( .C1(n6672), .C2(n6608), .A(n6604), .B(n6603), .ZN(U3048)
         );
  AOI22_X1 U7575 ( .A1(n6636), .A2(n6605), .B1(n6733), .B2(n6611), .ZN(n6607)
         );
  AOI22_X1 U7576 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6614), .B1(n6732), 
        .B2(n6613), .ZN(n6606) );
  OAI211_X1 U7577 ( .C1(n6640), .C2(n6608), .A(n6607), .B(n6606), .ZN(U3049)
         );
  AOI22_X1 U7578 ( .A1(n6740), .A2(n6612), .B1(n6739), .B2(n6611), .ZN(n6610)
         );
  AOI22_X1 U7579 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6614), .B1(n6738), 
        .B2(n6613), .ZN(n6609) );
  OAI211_X1 U7580 ( .C1(n6617), .C2(n6743), .A(n6610), .B(n6609), .ZN(U3050)
         );
  AOI22_X1 U7581 ( .A1(n6749), .A2(n6612), .B1(n6747), .B2(n6611), .ZN(n6616)
         );
  AOI22_X1 U7582 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6614), .B1(n6745), 
        .B2(n6613), .ZN(n6615) );
  OAI211_X1 U7583 ( .C1(n6617), .C2(n6754), .A(n6616), .B(n6615), .ZN(U3051)
         );
  AOI22_X1 U7584 ( .A1(n6692), .A2(n6644), .B1(n6618), .B2(n6635), .ZN(n6620)
         );
  AOI22_X1 U7585 ( .A1(n6704), .A2(n6643), .B1(n6693), .B2(n6645), .ZN(n6619)
         );
  OAI211_X1 U7586 ( .C1(n6631), .C2(n6621), .A(n6620), .B(n6619), .ZN(U3076)
         );
  INV_X1 U7587 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6625) );
  AOI22_X1 U7588 ( .A1(n6709), .A2(n6644), .B1(n6643), .B2(n6710), .ZN(n6624)
         );
  AOI22_X1 U7589 ( .A1(n6622), .A2(n6635), .B1(n6708), .B2(n6645), .ZN(n6623)
         );
  OAI211_X1 U7590 ( .C1(n6631), .C2(n6625), .A(n6624), .B(n6623), .ZN(U3077)
         );
  INV_X1 U7591 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U7592 ( .A1(n6714), .A2(n6644), .B1(n6643), .B2(n6716), .ZN(n6628)
         );
  AOI22_X1 U7593 ( .A1(n6626), .A2(n6635), .B1(n6715), .B2(n6645), .ZN(n6627)
         );
  OAI211_X1 U7594 ( .C1(n6631), .C2(n6629), .A(n6628), .B(n6627), .ZN(U3078)
         );
  AOI22_X1 U7595 ( .A1(n6721), .A2(n6644), .B1(n6630), .B2(n6635), .ZN(n6633)
         );
  INV_X1 U7596 ( .A(n6631), .ZN(n6646) );
  AOI22_X1 U7597 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6646), .B1(n6720), 
        .B2(n6645), .ZN(n6632) );
  OAI211_X1 U7598 ( .C1(n6634), .C2(n6639), .A(n6633), .B(n6632), .ZN(U3079)
         );
  AOI22_X1 U7599 ( .A1(n6733), .A2(n6644), .B1(n6636), .B2(n6635), .ZN(n6638)
         );
  AOI22_X1 U7600 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6646), .B1(n6732), 
        .B2(n6645), .ZN(n6637) );
  OAI211_X1 U7601 ( .C1(n6640), .C2(n6639), .A(n6638), .B(n6637), .ZN(U3081)
         );
  AOI22_X1 U7602 ( .A1(n6739), .A2(n6644), .B1(n6643), .B2(n6740), .ZN(n6642)
         );
  AOI22_X1 U7603 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6646), .B1(n6738), 
        .B2(n6645), .ZN(n6641) );
  OAI211_X1 U7604 ( .C1(n6743), .C2(n6649), .A(n6642), .B(n6641), .ZN(U3082)
         );
  AOI22_X1 U7605 ( .A1(n6747), .A2(n6644), .B1(n6643), .B2(n6749), .ZN(n6648)
         );
  AOI22_X1 U7606 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6646), .B1(n6745), 
        .B2(n6645), .ZN(n6647) );
  OAI211_X1 U7607 ( .C1(n6754), .C2(n6649), .A(n6648), .B(n6647), .ZN(U3083)
         );
  NOR2_X1 U7608 ( .A1(n6650), .A2(n6777), .ZN(n6682) );
  AOI22_X1 U7609 ( .A1(n6692), .A2(n6682), .B1(n6681), .B2(n6704), .ZN(n6662)
         );
  OAI21_X1 U7610 ( .B1(n6652), .B2(n6651), .A(n6703), .ZN(n6660) );
  AOI21_X1 U7611 ( .B1(n6654), .B2(n6653), .A(n6682), .ZN(n6659) );
  INV_X1 U7612 ( .A(n6659), .ZN(n6657) );
  AOI21_X1 U7613 ( .B1(n6934), .B2(n6658), .A(n6655), .ZN(n6656) );
  OAI21_X1 U7614 ( .B1(n6660), .B2(n6657), .A(n6656), .ZN(n6684) );
  OAI22_X1 U7615 ( .A1(n6660), .A2(n6659), .B1(n6658), .B2(n6937), .ZN(n6683)
         );
  AOI22_X1 U7616 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6684), .B1(n6693), 
        .B2(n6683), .ZN(n6661) );
  OAI211_X1 U7617 ( .C1(n6707), .C2(n6687), .A(n6662), .B(n6661), .ZN(U3108)
         );
  AOI22_X1 U7618 ( .A1(n6709), .A2(n6682), .B1(n6681), .B2(n6710), .ZN(n6664)
         );
  AOI22_X1 U7619 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6684), .B1(n6708), 
        .B2(n6683), .ZN(n6663) );
  OAI211_X1 U7620 ( .C1(n6713), .C2(n6687), .A(n6664), .B(n6663), .ZN(U3109)
         );
  AOI22_X1 U7621 ( .A1(n6714), .A2(n6682), .B1(n6681), .B2(n6716), .ZN(n6666)
         );
  AOI22_X1 U7622 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6684), .B1(n6715), 
        .B2(n6683), .ZN(n6665) );
  OAI211_X1 U7623 ( .C1(n6719), .C2(n6687), .A(n6666), .B(n6665), .ZN(U3110)
         );
  AOI22_X1 U7624 ( .A1(n6721), .A2(n6682), .B1(n6681), .B2(n6722), .ZN(n6668)
         );
  AOI22_X1 U7625 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6684), .B1(n6720), 
        .B2(n6683), .ZN(n6667) );
  OAI211_X1 U7626 ( .C1(n6725), .C2(n6687), .A(n6668), .B(n6667), .ZN(U3111)
         );
  INV_X1 U7627 ( .A(n6687), .ZN(n6676) );
  AOI22_X1 U7628 ( .A1(n6727), .A2(n6682), .B1(n6676), .B2(n6669), .ZN(n6671)
         );
  AOI22_X1 U7629 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6684), .B1(n6726), 
        .B2(n6683), .ZN(n6670) );
  OAI211_X1 U7630 ( .C1(n6672), .C2(n6679), .A(n6671), .B(n6670), .ZN(U3112)
         );
  AOI22_X1 U7631 ( .A1(n6733), .A2(n6682), .B1(n6681), .B2(n6734), .ZN(n6674)
         );
  AOI22_X1 U7632 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6684), .B1(n6732), 
        .B2(n6683), .ZN(n6673) );
  OAI211_X1 U7633 ( .C1(n6737), .C2(n6687), .A(n6674), .B(n6673), .ZN(U3113)
         );
  AOI22_X1 U7634 ( .A1(n6739), .A2(n6682), .B1(n6676), .B2(n6675), .ZN(n6678)
         );
  AOI22_X1 U7635 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6684), .B1(n6738), 
        .B2(n6683), .ZN(n6677) );
  OAI211_X1 U7636 ( .C1(n6680), .C2(n6679), .A(n6678), .B(n6677), .ZN(U3114)
         );
  AOI22_X1 U7637 ( .A1(n6747), .A2(n6682), .B1(n6681), .B2(n6749), .ZN(n6686)
         );
  AOI22_X1 U7638 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6684), .B1(n6745), 
        .B2(n6683), .ZN(n6685) );
  OAI211_X1 U7639 ( .C1(n6754), .C2(n6687), .A(n6686), .B(n6685), .ZN(U3115)
         );
  INV_X1 U7640 ( .A(n6688), .ZN(n6746) );
  AOI21_X1 U7641 ( .B1(n6690), .B2(n6689), .A(n6746), .ZN(n6698) );
  OAI22_X1 U7642 ( .A1(n6698), .A2(n6934), .B1(n6691), .B2(n6937), .ZN(n6744)
         );
  AOI22_X1 U7643 ( .A1(n6693), .A2(n6744), .B1(n6746), .B2(n6692), .ZN(n6706)
         );
  INV_X1 U7644 ( .A(n6694), .ZN(n6697) );
  OAI21_X1 U7645 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(n6699) );
  NAND2_X1 U7646 ( .A1(n6699), .A2(n6698), .ZN(n6701) );
  OAI211_X1 U7647 ( .C1(n6703), .C2(n6702), .A(n6701), .B(n6700), .ZN(n6750)
         );
  AOI22_X1 U7648 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6750), .B1(n6704), 
        .B2(n6748), .ZN(n6705) );
  OAI211_X1 U7649 ( .C1(n6707), .C2(n6753), .A(n6706), .B(n6705), .ZN(U3140)
         );
  AOI22_X1 U7650 ( .A1(n6709), .A2(n6746), .B1(n6708), .B2(n6744), .ZN(n6712)
         );
  AOI22_X1 U7651 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6750), .B1(n6710), 
        .B2(n6748), .ZN(n6711) );
  OAI211_X1 U7652 ( .C1(n6713), .C2(n6753), .A(n6712), .B(n6711), .ZN(U3141)
         );
  AOI22_X1 U7653 ( .A1(n6715), .A2(n6744), .B1(n6746), .B2(n6714), .ZN(n6718)
         );
  AOI22_X1 U7654 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6750), .B1(n6716), 
        .B2(n6748), .ZN(n6717) );
  OAI211_X1 U7655 ( .C1(n6719), .C2(n6753), .A(n6718), .B(n6717), .ZN(U3142)
         );
  AOI22_X1 U7656 ( .A1(n6721), .A2(n6746), .B1(n6720), .B2(n6744), .ZN(n6724)
         );
  AOI22_X1 U7657 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6750), .B1(n6722), 
        .B2(n6748), .ZN(n6723) );
  OAI211_X1 U7658 ( .C1(n6725), .C2(n6753), .A(n6724), .B(n6723), .ZN(U3143)
         );
  AOI22_X1 U7659 ( .A1(n6727), .A2(n6746), .B1(n6726), .B2(n6744), .ZN(n6730)
         );
  AOI22_X1 U7660 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6750), .B1(n6728), 
        .B2(n6748), .ZN(n6729) );
  OAI211_X1 U7661 ( .C1(n6731), .C2(n6753), .A(n6730), .B(n6729), .ZN(U3144)
         );
  AOI22_X1 U7662 ( .A1(n6733), .A2(n6746), .B1(n6732), .B2(n6744), .ZN(n6736)
         );
  AOI22_X1 U7663 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6750), .B1(n6734), 
        .B2(n6748), .ZN(n6735) );
  OAI211_X1 U7664 ( .C1(n6737), .C2(n6753), .A(n6736), .B(n6735), .ZN(U3145)
         );
  AOI22_X1 U7665 ( .A1(n6739), .A2(n6746), .B1(n6738), .B2(n6744), .ZN(n6742)
         );
  AOI22_X1 U7666 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6750), .B1(n6740), 
        .B2(n6748), .ZN(n6741) );
  OAI211_X1 U7667 ( .C1(n6743), .C2(n6753), .A(n6742), .B(n6741), .ZN(U3146)
         );
  AOI22_X1 U7668 ( .A1(n6747), .A2(n6746), .B1(n6745), .B2(n6744), .ZN(n6752)
         );
  AOI22_X1 U7669 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6750), .B1(n6749), 
        .B2(n6748), .ZN(n6751) );
  OAI211_X1 U7670 ( .C1(n6754), .C2(n6753), .A(n6752), .B(n6751), .ZN(U3147)
         );
  NAND2_X1 U7671 ( .A1(n6755), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6919) );
  INV_X1 U7672 ( .A(n6919), .ZN(n6760) );
  OAI22_X1 U7673 ( .A1(n6758), .A2(n6757), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6756), .ZN(n6911) );
  NOR3_X1 U7674 ( .A1(n6760), .A2(n6911), .A3(n6759), .ZN(n6766) );
  INV_X1 U7675 ( .A(n6766), .ZN(n6763) );
  OAI211_X1 U7676 ( .C1(n6764), .C2(n6763), .A(n6762), .B(n6761), .ZN(n6765)
         );
  OAI21_X1 U7677 ( .B1(n6766), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6765), 
        .ZN(n6771) );
  NAND2_X1 U7678 ( .A1(n6770), .A2(n6771), .ZN(n6767) );
  NAND2_X1 U7679 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  OAI21_X1 U7680 ( .B1(n6771), .B2(n6770), .A(n6769), .ZN(n6773) );
  NAND2_X1 U7681 ( .A1(n6776), .A2(n6777), .ZN(n6772) );
  NAND2_X1 U7682 ( .A1(n6773), .A2(n6772), .ZN(n6775) );
  OAI211_X1 U7683 ( .C1(n6777), .C2(n6776), .A(n6775), .B(n6774), .ZN(n6786)
         );
  NOR2_X1 U7684 ( .A1(MORE_REG_SCAN_IN), .A2(FLUSH_REG_SCAN_IN), .ZN(n6780) );
  OAI211_X1 U7685 ( .C1(n6781), .C2(n6780), .A(n6779), .B(n6778), .ZN(n6782)
         );
  NOR2_X1 U7686 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  AND3_X1 U7687 ( .A1(n6786), .A2(n6785), .A3(n6784), .ZN(n6801) );
  NAND2_X1 U7688 ( .A1(n6801), .A2(n6802), .ZN(n6787) );
  NAND2_X1 U7689 ( .A1(READY_N), .A2(n6932), .ZN(n6805) );
  NAND2_X1 U7690 ( .A1(n6787), .A2(n6805), .ZN(n6792) );
  NOR2_X1 U7691 ( .A1(n6788), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6938) );
  NAND4_X1 U7692 ( .A1(n6790), .A2(n6789), .A3(n6938), .A4(n6827), .ZN(n6791)
         );
  NAND2_X1 U7693 ( .A1(n6792), .A2(n6791), .ZN(n6903) );
  INV_X1 U7694 ( .A(n6903), .ZN(n6808) );
  AOI21_X1 U7695 ( .B1(READY_N), .B2(n6937), .A(n6808), .ZN(n6793) );
  NOR2_X1 U7696 ( .A1(n6793), .A2(n6809), .ZN(n6804) );
  AOI211_X1 U7697 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n6804), .ZN(n6799)
         );
  OAI211_X1 U7698 ( .C1(n6810), .C2(n6797), .A(n6809), .B(n6903), .ZN(n6798)
         );
  OAI211_X1 U7699 ( .C1(n6801), .C2(n6800), .A(n6799), .B(n6798), .ZN(U3148)
         );
  NOR2_X1 U7700 ( .A1(READY_N), .A2(n6809), .ZN(n6811) );
  AOI21_X1 U7701 ( .B1(n6906), .B2(n6811), .A(n6802), .ZN(n6807) );
  AOI21_X1 U7702 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6804), .A(n6803), .ZN(
        n6806) );
  OAI211_X1 U7703 ( .C1(n6808), .C2(n6807), .A(n6806), .B(n6805), .ZN(U3149)
         );
  NAND3_X1 U7704 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), 
        .A3(n6809), .ZN(n6813) );
  OAI211_X1 U7705 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6811), .A(n6902), .B(
        n6810), .ZN(n6812) );
  NAND2_X1 U7706 ( .A1(n6813), .A2(n6812), .ZN(U3150) );
  INV_X1 U7707 ( .A(n6901), .ZN(n6898) );
  AND2_X1 U7708 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6898), .ZN(U3151) );
  NOR2_X1 U7709 ( .A1(n6901), .A2(n6814), .ZN(U3152) );
  AND2_X1 U7710 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6898), .ZN(U3153) );
  AND2_X1 U7711 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6898), .ZN(U3154) );
  NOR2_X1 U7712 ( .A1(n6901), .A2(n6815), .ZN(U3155) );
  AND2_X1 U7713 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6898), .ZN(U3156) );
  AND2_X1 U7714 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6898), .ZN(U3157) );
  AND2_X1 U7715 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6898), .ZN(U3158) );
  AND2_X1 U7716 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6898), .ZN(U3159) );
  AND2_X1 U7717 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6898), .ZN(U3160) );
  AND2_X1 U7718 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6898), .ZN(U3161) );
  AND2_X1 U7719 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6898), .ZN(U3162) );
  AND2_X1 U7720 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6898), .ZN(U3163) );
  AND2_X1 U7721 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6898), .ZN(U3164) );
  AND2_X1 U7722 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6898), .ZN(U3165) );
  AND2_X1 U7723 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6898), .ZN(U3166) );
  AND2_X1 U7724 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6898), .ZN(U3167) );
  AND2_X1 U7725 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6898), .ZN(U3168) );
  NOR2_X1 U7726 ( .A1(n6901), .A2(n6816), .ZN(U3169) );
  AND2_X1 U7727 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6898), .ZN(U3170) );
  AND2_X1 U7728 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6898), .ZN(U3171) );
  AND2_X1 U7729 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6898), .ZN(U3172) );
  AND2_X1 U7730 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6898), .ZN(U3173) );
  AND2_X1 U7731 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6898), .ZN(U3174) );
  NOR2_X1 U7732 ( .A1(n6901), .A2(n6817), .ZN(U3175) );
  AND2_X1 U7733 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6898), .ZN(U3176) );
  AND2_X1 U7734 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6898), .ZN(U3177) );
  NOR2_X1 U7735 ( .A1(n6901), .A2(n6818), .ZN(U3178) );
  AND2_X1 U7736 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6898), .ZN(U3179) );
  AND2_X1 U7737 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6898), .ZN(U3180) );
  NAND2_X1 U7738 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6822) );
  NAND2_X1 U7739 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6828) );
  NAND2_X1 U7740 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n6829) );
  NAND2_X1 U7741 ( .A1(n6828), .A2(n6829), .ZN(n6820) );
  INV_X1 U7742 ( .A(NA_N), .ZN(n6819) );
  AOI221_X1 U7743 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6819), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6834) );
  AOI21_X1 U7744 ( .B1(n6830), .B2(n6820), .A(n6834), .ZN(n6821) );
  OAI221_X1 U7745 ( .B1(n6945), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6945), 
        .C2(n6822), .A(n6821), .ZN(U3181) );
  INV_X1 U7746 ( .A(n6828), .ZN(n6826) );
  INV_X1 U7747 ( .A(n6822), .ZN(n6823) );
  AOI21_X1 U7748 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6823), .ZN(n6825) );
  OAI211_X1 U7749 ( .C1(n6826), .C2(n6825), .A(n6824), .B(n6829), .ZN(U3182)
         );
  AOI221_X1 U7750 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6827), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6832) );
  OAI211_X1 U7751 ( .C1(n6830), .C2(n6829), .A(STATE_REG_0__SCAN_IN), .B(n6828), .ZN(n6831) );
  AOI21_X1 U7752 ( .B1(HOLD), .B2(n6832), .A(n6831), .ZN(n6835) );
  NAND4_X1 U7753 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .A3(
        READY_N), .A4(REQUESTPENDING_REG_SCAN_IN), .ZN(n6833) );
  OAI22_X1 U7754 ( .A1(n6835), .A2(n6834), .B1(NA_N), .B2(n6833), .ZN(U3183)
         );
  NAND2_X1 U7755 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6945), .ZN(n6891) );
  NOR2_X2 U7756 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6931), .ZN(n6889) );
  INV_X1 U7757 ( .A(n6945), .ZN(n6878) );
  AOI22_X1 U7758 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6878), .ZN(n6836) );
  OAI21_X1 U7759 ( .B1(n6921), .B2(n6891), .A(n6836), .ZN(U3184) );
  INV_X1 U7760 ( .A(n6891), .ZN(n6876) );
  INV_X1 U7761 ( .A(n6876), .ZN(n6883) );
  AOI22_X1 U7762 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6878), .ZN(n6837) );
  OAI21_X1 U7763 ( .B1(n6230), .B2(n6883), .A(n6837), .ZN(U3185) );
  AOI22_X1 U7764 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6878), .ZN(n6838) );
  OAI21_X1 U7765 ( .B1(n6839), .B2(n6883), .A(n6838), .ZN(U3186) );
  INV_X1 U7766 ( .A(n6889), .ZN(n6884) );
  OAI222_X1 U7767 ( .A1(n6883), .A2(n6841), .B1(n6840), .B2(n6945), .C1(n4566), 
        .C2(n6884), .ZN(U3187) );
  AOI22_X1 U7768 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6878), .ZN(n6842) );
  OAI21_X1 U7769 ( .B1(n4566), .B2(n6891), .A(n6842), .ZN(U3188) );
  OAI222_X1 U7770 ( .A1(n6883), .A2(n6844), .B1(n6843), .B2(n6945), .C1(n6846), 
        .C2(n6884), .ZN(U3189) );
  OAI222_X1 U7771 ( .A1(n6883), .A2(n6846), .B1(n6845), .B2(n6945), .C1(n6848), 
        .C2(n6884), .ZN(U3190) );
  AOI22_X1 U7772 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6878), .ZN(n6847) );
  OAI21_X1 U7773 ( .B1(n6848), .B2(n6883), .A(n6847), .ZN(U3191) );
  OAI222_X1 U7774 ( .A1(n6883), .A2(n6850), .B1(n6849), .B2(n6945), .C1(n6852), 
        .C2(n6884), .ZN(U3192) );
  AOI22_X1 U7775 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6878), .ZN(n6851) );
  OAI21_X1 U7776 ( .B1(n6852), .B2(n6891), .A(n6851), .ZN(U3193) );
  AOI22_X1 U7777 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6876), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6878), .ZN(n6853) );
  OAI21_X1 U7778 ( .B1(n6855), .B2(n6884), .A(n6853), .ZN(U3194) );
  OAI222_X1 U7779 ( .A1(n6883), .A2(n6855), .B1(n6854), .B2(n6945), .C1(n5385), 
        .C2(n6884), .ZN(U3195) );
  AOI22_X1 U7780 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6878), .ZN(n6856) );
  OAI21_X1 U7781 ( .B1(n5385), .B2(n6891), .A(n6856), .ZN(U3196) );
  AOI22_X1 U7782 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6876), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6878), .ZN(n6857) );
  OAI21_X1 U7783 ( .B1(n6858), .B2(n6884), .A(n6857), .ZN(U3197) );
  OAI222_X1 U7784 ( .A1(n6884), .A2(n5798), .B1(n6859), .B2(n6945), .C1(n6858), 
        .C2(n6883), .ZN(U3198) );
  AOI22_X1 U7785 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6878), .ZN(n6860) );
  OAI21_X1 U7786 ( .B1(n5798), .B2(n6891), .A(n6860), .ZN(U3199) );
  AOI22_X1 U7787 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6878), .ZN(n6861) );
  OAI21_X1 U7788 ( .B1(n6862), .B2(n6891), .A(n6861), .ZN(U3200) );
  AOI22_X1 U7789 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6931), .ZN(n6863) );
  OAI21_X1 U7790 ( .B1(n5790), .B2(n6891), .A(n6863), .ZN(U3201) );
  INV_X1 U7791 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U7792 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6931), .ZN(n6864) );
  OAI21_X1 U7793 ( .B1(n6865), .B2(n6891), .A(n6864), .ZN(U3202) );
  AOI22_X1 U7794 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6876), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6931), .ZN(n6866) );
  OAI21_X1 U7795 ( .B1(n6869), .B2(n6884), .A(n6866), .ZN(U3203) );
  OAI222_X1 U7796 ( .A1(n6883), .A2(n6869), .B1(n6868), .B2(n6945), .C1(n6867), 
        .C2(n6884), .ZN(U3204) );
  AOI22_X1 U7797 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6876), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6931), .ZN(n6870) );
  OAI21_X1 U7798 ( .B1(n6872), .B2(n6884), .A(n6870), .ZN(U3205) );
  AOI22_X1 U7799 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6931), .ZN(n6871) );
  OAI21_X1 U7800 ( .B1(n6872), .B2(n6891), .A(n6871), .ZN(U3206) );
  OAI222_X1 U7801 ( .A1(n6884), .A2(n6875), .B1(n6874), .B2(n6945), .C1(n6873), 
        .C2(n6883), .ZN(U3207) );
  AOI22_X1 U7802 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6876), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6931), .ZN(n6877) );
  OAI21_X1 U7803 ( .B1(n6880), .B2(n6884), .A(n6877), .ZN(U3208) );
  AOI22_X1 U7804 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6878), .ZN(n6879) );
  OAI21_X1 U7805 ( .B1(n6880), .B2(n6891), .A(n6879), .ZN(U3209) );
  OAI222_X1 U7806 ( .A1(n6883), .A2(n6882), .B1(n6881), .B2(n6945), .C1(n6886), 
        .C2(n6884), .ZN(U3210) );
  OAI222_X1 U7807 ( .A1(n6891), .A2(n6886), .B1(n6885), .B2(n6945), .C1(n6888), 
        .C2(n6884), .ZN(U3211) );
  AOI22_X1 U7808 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6931), .ZN(n6887) );
  OAI21_X1 U7809 ( .B1(n6888), .B2(n6891), .A(n6887), .ZN(U3212) );
  AOI22_X1 U7810 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6889), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6931), .ZN(n6890) );
  OAI21_X1 U7811 ( .B1(n6892), .B2(n6891), .A(n6890), .ZN(U3213) );
  MUX2_X1 U7812 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6945), .Z(U3445) );
  MUX2_X1 U7813 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6945), .Z(U3446) );
  AOI22_X1 U7814 ( .A1(n6945), .A2(n6894), .B1(n6893), .B2(n6931), .ZN(U3447)
         );
  INV_X1 U7815 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7816 ( .A1(n6945), .A2(n6896), .B1(n6895), .B2(n6931), .ZN(U3448)
         );
  INV_X1 U7817 ( .A(n6899), .ZN(n6897) );
  AOI21_X1 U7818 ( .B1(n6925), .B2(n6898), .A(n6897), .ZN(U3451) );
  OAI21_X1 U7819 ( .B1(n6901), .B2(n6900), .A(n6899), .ZN(U3452) );
  OAI221_X1 U7820 ( .B1(n6904), .B2(STATE2_REG_0__SCAN_IN), .C1(n6904), .C2(
        n6903), .A(n6902), .ZN(U3453) );
  AOI22_X1 U7821 ( .A1(n6908), .A2(n6907), .B1(n6906), .B2(n6905), .ZN(n6909)
         );
  INV_X1 U7822 ( .A(n6909), .ZN(n6910) );
  MUX2_X1 U7823 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6910), .S(n6916), 
        .Z(U3456) );
  INV_X1 U7824 ( .A(n6911), .ZN(n6913) );
  OAI22_X1 U7825 ( .A1(n6913), .A2(n6918), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6912), .ZN(n6915) );
  OAI22_X1 U7826 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6916), .B1(n6915), .B2(n6914), .ZN(n6917) );
  OAI21_X1 U7827 ( .B1(n6919), .B2(n6918), .A(n6917), .ZN(U3461) );
  NAND2_X1 U7828 ( .A1(n6920), .A2(n6921), .ZN(n6927) );
  NOR2_X1 U7829 ( .A1(n6923), .A2(n6921), .ZN(n6922) );
  AOI22_X1 U7830 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6923), .B1(
        REIP_REG_0__SCAN_IN), .B2(n6922), .ZN(n6924) );
  OAI221_X1 U7831 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6926), .C1(n6925), 
        .C2(n6927), .A(n6924), .ZN(U3468) );
  OAI21_X1 U7832 ( .B1(n6928), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6927), .ZN(
        n6929) );
  INV_X1 U7833 ( .A(n6929), .ZN(U3469) );
  NAND2_X1 U7834 ( .A1(n6931), .A2(W_R_N_REG_SCAN_IN), .ZN(n6930) );
  OAI21_X1 U7835 ( .B1(n6931), .B2(READREQUEST_REG_SCAN_IN), .A(n6930), .ZN(
        U3470) );
  OAI211_X1 U7836 ( .C1(READY_N), .C2(n6328), .A(n6934), .B(n6933), .ZN(n6935)
         );
  NOR2_X1 U7837 ( .A1(n6936), .A2(n6935), .ZN(n6944) );
  OR3_X1 U7838 ( .A1(n6939), .A2(n6938), .A3(n6937), .ZN(n6941) );
  AOI21_X1 U7839 ( .B1(n6941), .B2(STATE2_REG_0__SCAN_IN), .A(n6940), .ZN(
        n6943) );
  NAND2_X1 U7840 ( .A1(n6944), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6942) );
  OAI21_X1 U7841 ( .B1(n6944), .B2(n6943), .A(n6942), .ZN(U3472) );
  MUX2_X1 U7842 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6945), .Z(U3473) );
  NOR2_X2 U3895 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U3551 ( .A1(n6162), .A2(keyinput11), .B1(keyinput78), .B2(n5181), 
        .ZN(n4316) );
  NAND2_X1 U3555 ( .A1(n3294), .A2(n3504), .ZN(n3348) );
  NOR4_X1 U3557 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(DATAO_REG_11__SCAN_IN), 
        .A3(n4519), .A4(n5181), .ZN(n4525) );
  NAND2_X1 U3561 ( .A1(n3360), .A2(n3359), .ZN(n4794) );
  CLKBUF_X2 U3562 ( .A(n4290), .Z(n5774) );
  NAND2_X2 U3564 ( .A1(n3361), .A2(n4794), .ZN(n4722) );
  NAND2_X1 U3568 ( .A1(n5383), .A2(n3687), .ZN(n5574) );
  AND2_X1 U3569 ( .A1(n5311), .A2(n5187), .ZN(n6946) );
  AND2_X1 U3602 ( .A1(n6147), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5311) );
  OR2_X1 U3609 ( .A1(n5485), .A2(n6476), .ZN(n3095) );
  AND2_X2 U3617 ( .A1(n3780), .A2(n3539), .ZN(n3779) );
  AND4_X2 U3641 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), .ZN(n3130)
         );
  AND4_X2 U3726 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3131)
         );
  AND2_X4 U3776 ( .A1(n5159), .A2(n5158), .ZN(n5383) );
  NAND2_X2 U4045 ( .A1(n3641), .A2(n3640), .ZN(n3645) );
  NAND2_X1 U4051 ( .A1(n3345), .A2(n3344), .ZN(n6427) );
  CLKBUF_X1 U4154 ( .A(n3303), .Z(n5438) );
  CLKBUF_X1 U4364 ( .A(n3425), .Z(n3295) );
endmodule

