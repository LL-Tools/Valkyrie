

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474;

  INV_X2 U7176 ( .A(n10023), .ZN(n13687) );
  INV_X2 U7177 ( .A(n9828), .ZN(n13338) );
  BUF_X1 U7178 ( .A(n12131), .Z(n12229) );
  AND3_X1 U7179 ( .A1(n7712), .A2(n7711), .A3(n7710), .ZN(n13222) );
  AND2_X1 U7180 ( .A1(n14693), .A2(n14697), .ZN(n10243) );
  INV_X1 U7181 ( .A(n8544), .ZN(n8614) );
  INV_X1 U7182 ( .A(n12131), .ZN(n12228) );
  AND2_X1 U7183 ( .A1(n11076), .A2(n8598), .ZN(n7792) );
  INV_X1 U7184 ( .A(n11074), .ZN(n10616) );
  AND2_X1 U7185 ( .A1(n8466), .A2(n10962), .ZN(n10305) );
  NAND2_X1 U7186 ( .A1(n14894), .A2(n12315), .ZN(n6625) );
  INV_X1 U7187 ( .A(n12131), .ZN(n12236) );
  NAND2_X1 U7188 ( .A1(n6607), .A2(n8331), .ZN(n13016) );
  NAND2_X1 U7189 ( .A1(n10962), .A2(n9628), .ZN(n8471) );
  INV_X1 U7190 ( .A(n10023), .ZN(n13343) );
  NOR2_X2 U7191 ( .A1(n10881), .A2(n12148), .ZN(n10880) );
  OR2_X1 U7192 ( .A1(n12068), .A2(n9755), .ZN(n14640) );
  NAND2_X1 U7193 ( .A1(n8025), .A2(n7676), .ZN(n8028) );
  INV_X1 U7194 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9236) );
  OAI211_X1 U7195 ( .C1(n9962), .C2(n12054), .A(n9960), .B(n9961), .ZN(n10045)
         );
  XNOR2_X1 U7196 ( .A(n7145), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9726) );
  XNOR2_X1 U7197 ( .A(n9712), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14433) );
  AOI21_X1 U7198 ( .B1(n12911), .B2(n8170), .A(n8161), .ZN(n12919) );
  INV_X1 U7199 ( .A(n6457), .ZN(n14606) );
  INV_X1 U7200 ( .A(n11076), .ZN(n8030) );
  NOR2_X4 U7201 ( .A1(n8234), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8390) );
  OAI21_X2 U7202 ( .B1(n8594), .B2(n7438), .A(n8624), .ZN(n7437) );
  XNOR2_X2 U7203 ( .A(n6625), .B(n12319), .ZN(n14136) );
  NAND2_X2 U7204 ( .A1(n8216), .A2(n8237), .ZN(n10769) );
  NAND2_X1 U7205 ( .A1(n7715), .A2(n7714), .ZN(n8216) );
  INV_X4 U7206 ( .A(n8614), .ZN(n9165) );
  AND2_X4 U7207 ( .A1(n8431), .A2(n13988), .ZN(n8510) );
  AOI21_X2 U7208 ( .B1(n10722), .B2(n10721), .A(n10720), .ZN(n10725) );
  OAI22_X2 U7209 ( .A1(n10434), .A2(n10433), .B1(n10432), .B2(n10431), .ZN(
        n10722) );
  BUF_X4 U7210 ( .A(n8194), .Z(n6428) );
  INV_X1 U7211 ( .A(n8184), .ZN(n8194) );
  AOI211_X2 U7212 ( .C1(n14575), .C2(n15068), .A(n14352), .B(n14351), .ZN(
        n14579) );
  BUF_X4 U7213 ( .A(n12041), .Z(n6429) );
  INV_X1 U7214 ( .A(n11902), .ZN(n12041) );
  AND2_X1 U7215 ( .A1(n7229), .A2(n7230), .ZN(n7187) );
  NOR2_X1 U7216 ( .A1(n6754), .A2(n6753), .ZN(n6752) );
  OAI21_X1 U7217 ( .B1(n13637), .B2(n13795), .A(n7638), .ZN(n13862) );
  NOR2_X1 U7218 ( .A1(n14565), .A2(n6843), .ZN(n6842) );
  XNOR2_X1 U7219 ( .A(n12922), .B(n12921), .ZN(n13145) );
  OR2_X1 U7220 ( .A1(n13597), .A2(n6916), .ZN(n6912) );
  OR2_X1 U7221 ( .A1(n13863), .A2(n7637), .ZN(n6621) );
  OR2_X1 U7222 ( .A1(n8925), .A2(n8924), .ZN(n6984) );
  NAND2_X1 U7223 ( .A1(n13332), .A2(n13331), .ZN(n13361) );
  NAND2_X1 U7224 ( .A1(n6906), .A2(n13591), .ZN(n13749) );
  XNOR2_X1 U7225 ( .A(n13333), .B(n7316), .ZN(n13332) );
  NAND2_X1 U7226 ( .A1(n14090), .A2(n14089), .ZN(n14088) );
  NAND2_X1 U7227 ( .A1(n13444), .A2(n6609), .ZN(n13333) );
  OAI21_X1 U7228 ( .B1(n14116), .B2(n7030), .A(n7028), .ZN(n14090) );
  NAND2_X1 U7229 ( .A1(n12337), .A2(n12336), .ZN(n14116) );
  NAND2_X1 U7230 ( .A1(n9111), .A2(n9110), .ZN(n13871) );
  AND2_X1 U7231 ( .A1(n13832), .A2(n13582), .ZN(n13810) );
  NAND2_X1 U7232 ( .A1(n9060), .A2(n9059), .ZN(n13955) );
  NOR2_X1 U7233 ( .A1(n7016), .A2(n7015), .ZN(n7014) );
  NAND2_X1 U7234 ( .A1(n11944), .A2(n11943), .ZN(n14600) );
  NAND2_X1 U7235 ( .A1(n8998), .A2(n8997), .ZN(n13964) );
  NAND2_X1 U7236 ( .A1(n8983), .A2(n8982), .ZN(n13753) );
  AND2_X1 U7237 ( .A1(n12471), .A2(n12472), .ZN(n12632) );
  OAI21_X1 U7238 ( .B1(n11677), .B2(n11676), .A(n11679), .ZN(n11685) );
  AND2_X1 U7239 ( .A1(n6437), .A2(n6835), .ZN(n14463) );
  OAI21_X1 U7240 ( .B1(n11414), .B2(n11356), .A(n11357), .ZN(n11677) );
  NAND2_X1 U7241 ( .A1(n7385), .A2(n11471), .ZN(n11760) );
  NAND2_X1 U7242 ( .A1(n8909), .A2(n8908), .ZN(n13920) );
  XNOR2_X1 U7243 ( .A(n12268), .B(n12270), .ZN(n12272) );
  OAI21_X1 U7244 ( .B1(n6820), .B2(n10725), .A(n6819), .ZN(n11428) );
  AOI21_X1 U7245 ( .B1(n10949), .B2(n7035), .A(n7034), .ZN(n12268) );
  NAND2_X1 U7246 ( .A1(n6668), .A2(n6666), .ZN(n11601) );
  OR2_X1 U7247 ( .A1(n10744), .A2(n12139), .ZN(n10881) );
  NAND2_X1 U7248 ( .A1(n8673), .A2(n8672), .ZN(n10723) );
  NAND2_X1 U7249 ( .A1(n8653), .A2(n8652), .ZN(n10552) );
  NAND2_X1 U7250 ( .A1(n6866), .A2(n10271), .ZN(n12132) );
  OAI21_X2 U7251 ( .B1(n9630), .B2(n10308), .A(n13841), .ZN(n9631) );
  INV_X2 U7252 ( .A(n13844), .ZN(n6430) );
  NAND2_X1 U7253 ( .A1(n10235), .A2(n10234), .ZN(n14067) );
  INV_X1 U7254 ( .A(n12122), .ZN(n14153) );
  NAND3_X1 U7255 ( .A1(n10241), .A2(n10239), .A3(n6503), .ZN(n14152) );
  AND3_X1 U7256 ( .A1(n9858), .A2(n9857), .A3(n9856), .ZN(n15053) );
  NAND2_X1 U7257 ( .A1(n6997), .A2(n6996), .ZN(n10684) );
  NAND4_X1 U7258 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(n13488)
         );
  INV_X1 U7259 ( .A(n13214), .ZN(n10712) );
  INV_X4 U7260 ( .A(n12037), .ZN(n12059) );
  OR2_X1 U7261 ( .A1(n7941), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U7262 ( .A1(n6990), .A2(n8509), .ZN(n10053) );
  NAND2_X1 U7263 ( .A1(n9378), .A2(n9278), .ZN(n9736) );
  NAND4_X1 U7264 ( .A1(n8480), .A2(n8479), .A3(n8478), .A4(n8477), .ZN(n13489)
         );
  INV_X1 U7265 ( .A(n9673), .ZN(n10541) );
  AND2_X2 U7266 ( .A1(n10615), .A2(n10893), .ZN(n11074) );
  NAND2_X1 U7267 ( .A1(n7704), .A2(n6435), .ZN(n6608) );
  MUX2_X1 U7268 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7703), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n7704) );
  NAND2_X1 U7269 ( .A1(n14700), .A2(n9491), .ZN(n9958) );
  AND2_X2 U7270 ( .A1(n7686), .A2(n7685), .ZN(n8195) );
  XNOR2_X1 U7271 ( .A(n8455), .B(n8454), .ZN(n8482) );
  NAND2_X1 U7272 ( .A1(n6640), .A2(n6639), .ZN(n14697) );
  INV_X1 U7273 ( .A(n9726), .ZN(n14693) );
  AOI21_X1 U7274 ( .B1(n8503), .B2(n6846), .A(n8502), .ZN(n8527) );
  NAND2_X1 U7275 ( .A1(n8464), .A2(n8463), .ZN(n10962) );
  INV_X1 U7276 ( .A(n10304), .ZN(n9628) );
  OR2_X1 U7277 ( .A1(n9274), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U7278 ( .A1(n7039), .A2(n9725), .ZN(n14700) );
  NAND2_X1 U7279 ( .A1(n6435), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U7280 ( .A(n7590), .B(n9365), .ZN(n9491) );
  OR2_X1 U7281 ( .A1(n9364), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U7282 ( .A1(n13299), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7682) );
  OR2_X1 U7283 ( .A1(n7702), .A2(n7699), .ZN(n6435) );
  INV_X2 U7284 ( .A(n8598), .ZN(n9040) );
  NOR2_X1 U7285 ( .A1(n8028), .A2(n6529), .ZN(n7683) );
  AND2_X1 U7286 ( .A1(n7512), .A2(n7674), .ZN(n7511) );
  AND4_X1 U7287 ( .A1(n6597), .A2(n7670), .A3(n6596), .A4(n6664), .ZN(n7756)
         );
  AND4_X1 U7288 ( .A1(n6776), .A2(n6775), .A3(n7675), .A4(n7924), .ZN(n6774)
         );
  AND4_X1 U7289 ( .A1(n6777), .A2(n7833), .A3(n7779), .A4(n7671), .ZN(n7672)
         );
  INV_X1 U7290 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7696) );
  INV_X1 U7291 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7697) );
  INV_X1 U7292 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7833) );
  NOR2_X1 U7293 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n6597) );
  INV_X4 U7294 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7295 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n6775) );
  INV_X1 U7296 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7924) );
  NOR2_X1 U7297 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n6776) );
  NOR2_X1 U7298 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n6777) );
  NOR2_X1 U7299 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9568) );
  NOR2_X1 U7300 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7512) );
  INV_X1 U7301 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8599) );
  INV_X1 U7302 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8648) );
  INV_X4 U7303 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X4 U7304 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7305 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8837) );
  INV_X1 U7306 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7670) );
  NAND2_X4 U7307 ( .A1(n10420), .A2(n10419), .ZN(n10859) );
  INV_X2 U7308 ( .A(n7721), .ZN(n7770) );
  NAND2_X2 U7309 ( .A1(n7687), .A2(n7686), .ZN(n7744) );
  XNOR2_X2 U7310 ( .A(n7684), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7686) );
  INV_X1 U7311 ( .A(n8030), .ZN(n6431) );
  INV_X2 U7312 ( .A(n6431), .ZN(n6432) );
  INV_X1 U7313 ( .A(n6431), .ZN(n6433) );
  AND2_X2 U7314 ( .A1(n8431), .A2(n8434), .ZN(n9160) );
  INV_X4 U7315 ( .A(n11950), .ZN(n8598) );
  BUF_X2 U7316 ( .A(n10697), .Z(n6434) );
  OAI211_X2 U7317 ( .C1(n9393), .C2(n9453), .A(n8488), .B(n8487), .ZN(n9644)
         );
  INV_X1 U7318 ( .A(n13608), .ZN(n7642) );
  NAND2_X1 U7319 ( .A1(n6614), .A2(n8784), .ZN(n8785) );
  NAND2_X1 U7320 ( .A1(n7084), .A2(n7087), .ZN(n6615) );
  AND2_X1 U7321 ( .A1(n13225), .A2(n12895), .ZN(n8384) );
  INV_X1 U7322 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7671) );
  INV_X1 U7323 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6596) );
  AND2_X1 U7324 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  NOR2_X1 U7325 ( .A1(n7018), .A2(n7017), .ZN(n7015) );
  INV_X1 U7326 ( .A(n13748), .ZN(n7016) );
  INV_X1 U7327 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8414) );
  INV_X1 U7328 ( .A(n14697), .ZN(n9727) );
  NOR2_X1 U7329 ( .A1(n12816), .A2(n12817), .ZN(n12818) );
  INV_X1 U7330 ( .A(n15215), .ZN(n14859) );
  NAND2_X1 U7331 ( .A1(n6603), .A2(n6604), .ZN(n7702) );
  INV_X1 U7332 ( .A(n7522), .ZN(n6604) );
  XNOR2_X1 U7333 ( .A(n8211), .B(P3_IR_REG_20__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U7334 ( .A1(n8028), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U7335 ( .A1(n9393), .A2(n8598), .ZN(n8749) );
  NAND2_X2 U7336 ( .A1(n9727), .A2(n14693), .ZN(n12037) );
  NAND2_X1 U7337 ( .A1(n9958), .A2(n8598), .ZN(n11902) );
  NAND2_X1 U7338 ( .A1(n14688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7145) );
  AND2_X1 U7339 ( .A1(n7072), .A2(n12158), .ZN(n7071) );
  INV_X1 U7340 ( .A(n12182), .ZN(n7423) );
  INV_X1 U7341 ( .A(n12183), .ZN(n7422) );
  NAND2_X1 U7342 ( .A1(n8782), .A2(n6486), .ZN(n7529) );
  OAI21_X1 U7343 ( .B1(n8763), .B2(n8762), .A(n6533), .ZN(n6977) );
  AOI21_X1 U7344 ( .B1(n8763), .B2(n8762), .A(n8761), .ZN(n6976) );
  INV_X1 U7345 ( .A(n12186), .ZN(n7416) );
  INV_X1 U7346 ( .A(n8981), .ZN(n7484) );
  OAI21_X1 U7347 ( .B1(n8878), .B2(n7082), .A(n7668), .ZN(n7081) );
  INV_X1 U7348 ( .A(n12715), .ZN(n6804) );
  OR2_X1 U7349 ( .A1(n9234), .A2(n8471), .ZN(n8472) );
  NAND2_X1 U7350 ( .A1(n7212), .A2(n8207), .ZN(n7211) );
  INV_X1 U7351 ( .A(n7215), .ZN(n7212) );
  AOI21_X1 U7352 ( .B1(n7221), .B2(n7217), .A(n7216), .ZN(n7215) );
  INV_X1 U7353 ( .A(n8381), .ZN(n7216) );
  INV_X1 U7354 ( .A(n7685), .ZN(n7687) );
  NAND2_X1 U7355 ( .A1(n6701), .A2(n6493), .ZN(n6700) );
  INV_X1 U7356 ( .A(n12701), .ZN(n6701) );
  NAND2_X1 U7357 ( .A1(n6705), .A2(n11152), .ZN(n6702) );
  NOR2_X1 U7358 ( .A1(n12734), .A2(n6560), .ZN(n11196) );
  NAND2_X1 U7359 ( .A1(n7365), .A2(n7364), .ZN(n7363) );
  NAND2_X1 U7360 ( .A1(n11393), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7364) );
  INV_X1 U7361 ( .A(n12773), .ZN(n7264) );
  AND2_X1 U7362 ( .A1(n7517), .A2(n6476), .ZN(n7516) );
  NAND2_X1 U7363 ( .A1(n7518), .A2(n12952), .ZN(n7517) );
  AND2_X1 U7364 ( .A1(n8364), .A2(n8365), .ZN(n8362) );
  NAND2_X1 U7365 ( .A1(n8111), .A2(n8110), .ZN(n8126) );
  INV_X1 U7366 ( .A(n8112), .ZN(n8111) );
  OR2_X1 U7367 ( .A1(n13269), .A2(n12682), .ZN(n8331) );
  OR2_X1 U7368 ( .A1(n12687), .A2(n14846), .ZN(n8296) );
  INV_X1 U7369 ( .A(n11046), .ZN(n6671) );
  OR2_X1 U7370 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7699) );
  INV_X1 U7371 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U7372 ( .A1(n8089), .A2(n8088), .ZN(n8091) );
  OR2_X1 U7373 ( .A1(n8052), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8053) );
  INV_X1 U7374 ( .A(n7020), .ZN(n7017) );
  AOI21_X1 U7375 ( .B1(n7641), .B2(n11866), .A(n6482), .ZN(n7640) );
  AND2_X1 U7376 ( .A1(n6741), .A2(n7641), .ZN(n6739) );
  NOR2_X1 U7377 ( .A1(n7118), .A2(n11863), .ZN(n7117) );
  INV_X1 U7378 ( .A(n7119), .ZN(n7118) );
  AOI21_X1 U7379 ( .B1(n13666), .B2(n13678), .A(n13634), .ZN(n13648) );
  INV_X1 U7380 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7546) );
  NOR2_X1 U7381 ( .A1(n8714), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8743) );
  OR2_X1 U7382 ( .A1(n8670), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8714) );
  INV_X1 U7383 ( .A(n12396), .ZN(n7571) );
  OR2_X1 U7384 ( .A1(n14107), .A2(n7577), .ZN(n7576) );
  INV_X1 U7385 ( .A(n6864), .ZN(n6861) );
  OR2_X1 U7386 ( .A1(n12308), .A2(n12306), .ZN(n12174) );
  XNOR2_X1 U7387 ( .A(n14152), .B(n14067), .ZN(n12004) );
  INV_X1 U7388 ( .A(n15002), .ZN(n9955) );
  XNOR2_X1 U7389 ( .A(n14155), .B(n10045), .ZN(n12113) );
  NAND2_X1 U7390 ( .A1(n14295), .A2(n7391), .ZN(n7390) );
  NOR2_X1 U7391 ( .A1(n14296), .A2(n7392), .ZN(n7391) );
  INV_X1 U7392 ( .A(n14294), .ZN(n7392) );
  INV_X1 U7393 ( .A(n9298), .ZN(n7279) );
  NAND2_X1 U7394 ( .A1(n7470), .A2(SI_14_), .ZN(n7473) );
  NAND2_X1 U7395 ( .A1(n8711), .A2(n9304), .ZN(n8736) );
  NAND2_X1 U7396 ( .A1(n7083), .A2(n8710), .ZN(n8738) );
  INV_X1 U7397 ( .A(n8499), .ZN(n6846) );
  XNOR2_X1 U7398 ( .A(n8529), .B(SI_2_), .ZN(n8528) );
  XNOR2_X1 U7399 ( .A(n14719), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14760) );
  OR2_X1 U7400 ( .A1(n10415), .A2(n10414), .ZN(n10420) );
  OAI21_X1 U7401 ( .B1(n12578), .B2(n12484), .A(n12486), .ZN(n12586) );
  NAND2_X1 U7402 ( .A1(n10858), .A2(n7176), .ZN(n10988) );
  AND2_X1 U7403 ( .A1(n7177), .A2(n10857), .ZN(n7176) );
  INV_X1 U7404 ( .A(n14861), .ZN(n12636) );
  AOI21_X1 U7405 ( .B1(n7148), .B2(n7151), .A(n6561), .ZN(n7146) );
  INV_X1 U7406 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8389) );
  INV_X1 U7407 ( .A(n8388), .ZN(n7229) );
  INV_X1 U7408 ( .A(n8199), .ZN(n8100) );
  NAND2_X1 U7409 ( .A1(n7685), .A2(n12417), .ZN(n8184) );
  OR2_X1 U7410 ( .A1(n8199), .A2(n11079), .ZN(n7708) );
  NAND2_X1 U7411 ( .A1(n8403), .A2(n8402), .ZN(n10394) );
  INV_X2 U7412 ( .A(n8195), .ZN(n8060) );
  XNOR2_X1 U7413 ( .A(n11196), .B(n7232), .ZN(n11173) );
  OR2_X1 U7414 ( .A1(n11173), .A2(n11161), .ZN(n6708) );
  NAND2_X1 U7415 ( .A1(n6994), .A2(n6993), .ZN(n7263) );
  INV_X1 U7416 ( .A(n11199), .ZN(n6993) );
  OR2_X1 U7417 ( .A1(n12729), .A2(n6573), .ZN(n7371) );
  OR2_X1 U7418 ( .A1(n11185), .A2(n11184), .ZN(n7365) );
  NOR2_X1 U7419 ( .A1(n11395), .A2(n7880), .ZN(n11718) );
  NAND2_X1 U7420 ( .A1(n6983), .A2(n6982), .ZN(n12747) );
  INV_X1 U7421 ( .A(n11720), .ZN(n6982) );
  INV_X1 U7422 ( .A(n7367), .ZN(n7366) );
  AOI21_X1 U7423 ( .B1(n12819), .B2(n12832), .A(n12842), .ZN(n7367) );
  OR2_X1 U7424 ( .A1(n12818), .A2(n12819), .ZN(n6660) );
  XNOR2_X1 U7425 ( .A(n12464), .B(n12677), .ZN(n12921) );
  NAND2_X1 U7426 ( .A1(n12960), .A2(n12447), .ZN(n12947) );
  OR2_X1 U7427 ( .A1(n12967), .A2(n12527), .ZN(n12447) );
  XNOR2_X1 U7428 ( .A(n12954), .B(n12679), .ZN(n12952) );
  OR2_X1 U7429 ( .A1(n12643), .A2(n13059), .ZN(n8322) );
  OAI21_X1 U7430 ( .B1(n13115), .B2(n7199), .A(n7197), .ZN(n13086) );
  INV_X1 U7431 ( .A(n7200), .ZN(n7199) );
  AOI21_X1 U7432 ( .B1(n7200), .B2(n7202), .A(n7198), .ZN(n7197) );
  NAND2_X1 U7433 ( .A1(n7205), .A2(n7206), .ZN(n7204) );
  INV_X1 U7434 ( .A(n13115), .ZN(n7205) );
  INV_X1 U7435 ( .A(n10416), .ZN(n10893) );
  AND2_X1 U7436 ( .A1(n11076), .A2(n11950), .ZN(n7721) );
  OR2_X1 U7437 ( .A1(n7683), .A2(n13298), .ZN(n7684) );
  NAND2_X1 U7438 ( .A1(n6950), .A2(n8122), .ZN(n8134) );
  INV_X1 U7439 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7676) );
  INV_X1 U7440 ( .A(n6941), .ZN(n6940) );
  OAI21_X1 U7441 ( .B1(n8005), .B2(n6942), .A(n8022), .ZN(n6941) );
  NAND2_X1 U7442 ( .A1(n7247), .A2(n7245), .ZN(n8006) );
  AOI21_X1 U7443 ( .B1(n7249), .B2(n7251), .A(n7246), .ZN(n7245) );
  NAND2_X1 U7444 ( .A1(n6924), .A2(n7249), .ZN(n7247) );
  INV_X1 U7445 ( .A(n8003), .ZN(n7246) );
  INV_X1 U7446 ( .A(n7331), .ZN(n6823) );
  AOI21_X1 U7447 ( .B1(n7333), .B2(n7332), .A(n11406), .ZN(n7331) );
  INV_X1 U7448 ( .A(n10724), .ZN(n7332) );
  AND2_X1 U7449 ( .A1(n9232), .A2(n8466), .ZN(n9633) );
  NAND2_X1 U7450 ( .A1(n9192), .A2(n7493), .ZN(n7492) );
  INV_X1 U7451 ( .A(n7494), .ZN(n7493) );
  XNOR2_X1 U7452 ( .A(n11263), .B(n11275), .ZN(n15159) );
  NOR2_X1 U7453 ( .A1(n13619), .A2(n7019), .ZN(n7018) );
  INV_X1 U7454 ( .A(n13617), .ZN(n7019) );
  OR2_X1 U7455 ( .A1(n13763), .A2(n13618), .ZN(n7020) );
  NAND2_X1 U7456 ( .A1(n13778), .A2(n13775), .ZN(n7635) );
  NAND2_X1 U7457 ( .A1(n6922), .A2(n11355), .ZN(n11414) );
  NAND2_X1 U7458 ( .A1(n11354), .A2(n11353), .ZN(n6922) );
  NAND2_X1 U7459 ( .A1(n10356), .A2(n6451), .ZN(n7652) );
  NAND2_X1 U7460 ( .A1(n6749), .A2(n10100), .ZN(n6748) );
  NOR2_X1 U7461 ( .A1(n10327), .A2(n6750), .ZN(n6749) );
  INV_X1 U7462 ( .A(n10099), .ZN(n6750) );
  AOI21_X1 U7463 ( .B1(n10331), .B2(n7005), .A(n6525), .ZN(n7004) );
  INV_X1 U7464 ( .A(n10102), .ZN(n7005) );
  NAND2_X1 U7465 ( .A1(n9946), .A2(n9945), .ZN(n10026) );
  OR2_X1 U7466 ( .A1(n9841), .A2(n6725), .ZN(n6724) );
  AND2_X1 U7467 ( .A1(n9670), .A2(n9669), .ZN(n13795) );
  BUF_X1 U7468 ( .A(n8749), .Z(n9152) );
  INV_X2 U7469 ( .A(n9393), .ZN(n8906) );
  NAND2_X1 U7470 ( .A1(n8482), .A2(n11035), .ZN(n10540) );
  NAND2_X1 U7471 ( .A1(n6620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6619) );
  AND2_X1 U7472 ( .A1(n14005), .A2(n7570), .ZN(n7569) );
  OR2_X1 U7473 ( .A1(n14126), .A2(n7571), .ZN(n7570) );
  AOI21_X1 U7474 ( .B1(n7573), .B2(n7575), .A(n7025), .ZN(n7024) );
  INV_X1 U7475 ( .A(n14082), .ZN(n7025) );
  INV_X1 U7476 ( .A(n7573), .ZN(n7026) );
  NAND2_X1 U7477 ( .A1(n10633), .A2(n10632), .ZN(n7552) );
  AND4_X1 U7478 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n12409) );
  AND2_X1 U7479 ( .A1(n11969), .A2(n11968), .ZN(n14297) );
  NAND2_X1 U7480 ( .A1(n7595), .A2(n6522), .ZN(n7592) );
  NAND2_X1 U7481 ( .A1(n9727), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7595) );
  INV_X1 U7482 ( .A(n14285), .ZN(n6856) );
  NAND2_X1 U7483 ( .A1(n14283), .A2(n7618), .ZN(n14345) );
  NOR2_X1 U7484 ( .A1(n14344), .A2(n7619), .ZN(n7618) );
  INV_X1 U7485 ( .A(n14282), .ZN(n7619) );
  OAI21_X1 U7486 ( .B1(n7401), .B2(n7136), .A(n7134), .ZN(n14372) );
  NOR2_X1 U7487 ( .A1(n7135), .A2(n6487), .ZN(n7134) );
  NOR2_X1 U7488 ( .A1(n14448), .A2(n7622), .ZN(n7621) );
  AOI21_X1 U7489 ( .B1(n14448), .B2(n7131), .A(n6519), .ZN(n7130) );
  INV_X1 U7490 ( .A(n14298), .ZN(n7131) );
  OR2_X1 U7491 ( .A1(n14453), .A2(n7132), .ZN(n7129) );
  OR2_X1 U7492 ( .A1(n14464), .A2(n14471), .ZN(n14298) );
  NOR2_X1 U7493 ( .A1(n14475), .A2(n6836), .ZN(n6835) );
  INV_X1 U7494 ( .A(n6837), .ZN(n6836) );
  OR2_X1 U7495 ( .A1(n14474), .A2(n14473), .ZN(n14270) );
  AND2_X1 U7496 ( .A1(n7599), .A2(n6874), .ZN(n6873) );
  AOI21_X1 U7497 ( .B1(n7600), .B2(n7602), .A(n6516), .ZN(n7599) );
  NAND2_X1 U7498 ( .A1(n7600), .A2(n6875), .ZN(n6874) );
  OR2_X1 U7499 ( .A1(n14263), .A2(n14287), .ZN(n14266) );
  NAND2_X1 U7500 ( .A1(n10823), .A2(n10822), .ZN(n12148) );
  INV_X1 U7501 ( .A(n12004), .ZN(n10251) );
  NAND2_X1 U7502 ( .A1(n6851), .A2(n10226), .ZN(n10460) );
  NAND2_X1 U7503 ( .A1(n10223), .A2(n12001), .ZN(n6851) );
  INV_X1 U7504 ( .A(n14155), .ZN(n10201) );
  INV_X2 U7505 ( .A(n12054), .ZN(n12023) );
  INV_X1 U7506 ( .A(n15079), .ZN(n14936) );
  NOR2_X1 U7507 ( .A1(n9380), .A2(n9738), .ZN(n10191) );
  AND3_X1 U7508 ( .A1(n7277), .A2(n7386), .A3(n7387), .ZN(n7276) );
  NAND2_X2 U7509 ( .A1(n7000), .A2(n6998), .ZN(n11950) );
  NAND2_X1 U7510 ( .A1(n6999), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U7511 ( .A1(n7002), .A2(n7001), .ZN(n7000) );
  NAND3_X1 U7512 ( .A1(n7696), .A2(n7697), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6999) );
  XNOR2_X1 U7513 ( .A(n6867), .B(n8623), .ZN(n10270) );
  NAND2_X1 U7514 ( .A1(n7436), .A2(n8597), .ZN(n6867) );
  NAND2_X1 U7515 ( .A1(n8595), .A2(n8594), .ZN(n7436) );
  AND2_X1 U7516 ( .A1(n7357), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14763) );
  INV_X1 U7517 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7357) );
  AOI21_X1 U7518 ( .B1(n14947), .B2(n14948), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n7348) );
  AOI21_X1 U7519 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14738), .A(n14737), .ZN(
        n14755) );
  NOR2_X1 U7520 ( .A1(n14796), .A2(n14795), .ZN(n14737) );
  AND2_X1 U7521 ( .A1(n6771), .A2(n6770), .ZN(n14826) );
  INV_X1 U7522 ( .A(n14819), .ZN(n6771) );
  NAND2_X1 U7523 ( .A1(n14806), .A2(n14822), .ZN(n6770) );
  NAND2_X1 U7524 ( .A1(n12937), .A2(n6679), .ZN(n13149) );
  NAND2_X1 U7525 ( .A1(n6680), .A2(n15201), .ZN(n6679) );
  NAND2_X1 U7526 ( .A1(n12043), .A2(n12042), .ZN(n14576) );
  AND4_X1 U7527 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n12122) );
  NOR2_X1 U7528 ( .A1(n14947), .A2(n14948), .ZN(n14946) );
  XNOR2_X1 U7529 ( .A(n14826), .B(n14825), .ZN(n14824) );
  AND2_X1 U7530 ( .A1(n8517), .A2(n8516), .ZN(n8523) );
  OAI21_X1 U7531 ( .B1(n12112), .B2(n7414), .A(n7413), .ZN(n7412) );
  INV_X1 U7532 ( .A(n7655), .ZN(n7414) );
  NAND2_X1 U7533 ( .A1(n10515), .A2(n14155), .ZN(n12114) );
  NOR2_X1 U7534 ( .A1(n6527), .A2(n7062), .ZN(n7061) );
  NOR2_X1 U7535 ( .A1(n7063), .A2(n12130), .ZN(n7062) );
  NAND2_X1 U7536 ( .A1(n7431), .A2(n12133), .ZN(n7430) );
  INV_X1 U7537 ( .A(n12138), .ZN(n7068) );
  INV_X1 U7538 ( .A(n12142), .ZN(n12145) );
  NAND2_X1 U7539 ( .A1(n7045), .A2(n7432), .ZN(n12169) );
  NAND2_X1 U7540 ( .A1(n7433), .A2(n12163), .ZN(n7432) );
  NOR2_X1 U7541 ( .A1(n7423), .A2(n7422), .ZN(n7421) );
  AOI21_X1 U7542 ( .B1(n7423), .B2(n7422), .A(n7420), .ZN(n7419) );
  NAND2_X1 U7543 ( .A1(n8803), .A2(n8804), .ZN(n8802) );
  INV_X1 U7544 ( .A(n7538), .ZN(n7537) );
  OAI21_X1 U7545 ( .B1(n7540), .B2(n6465), .A(n8849), .ZN(n7538) );
  AOI21_X1 U7546 ( .B1(n7427), .B2(n7048), .A(n7047), .ZN(n7046) );
  AOI21_X1 U7547 ( .B1(n12204), .B2(n7049), .A(n6536), .ZN(n7048) );
  NOR2_X1 U7548 ( .A1(n7049), .A2(n12204), .ZN(n7047) );
  INV_X1 U7549 ( .A(n12205), .ZN(n7411) );
  NAND2_X1 U7550 ( .A1(n12217), .A2(n7052), .ZN(n7051) );
  INV_X1 U7551 ( .A(n12216), .ZN(n7052) );
  NAND2_X1 U7552 ( .A1(n7535), .A2(n6484), .ZN(n7534) );
  AND2_X1 U7553 ( .A1(n6957), .A2(n9006), .ZN(n6956) );
  INV_X1 U7554 ( .A(n6549), .ZN(n6957) );
  NAND2_X1 U7555 ( .A1(n9007), .A2(n6549), .ZN(n6955) );
  INV_X1 U7556 ( .A(n9189), .ZN(n7497) );
  INV_X1 U7557 ( .A(n9190), .ZN(n7496) );
  NOR2_X1 U7558 ( .A1(n7304), .A2(n6918), .ZN(n6917) );
  INV_X1 U7559 ( .A(n13599), .ZN(n6918) );
  INV_X1 U7560 ( .A(n7305), .ZN(n7304) );
  NAND2_X1 U7561 ( .A1(n12227), .A2(n7057), .ZN(n7056) );
  INV_X1 U7562 ( .A(n12226), .ZN(n7057) );
  NOR2_X1 U7563 ( .A1(n12241), .A2(n14312), .ZN(n7095) );
  NOR2_X1 U7564 ( .A1(n14361), .A2(n7098), .ZN(n12066) );
  NOR2_X1 U7565 ( .A1(n14394), .A2(n7132), .ZN(n7099) );
  AND2_X1 U7566 ( .A1(n14379), .A2(n14306), .ZN(n7139) );
  INV_X1 U7567 ( .A(n7443), .ZN(n7441) );
  NAND2_X1 U7568 ( .A1(n7481), .A2(n7479), .ZN(n9037) );
  AOI21_X1 U7569 ( .B1(n7482), .B2(n7484), .A(n7480), .ZN(n7479) );
  INV_X1 U7570 ( .A(n9019), .ZN(n7480) );
  AOI21_X1 U7571 ( .B1(n7080), .B2(n7082), .A(n7078), .ZN(n7077) );
  INV_X1 U7572 ( .A(n7081), .ZN(n7080) );
  NAND2_X1 U7573 ( .A1(n7079), .A2(n8880), .ZN(n8928) );
  NAND2_X1 U7574 ( .A1(n8739), .A2(n9322), .ZN(n8765) );
  OAI21_X1 U7575 ( .B1(n8528), .B2(n7468), .A(n8551), .ZN(n7467) );
  INV_X1 U7576 ( .A(n8531), .ZN(n7468) );
  OAI21_X1 U7577 ( .B1(n14768), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14718), .ZN(
        n14719) );
  NAND2_X1 U7578 ( .A1(n6951), .A2(n7167), .ZN(n7159) );
  AND2_X1 U7579 ( .A1(n7169), .A2(n7160), .ZN(n6951) );
  INV_X1 U7580 ( .A(n11238), .ZN(n6714) );
  NOR2_X1 U7581 ( .A1(n11237), .A2(n6490), .ZN(n11139) );
  NAND2_X1 U7582 ( .A1(n6800), .A2(n6804), .ZN(n6799) );
  INV_X1 U7583 ( .A(n6801), .ZN(n6800) );
  AOI21_X1 U7584 ( .B1(n7663), .B2(n11115), .A(n6802), .ZN(n6801) );
  INV_X1 U7585 ( .A(n12716), .ZN(n6802) );
  NAND2_X1 U7586 ( .A1(n12698), .A2(n6497), .ZN(n6798) );
  NAND2_X1 U7587 ( .A1(n7263), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U7588 ( .A1(n11393), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7262) );
  OR2_X1 U7589 ( .A1(n13133), .A2(n12907), .ZN(n8381) );
  OR2_X1 U7590 ( .A1(n13170), .A2(n13020), .ZN(n8340) );
  OAI21_X1 U7591 ( .B1(n12428), .B2(n6684), .A(n6682), .ZN(n6687) );
  INV_X1 U7592 ( .A(n6683), .ZN(n6682) );
  OAI21_X1 U7593 ( .B1(n6685), .B2(n6684), .A(n12431), .ZN(n6683) );
  INV_X1 U7594 ( .A(n12429), .ZN(n6684) );
  INV_X1 U7595 ( .A(n8273), .ZN(n7195) );
  INV_X1 U7596 ( .A(n7194), .ZN(n7193) );
  OAI21_X1 U7597 ( .B1(n11441), .B2(n7195), .A(n11047), .ZN(n7194) );
  OAI21_X1 U7598 ( .B1(n11042), .B2(n6459), .A(n11597), .ZN(n6667) );
  AND3_X1 U7599 ( .A1(n7784), .A2(n7783), .A3(n7782), .ZN(n11040) );
  NAND2_X1 U7600 ( .A1(n6601), .A2(n6600), .ZN(n11012) );
  OR2_X1 U7601 ( .A1(n7743), .A2(n11013), .ZN(n6601) );
  INV_X1 U7602 ( .A(n8259), .ZN(n6602) );
  NAND2_X1 U7603 ( .A1(n8400), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U7604 ( .A1(n7922), .A2(n7921), .ZN(n7923) );
  INV_X1 U7605 ( .A(n7885), .ZN(n7234) );
  INV_X1 U7606 ( .A(n7845), .ZN(n6948) );
  AND2_X1 U7607 ( .A1(n7242), .A2(n7807), .ZN(n7241) );
  INV_X1 U7608 ( .A(n7810), .ZN(n7242) );
  NAND2_X1 U7609 ( .A1(n14882), .A2(n6464), .ZN(n6828) );
  INV_X1 U7610 ( .A(n11818), .ZN(n6826) );
  NAND2_X1 U7611 ( .A1(n6975), .A2(n6973), .ZN(n6972) );
  INV_X1 U7612 ( .A(n9547), .ZN(n6902) );
  NOR2_X1 U7613 ( .A1(n6895), .A2(n6901), .ZN(n6894) );
  AND2_X1 U7614 ( .A1(n9807), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6901) );
  INV_X1 U7615 ( .A(n6897), .ZN(n6895) );
  NOR2_X1 U7616 ( .A1(n13660), .A2(n13871), .ZN(n7124) );
  AND2_X1 U7617 ( .A1(n7124), .A2(n7123), .ZN(n7122) );
  INV_X1 U7618 ( .A(n13600), .ZN(n7303) );
  INV_X1 U7619 ( .A(n6917), .ZN(n6916) );
  NAND2_X1 U7620 ( .A1(n6917), .A2(n6915), .ZN(n6914) );
  INV_X1 U7621 ( .A(n6919), .ZN(n6915) );
  AND2_X1 U7622 ( .A1(n13685), .A2(n6543), .ZN(n7634) );
  INV_X1 U7623 ( .A(n7312), .ZN(n7311) );
  AOI21_X1 U7624 ( .B1(n7312), .B2(n7310), .A(n7309), .ZN(n7308) );
  AND2_X1 U7625 ( .A1(n13594), .A2(n7313), .ZN(n7312) );
  INV_X1 U7626 ( .A(n7291), .ZN(n7290) );
  OAI21_X1 U7627 ( .B1(n13809), .B2(n7292), .A(n13585), .ZN(n7291) );
  INV_X1 U7628 ( .A(n13584), .ZN(n7292) );
  AOI21_X1 U7629 ( .B1(n11861), .B2(n6742), .A(n6517), .ZN(n6741) );
  INV_X1 U7630 ( .A(n11696), .ZN(n6742) );
  AND2_X1 U7631 ( .A1(n11420), .A2(n11344), .ZN(n7648) );
  INV_X1 U7632 ( .A(n10935), .ZN(n10933) );
  NAND2_X1 U7633 ( .A1(n10347), .A2(n10546), .ZN(n6909) );
  NOR2_X1 U7634 ( .A1(n10357), .A2(n7297), .ZN(n7296) );
  INV_X1 U7635 ( .A(n10349), .ZN(n7297) );
  NAND2_X1 U7636 ( .A1(n13797), .A2(n13566), .ZN(n13798) );
  AND2_X1 U7637 ( .A1(n8482), .A2(n8481), .ZN(n9665) );
  NOR2_X1 U7638 ( .A1(n8450), .A2(n8443), .ZN(n7649) );
  INV_X1 U7639 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8442) );
  AND2_X1 U7640 ( .A1(n8445), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6989) );
  INV_X1 U7641 ( .A(n8443), .ZN(n8446) );
  INV_X1 U7642 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9235) );
  INV_X1 U7643 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U7644 ( .A1(n12269), .A2(n12270), .ZN(n6638) );
  INV_X1 U7645 ( .A(n10953), .ZN(n7586) );
  NAND2_X1 U7646 ( .A1(n9755), .A2(n10923), .ZN(n7038) );
  NAND2_X1 U7647 ( .A1(n12086), .A2(n12076), .ZN(n12098) );
  AOI21_X1 U7648 ( .B1(n14416), .B2(n7403), .A(n6477), .ZN(n7402) );
  INV_X1 U7649 ( .A(n14302), .ZN(n7403) );
  NOR2_X1 U7650 ( .A1(n14430), .A2(n7128), .ZN(n7127) );
  INV_X1 U7651 ( .A(n7130), .ZN(n7128) );
  NOR2_X1 U7652 ( .A1(n14633), .A2(n6838), .ZN(n6837) );
  INV_X1 U7653 ( .A(n6839), .ZN(n6838) );
  NOR2_X1 U7654 ( .A1(n14547), .A2(n14905), .ZN(n6841) );
  NAND2_X1 U7655 ( .A1(n10817), .A2(n10816), .ZN(n10819) );
  INV_X1 U7656 ( .A(n14397), .ZN(n7138) );
  INV_X1 U7657 ( .A(n14306), .ZN(n7137) );
  NAND2_X1 U7658 ( .A1(n14397), .A2(n7139), .ZN(n14378) );
  NAND2_X1 U7659 ( .A1(n6437), .A2(n6837), .ZN(n14493) );
  NOR2_X1 U7660 ( .A1(n10273), .A2(n12132), .ZN(n10495) );
  INV_X1 U7661 ( .A(n9736), .ZN(n9738) );
  INV_X1 U7662 ( .A(n7489), .ZN(n7488) );
  AOI21_X1 U7663 ( .B1(n7489), .B2(n7487), .A(n7486), .ZN(n7485) );
  INV_X1 U7664 ( .A(n9123), .ZN(n7486) );
  INV_X1 U7665 ( .A(n9131), .ZN(n7487) );
  NAND2_X1 U7666 ( .A1(n9150), .A2(n9082), .ZN(n9132) );
  OR2_X1 U7667 ( .A1(n9148), .A2(n9147), .ZN(n9150) );
  AND3_X1 U7668 ( .A1(n9568), .A2(n9258), .A3(n9257), .ZN(n7387) );
  NOR2_X1 U7669 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n9257) );
  AND2_X1 U7670 ( .A1(n9259), .A2(n9260), .ZN(n7386) );
  AND2_X1 U7671 ( .A1(n7446), .A2(n7444), .ZN(n7443) );
  NAND2_X1 U7672 ( .A1(n7448), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U7673 ( .A1(n7449), .A2(n7445), .ZN(n7444) );
  INV_X1 U7674 ( .A(n9055), .ZN(n7447) );
  XNOR2_X1 U7675 ( .A(n9037), .B(SI_24_), .ZN(n9034) );
  XNOR2_X1 U7676 ( .A(n9012), .B(n9014), .ZN(n8992) );
  NOR2_X1 U7677 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9357) );
  XNOR2_X1 U7678 ( .A(n8953), .B(SI_20_), .ZN(n8952) );
  NAND2_X1 U7679 ( .A1(n8900), .A2(n8929), .ZN(n6613) );
  XNOR2_X1 U7680 ( .A(n8928), .B(SI_18_), .ZN(n8900) );
  NAND2_X1 U7681 ( .A1(n8831), .A2(n8830), .ZN(n8851) );
  OAI21_X1 U7682 ( .B1(n8785), .B2(n7472), .A(n7471), .ZN(n8831) );
  NOR2_X1 U7683 ( .A1(n7474), .A2(SI_14_), .ZN(n7472) );
  NAND2_X1 U7684 ( .A1(n6453), .A2(n7474), .ZN(n7471) );
  AND2_X1 U7685 ( .A1(n8852), .A2(n8834), .ZN(n8850) );
  NAND2_X1 U7686 ( .A1(n8713), .A2(n8736), .ZN(n8737) );
  NAND2_X1 U7687 ( .A1(n7452), .A2(n7453), .ZN(n8708) );
  AOI21_X1 U7688 ( .B1(n7455), .B2(n7457), .A(n6532), .ZN(n7453) );
  NAND2_X1 U7689 ( .A1(n7437), .A2(n6441), .ZN(n7096) );
  INV_X1 U7690 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7272) );
  XNOR2_X1 U7691 ( .A(n8500), .B(SI_1_), .ZN(n8499) );
  XNOR2_X1 U7692 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n6756) );
  AOI21_X1 U7693 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14732), .A(n14731), .ZN(
        n14756) );
  NOR2_X1 U7694 ( .A1(n7159), .A2(n12443), .ZN(n7157) );
  INV_X1 U7695 ( .A(n7159), .ZN(n7158) );
  INV_X1 U7696 ( .A(n12654), .ZN(n7167) );
  NOR2_X1 U7697 ( .A1(n12511), .A2(n12678), .ZN(n7166) );
  AOI21_X1 U7698 ( .B1(n7152), .B2(n7150), .A(n7149), .ZN(n7148) );
  INV_X1 U7699 ( .A(n7154), .ZN(n7150) );
  INV_X1 U7700 ( .A(n12615), .ZN(n7149) );
  INV_X1 U7701 ( .A(n7152), .ZN(n7151) );
  AOI21_X1 U7702 ( .B1(n7180), .B2(n7179), .A(n6565), .ZN(n7178) );
  INV_X1 U7703 ( .A(n12607), .ZN(n7179) );
  OAI211_X1 U7704 ( .C1(n7770), .C2(SI_2_), .A(n7728), .B(n7727), .ZN(n10576)
         );
  OR2_X1 U7705 ( .A1(n7170), .A2(n12570), .ZN(n7169) );
  INV_X1 U7706 ( .A(n7172), .ZN(n7170) );
  NAND2_X1 U7707 ( .A1(n7172), .A2(n12507), .ZN(n7171) );
  NAND2_X1 U7708 ( .A1(n11649), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U7709 ( .A1(n7383), .A2(n7384), .ZN(n7382) );
  XNOR2_X1 U7710 ( .A(n11258), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n11239) );
  NOR2_X1 U7711 ( .A1(n11244), .A2(n6489), .ZN(n11124) );
  NAND2_X1 U7712 ( .A1(n6704), .A2(n6698), .ZN(n6697) );
  AND2_X1 U7713 ( .A1(n11142), .A2(n12700), .ZN(n6698) );
  NAND2_X1 U7714 ( .A1(n6702), .A2(n6700), .ZN(n12732) );
  NAND2_X1 U7715 ( .A1(n6463), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U7716 ( .A1(n6708), .A2(n6495), .ZN(n6994) );
  XNOR2_X1 U7717 ( .A(n7261), .B(n11394), .ZN(n11388) );
  NOR2_X1 U7718 ( .A1(n11388), .A2(n7879), .ZN(n11705) );
  OR2_X1 U7719 ( .A1(n11718), .A2(n11719), .ZN(n6983) );
  INV_X1 U7720 ( .A(n7363), .ZN(n11716) );
  NAND2_X1 U7721 ( .A1(n6710), .A2(n6709), .ZN(n12752) );
  INV_X1 U7722 ( .A(n11707), .ZN(n6709) );
  OAI21_X1 U7723 ( .B1(n12754), .B2(n12771), .A(n6719), .ZN(n12755) );
  NAND2_X1 U7724 ( .A1(n6711), .A2(n12809), .ZN(n6712) );
  OR2_X1 U7725 ( .A1(n8370), .A2(n7219), .ZN(n7218) );
  INV_X1 U7726 ( .A(n8371), .ZN(n7219) );
  INV_X1 U7727 ( .A(n8169), .ZN(n12457) );
  AOI21_X1 U7728 ( .B1(n7516), .B2(n7669), .A(n6537), .ZN(n7514) );
  INV_X1 U7729 ( .A(n7516), .ZN(n7515) );
  NOR2_X1 U7730 ( .A1(n12917), .A2(n12921), .ZN(n12918) );
  NAND2_X1 U7731 ( .A1(n6606), .A2(n8365), .ZN(n12922) );
  NAND2_X1 U7732 ( .A1(n12931), .A2(n8364), .ZN(n6606) );
  INV_X1 U7733 ( .A(n12678), .ZN(n12948) );
  OAI21_X1 U7734 ( .B1(n8087), .B2(n7209), .A(n7207), .ZN(n12951) );
  INV_X1 U7735 ( .A(n7208), .ZN(n7207) );
  OAI21_X1 U7736 ( .B1(n6458), .B2(n7209), .A(n12952), .ZN(n7208) );
  INV_X1 U7737 ( .A(n8356), .ZN(n7209) );
  NOR2_X1 U7738 ( .A1(n12977), .A2(n7502), .ZN(n7501) );
  NAND2_X1 U7739 ( .A1(n7500), .A2(n7498), .ZN(n12960) );
  NOR2_X1 U7740 ( .A1(n7503), .A2(n8104), .ZN(n7498) );
  OR2_X1 U7741 ( .A1(n12974), .A2(n12965), .ZN(n8352) );
  NAND2_X1 U7742 ( .A1(n8087), .A2(n6458), .ZN(n12966) );
  XNOR2_X1 U7743 ( .A(n12974), .B(n12988), .ZN(n12977) );
  OAI21_X1 U7744 ( .B1(n13016), .B2(n7226), .A(n7222), .ZN(n12998) );
  AOI21_X1 U7745 ( .B1(n7225), .B2(n7224), .A(n7223), .ZN(n7222) );
  INV_X1 U7746 ( .A(n8336), .ZN(n7224) );
  INV_X1 U7747 ( .A(n8340), .ZN(n7223) );
  AND2_X1 U7748 ( .A1(n12441), .A2(n12440), .ZN(n7520) );
  OR2_X1 U7749 ( .A1(n12605), .A2(n13028), .ZN(n8336) );
  AND2_X1 U7750 ( .A1(n8331), .A2(n8332), .ZN(n13026) );
  NAND2_X1 U7751 ( .A1(n13060), .A2(n8018), .ZN(n13040) );
  AND4_X1 U7752 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .ZN(n13059)
         );
  AND4_X1 U7753 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n7996), .ZN(n13075)
         );
  AND4_X1 U7754 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n13085)
         );
  AOI21_X1 U7755 ( .B1(n7203), .B2(n8302), .A(n7201), .ZN(n7200) );
  INV_X1 U7756 ( .A(n8305), .ZN(n7201) );
  NAND2_X1 U7757 ( .A1(n6681), .A2(n12429), .ZN(n13098) );
  NAND2_X1 U7758 ( .A1(n12428), .A2(n6685), .ZN(n6681) );
  OR2_X1 U7759 ( .A1(n7918), .A2(n7917), .ZN(n7919) );
  NAND2_X1 U7760 ( .A1(n14851), .A2(n7915), .ZN(n7920) );
  AND4_X1 U7761 ( .A1(n7946), .A2(n7945), .A3(n7944), .A4(n7943), .ZN(n13119)
         );
  AOI21_X1 U7762 ( .B1(n7507), .B2(n7506), .A(n6471), .ZN(n7505) );
  INV_X1 U7763 ( .A(n12422), .ZN(n7506) );
  NAND2_X1 U7764 ( .A1(n7504), .A2(n7507), .ZN(n15193) );
  NAND2_X1 U7765 ( .A1(n11601), .A2(n12422), .ZN(n7504) );
  AOI21_X1 U7766 ( .B1(n7193), .B2(n7195), .A(n7191), .ZN(n7190) );
  INV_X1 U7767 ( .A(n8277), .ZN(n7191) );
  AND2_X1 U7768 ( .A1(n8273), .A2(n8272), .ZN(n11441) );
  NAND3_X1 U7769 ( .A1(n11076), .A2(n11118), .A3(n11074), .ZN(n14857) );
  OR2_X1 U7770 ( .A1(n13213), .A2(n10626), .ZN(n13219) );
  NAND2_X1 U7771 ( .A1(n8139), .A2(n8138), .ZN(n12464) );
  INV_X1 U7772 ( .A(n12421), .ZN(n15282) );
  AND2_X1 U7773 ( .A1(n10402), .A2(n11074), .ZN(n15215) );
  INV_X1 U7774 ( .A(n15218), .ZN(n14854) );
  XNOR2_X1 U7775 ( .A(n8391), .B(n8392), .ZN(n11073) );
  NAND2_X1 U7776 ( .A1(n8165), .A2(n8164), .ZN(n8177) );
  OR2_X1 U7777 ( .A1(n8163), .A2(n8162), .ZN(n8165) );
  NAND2_X1 U7778 ( .A1(n8136), .A2(n8135), .ZN(n8151) );
  OR2_X1 U7779 ( .A1(n8134), .A2(n8133), .ZN(n8136) );
  AND2_X1 U7780 ( .A1(n8389), .A2(n8392), .ZN(n7183) );
  OR2_X1 U7781 ( .A1(n8092), .A2(n11745), .ZN(n8106) );
  NAND2_X1 U7782 ( .A1(n7253), .A2(n7252), .ZN(n8089) );
  AOI21_X1 U7783 ( .B1(n7255), .B2(n7257), .A(n6583), .ZN(n7252) );
  NAND2_X1 U7784 ( .A1(n6944), .A2(n6943), .ZN(n7253) );
  INV_X1 U7785 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8209) );
  OAI21_X1 U7786 ( .B1(n8051), .B2(n6945), .A(n8053), .ZN(n8066) );
  XNOR2_X1 U7787 ( .A(n8052), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8051) );
  INV_X1 U7788 ( .A(n8019), .ZN(n6942) );
  NAND2_X1 U7789 ( .A1(n8020), .A2(n8019), .ZN(n8023) );
  AND2_X1 U7790 ( .A1(n8041), .A2(n8021), .ZN(n8022) );
  NAND2_X1 U7791 ( .A1(n8006), .A2(n8005), .ZN(n8020) );
  NAND2_X1 U7792 ( .A1(n7970), .A2(n7969), .ZN(n6924) );
  NAND2_X1 U7793 ( .A1(n7968), .A2(n7967), .ZN(n7970) );
  NAND2_X1 U7794 ( .A1(n7923), .A2(n9902), .ZN(n7271) );
  NAND2_X1 U7795 ( .A1(n6935), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6934) );
  INV_X1 U7796 ( .A(n7923), .ZN(n6935) );
  INV_X1 U7797 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7673) );
  AND2_X1 U7798 ( .A1(n7885), .A2(n7867), .ZN(n7868) );
  INV_X1 U7799 ( .A(n7865), .ZN(n7237) );
  AND2_X1 U7800 ( .A1(n7865), .A2(n7847), .ZN(n7848) );
  NAND2_X1 U7801 ( .A1(n7846), .A2(n7845), .ZN(n7849) );
  NAND2_X1 U7802 ( .A1(n7849), .A2(n7848), .ZN(n7866) );
  AND2_X1 U7803 ( .A1(n7845), .A2(n7827), .ZN(n7828) );
  OAI21_X1 U7804 ( .B1(n7808), .B2(n7240), .A(n7238), .ZN(n7846) );
  INV_X1 U7805 ( .A(n7239), .ZN(n7238) );
  OAI21_X1 U7806 ( .B1(n7241), .B2(n7240), .A(n7828), .ZN(n7239) );
  INV_X1 U7807 ( .A(n7825), .ZN(n7240) );
  NAND2_X1 U7808 ( .A1(n7808), .A2(n7241), .ZN(n7826) );
  NAND2_X1 U7809 ( .A1(n7796), .A2(n7795), .ZN(n7806) );
  CLKBUF_X1 U7810 ( .A(n7756), .Z(n7757) );
  NAND2_X1 U7811 ( .A1(n6925), .A2(n7736), .ZN(n7752) );
  INV_X1 U7812 ( .A(n7726), .ZN(n7524) );
  INV_X1 U7813 ( .A(n6828), .ZN(n6827) );
  NOR2_X1 U7814 ( .A1(n7326), .A2(n13435), .ZN(n7322) );
  XNOR2_X1 U7815 ( .A(n9828), .B(n10684), .ZN(n9920) );
  AOI21_X1 U7816 ( .B1(n7326), .B2(n13453), .A(n7325), .ZN(n7324) );
  INV_X1 U7817 ( .A(n13323), .ZN(n7325) );
  NOR2_X1 U7818 ( .A1(n7327), .A2(n13368), .ZN(n7326) );
  INV_X1 U7819 ( .A(n7329), .ZN(n7327) );
  NAND2_X1 U7820 ( .A1(n13387), .A2(n6817), .ZN(n13329) );
  NAND2_X1 U7821 ( .A1(n13326), .A2(n6818), .ZN(n6817) );
  INV_X1 U7822 ( .A(n13327), .ZN(n6818) );
  INV_X1 U7823 ( .A(n7335), .ZN(n7334) );
  XNOR2_X1 U7824 ( .A(n9828), .B(n9644), .ZN(n9685) );
  XNOR2_X1 U7825 ( .A(n9828), .B(n10053), .ZN(n9681) );
  NAND2_X1 U7826 ( .A1(n13398), .A2(n6830), .ZN(n13460) );
  NOR2_X1 U7827 ( .A1(n13463), .A2(n13341), .ZN(n6830) );
  NAND2_X1 U7828 ( .A1(n8790), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8819) );
  AND2_X1 U7829 ( .A1(n11821), .A2(n11820), .ZN(n13306) );
  AND2_X1 U7830 ( .A1(n9188), .A2(n9169), .ZN(n9187) );
  NAND2_X1 U7831 ( .A1(n10962), .A2(n10304), .ZN(n9231) );
  INV_X1 U7832 ( .A(n8536), .ZN(n9094) );
  NOR2_X1 U7833 ( .A1(n13511), .A2(n6884), .ZN(n9595) );
  NOR2_X1 U7834 ( .A1(n6886), .A2(n6885), .ZN(n6884) );
  AOI21_X1 U7835 ( .B1(n9436), .B2(n9406), .A(n9405), .ZN(n9543) );
  NAND2_X1 U7836 ( .A1(n6902), .A2(n6898), .ZN(n6897) );
  INV_X1 U7837 ( .A(n9548), .ZN(n6898) );
  OR2_X1 U7838 ( .A1(n15131), .A2(n6899), .ZN(n6896) );
  NAND2_X1 U7839 ( .A1(n6902), .A2(n6900), .ZN(n6899) );
  INV_X1 U7840 ( .A(n15130), .ZN(n6900) );
  NAND2_X1 U7841 ( .A1(n13525), .A2(n11262), .ZN(n11263) );
  NAND2_X1 U7842 ( .A1(n6891), .A2(n13550), .ZN(n6890) );
  INV_X1 U7843 ( .A(n13533), .ZN(n6891) );
  NAND2_X1 U7844 ( .A1(n6890), .A2(n6889), .ZN(n6888) );
  INV_X1 U7845 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6889) );
  NOR2_X1 U7846 ( .A1(n13649), .A2(n7009), .ZN(n7008) );
  NOR2_X1 U7847 ( .A1(n13660), .A2(n7010), .ZN(n7009) );
  OR2_X1 U7848 ( .A1(n7010), .A2(n13640), .ZN(n7639) );
  NAND2_X1 U7849 ( .A1(n13670), .A2(n7124), .ZN(n13658) );
  NAND2_X1 U7850 ( .A1(n13686), .A2(n13600), .ZN(n7307) );
  NAND2_X1 U7851 ( .A1(n13700), .A2(n13599), .ZN(n13686) );
  NAND2_X1 U7852 ( .A1(n6735), .A2(n13627), .ZN(n13697) );
  OAI21_X1 U7853 ( .B1(n7012), .B2(n6733), .A(n6731), .ZN(n6735) );
  AOI21_X1 U7854 ( .B1(n7014), .B2(n7017), .A(n6518), .ZN(n7011) );
  OR2_X1 U7855 ( .A1(n13749), .A2(n13748), .ZN(n13751) );
  NOR2_X1 U7856 ( .A1(n13798), .A2(n13915), .ZN(n13783) );
  NAND2_X1 U7857 ( .A1(n13783), .A2(n13975), .ZN(n13761) );
  NAND2_X1 U7858 ( .A1(n6907), .A2(n13589), .ZN(n13760) );
  OAI21_X1 U7859 ( .B1(n13792), .B2(n13613), .A(n13615), .ZN(n13778) );
  NAND2_X1 U7860 ( .A1(n13810), .A2(n13809), .ZN(n13808) );
  OAI21_X1 U7861 ( .B1(n11865), .B2(n7300), .A(n7298), .ZN(n13832) );
  INV_X1 U7862 ( .A(n7299), .ZN(n7298) );
  OAI21_X1 U7863 ( .B1(n7301), .B2(n7300), .A(n13834), .ZN(n7299) );
  INV_X1 U7864 ( .A(n13579), .ZN(n7300) );
  NAND2_X1 U7865 ( .A1(n6531), .A2(n11360), .ZN(n13824) );
  NAND2_X1 U7866 ( .A1(n6740), .A2(n6741), .ZN(n13605) );
  OR2_X1 U7867 ( .A1(n11697), .A2(n11688), .ZN(n6740) );
  AND2_X1 U7868 ( .A1(n11866), .A2(n11864), .ZN(n7301) );
  NAND2_X1 U7869 ( .A1(n6921), .A2(n11688), .ZN(n11865) );
  INV_X1 U7870 ( .A(n11862), .ZN(n6921) );
  NAND2_X1 U7871 ( .A1(n11668), .A2(n11667), .ZN(n11695) );
  NAND2_X1 U7872 ( .A1(n11345), .A2(n7648), .ZN(n11418) );
  NAND2_X1 U7873 ( .A1(n10933), .A2(n10929), .ZN(n11345) );
  NAND2_X1 U7874 ( .A1(n10928), .A2(n10927), .ZN(n11354) );
  NAND2_X1 U7875 ( .A1(n10926), .A2(n10925), .ZN(n10928) );
  INV_X1 U7876 ( .A(n6909), .ZN(n6911) );
  NAND2_X1 U7877 ( .A1(n7652), .A2(n7651), .ZN(n10692) );
  AND2_X1 U7878 ( .A1(n10548), .A2(n10553), .ZN(n7651) );
  NAND2_X1 U7879 ( .A1(n10350), .A2(n7296), .ZN(n10547) );
  NAND2_X1 U7880 ( .A1(n6748), .A2(n6746), .ZN(n10356) );
  NOR2_X1 U7881 ( .A1(n10352), .A2(n6747), .ZN(n6746) );
  INV_X1 U7882 ( .A(n7004), .ZN(n6747) );
  NAND2_X1 U7883 ( .A1(n10029), .A2(n10028), .ZN(n10100) );
  XNOR2_X1 U7884 ( .A(n9944), .B(n10684), .ZN(n9843) );
  NAND2_X1 U7885 ( .A1(n9847), .A2(n10057), .ZN(n9940) );
  NAND2_X1 U7886 ( .A1(n7630), .A2(n9800), .ZN(n9841) );
  NAND2_X1 U7887 ( .A1(n9795), .A2(n9794), .ZN(n6905) );
  NOR2_X1 U7888 ( .A1(n9797), .A2(n10053), .ZN(n9847) );
  OR2_X1 U7889 ( .A1(n9666), .A2(n9662), .ZN(n9795) );
  NOR2_X1 U7890 ( .A1(n13491), .A2(n9673), .ZN(n9667) );
  INV_X1 U7891 ( .A(n13795), .ZN(n13822) );
  NAND2_X1 U7892 ( .A1(n10049), .A2(n9673), .ZN(n9797) );
  OR2_X1 U7893 ( .A1(n13687), .A2(n9628), .ZN(n9659) );
  XNOR2_X1 U7894 ( .A(n10305), .B(n8482), .ZN(n7315) );
  MUX2_X1 U7895 ( .A(n8484), .B(n14003), .S(n9393), .Z(n9673) );
  OR2_X1 U7896 ( .A1(n14694), .A2(n9089), .ZN(n9091) );
  AND2_X1 U7897 ( .A1(n6751), .A2(n13651), .ZN(n13867) );
  NAND2_X1 U7898 ( .A1(n9045), .A2(n9044), .ZN(n13705) );
  NAND2_X1 U7899 ( .A1(n8957), .A2(n8956), .ZN(n13763) );
  XNOR2_X1 U7900 ( .A(n8428), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U7901 ( .A1(n13981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8428) );
  XNOR2_X1 U7902 ( .A(n8430), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U7903 ( .A1(n8429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U7904 ( .A1(n7545), .A2(n7544), .ZN(n8468) );
  AND2_X1 U7905 ( .A1(n6545), .A2(n8453), .ZN(n7544) );
  INV_X1 U7906 ( .A(n8456), .ZN(n7545) );
  NAND2_X1 U7907 ( .A1(n8464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8458) );
  AND2_X1 U7908 ( .A1(n8743), .A2(n8742), .ZN(n8746) );
  NAND2_X1 U7909 ( .A1(n14116), .A2(n14117), .ZN(n7033) );
  AOI21_X1 U7910 ( .B1(n7569), .B2(n7571), .A(n6512), .ZN(n7568) );
  NAND2_X1 U7911 ( .A1(n14088), .A2(n6569), .ZN(n14026) );
  AND2_X1 U7912 ( .A1(n6634), .A2(n6638), .ZN(n14908) );
  NAND2_X1 U7913 ( .A1(n12272), .A2(n12271), .ZN(n6634) );
  OR2_X1 U7914 ( .A1(n12286), .A2(n7558), .ZN(n7557) );
  INV_X1 U7915 ( .A(n12290), .ZN(n7558) );
  NAND2_X1 U7916 ( .A1(n10635), .A2(n7549), .ZN(n6631) );
  INV_X1 U7917 ( .A(n14052), .ZN(n7583) );
  NOR2_X1 U7918 ( .A1(n7583), .A2(n7584), .ZN(n7582) );
  INV_X1 U7919 ( .A(n14137), .ZN(n7584) );
  AOI21_X1 U7920 ( .B1(n7574), .B2(n7577), .A(n6509), .ZN(n7573) );
  INV_X1 U7921 ( .A(n14117), .ZN(n7029) );
  NOR2_X1 U7922 ( .A1(n14018), .A2(n7032), .ZN(n7031) );
  INV_X1 U7923 ( .A(n12344), .ZN(n7032) );
  AND2_X1 U7924 ( .A1(n12032), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12034) );
  AND2_X1 U7925 ( .A1(n14920), .A2(n14918), .ZN(n12286) );
  OR2_X1 U7926 ( .A1(n10038), .A2(n10037), .ZN(n7581) );
  OR2_X1 U7927 ( .A1(n11996), .A2(n11995), .ZN(n11998) );
  NOR2_X1 U7928 ( .A1(n10635), .A2(n7549), .ZN(n6630) );
  AND2_X1 U7929 ( .A1(n12235), .A2(n12234), .ZN(n12239) );
  OR2_X1 U7930 ( .A1(n12233), .A2(n12232), .ZN(n12234) );
  NAND2_X1 U7931 ( .A1(n7089), .A2(n12248), .ZN(n7088) );
  NAND2_X1 U7932 ( .A1(n12244), .A2(n12245), .ZN(n7089) );
  NAND2_X1 U7933 ( .A1(n7091), .A2(n7090), .ZN(n12243) );
  OR2_X1 U7934 ( .A1(n12084), .A2(n12085), .ZN(n7090) );
  NAND2_X1 U7935 ( .A1(n7092), .A2(n12092), .ZN(n7091) );
  AND4_X1 U7936 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n10225)
         );
  OAI21_X1 U7937 ( .B1(n12037), .B2(n9476), .A(n9872), .ZN(n6649) );
  NOR2_X1 U7938 ( .A1(n14329), .A2(n14321), .ZN(n14314) );
  OR2_X1 U7939 ( .A1(n14384), .A2(n14583), .ZN(n14363) );
  NAND2_X1 U7940 ( .A1(n14375), .A2(n14280), .ZN(n14362) );
  OR2_X1 U7941 ( .A1(n7627), .A2(n7625), .ZN(n7624) );
  INV_X1 U7942 ( .A(n14279), .ZN(n7625) );
  NOR2_X1 U7943 ( .A1(n7626), .A2(n6881), .ZN(n6880) );
  INV_X1 U7944 ( .A(n14276), .ZN(n6881) );
  NAND2_X1 U7945 ( .A1(n7628), .A2(n14279), .ZN(n7626) );
  OAI21_X1 U7946 ( .B1(n14429), .B2(n6879), .A(n6877), .ZN(n14375) );
  INV_X1 U7947 ( .A(n6878), .ZN(n6877) );
  OAI21_X1 U7948 ( .B1(n6880), .B2(n6879), .A(n14376), .ZN(n6878) );
  INV_X1 U7949 ( .A(n7624), .ZN(n6879) );
  AND2_X1 U7950 ( .A1(n14394), .A2(n14277), .ZN(n7627) );
  NAND2_X1 U7951 ( .A1(n7401), .A2(n7399), .ZN(n14397) );
  NAND2_X1 U7952 ( .A1(n6475), .A2(n7628), .ZN(n14417) );
  NAND2_X1 U7953 ( .A1(n14303), .A2(n14302), .ZN(n14412) );
  NOR2_X1 U7954 ( .A1(n14271), .A2(n6438), .ZN(n7389) );
  INV_X1 U7955 ( .A(n14679), .ZN(n14464) );
  NAND2_X1 U7956 ( .A1(n14270), .A2(n7623), .ZN(n14458) );
  AND2_X1 U7957 ( .A1(n14271), .A2(n14269), .ZN(n7623) );
  NAND2_X1 U7958 ( .A1(n6868), .A2(n6869), .ZN(n14474) );
  AOI21_X1 U7959 ( .B1(n6870), .B2(n7601), .A(n6442), .ZN(n6869) );
  NOR2_X1 U7960 ( .A1(n7143), .A2(n14529), .ZN(n7142) );
  INV_X1 U7961 ( .A(n14289), .ZN(n7143) );
  NAND2_X1 U7962 ( .A1(n7141), .A2(n7140), .ZN(n14503) );
  AND2_X1 U7963 ( .A1(n14501), .A2(n14292), .ZN(n7140) );
  NAND2_X1 U7964 ( .A1(n14266), .A2(n14265), .ZN(n14530) );
  NAND2_X1 U7965 ( .A1(n14530), .A2(n14529), .ZN(n14528) );
  NAND2_X1 U7966 ( .A1(n6858), .A2(n6857), .ZN(n14263) );
  AOI21_X1 U7967 ( .B1(n6860), .B2(n12015), .A(n6859), .ZN(n6858) );
  NOR2_X1 U7968 ( .A1(n7615), .A2(n6861), .ZN(n6860) );
  INV_X1 U7969 ( .A(n12019), .ZN(n14287) );
  NAND2_X1 U7970 ( .A1(n11766), .A2(n11765), .ZN(n12308) );
  AND2_X1 U7971 ( .A1(n12174), .A2(n12165), .ZN(n12172) );
  NOR2_X1 U7972 ( .A1(n12172), .A2(n7617), .ZN(n7616) );
  INV_X1 U7973 ( .A(n11767), .ZN(n7617) );
  NAND2_X1 U7974 ( .A1(n6862), .A2(n6864), .ZN(n11485) );
  NAND2_X1 U7975 ( .A1(n6863), .A2(n11531), .ZN(n6862) );
  INV_X1 U7976 ( .A(n11484), .ZN(n6863) );
  NAND2_X1 U7977 ( .A1(n11485), .A2(n12018), .ZN(n11768) );
  NAND2_X1 U7978 ( .A1(n11465), .A2(n11464), .ZN(n11533) );
  NAND2_X1 U7979 ( .A1(n10877), .A2(n7407), .ZN(n11336) );
  NOR2_X1 U7980 ( .A1(n10839), .A2(n7408), .ZN(n7407) );
  INV_X1 U7981 ( .A(n10824), .ZN(n7408) );
  OR2_X1 U7982 ( .A1(n12010), .A2(n6855), .ZN(n6854) );
  INV_X1 U7983 ( .A(n10837), .ZN(n6855) );
  NAND2_X1 U7984 ( .A1(n10819), .A2(n7409), .ZN(n10877) );
  NOR2_X1 U7985 ( .A1(n12011), .A2(n7410), .ZN(n7409) );
  INV_X1 U7986 ( .A(n10818), .ZN(n7410) );
  INV_X1 U7987 ( .A(n14909), .ZN(n11751) );
  NAND2_X1 U7988 ( .A1(n10743), .A2(n12010), .ZN(n10838) );
  OAI21_X1 U7989 ( .B1(n7605), .B2(n10460), .A(n6849), .ZN(n10492) );
  OR2_X1 U7990 ( .A1(n10231), .A2(n7606), .ZN(n7605) );
  NOR2_X1 U7991 ( .A1(n6850), .A2(n12005), .ZN(n6849) );
  NOR2_X1 U7992 ( .A1(n7607), .A2(n7606), .ZN(n6850) );
  INV_X1 U7993 ( .A(n12005), .ZN(n10279) );
  INV_X1 U7994 ( .A(n10460), .ZN(n7610) );
  NAND2_X1 U7995 ( .A1(n10463), .A2(n15073), .ZN(n10462) );
  AND2_X1 U7996 ( .A1(n12118), .A2(n12119), .ZN(n12116) );
  NAND2_X1 U7997 ( .A1(n10197), .A2(n10196), .ZN(n10223) );
  AND2_X1 U7998 ( .A1(n9871), .A2(n9895), .ZN(n15007) );
  OAI21_X1 U7999 ( .B1(n9705), .B2(P1_D_REG_0__SCAN_IN), .A(n9693), .ZN(n10203) );
  NAND2_X1 U8000 ( .A1(n11894), .A2(n11893), .ZN(n14251) );
  INV_X1 U8001 ( .A(n14566), .ZN(n6844) );
  NAND2_X1 U8002 ( .A1(n11963), .A2(n11962), .ZN(n14475) );
  INV_X1 U8003 ( .A(n15072), .ZN(n15062) );
  AND2_X1 U8004 ( .A1(n9370), .A2(n7612), .ZN(n7611) );
  INV_X1 U8005 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7612) );
  NOR2_X1 U8006 ( .A1(n9086), .A2(n7490), .ZN(n7489) );
  INV_X1 U8007 ( .A(n9084), .ZN(n7490) );
  INV_X1 U8008 ( .A(n14688), .ZN(n6642) );
  NOR2_X1 U8009 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6641) );
  NAND2_X1 U8010 ( .A1(n9371), .A2(n9370), .ZN(n7041) );
  AND2_X1 U8011 ( .A1(n7279), .A2(n9270), .ZN(n7275) );
  OAI21_X1 U8012 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9075) );
  NAND2_X1 U8013 ( .A1(n7075), .A2(n8981), .ZN(n9012) );
  NAND2_X1 U8014 ( .A1(n8979), .A2(n8978), .ZN(n7075) );
  NAND2_X1 U8015 ( .A1(n9371), .A2(n7036), .ZN(n9361) );
  NOR2_X1 U8016 ( .A1(n7037), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7036) );
  INV_X1 U8017 ( .A(n8992), .ZN(n11951) );
  NAND2_X1 U8018 ( .A1(n7476), .A2(n7478), .ZN(n8829) );
  NAND2_X1 U8019 ( .A1(n7473), .A2(n7477), .ZN(n7476) );
  XNOR2_X1 U8020 ( .A(n8552), .B(n8550), .ZN(n10111) );
  INV_X1 U8021 ( .A(n8528), .ZN(n7465) );
  OAI21_X1 U8022 ( .B1(n15464), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6479), .ZN(
        n7107) );
  NAND2_X1 U8023 ( .A1(n14723), .A2(n14722), .ZN(n14778) );
  OR2_X1 U8024 ( .A1(n14774), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U8025 ( .A1(n7105), .A2(n14783), .ZN(n14784) );
  NAND2_X1 U8026 ( .A1(n15467), .A2(n15468), .ZN(n7105) );
  NAND2_X1 U8027 ( .A1(n7361), .A2(n14790), .ZN(n14791) );
  NAND2_X1 U8028 ( .A1(n14817), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7361) );
  OAI21_X1 U8029 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14736), .A(n14735), .ZN(
        n14796) );
  OR2_X1 U8030 ( .A1(n14952), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7114) );
  OAI22_X1 U8031 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14740), .B1(n14755), 
        .B2(n14739), .ZN(n14752) );
  NOR2_X1 U8032 ( .A1(n6767), .A2(n6766), .ZN(n6764) );
  NAND2_X1 U8033 ( .A1(n10631), .A2(n7660), .ZN(n10633) );
  OR2_X1 U8034 ( .A1(n10630), .A2(n10629), .ZN(n7660) );
  AND2_X1 U8035 ( .A1(n10577), .A2(n10422), .ZN(n10427) );
  AND3_X1 U8036 ( .A1(n8103), .A2(n8102), .A3(n8101), .ZN(n12978) );
  NAND2_X1 U8037 ( .A1(n8109), .A2(n8108), .ZN(n12954) );
  NAND2_X1 U8038 ( .A1(n12483), .A2(n12482), .ZN(n12578) );
  OR2_X1 U8039 ( .A1(n12586), .A2(n12585), .ZN(n12587) );
  NAND2_X1 U8040 ( .A1(n8095), .A2(n8094), .ZN(n12967) );
  NAND2_X1 U8041 ( .A1(n10711), .A2(n10710), .ZN(n10858) );
  OR2_X1 U8042 ( .A1(n10714), .A2(n10713), .ZN(n12656) );
  AND2_X1 U8043 ( .A1(n7927), .A2(n7926), .ZN(n12621) );
  NAND2_X1 U8044 ( .A1(n10579), .A2(n10580), .ZN(n10711) );
  NAND2_X1 U8045 ( .A1(n10399), .A2(n11070), .ZN(n12674) );
  XNOR2_X1 U8046 ( .A(n8236), .B(n8389), .ZN(n10777) );
  NAND2_X1 U8047 ( .A1(n7188), .A2(n7187), .ZN(n7186) );
  NAND2_X1 U8048 ( .A1(n8213), .A2(n8212), .ZN(n7188) );
  NAND2_X1 U8049 ( .A1(n8119), .A2(n8118), .ZN(n12679) );
  NAND4_X1 U8050 ( .A1(n7732), .A2(n7731), .A3(n7730), .A4(n7729), .ZN(n12691)
         );
  OR2_X1 U8051 ( .A1(n8060), .A2(n11090), .ZN(n7730) );
  AOI21_X1 U8052 ( .B1(n12723), .B2(n11153), .A(n12724), .ZN(n12729) );
  XNOR2_X1 U8053 ( .A(n7371), .B(n11172), .ZN(n11154) );
  NOR2_X1 U8054 ( .A1(n11386), .A2(n11385), .ZN(n11710) );
  NAND2_X1 U8055 ( .A1(n12770), .A2(n6559), .ZN(n12775) );
  XNOR2_X1 U8056 ( .A(n12810), .B(n12809), .ZN(n12783) );
  NOR2_X1 U8057 ( .A1(n12783), .A2(n12782), .ZN(n12808) );
  AOI21_X1 U8058 ( .B1(n6661), .B2(n6660), .A(n12850), .ZN(n12833) );
  NOR2_X1 U8059 ( .A1(n7369), .A2(n7368), .ZN(n6661) );
  OAI211_X1 U8060 ( .C1(n12843), .C2(n12892), .A(n6653), .B(n6652), .ZN(n6651)
         );
  AOI21_X1 U8061 ( .B1(n12859), .B2(n12842), .A(n6654), .ZN(n6653) );
  INV_X1 U8062 ( .A(n12841), .ZN(n6652) );
  AOI21_X1 U8063 ( .B1(n12863), .B2(n12862), .A(n12861), .ZN(n12872) );
  OR2_X1 U8064 ( .A1(n11144), .A2(n11143), .ZN(n12892) );
  NAND2_X1 U8065 ( .A1(n6809), .A2(n6579), .ZN(n7376) );
  NAND2_X1 U8066 ( .A1(n6810), .A2(n12890), .ZN(n6809) );
  NAND2_X1 U8067 ( .A1(n12887), .A2(n12886), .ZN(n7377) );
  XNOR2_X1 U8068 ( .A(n7379), .B(n12885), .ZN(n7378) );
  NAND2_X1 U8069 ( .A1(n12856), .A2(n12882), .ZN(n7379) );
  NAND2_X1 U8070 ( .A1(n8125), .A2(n8124), .ZN(n12942) );
  NAND2_X1 U8071 ( .A1(n8182), .A2(n8181), .ZN(n13225) );
  NOR2_X1 U8072 ( .A1(n13149), .A2(n6483), .ZN(n13239) );
  NAND2_X1 U8073 ( .A1(n8032), .A2(n8031), .ZN(n13269) );
  NAND2_X1 U8074 ( .A1(n7940), .A2(n7939), .ZN(n13289) );
  OR2_X1 U8075 ( .A1(n15295), .A2(n15281), .ZN(n13294) );
  AND2_X1 U8076 ( .A1(n10377), .A2(n10376), .ZN(n13296) );
  INV_X1 U8077 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U8078 ( .A1(n8789), .A2(n8788), .ZN(n14887) );
  NAND2_X1 U8079 ( .A1(n11819), .A2(n11818), .ZN(n6829) );
  NAND2_X1 U8080 ( .A1(n6829), .A2(n6827), .ZN(n14880) );
  AOI21_X1 U8081 ( .B1(n6436), .B2(n13463), .A(n7343), .ZN(n7342) );
  INV_X1 U8082 ( .A(n13374), .ZN(n7343) );
  NOR2_X1 U8083 ( .A1(n11428), .A2(n6988), .ZN(n11554) );
  AND2_X1 U8084 ( .A1(n11429), .A2(n11430), .ZN(n6988) );
  OAI21_X1 U8085 ( .B1(n13361), .B2(n6831), .A(n7317), .ZN(n13397) );
  INV_X1 U8086 ( .A(n13427), .ZN(n6831) );
  NAND2_X1 U8087 ( .A1(n13397), .A2(n13399), .ZN(n13398) );
  NAND2_X1 U8088 ( .A1(n8861), .A2(n8860), .ZN(n13930) );
  OAI21_X1 U8089 ( .B1(n11554), .B2(n11553), .A(n11552), .ZN(n11819) );
  NAND2_X1 U8090 ( .A1(n8603), .A2(n8602), .ZN(n10334) );
  NOR2_X1 U8091 ( .A1(n9595), .A2(n9594), .ZN(n9593) );
  OR2_X1 U8092 ( .A1(n15131), .A2(n15130), .ZN(n15132) );
  NAND2_X1 U8093 ( .A1(n13526), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U8094 ( .A1(n6448), .A2(n10023), .ZN(n13856) );
  XNOR2_X1 U8095 ( .A(n13603), .B(n7007), .ZN(n13865) );
  AND2_X1 U8096 ( .A1(n13856), .A2(n13858), .ZN(n13940) );
  OAI21_X1 U8097 ( .B1(n13865), .B2(n15182), .A(n6923), .ZN(n13947) );
  NOR2_X1 U8098 ( .A1(n13862), .A2(n6621), .ZN(n6923) );
  AND2_X1 U8099 ( .A1(n13864), .A2(n15179), .ZN(n7637) );
  NAND2_X1 U8100 ( .A1(n8752), .A2(n8751), .ZN(n13847) );
  NAND2_X1 U8101 ( .A1(n10954), .A2(n10953), .ZN(n11058) );
  NAND2_X1 U8102 ( .A1(n10949), .A2(n10948), .ZN(n10954) );
  OAI21_X1 U8103 ( .B1(n12389), .B2(n6646), .A(n6643), .ZN(n6647) );
  INV_X1 U8104 ( .A(n14126), .ZN(n6646) );
  AND2_X1 U8105 ( .A1(n6644), .A2(n12396), .ZN(n6643) );
  NAND2_X1 U8106 ( .A1(n14126), .A2(n6645), .ZN(n6644) );
  INV_X1 U8107 ( .A(n14005), .ZN(n7027) );
  NAND2_X1 U8108 ( .A1(n10123), .A2(n10122), .ZN(n10631) );
  NOR2_X1 U8109 ( .A1(n9870), .A2(n9869), .ZN(n10038) );
  NAND2_X1 U8110 ( .A1(n12031), .A2(n12030), .ZN(n14443) );
  NAND2_X1 U8111 ( .A1(n6633), .A2(n7554), .ZN(n14036) );
  AOI21_X1 U8112 ( .B1(n7557), .B2(n7560), .A(n7555), .ZN(n7554) );
  OAI21_X1 U8113 ( .B1(n6637), .B2(n12272), .A(n6635), .ZN(n6633) );
  INV_X1 U8114 ( .A(n14037), .ZN(n7555) );
  NAND2_X1 U8115 ( .A1(n11994), .A2(n11993), .ZN(n14637) );
  NAND2_X1 U8116 ( .A1(n14098), .A2(n14097), .ZN(n14893) );
  NAND2_X1 U8117 ( .A1(n9746), .A2(n9745), .ZN(n14133) );
  NAND2_X1 U8118 ( .A1(n7592), .A2(n9726), .ZN(n7593) );
  NAND2_X1 U8119 ( .A1(n12059), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7594) );
  OAI21_X1 U8120 ( .B1(n14694), .B2(n11902), .A(n11901), .ZN(n14261) );
  XNOR2_X1 U8121 ( .A(n14313), .B(n14312), .ZN(n14567) );
  NAND2_X1 U8122 ( .A1(n14345), .A2(n14285), .ZN(n14338) );
  INV_X1 U8123 ( .A(n15012), .ZN(n14546) );
  NAND2_X1 U8124 ( .A1(n7133), .A2(n10250), .ZN(n10252) );
  INV_X1 U8125 ( .A(n15018), .ZN(n14537) );
  NAND2_X1 U8126 ( .A1(n14700), .A2(n6467), .ZN(n9960) );
  OR2_X1 U8127 ( .A1(n11902), .A2(n9291), .ZN(n9961) );
  NAND3_X1 U8128 ( .A1(n7611), .A2(n9371), .A3(n7144), .ZN(n14688) );
  INV_X1 U8129 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7144) );
  INV_X1 U8130 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14764) );
  XNOR2_X1 U8131 ( .A(n14765), .B(n7102), .ZN(n15473) );
  XNOR2_X1 U8132 ( .A(n14791), .B(n14792), .ZN(n14818) );
  NOR2_X1 U8133 ( .A1(n7348), .A2(n14946), .ZN(n14953) );
  NAND2_X1 U8134 ( .A1(n7353), .A2(n7352), .ZN(n7351) );
  NAND2_X1 U8135 ( .A1(n14797), .A2(n14959), .ZN(n7352) );
  INV_X1 U8136 ( .A(n14956), .ZN(n7353) );
  NAND2_X1 U8137 ( .A1(n14800), .A2(n6501), .ZN(n6763) );
  NAND2_X1 U8138 ( .A1(n7351), .A2(n6764), .ZN(n6758) );
  AOI21_X1 U8139 ( .B1(n7351), .B2(n6760), .A(n6759), .ZN(n14967) );
  NAND2_X1 U8140 ( .A1(n6762), .A2(n6761), .ZN(n6760) );
  OAI21_X1 U8141 ( .B1(n6762), .B2(n7103), .A(n6763), .ZN(n6759) );
  INV_X1 U8142 ( .A(n6764), .ZN(n6761) );
  OAI21_X1 U8143 ( .B1(n14824), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6480), .ZN(
        n6769) );
  AOI21_X1 U8144 ( .B1(n12106), .B2(n12105), .A(n7065), .ZN(n7655) );
  INV_X1 U8145 ( .A(n12107), .ZN(n7065) );
  OAI21_X1 U8146 ( .B1(n7667), .B2(n12121), .A(n12120), .ZN(n12126) );
  AND2_X1 U8147 ( .A1(n7412), .A2(n12113), .ZN(n7667) );
  INV_X1 U8148 ( .A(n12129), .ZN(n7063) );
  INV_X1 U8149 ( .A(n12130), .ZN(n7064) );
  NOR2_X1 U8150 ( .A1(n6991), .A2(n6980), .ZN(n6978) );
  INV_X1 U8151 ( .A(n8591), .ZN(n6980) );
  NOR2_X1 U8152 ( .A1(n7068), .A2(n12136), .ZN(n7067) );
  NAND2_X1 U8153 ( .A1(n6462), .A2(n6968), .ZN(n6967) );
  NAND2_X1 U8154 ( .A1(n6970), .A2(n6969), .ZN(n6968) );
  INV_X1 U8155 ( .A(n8638), .ZN(n6970) );
  INV_X1 U8156 ( .A(n8637), .ZN(n6969) );
  AOI21_X1 U8157 ( .B1(n6962), .B2(n6967), .A(n6452), .ZN(n6960) );
  NAND2_X1 U8158 ( .A1(n6460), .A2(n7548), .ZN(n7547) );
  NAND2_X1 U8159 ( .A1(n6462), .A2(n6965), .ZN(n6964) );
  AND2_X1 U8160 ( .A1(n8638), .A2(n8637), .ZN(n6965) );
  NOR2_X1 U8161 ( .A1(n12154), .A2(n12151), .ZN(n7074) );
  NAND2_X1 U8162 ( .A1(n7426), .A2(n12149), .ZN(n7425) );
  NAND2_X1 U8163 ( .A1(n12154), .A2(n12151), .ZN(n7073) );
  NAND2_X1 U8164 ( .A1(n7074), .A2(n7073), .ZN(n7072) );
  INV_X1 U8165 ( .A(n7043), .ZN(n12177) );
  OAI21_X1 U8166 ( .B1(n12169), .B2(n6526), .A(n7044), .ZN(n7043) );
  NAND2_X1 U8167 ( .A1(n12176), .A2(n12175), .ZN(n7044) );
  NAND2_X1 U8168 ( .A1(n7542), .A2(n7541), .ZN(n7540) );
  INV_X1 U8169 ( .A(n8827), .ZN(n7542) );
  INV_X1 U8170 ( .A(n8826), .ZN(n7541) );
  OAI21_X1 U8171 ( .B1(n7417), .B2(n12181), .A(n7415), .ZN(n12189) );
  AOI21_X1 U8172 ( .B1(n7419), .B2(n6502), .A(n7416), .ZN(n7415) );
  NAND2_X1 U8173 ( .A1(n7418), .A2(n7419), .ZN(n7417) );
  NAND2_X1 U8174 ( .A1(n8808), .A2(n8807), .ZN(n6959) );
  AND2_X1 U8175 ( .A1(n8826), .A2(n8827), .ZN(n7543) );
  INV_X1 U8176 ( .A(n8896), .ZN(n7527) );
  INV_X1 U8177 ( .A(n8947), .ZN(n7526) );
  OAI22_X1 U8178 ( .A1(n12206), .A2(n6449), .B1(n12207), .B2(n7411), .ZN(
        n12210) );
  INV_X1 U8179 ( .A(n8991), .ZN(n7535) );
  NAND2_X1 U8180 ( .A1(n7054), .A2(n12216), .ZN(n7053) );
  AND2_X1 U8181 ( .A1(n9055), .A2(SI_26_), .ZN(n7451) );
  INV_X1 U8182 ( .A(n7483), .ZN(n7482) );
  OAI21_X1 U8183 ( .B1(n8978), .B2(n7484), .A(n9011), .ZN(n7483) );
  INV_X1 U8184 ( .A(n8880), .ZN(n7082) );
  INV_X1 U8185 ( .A(n8934), .ZN(n7078) );
  AND2_X1 U8186 ( .A1(n7460), .A2(n7085), .ZN(n7084) );
  NAND2_X1 U8187 ( .A1(n7086), .A2(n8710), .ZN(n7085) );
  INV_X1 U8188 ( .A(n8707), .ZN(n7086) );
  INV_X1 U8189 ( .A(n8710), .ZN(n7087) );
  INV_X1 U8190 ( .A(n7659), .ZN(n7459) );
  NAND2_X1 U8191 ( .A1(n8708), .A2(n7084), .ZN(n6616) );
  NAND2_X1 U8192 ( .A1(n11141), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6707) );
  OAI21_X1 U8193 ( .B1(n6981), .B2(n6796), .A(n6586), .ZN(n6795) );
  INV_X1 U8194 ( .A(n12782), .ZN(n6796) );
  INV_X1 U8195 ( .A(n6981), .ZN(n6793) );
  OR2_X1 U8196 ( .A1(n7914), .A2(n14844), .ZN(n7916) );
  AND2_X1 U8197 ( .A1(n10771), .A2(n10912), .ZN(n6674) );
  NAND2_X1 U8198 ( .A1(n9053), .A2(n9054), .ZN(n6974) );
  NAND2_X1 U8199 ( .A1(n6954), .A2(n6953), .ZN(n9032) );
  AOI21_X1 U8200 ( .B1(n6956), .B2(n6955), .A(n6562), .ZN(n6953) );
  INV_X1 U8201 ( .A(n9054), .ZN(n6975) );
  INV_X1 U8202 ( .A(n9053), .ZN(n6973) );
  NAND2_X1 U8203 ( .A1(n13748), .A2(n13593), .ZN(n7313) );
  INV_X1 U8204 ( .A(n13595), .ZN(n7309) );
  INV_X1 U8205 ( .A(n13593), .ZN(n7310) );
  INV_X1 U8206 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8408) );
  INV_X1 U8207 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8409) );
  AOI21_X1 U8208 ( .B1(n9056), .B2(n7451), .A(n7450), .ZN(n7449) );
  INV_X1 U8209 ( .A(n9074), .ZN(n7450) );
  INV_X1 U8210 ( .A(n7451), .ZN(n7445) );
  AOI21_X1 U8211 ( .B1(n9056), .B2(n9055), .A(SI_26_), .ZN(n7448) );
  NAND2_X1 U8212 ( .A1(n8828), .A2(n7477), .ZN(n7474) );
  AND2_X1 U8213 ( .A1(n7666), .A2(n6618), .ZN(n7464) );
  NAND2_X1 U8214 ( .A1(n8737), .A2(n8736), .ZN(n6618) );
  INV_X1 U8215 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U8216 ( .B1(n8665), .B2(n7457), .A(n8689), .ZN(n7456) );
  INV_X1 U8217 ( .A(n8668), .ZN(n7457) );
  OAI21_X1 U8218 ( .B1(n11950), .B2(n6848), .A(n6847), .ZN(n8500) );
  NAND2_X1 U8219 ( .A1(n11950), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6847) );
  AOI21_X1 U8220 ( .B1(n12474), .B2(n7154), .A(n7153), .ZN(n7152) );
  INV_X1 U8221 ( .A(n12614), .ZN(n7153) );
  INV_X1 U8222 ( .A(n12497), .ZN(n7182) );
  NAND2_X1 U8223 ( .A1(n12468), .A2(n6492), .ZN(n12472) );
  INV_X1 U8224 ( .A(n12469), .ZN(n7175) );
  NAND2_X1 U8225 ( .A1(n12509), .A2(n12964), .ZN(n7172) );
  INV_X1 U8226 ( .A(n12508), .ZN(n7160) );
  NAND2_X1 U8227 ( .A1(n7168), .A2(n7174), .ZN(n7161) );
  INV_X1 U8228 ( .A(n11252), .ZN(n6791) );
  NAND2_X1 U8229 ( .A1(n7382), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7381) );
  NOR2_X1 U8230 ( .A1(n11139), .A2(n11138), .ZN(n11140) );
  OR2_X1 U8231 ( .A1(n12764), .A2(n6718), .ZN(n7265) );
  NAND2_X1 U8232 ( .A1(n6657), .A2(n6588), .ZN(n12798) );
  NAND2_X1 U8233 ( .A1(n6797), .A2(n12837), .ZN(n12839) );
  NAND2_X1 U8234 ( .A1(n6794), .A2(n6792), .ZN(n6797) );
  NAND2_X1 U8235 ( .A1(n12783), .A2(n6793), .ZN(n6792) );
  INV_X1 U8236 ( .A(n6795), .ZN(n6794) );
  NAND2_X1 U8237 ( .A1(n7259), .A2(n6589), .ZN(n6695) );
  OR2_X1 U8238 ( .A1(n12942), .A2(n12948), .ZN(n8364) );
  INV_X1 U8239 ( .A(n8098), .ZN(n8097) );
  OR2_X1 U8240 ( .A1(n12967), .A2(n12978), .ZN(n8353) );
  OR2_X1 U8241 ( .A1(n12996), .A2(n13004), .ZN(n8344) );
  NAND2_X1 U8242 ( .A1(n13017), .A2(n8336), .ZN(n7227) );
  NAND2_X1 U8243 ( .A1(n8057), .A2(n8056), .ZN(n8070) );
  INV_X1 U8244 ( .A(n8058), .ZN(n8057) );
  NAND2_X1 U8245 ( .A1(n13018), .A2(n13017), .ZN(n7521) );
  NAND2_X1 U8246 ( .A1(n8034), .A2(n8033), .ZN(n8045) );
  NOR2_X1 U8247 ( .A1(n12430), .A2(n6686), .ZN(n6685) );
  INV_X1 U8248 ( .A(n12427), .ZN(n6686) );
  NAND2_X1 U8249 ( .A1(n11600), .A2(n12422), .ZN(n7509) );
  OR2_X1 U8250 ( .A1(n15213), .A2(n11024), .ZN(n8266) );
  NAND2_X1 U8251 ( .A1(n8252), .A2(n8251), .ZN(n10895) );
  INV_X1 U8252 ( .A(n10762), .ZN(n10771) );
  NAND2_X1 U8253 ( .A1(n13257), .A2(n13004), .ZN(n12445) );
  NAND2_X1 U8254 ( .A1(n6599), .A2(n8280), .ZN(n15192) );
  NAND2_X1 U8255 ( .A1(n7189), .A2(n6481), .ZN(n6599) );
  INV_X1 U8256 ( .A(n8282), .ZN(n6598) );
  INV_X1 U8257 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7523) );
  AOI21_X1 U8258 ( .B1(n8053), .B2(n6945), .A(n7256), .ZN(n6943) );
  INV_X1 U8259 ( .A(n8067), .ZN(n7257) );
  NAND2_X1 U8260 ( .A1(n6939), .A2(n6937), .ZN(n8052) );
  AOI21_X1 U8261 ( .B1(n6940), .B2(n6942), .A(n6938), .ZN(n6937) );
  INV_X1 U8262 ( .A(n8041), .ZN(n6938) );
  INV_X1 U8263 ( .A(n7250), .ZN(n7249) );
  OAI21_X1 U8264 ( .B1(n7983), .B2(n7251), .A(n8001), .ZN(n7250) );
  INV_X1 U8265 ( .A(n7984), .ZN(n7251) );
  OAI21_X1 U8266 ( .B1(n7271), .B2(n6930), .A(n7949), .ZN(n6928) );
  OAI22_X1 U8267 ( .A1(n9191), .A2(n7495), .B1(n9194), .B2(n9193), .ZN(n7494)
         );
  NAND2_X1 U8268 ( .A1(n7497), .A2(n7496), .ZN(n7495) );
  AND2_X1 U8269 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  AND2_X1 U8270 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n9113), .ZN(n9135) );
  INV_X1 U8271 ( .A(n6732), .ZN(n6731) );
  OAI21_X1 U8272 ( .B1(n7011), .B2(n6733), .A(n6727), .ZN(n6732) );
  AND2_X1 U8273 ( .A1(n6728), .A2(n13712), .ZN(n6727) );
  OR2_X1 U8274 ( .A1(n6733), .A2(n6729), .ZN(n6728) );
  INV_X1 U8275 ( .A(n13624), .ZN(n6733) );
  NOR2_X1 U8276 ( .A1(n13628), .A2(n6920), .ZN(n6919) );
  INV_X1 U8277 ( .A(n13596), .ZN(n6920) );
  NOR2_X1 U8278 ( .A1(n8885), .A2(n15444), .ZN(n8910) );
  NOR2_X1 U8279 ( .A1(n14887), .A2(n11678), .ZN(n7119) );
  INV_X1 U8280 ( .A(n11347), .ZN(n7645) );
  NOR2_X1 U8281 ( .A1(n8605), .A2(n8604), .ZN(n8629) );
  INV_X1 U8282 ( .A(n9842), .ZN(n6725) );
  NOR2_X1 U8283 ( .A1(n13649), .A2(n13795), .ZN(n6755) );
  NOR2_X1 U8284 ( .A1(n8646), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8649) );
  INV_X1 U8285 ( .A(n12369), .ZN(n7577) );
  AND2_X1 U8286 ( .A1(n12105), .A2(n9736), .ZN(n10039) );
  AND2_X1 U8287 ( .A1(n12074), .A2(n12073), .ZN(n12078) );
  OR2_X1 U8288 ( .A1(n12072), .A2(n14433), .ZN(n12073) );
  NAND2_X1 U8289 ( .A1(n7059), .A2(n12226), .ZN(n7058) );
  NAND2_X1 U8290 ( .A1(n12075), .A2(n12078), .ZN(n12086) );
  XNOR2_X1 U8291 ( .A(n7093), .B(n14433), .ZN(n7092) );
  NOR2_X1 U8292 ( .A1(n12067), .A2(n7094), .ZN(n7093) );
  NAND2_X1 U8293 ( .A1(n6470), .A2(n7095), .ZN(n7094) );
  INV_X1 U8294 ( .A(n7139), .ZN(n7136) );
  NOR2_X1 U8295 ( .A1(n14432), .A2(n14600), .ZN(n7284) );
  NOR2_X1 U8296 ( .A1(n7400), .A2(n14394), .ZN(n7399) );
  INV_X1 U8297 ( .A(n7402), .ZN(n7400) );
  INV_X1 U8298 ( .A(n14272), .ZN(n7622) );
  INV_X1 U8299 ( .A(n14265), .ZN(n6875) );
  INV_X1 U8300 ( .A(n14267), .ZN(n7602) );
  NOR2_X1 U8301 ( .A1(n14637), .A2(n14535), .ZN(n6839) );
  INV_X1 U8302 ( .A(n7616), .ZN(n7615) );
  INV_X1 U8303 ( .A(n7613), .ZN(n6859) );
  AOI21_X1 U8304 ( .B1(n7616), .B2(n7614), .A(n6508), .ZN(n7613) );
  NOR2_X1 U8305 ( .A1(n12308), .A2(n11770), .ZN(n7281) );
  AOI21_X1 U8306 ( .B1(n11531), .B2(n6865), .A(n6513), .ZN(n6864) );
  INV_X1 U8307 ( .A(n11483), .ZN(n6865) );
  NAND2_X1 U8308 ( .A1(n10201), .A2(n10045), .ZN(n12115) );
  INV_X1 U8309 ( .A(n7038), .ZN(n12105) );
  NAND2_X1 U8310 ( .A1(n7285), .A2(n14606), .ZN(n14432) );
  NOR2_X1 U8311 ( .A1(n7441), .A2(n9076), .ZN(n7440) );
  INV_X1 U8312 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9262) );
  INV_X1 U8313 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9261) );
  NOR2_X1 U8314 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n9367) );
  NOR2_X1 U8315 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9269) );
  INV_X1 U8316 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7694) );
  NAND2_X1 U8317 ( .A1(n8955), .A2(n8954), .ZN(n8979) );
  OR2_X1 U8318 ( .A1(n8953), .A2(n10185), .ZN(n8954) );
  NAND2_X1 U8319 ( .A1(n8952), .A2(n8951), .ZN(n8955) );
  AND2_X1 U8320 ( .A1(n8880), .A2(n8856), .ZN(n8878) );
  AOI21_X1 U8321 ( .B1(n7464), .B2(n7462), .A(n7461), .ZN(n7460) );
  INV_X1 U8322 ( .A(n8765), .ZN(n7461) );
  INV_X1 U8323 ( .A(n8736), .ZN(n7462) );
  INV_X1 U8324 ( .A(n7464), .ZN(n7463) );
  OR2_X1 U8325 ( .A1(n9350), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9570) );
  INV_X1 U8326 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9325) );
  INV_X1 U8327 ( .A(n7467), .ZN(n7466) );
  NAND2_X1 U8328 ( .A1(n14716), .A2(n7358), .ZN(n14717) );
  NAND2_X1 U8329 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7359), .ZN(n7358) );
  OAI21_X1 U8330 ( .B1(n14760), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14720), .ZN(
        n14721) );
  XNOR2_X1 U8331 ( .A(n14721), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U8332 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14725), .B1(n14778), .B2(
        n14724), .ZN(n14726) );
  OR2_X1 U8333 ( .A1(n14725), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14724) );
  OAI21_X1 U8334 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14730), .A(n14729), .ZN(
        n14787) );
  INV_X1 U8335 ( .A(n10039), .ZN(n12361) );
  NOR2_X1 U8336 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7764) );
  NAND2_X1 U8337 ( .A1(n10988), .A2(n10987), .ZN(n10989) );
  INV_X1 U8338 ( .A(n11040), .ZN(n11024) );
  NAND2_X1 U8339 ( .A1(n7993), .A2(n7992), .ZN(n8012) );
  INV_X1 U8340 ( .A(n7994), .ZN(n7993) );
  INV_X1 U8341 ( .A(n7161), .ZN(n12595) );
  OR2_X1 U8342 ( .A1(n12558), .A2(n14858), .ZN(n7154) );
  NAND2_X1 U8343 ( .A1(n7161), .A2(n7160), .ZN(n7173) );
  NAND2_X1 U8344 ( .A1(n7959), .A2(n7958), .ZN(n7975) );
  INV_X1 U8345 ( .A(n7960), .ZN(n7959) );
  NOR2_X1 U8346 ( .A1(n7270), .A2(n8384), .ZN(n8231) );
  AOI21_X1 U8347 ( .B1(n7213), .B2(n6445), .A(n7210), .ZN(n8208) );
  NAND2_X1 U8348 ( .A1(n6538), .A2(n7211), .ZN(n7210) );
  AND2_X1 U8349 ( .A1(n8202), .A2(n8189), .ZN(n12895) );
  OR2_X1 U8350 ( .A1(n7704), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6816) );
  NOR2_X1 U8351 ( .A1(n6815), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6814) );
  NOR2_X1 U8352 ( .A1(n11095), .A2(n6789), .ZN(n6780) );
  INV_X1 U8353 ( .A(n11295), .ZN(n6789) );
  AOI21_X1 U8354 ( .B1(n11578), .B2(n11294), .A(n11577), .ZN(n6786) );
  NAND2_X1 U8355 ( .A1(n6717), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11584) );
  INV_X1 U8356 ( .A(n11582), .ZN(n6717) );
  NAND2_X1 U8357 ( .A1(n6716), .A2(n6714), .ZN(n6713) );
  INV_X1 U8358 ( .A(n11239), .ZN(n6716) );
  NAND2_X1 U8359 ( .A1(n6791), .A2(n6784), .ZN(n6783) );
  INV_X1 U8360 ( .A(n11253), .ZN(n6784) );
  AOI21_X1 U8361 ( .B1(n7381), .B2(n11245), .A(n11246), .ZN(n11244) );
  NAND2_X1 U8362 ( .A1(n7380), .A2(n11245), .ZN(n11587) );
  INV_X1 U8363 ( .A(n7381), .ZN(n7380) );
  NOR2_X1 U8364 ( .A1(n11124), .A2(n11138), .ZN(n11125) );
  NAND2_X1 U8365 ( .A1(n12701), .A2(n12699), .ZN(n6703) );
  NAND2_X1 U8366 ( .A1(n6790), .A2(n11208), .ZN(n12696) );
  NAND2_X1 U8367 ( .A1(n6782), .A2(n6781), .ZN(n6790) );
  AND2_X1 U8368 ( .A1(n6783), .A2(n11100), .ZN(n6781) );
  NOR2_X1 U8369 ( .A1(n11126), .A2(n11142), .ZN(n12727) );
  OAI21_X1 U8370 ( .B1(n12698), .B2(n11115), .A(n7663), .ZN(n12717) );
  NAND2_X1 U8371 ( .A1(n6798), .A2(n6799), .ZN(n12719) );
  NAND2_X1 U8372 ( .A1(n6803), .A2(n7662), .ZN(n11192) );
  NAND2_X1 U8373 ( .A1(n6798), .A2(n6450), .ZN(n6803) );
  XNOR2_X1 U8374 ( .A(n7363), .B(n11394), .ZN(n11395) );
  OR2_X1 U8375 ( .A1(n11705), .A2(n11706), .ZN(n6710) );
  INV_X1 U8376 ( .A(n7261), .ZN(n11704) );
  INV_X1 U8377 ( .A(n7375), .ZN(n7372) );
  INV_X1 U8378 ( .A(n6656), .ZN(n12763) );
  NAND2_X1 U8379 ( .A1(n7373), .A2(n6656), .ZN(n6659) );
  OR2_X1 U8380 ( .A1(n7954), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U8381 ( .A1(n6696), .A2(n6695), .ZN(n12829) );
  NAND2_X1 U8382 ( .A1(n6691), .A2(n7368), .ZN(n6696) );
  NAND2_X1 U8383 ( .A1(n7259), .A2(n7258), .ZN(n6691) );
  OAI21_X1 U8384 ( .B1(n12849), .B2(n14805), .A(n12836), .ZN(n6654) );
  NAND2_X1 U8385 ( .A1(n6692), .A2(n6695), .ZN(n12863) );
  AOI21_X1 U8386 ( .B1(n6690), .B2(n7368), .A(n6689), .ZN(n6692) );
  INV_X1 U8387 ( .A(n6693), .ZN(n6689) );
  AOI21_X1 U8388 ( .B1(n7368), .B2(n12827), .A(n13191), .ZN(n6693) );
  NAND2_X1 U8389 ( .A1(n6694), .A2(n7368), .ZN(n12862) );
  NAND2_X1 U8390 ( .A1(n7259), .A2(n7258), .ZN(n6694) );
  NOR2_X1 U8391 ( .A1(n12677), .A2(n12464), .ZN(n12448) );
  NOR2_X1 U8392 ( .A1(n12946), .A2(n7669), .ZN(n12932) );
  NOR2_X1 U8393 ( .A1(n12947), .A2(n12952), .ZN(n12946) );
  OR2_X1 U8394 ( .A1(n8070), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8081) );
  AND2_X1 U8395 ( .A1(n8340), .A2(n8341), .ZN(n13011) );
  NAND2_X1 U8396 ( .A1(n7521), .A2(n12440), .ZN(n13001) );
  NAND2_X1 U8397 ( .A1(n13040), .A2(n6564), .ZN(n6607) );
  NAND2_X1 U8398 ( .A1(n8336), .A2(n8337), .ZN(n13017) );
  NAND2_X1 U8399 ( .A1(n13056), .A2(n13057), .ZN(n7519) );
  AND2_X1 U8400 ( .A1(n8322), .A2(n8325), .ZN(n13047) );
  NAND2_X1 U8401 ( .A1(n8319), .A2(n13041), .ZN(n13057) );
  NAND2_X1 U8402 ( .A1(n6687), .A2(n7510), .ZN(n12433) );
  AOI21_X1 U8403 ( .B1(n13097), .B2(n12431), .A(n6514), .ZN(n7510) );
  NAND2_X1 U8404 ( .A1(n7929), .A2(n7928), .ZN(n7941) );
  INV_X1 U8405 ( .A(n7930), .ZN(n7929) );
  OR2_X1 U8406 ( .A1(n15197), .A2(n12636), .ZN(n14842) );
  AND3_X1 U8407 ( .A1(n7913), .A2(n7912), .A3(n7911), .ZN(n14846) );
  INV_X1 U8408 ( .A(n12426), .ZN(n14844) );
  NOR2_X1 U8409 ( .A1(n7877), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7895) );
  AND2_X1 U8410 ( .A1(n14842), .A2(n8290), .ZN(n14850) );
  AND3_X1 U8411 ( .A1(n7894), .A2(n7893), .A3(n7892), .ZN(n14861) );
  OR2_X1 U8412 ( .A1(n7859), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U8413 ( .A1(n12423), .A2(n12422), .ZN(n15195) );
  NAND2_X1 U8414 ( .A1(n6670), .A2(n6669), .ZN(n6668) );
  NOR2_X1 U8415 ( .A1(n11043), .A2(n6459), .ZN(n6669) );
  OR2_X1 U8416 ( .A1(n11601), .A2(n11600), .ZN(n12423) );
  NOR2_X1 U8417 ( .A1(n7803), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7818) );
  AND2_X1 U8418 ( .A1(n7818), .A2(n11736), .ZN(n7839) );
  NAND2_X1 U8419 ( .A1(n6672), .A2(n11046), .ZN(n11599) );
  OAI21_X1 U8420 ( .B1(n11044), .B2(n11043), .A(n11042), .ZN(n6672) );
  OR2_X1 U8421 ( .A1(n7786), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U8422 ( .A1(n10763), .A2(n10762), .ZN(n6605) );
  NAND2_X1 U8423 ( .A1(n10597), .A2(n10596), .ZN(n15218) );
  NAND2_X1 U8424 ( .A1(n8155), .A2(n8154), .ZN(n13139) );
  NAND2_X1 U8425 ( .A1(n8044), .A2(n8043), .ZN(n12605) );
  INV_X1 U8426 ( .A(n15281), .ZN(n15287) );
  OR2_X1 U8427 ( .A1(n10389), .A2(n10610), .ZN(n10591) );
  AND2_X1 U8428 ( .A1(n10394), .A2(n13295), .ZN(n11070) );
  INV_X1 U8429 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7763) );
  INV_X1 U8430 ( .A(n8178), .ZN(n7267) );
  INV_X1 U8431 ( .A(n7269), .ZN(n7268) );
  OAI21_X1 U8432 ( .B1(n8151), .B2(n8150), .A(n8152), .ZN(n8163) );
  NAND2_X1 U8433 ( .A1(n6779), .A2(n6778), .ZN(n8400) );
  INV_X1 U8434 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8435 ( .A1(n8106), .A2(n6949), .ZN(n8121) );
  AND2_X1 U8436 ( .A1(n8019), .A2(n8004), .ZN(n8005) );
  OAI21_X1 U8437 ( .B1(n6932), .B2(n6929), .A(n6927), .ZN(n7968) );
  NAND2_X1 U8438 ( .A1(n7947), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6929) );
  INV_X1 U8439 ( .A(n6934), .ZN(n6932) );
  INV_X1 U8440 ( .A(n6928), .ZN(n6927) );
  NAND2_X1 U8441 ( .A1(n7903), .A2(n7902), .ZN(n7906) );
  AND2_X1 U8442 ( .A1(n7921), .A2(n7904), .ZN(n7905) );
  NAND2_X1 U8443 ( .A1(n7906), .A2(n7905), .ZN(n7922) );
  AND2_X1 U8444 ( .A1(n7233), .A2(n6947), .ZN(n6946) );
  NAND2_X1 U8445 ( .A1(n7235), .A2(n6948), .ZN(n6947) );
  AOI21_X1 U8446 ( .B1(n7235), .B2(n7237), .A(n7234), .ZN(n7233) );
  AND2_X1 U8447 ( .A1(n7902), .A2(n7887), .ZN(n7888) );
  NAND2_X1 U8448 ( .A1(n7889), .A2(n7888), .ZN(n7903) );
  OR2_X1 U8449 ( .A1(n7813), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U8450 ( .A1(n7775), .A2(n7774), .ZN(n7794) );
  NOR2_X1 U8451 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U8452 ( .A1(n11120), .A2(n7244), .ZN(n7726) );
  NAND2_X1 U8453 ( .A1(n6926), .A2(n7724), .ZN(n7735) );
  XNOR2_X1 U8454 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7723) );
  AND2_X1 U8455 ( .A1(n8438), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7722) );
  INV_X1 U8456 ( .A(n10071), .ZN(n7338) );
  INV_X1 U8457 ( .A(n13464), .ZN(n13640) );
  OR2_X1 U8458 ( .A1(n11004), .A2(n11005), .ZN(n7335) );
  AND2_X1 U8459 ( .A1(n8696), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8718) );
  XNOR2_X1 U8460 ( .A(n13920), .B(n13338), .ZN(n6611) );
  NAND2_X1 U8461 ( .A1(n6611), .A2(n13322), .ZN(n13323) );
  NAND2_X1 U8462 ( .A1(n13320), .A2(n7330), .ZN(n7329) );
  INV_X1 U8463 ( .A(n13321), .ZN(n7330) );
  OR2_X1 U8464 ( .A1(n13454), .A2(n13453), .ZN(n7328) );
  INV_X1 U8465 ( .A(n13347), .ZN(n7344) );
  NAND2_X1 U8466 ( .A1(n8718), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8753) );
  INV_X1 U8467 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11435) );
  OAI22_X1 U8468 ( .A1(n11819), .A2(n6523), .B1(n6824), .B2(n6444), .ZN(n13406) );
  AOI21_X1 U8469 ( .B1(n6827), .B2(n6826), .A(n6825), .ZN(n6824) );
  INV_X1 U8470 ( .A(n13311), .ZN(n6825) );
  NAND2_X1 U8471 ( .A1(n13406), .A2(n13407), .ZN(n13405) );
  NAND2_X1 U8472 ( .A1(n13333), .A2(n13334), .ZN(n7656) );
  NOR2_X1 U8473 ( .A1(n9022), .A2(n13431), .ZN(n9046) );
  NAND2_X1 U8474 ( .A1(n10725), .A2(n10724), .ZN(n11003) );
  OR2_X1 U8475 ( .A1(n8655), .A2(n8654), .ZN(n8674) );
  NOR2_X1 U8476 ( .A1(n8674), .A2(n10729), .ZN(n8696) );
  INV_X1 U8477 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10729) );
  OR2_X1 U8478 ( .A1(n8753), .A2(n11435), .ZN(n8775) );
  NAND2_X1 U8479 ( .A1(n8958), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8984) );
  AND2_X1 U8480 ( .A1(n9633), .A2(n9247), .ZN(n13570) );
  XNOR2_X1 U8481 ( .A(n10334), .B(n9828), .ZN(n10261) );
  INV_X1 U8482 ( .A(n8819), .ZN(n8818) );
  AND2_X1 U8483 ( .A1(n9633), .A2(n9248), .ZN(n13464) );
  INV_X1 U8485 ( .A(n9160), .ZN(n9114) );
  NAND3_X1 U8486 ( .A1(n8437), .A2(n8436), .A3(n8435), .ZN(n9211) );
  AND2_X1 U8487 ( .A1(n8433), .A2(n8432), .ZN(n8437) );
  AND2_X1 U8488 ( .A1(n6896), .A2(n6894), .ZN(n9813) );
  NAND2_X1 U8489 ( .A1(n6896), .A2(n6496), .ZN(n9907) );
  OR2_X1 U8490 ( .A1(n9910), .A2(n9909), .ZN(n6893) );
  AND2_X1 U8491 ( .A1(n6893), .A2(n6892), .ZN(n9997) );
  NAND2_X1 U8492 ( .A1(n9994), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8493 ( .A1(n9997), .A2(n9996), .ZN(n10176) );
  AOI21_X1 U8494 ( .B1(n10176), .B2(n10174), .A(n10175), .ZN(n11259) );
  NOR2_X1 U8495 ( .A1(n13565), .A2(n7121), .ZN(n7120) );
  INV_X1 U8496 ( .A(n7122), .ZN(n7121) );
  AND2_X1 U8497 ( .A1(n13670), .A2(n7122), .ZN(n13641) );
  AND2_X1 U8498 ( .A1(n6914), .A2(n7302), .ZN(n6913) );
  AOI21_X1 U8499 ( .B1(n7305), .B2(n7303), .A(n6500), .ZN(n7302) );
  AND2_X1 U8500 ( .A1(n9135), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13642) );
  NAND2_X1 U8501 ( .A1(n13670), .A2(n13357), .ZN(n13671) );
  NOR2_X1 U8502 ( .A1(n13678), .A2(n7306), .ZN(n7305) );
  INV_X1 U8503 ( .A(n13601), .ZN(n7306) );
  NAND2_X1 U8504 ( .A1(n7632), .A2(n7631), .ZN(n13666) );
  AOI21_X1 U8505 ( .B1(n7634), .B2(n6440), .A(n6472), .ZN(n7631) );
  NAND2_X1 U8506 ( .A1(n6730), .A2(n13624), .ZN(n13715) );
  NAND2_X1 U8507 ( .A1(n7012), .A2(n6734), .ZN(n6730) );
  NOR2_X1 U8508 ( .A1(n6726), .A2(n13622), .ZN(n6734) );
  INV_X1 U8509 ( .A(n7011), .ZN(n6726) );
  AOI21_X1 U8510 ( .B1(n7290), .B2(n7292), .A(n7289), .ZN(n7288) );
  NAND2_X1 U8511 ( .A1(n13810), .A2(n7290), .ZN(n7287) );
  INV_X1 U8512 ( .A(n13586), .ZN(n7289) );
  NAND2_X1 U8513 ( .A1(n6738), .A2(n6736), .ZN(n13805) );
  AOI21_X1 U8514 ( .B1(n6739), .B2(n11688), .A(n6737), .ZN(n6736) );
  INV_X1 U8515 ( .A(n7640), .ZN(n6737) );
  NAND2_X1 U8516 ( .A1(n11360), .A2(n7119), .ZN(n11689) );
  NAND2_X1 U8517 ( .A1(n6720), .A2(n11358), .ZN(n11668) );
  OAI21_X1 U8518 ( .B1(n10933), .B2(n7647), .A(n7644), .ZN(n6720) );
  AOI21_X1 U8519 ( .B1(n7648), .B2(n7646), .A(n7645), .ZN(n7644) );
  INV_X1 U8520 ( .A(n7648), .ZN(n7647) );
  NAND2_X1 U8521 ( .A1(n11360), .A2(n11359), .ZN(n11672) );
  AOI21_X1 U8522 ( .B1(n7293), .B2(n6909), .A(n6491), .ZN(n6908) );
  NOR2_X1 U8523 ( .A1(n10559), .A2(n10723), .ZN(n10697) );
  NAND2_X1 U8524 ( .A1(n7126), .A2(n7125), .ZN(n10559) );
  NAND2_X1 U8525 ( .A1(n10348), .A2(n10347), .ZN(n10350) );
  NAND2_X1 U8526 ( .A1(n10096), .A2(n10311), .ZN(n10338) );
  AND2_X1 U8527 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8583) );
  NAND2_X1 U8528 ( .A1(n9021), .A2(n9020), .ZN(n13888) );
  AND2_X1 U8529 ( .A1(n11345), .A2(n11344), .ZN(n11419) );
  AOI21_X1 U8530 ( .B1(n9606), .B2(n11807), .A(n14002), .ZN(n15167) );
  AOI21_X1 U8531 ( .B1(n8881), .B2(n8448), .A(n8447), .ZN(n8449) );
  AOI21_X1 U8532 ( .B1(n8446), .B2(n6989), .A(n7658), .ZN(n8447) );
  NAND2_X1 U8533 ( .A1(n8452), .A2(n6505), .ZN(n6744) );
  INV_X1 U8534 ( .A(n8450), .ZN(n6745) );
  OR2_X1 U8535 ( .A1(n9241), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U8536 ( .A1(n6578), .A2(n9235), .ZN(n9241) );
  OAI21_X1 U8537 ( .B1(n8468), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8470) );
  AND2_X1 U8538 ( .A1(n8421), .A2(n7347), .ZN(n7346) );
  NAND2_X1 U8539 ( .A1(n7650), .A2(n8421), .ZN(n8881) );
  OR2_X1 U8540 ( .A1(n8770), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8814) );
  OR2_X1 U8541 ( .A1(n8836), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8646) );
  INV_X1 U8542 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8438) );
  INV_X1 U8543 ( .A(n12388), .ZN(n6645) );
  AOI21_X1 U8544 ( .B1(n6638), .B2(n6636), .A(n7556), .ZN(n6635) );
  INV_X1 U8545 ( .A(n12271), .ZN(n6636) );
  INV_X1 U8546 ( .A(n7557), .ZN(n7556) );
  INV_X1 U8547 ( .A(n6638), .ZN(n6637) );
  NOR2_X1 U8548 ( .A1(n11773), .A2(n11772), .ZN(n11791) );
  AND2_X1 U8549 ( .A1(n7587), .A2(n10948), .ZN(n7035) );
  INV_X1 U8550 ( .A(n7585), .ZN(n7034) );
  AOI21_X1 U8551 ( .B1(n7587), .B2(n7586), .A(n6524), .ZN(n7585) );
  OR2_X1 U8552 ( .A1(n11477), .A2(n11476), .ZN(n11488) );
  NAND2_X1 U8553 ( .A1(n14106), .A2(n14107), .ZN(n14105) );
  NOR2_X1 U8554 ( .A1(n10828), .A2(n15349), .ZN(n10843) );
  AND2_X1 U8555 ( .A1(n10843), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11329) );
  OAI21_X1 U8556 ( .B1(n6630), .B2(n6631), .A(n6628), .ZN(n6627) );
  INV_X1 U8557 ( .A(n14061), .ZN(n6628) );
  NAND2_X1 U8558 ( .A1(n14136), .A2(n14137), .ZN(n14135) );
  AND4_X1 U8559 ( .A1(n11494), .A2(n11493), .A3(n11492), .A4(n11491), .ZN(
        n12306) );
  NOR2_X1 U8560 ( .A1(n14576), .A2(n14363), .ZN(n14353) );
  NAND2_X1 U8561 ( .A1(n14404), .A2(n14668), .ZN(n14384) );
  AND2_X1 U8562 ( .A1(n7284), .A2(n6832), .ZN(n14404) );
  INV_X1 U8563 ( .A(n7284), .ZN(n14419) );
  NAND2_X1 U8564 ( .A1(n7401), .A2(n7402), .ZN(n14395) );
  AND2_X1 U8565 ( .A1(n11984), .A2(n11905), .ZN(n12032) );
  NAND2_X1 U8566 ( .A1(n6437), .A2(n14647), .ZN(n14531) );
  INV_X1 U8567 ( .A(n7281), .ZN(n11799) );
  NAND3_X1 U8568 ( .A1(n10880), .A2(n6443), .A3(n7282), .ZN(n11770) );
  NAND2_X1 U8569 ( .A1(n10880), .A2(n6841), .ZN(n11537) );
  NAND2_X1 U8570 ( .A1(n10880), .A2(n10842), .ZN(n11327) );
  AOI21_X1 U8571 ( .B1(n6439), .B2(n6855), .A(n6515), .ZN(n6853) );
  NAND2_X1 U8572 ( .A1(n10819), .A2(n10818), .ZN(n10875) );
  NAND2_X1 U8573 ( .A1(n10495), .A2(n10494), .ZN(n10744) );
  NAND2_X1 U8574 ( .A1(n7404), .A2(n7406), .ZN(n7133) );
  NOR2_X1 U8575 ( .A1(n10249), .A2(n7405), .ZN(n7404) );
  INV_X1 U8576 ( .A(n12118), .ZN(n7405) );
  NAND2_X1 U8577 ( .A1(n6834), .A2(n6833), .ZN(n10273) );
  INV_X1 U8578 ( .A(n10462), .ZN(n6834) );
  AND2_X1 U8579 ( .A1(n7273), .A2(n15001), .ZN(n10463) );
  NAND2_X1 U8580 ( .A1(n15001), .A2(n10515), .ZN(n10206) );
  NAND2_X1 U8581 ( .A1(n9957), .A2(n9956), .ZN(n10195) );
  NAND2_X1 U8582 ( .A1(n9757), .A2(n15006), .ZN(n14998) );
  NAND2_X1 U8583 ( .A1(n14998), .A2(n7066), .ZN(n12106) );
  OR2_X1 U8584 ( .A1(n9757), .A2(n15006), .ZN(n7066) );
  NOR2_X1 U8585 ( .A1(n7138), .A2(n7137), .ZN(n14380) );
  NOR2_X1 U8586 ( .A1(n7388), .A2(n6438), .ZN(n14454) );
  INV_X1 U8587 ( .A(n7390), .ZN(n7388) );
  INV_X1 U8588 ( .A(n14463), .ZN(n14476) );
  INV_X1 U8589 ( .A(n10242), .ZN(n15068) );
  NAND2_X1 U8590 ( .A1(n12075), .A2(n9713), .ZN(n15072) );
  XNOR2_X1 U8591 ( .A(n9127), .B(n9126), .ZN(n11892) );
  OAI21_X1 U8592 ( .B1(n9132), .B2(n7488), .A(n7485), .ZN(n9127) );
  XNOR2_X1 U8593 ( .A(n9132), .B(n9131), .ZN(n13987) );
  NAND2_X1 U8594 ( .A1(n7442), .A2(n7443), .ZN(n9109) );
  XNOR2_X1 U8595 ( .A(n9277), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U8596 ( .A1(n7275), .A2(n7276), .ZN(n9364) );
  AND2_X1 U8597 ( .A1(n9360), .A2(n9359), .ZN(n9755) );
  INV_X1 U8598 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9355) );
  AND2_X1 U8599 ( .A1(n6478), .A2(n7435), .ZN(n7434) );
  INV_X1 U8600 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7435) );
  XNOR2_X1 U8601 ( .A(n6612), .B(n8905), .ZN(n11961) );
  NAND2_X1 U8602 ( .A1(n6613), .A2(n8902), .ZN(n6612) );
  NAND2_X1 U8603 ( .A1(n7473), .A2(n7478), .ZN(n8810) );
  AND2_X1 U8604 ( .A1(n10061), .A2(n9901), .ZN(n11473) );
  OAI21_X1 U8605 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8764) );
  NAND2_X1 U8606 ( .A1(n7454), .A2(n8668), .ZN(n8690) );
  NAND2_X1 U8607 ( .A1(n8666), .A2(n8665), .ZN(n7454) );
  AND2_X1 U8608 ( .A1(n7097), .A2(n7096), .ZN(n8642) );
  NAND2_X1 U8609 ( .A1(n9281), .A2(n7591), .ZN(n9298) );
  AND2_X1 U8610 ( .A1(n9263), .A2(n7272), .ZN(n7591) );
  NAND2_X1 U8611 ( .A1(n7356), .A2(n7354), .ZN(n14762) );
  NAND2_X1 U8612 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7355), .ZN(n7354) );
  NAND2_X1 U8613 ( .A1(n14763), .A2(n6756), .ZN(n7356) );
  INV_X1 U8614 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7355) );
  XNOR2_X1 U8615 ( .A(n14717), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14768) );
  NOR2_X1 U8616 ( .A1(n14772), .A2(n14773), .ZN(n14776) );
  NAND2_X1 U8617 ( .A1(n6757), .A2(n14780), .ZN(n14782) );
  NAND2_X1 U8618 ( .A1(n14815), .A2(n14814), .ZN(n6757) );
  INV_X1 U8619 ( .A(n7107), .ZN(n14777) );
  INV_X1 U8620 ( .A(n6772), .ZN(n14788) );
  OAI21_X1 U8621 ( .B1(n14816), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6473), .ZN(
        n6772) );
  OAI21_X1 U8622 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14734), .A(n14733), .ZN(
        n14794) );
  NAND2_X1 U8623 ( .A1(n7348), .A2(n7113), .ZN(n7109) );
  INV_X1 U8624 ( .A(n7111), .ZN(n7110) );
  OAI21_X1 U8625 ( .B1(n7114), .B2(n7112), .A(n14957), .ZN(n7111) );
  INV_X1 U8626 ( .A(n6765), .ZN(n6762) );
  AOI21_X1 U8627 ( .B1(n7103), .B2(n6766), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n6765) );
  NAND2_X1 U8628 ( .A1(n12502), .A2(n7158), .ZN(n7155) );
  NAND2_X1 U8629 ( .A1(n8080), .A2(n8079), .ZN(n12974) );
  NAND2_X1 U8630 ( .A1(n10427), .A2(n10425), .ZN(n10578) );
  NAND2_X1 U8631 ( .A1(n12606), .A2(n12497), .ZN(n12551) );
  NAND2_X1 U8632 ( .A1(n7173), .A2(n12507), .ZN(n12569) );
  NAND2_X1 U8633 ( .A1(n12608), .A2(n12607), .ZN(n12606) );
  INV_X1 U8634 ( .A(n12682), .ZN(n13049) );
  NAND2_X1 U8635 ( .A1(n12587), .A2(n12489), .ZN(n12647) );
  INV_X1 U8636 ( .A(n12659), .ZN(n12668) );
  OR2_X1 U8637 ( .A1(n10589), .A2(n10404), .ZN(n12666) );
  INV_X1 U8638 ( .A(n7162), .ZN(n12653) );
  AOI21_X1 U8639 ( .B1(n7173), .B2(n7164), .A(n7163), .ZN(n7162) );
  INV_X1 U8640 ( .A(n7171), .ZN(n7164) );
  INV_X1 U8641 ( .A(n7169), .ZN(n7163) );
  NAND2_X1 U8642 ( .A1(n12479), .A2(n12478), .ZN(n12664) );
  NAND2_X1 U8643 ( .A1(n7147), .A2(n7146), .ZN(n12479) );
  INV_X1 U8644 ( .A(n12652), .ZN(n12672) );
  AND2_X1 U8645 ( .A1(n8202), .A2(n8174), .ZN(n12907) );
  NAND2_X1 U8646 ( .A1(n8132), .A2(n8131), .ZN(n12678) );
  INV_X1 U8647 ( .A(n12978), .ZN(n12527) );
  OAI211_X1 U8648 ( .C1(n8184), .C2(n13251), .A(n8086), .B(n8085), .ZN(n12988)
         );
  INV_X1 U8649 ( .A(n13028), .ZN(n12681) );
  INV_X1 U8650 ( .A(n13059), .ZN(n12683) );
  OR2_X1 U8651 ( .A1(n8184), .A2(n7705), .ZN(n7707) );
  NAND4_X1 U8652 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n13213)
         );
  OR2_X1 U8653 ( .A1(n8060), .A2(n11084), .ZN(n7689) );
  AND2_X1 U8654 ( .A1(n6788), .A2(n6787), .ZN(n11576) );
  INV_X1 U8655 ( .A(n11294), .ZN(n6788) );
  NAND2_X1 U8656 ( .A1(n11618), .A2(n11295), .ZN(n6787) );
  NAND2_X1 U8657 ( .A1(n7382), .A2(n11245), .ZN(n11585) );
  NAND2_X1 U8658 ( .A1(n6786), .A2(n6785), .ZN(n11581) );
  NAND2_X1 U8659 ( .A1(n6782), .A2(n6783), .ZN(n11255) );
  NAND2_X1 U8660 ( .A1(n11127), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n12723) );
  AOI21_X1 U8661 ( .B1(n12730), .B2(n11171), .A(n6992), .ZN(n12734) );
  INV_X1 U8662 ( .A(n6594), .ZN(n6992) );
  INV_X1 U8663 ( .A(n6708), .ZN(n11197) );
  AOI21_X1 U8664 ( .B1(n11192), .B2(n11191), .A(n11190), .ZN(n11384) );
  INV_X1 U8665 ( .A(n6994), .ZN(n11200) );
  INV_X1 U8666 ( .A(n7263), .ZN(n11387) );
  INV_X1 U8667 ( .A(n7371), .ZN(n11180) );
  INV_X1 U8668 ( .A(n7365), .ZN(n11392) );
  INV_X1 U8669 ( .A(n6983), .ZN(n11721) );
  NOR2_X1 U8670 ( .A1(n11710), .A2(n6808), .ZN(n11713) );
  AND2_X1 U8671 ( .A1(n11711), .A2(n11717), .ZN(n6808) );
  NAND2_X1 U8672 ( .A1(n11713), .A2(n11712), .ZN(n12743) );
  INV_X1 U8673 ( .A(n12752), .ZN(n12751) );
  INV_X1 U8674 ( .A(n6710), .ZN(n11708) );
  NAND2_X1 U8675 ( .A1(n12743), .A2(n6805), .ZN(n12770) );
  NOR2_X1 U8676 ( .A1(n6807), .A2(n6806), .ZN(n6805) );
  INV_X1 U8677 ( .A(n12742), .ZN(n6806) );
  INV_X1 U8678 ( .A(n12741), .ZN(n6807) );
  NAND2_X1 U8679 ( .A1(n6712), .A2(n12787), .ZN(n12789) );
  INV_X1 U8680 ( .A(n6660), .ZN(n12831) );
  AND2_X1 U8681 ( .A1(n7260), .A2(n12787), .ZN(n12807) );
  NOR2_X1 U8682 ( .A1(n12808), .A2(n6981), .ZN(n12838) );
  INV_X1 U8683 ( .A(n12881), .ZN(n12859) );
  NAND2_X1 U8684 ( .A1(n8168), .A2(n8167), .ZN(n13133) );
  NAND2_X1 U8685 ( .A1(n7214), .A2(n7217), .ZN(n12460) );
  NAND2_X1 U8686 ( .A1(n13145), .A2(n15201), .ZN(n12923) );
  NAND2_X1 U8687 ( .A1(n12966), .A2(n8356), .ZN(n12953) );
  NAND2_X1 U8688 ( .A1(n8055), .A2(n8054), .ZN(n13170) );
  NAND2_X1 U8689 ( .A1(n13040), .A2(n8322), .ZN(n13037) );
  NAND2_X1 U8690 ( .A1(n13096), .A2(n12431), .ZN(n13083) );
  NAND2_X1 U8691 ( .A1(n7196), .A2(n7200), .ZN(n13088) );
  NAND2_X1 U8692 ( .A1(n13115), .A2(n7203), .ZN(n7196) );
  NAND2_X1 U8693 ( .A1(n7204), .A2(n7203), .ZN(n13111) );
  NAND2_X1 U8694 ( .A1(n7204), .A2(n8215), .ZN(n13109) );
  NAND2_X1 U8695 ( .A1(n15248), .A2(n14860), .ZN(n13125) );
  NAND2_X1 U8696 ( .A1(n12428), .A2(n12427), .ZN(n13117) );
  INV_X1 U8697 ( .A(n13107), .ZN(n15206) );
  NAND2_X1 U8698 ( .A1(n7189), .A2(n7190), .ZN(n11595) );
  AND3_X1 U8699 ( .A1(n7858), .A2(n7857), .A3(n7856), .ZN(n12421) );
  NAND2_X1 U8700 ( .A1(n7192), .A2(n8273), .ZN(n11037) );
  NAND2_X1 U8701 ( .A1(n11304), .A2(n11441), .ZN(n7192) );
  AND2_X1 U8702 ( .A1(n10417), .A2(n12878), .ZN(n15232) );
  INV_X1 U8703 ( .A(n15234), .ZN(n15244) );
  NOR2_X1 U8704 ( .A1(n10917), .A2(n15281), .ZN(n13107) );
  AND2_X2 U8705 ( .A1(n10657), .A2(n10623), .ZN(n15308) );
  NAND2_X1 U8706 ( .A1(n15308), .A2(n15287), .ZN(n13210) );
  NAND2_X1 U8707 ( .A1(n8193), .A2(n8192), .ZN(n13229) );
  INV_X1 U8708 ( .A(n12621), .ZN(n13293) );
  AND2_X1 U8709 ( .A1(n11073), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13295) );
  INV_X1 U8710 ( .A(n13295), .ZN(n11882) );
  AOI21_X1 U8711 ( .B1(n7269), .B2(n7267), .A(n6595), .ZN(n7266) );
  INV_X1 U8712 ( .A(n7686), .ZN(n12417) );
  MUX2_X1 U8713 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8393), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8394) );
  NAND2_X1 U8714 ( .A1(n8398), .A2(n8397), .ZN(n10908) );
  NAND2_X1 U8715 ( .A1(n8106), .A2(n8093), .ZN(n8105) );
  NAND2_X1 U8716 ( .A1(n7254), .A2(n8067), .ZN(n8078) );
  NAND2_X1 U8717 ( .A1(n8066), .A2(n8065), .ZN(n7254) );
  INV_X1 U8718 ( .A(n10777), .ZN(n10615) );
  XNOR2_X1 U8719 ( .A(n8210), .B(n8209), .ZN(n10416) );
  INV_X1 U8720 ( .A(n10617), .ZN(n10417) );
  NAND2_X1 U8721 ( .A1(n6936), .A2(n6940), .ZN(n8042) );
  OR2_X1 U8722 ( .A1(n8006), .A2(n6942), .ZN(n6936) );
  NAND2_X1 U8723 ( .A1(n7248), .A2(n7984), .ZN(n8002) );
  INV_X1 U8724 ( .A(SI_16_), .ZN(n9655) );
  INV_X1 U8725 ( .A(SI_15_), .ZN(n9604) );
  NAND2_X1 U8726 ( .A1(n6933), .A2(n7271), .ZN(n7948) );
  NAND2_X1 U8727 ( .A1(n6934), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6933) );
  INV_X1 U8728 ( .A(SI_13_), .ZN(n9375) );
  NAND2_X1 U8729 ( .A1(n6934), .A2(n7271), .ZN(n7936) );
  XNOR2_X1 U8730 ( .A(n7925), .B(n7924), .ZN(n12771) );
  INV_X1 U8731 ( .A(SI_12_), .ZN(n9322) );
  INV_X1 U8732 ( .A(SI_11_), .ZN(n9304) );
  OR2_X1 U8733 ( .A1(n7874), .A2(n7873), .ZN(n11393) );
  OAI21_X1 U8734 ( .B1(n7849), .B2(n7237), .A(n7235), .ZN(n7886) );
  NAND2_X1 U8735 ( .A1(n7866), .A2(n7865), .ZN(n7869) );
  NAND2_X1 U8736 ( .A1(n7826), .A2(n7825), .ZN(n7829) );
  NAND2_X1 U8737 ( .A1(n7808), .A2(n7807), .ZN(n7811) );
  OR2_X1 U8738 ( .A1(n7781), .A2(n7780), .ZN(n11222) );
  NAND2_X1 U8739 ( .A1(n7759), .A2(n7760), .ZN(n11258) );
  OAI211_X1 U8740 ( .C1(n11120), .C2(n7370), .A(n7726), .B(n7243), .ZN(n11299)
         );
  NAND2_X1 U8741 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7370) );
  NAND2_X1 U8742 ( .A1(n13298), .A2(n7244), .ZN(n7243) );
  NAND2_X1 U8743 ( .A1(n6665), .A2(n6662), .ZN(n11629) );
  NAND2_X1 U8744 ( .A1(n6664), .A2(n6663), .ZN(n6662) );
  OAI21_X1 U8745 ( .B1(n10072), .B2(n7337), .A(n7336), .ZN(n10434) );
  NAND2_X1 U8746 ( .A1(n7339), .A2(n7340), .ZN(n7336) );
  NAND2_X1 U8747 ( .A1(n7338), .A2(n7340), .ZN(n7337) );
  NAND2_X1 U8748 ( .A1(n10261), .A2(n10262), .ZN(n7340) );
  NAND2_X1 U8749 ( .A1(n13351), .A2(n13350), .ZN(n6979) );
  NAND2_X1 U8750 ( .A1(n13460), .A2(n6436), .ZN(n13375) );
  AND2_X1 U8751 ( .A1(n11003), .A2(n7333), .ZN(n11407) );
  NAND2_X1 U8752 ( .A1(n13323), .A2(n6610), .ZN(n13368) );
  OR2_X1 U8753 ( .A1(n6611), .A2(n13322), .ZN(n6610) );
  NAND2_X1 U8754 ( .A1(n7328), .A2(n7329), .ZN(n13369) );
  NAND2_X1 U8755 ( .A1(n7320), .A2(n6617), .ZN(n13389) );
  AOI21_X1 U8756 ( .B1(n7324), .B2(n7322), .A(n7321), .ZN(n7320) );
  INV_X1 U8757 ( .A(n13436), .ZN(n7321) );
  NOR2_X1 U8758 ( .A1(n10072), .A2(n10071), .ZN(n10140) );
  NAND2_X1 U8759 ( .A1(n13428), .A2(n13427), .ZN(n13426) );
  NAND2_X1 U8760 ( .A1(n7656), .A2(n13361), .ZN(n13428) );
  NOR2_X1 U8761 ( .A1(n9929), .A2(n9928), .ZN(n10068) );
  NOR2_X1 U8762 ( .A1(n9667), .A2(n6507), .ZN(n9648) );
  NAND2_X1 U8763 ( .A1(n7319), .A2(n7324), .ZN(n13438) );
  NAND2_X1 U8764 ( .A1(n13454), .A2(n7326), .ZN(n7319) );
  XNOR2_X1 U8765 ( .A(n13329), .B(n13328), .ZN(n13446) );
  NAND2_X1 U8766 ( .A1(n13446), .A2(n13445), .ZN(n13444) );
  NAND2_X1 U8767 ( .A1(n6821), .A2(n7333), .ZN(n6820) );
  NAND2_X1 U8768 ( .A1(n6821), .A2(n6823), .ZN(n6819) );
  INV_X1 U8769 ( .A(n11409), .ZN(n6821) );
  AOI21_X1 U8770 ( .B1(n6822), .B2(n7333), .A(n6823), .ZN(n11408) );
  INV_X1 U8771 ( .A(n10725), .ZN(n6822) );
  AOI21_X1 U8772 ( .B1(n9682), .B2(n9681), .A(n9825), .ZN(n9689) );
  NAND2_X1 U8773 ( .A1(n13416), .A2(n13319), .ZN(n13454) );
  NAND2_X1 U8774 ( .A1(n13398), .A2(n13342), .ZN(n13462) );
  AOI21_X1 U8775 ( .B1(n7492), .B2(n9195), .A(n9201), .ZN(n9202) );
  OR2_X1 U8776 ( .A1(n9094), .A2(n8537), .ZN(n8539) );
  OR2_X1 U8777 ( .A1(n8962), .A2(n8476), .ZN(n8479) );
  CLKBUF_X1 U8778 ( .A(n9211), .Z(n13491) );
  NAND2_X1 U8779 ( .A1(n6883), .A2(n9402), .ZN(n9436) );
  OR2_X1 U8780 ( .A1(n9593), .A2(n9433), .ZN(n6883) );
  NAND2_X1 U8781 ( .A1(n6896), .A2(n6897), .ZN(n9805) );
  INV_X1 U8782 ( .A(n6893), .ZN(n9993) );
  XNOR2_X1 U8783 ( .A(n11261), .B(n11273), .ZN(n13526) );
  NAND2_X1 U8784 ( .A1(n15157), .A2(n11264), .ZN(n11268) );
  NAND2_X1 U8785 ( .A1(n11268), .A2(n11267), .ZN(n11506) );
  NAND2_X1 U8786 ( .A1(n11506), .A2(n6882), .ZN(n11507) );
  OR2_X1 U8787 ( .A1(n11511), .A2(n11858), .ZN(n6882) );
  NAND2_X1 U8788 ( .A1(n11507), .A2(n11508), .ZN(n13532) );
  NOR2_X1 U8789 ( .A1(n6888), .A2(n13546), .ZN(n13547) );
  NAND2_X1 U8790 ( .A1(n6887), .A2(n6890), .ZN(n13534) );
  AND2_X1 U8791 ( .A1(n6888), .A2(n6887), .ZN(n13548) );
  AND2_X1 U8792 ( .A1(n7639), .A2(n6592), .ZN(n7638) );
  XNOR2_X1 U8793 ( .A(n7008), .B(n7007), .ZN(n13637) );
  NAND2_X1 U8794 ( .A1(n7307), .A2(n13601), .ZN(n13679) );
  NAND2_X1 U8795 ( .A1(n7307), .A2(n7305), .ZN(n13873) );
  INV_X1 U8796 ( .A(n7633), .ZN(n13682) );
  AOI21_X1 U8797 ( .B1(n13697), .B2(n13628), .A(n6440), .ZN(n7633) );
  NAND2_X1 U8798 ( .A1(n7012), .A2(n7011), .ZN(n13739) );
  NAND2_X1 U8799 ( .A1(n13751), .A2(n13593), .ZN(n13729) );
  NAND2_X1 U8800 ( .A1(n7013), .A2(n7020), .ZN(n13745) );
  NAND2_X1 U8801 ( .A1(n7635), .A2(n7018), .ZN(n7013) );
  NAND2_X1 U8802 ( .A1(n7635), .A2(n13617), .ZN(n13769) );
  NAND2_X1 U8803 ( .A1(n8936), .A2(n8935), .ZN(n13915) );
  NAND2_X1 U8804 ( .A1(n13808), .A2(n13584), .ZN(n13791) );
  NAND2_X1 U8805 ( .A1(n8884), .A2(n8883), .ZN(n13925) );
  NAND2_X1 U8806 ( .A1(n13580), .A2(n13579), .ZN(n13833) );
  NAND2_X1 U8807 ( .A1(n7643), .A2(n13608), .ZN(n13820) );
  NAND2_X1 U8808 ( .A1(n13605), .A2(n13604), .ZN(n7643) );
  NAND2_X1 U8809 ( .A1(n11865), .A2(n7301), .ZN(n13580) );
  NAND2_X1 U8810 ( .A1(n11865), .A2(n11864), .ZN(n11867) );
  NAND2_X1 U8811 ( .A1(n8840), .A2(n8839), .ZN(n13607) );
  NAND2_X1 U8812 ( .A1(n11697), .A2(n11696), .ZN(n11853) );
  NAND2_X1 U8813 ( .A1(n6910), .A2(n7293), .ZN(n10702) );
  NAND2_X1 U8814 ( .A1(n10547), .A2(n10546), .ZN(n10549) );
  NAND2_X1 U8815 ( .A1(n10348), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U8816 ( .A1(n7652), .A2(n10553), .ZN(n10555) );
  NAND2_X1 U8817 ( .A1(n10356), .A2(n10355), .ZN(n10550) );
  NAND2_X1 U8818 ( .A1(n6748), .A2(n7004), .ZN(n10353) );
  NAND2_X1 U8819 ( .A1(n7006), .A2(n10102), .ZN(n10332) );
  NAND2_X1 U8820 ( .A1(n10100), .A2(n10099), .ZN(n7006) );
  NAND2_X1 U8821 ( .A1(n13844), .A2(n10309), .ZN(n13816) );
  AOI22_X1 U8822 ( .A1(n8907), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8906), .B2(
        n13505), .ZN(n6996) );
  NAND2_X1 U8823 ( .A1(n10111), .A2(n8786), .ZN(n6997) );
  OR2_X1 U8824 ( .A1(n8749), .A2(n9313), .ZN(n8487) );
  INV_X1 U8825 ( .A(n13850), .ZN(n13766) );
  INV_X1 U8826 ( .A(n13835), .ZN(n13848) );
  NAND2_X1 U8827 ( .A1(n9629), .A2(n15176), .ZN(n13841) );
  NAND2_X1 U8828 ( .A1(n8695), .A2(n8694), .ZN(n11010) );
  INV_X1 U8829 ( .A(n13912), .ZN(n13899) );
  AND2_X2 U8830 ( .A1(n9660), .A2(n9767), .ZN(n15190) );
  INV_X1 U8831 ( .A(n13866), .ZN(n6754) );
  NOR2_X1 U8832 ( .A1(n13868), .A2(n15182), .ZN(n6753) );
  INV_X1 U8833 ( .A(n13753), .ZN(n13970) );
  NAND2_X1 U8834 ( .A1(n8817), .A2(n8816), .ZN(n11863) );
  NAND2_X1 U8835 ( .A1(n8717), .A2(n8716), .ZN(n11412) );
  INV_X1 U8836 ( .A(n10684), .ZN(n10057) );
  AOI22_X1 U8837 ( .A1(n8907), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9415), .B2(
        n8906), .ZN(n6990) );
  INV_X1 U8838 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8426) );
  INV_X1 U8839 ( .A(n8431), .ZN(n13986) );
  NAND2_X1 U8840 ( .A1(n6744), .A2(n8449), .ZN(n13996) );
  INV_X1 U8841 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U8842 ( .A1(n8468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8455) );
  INV_X1 U8843 ( .A(n8466), .ZN(n11035) );
  INV_X1 U8844 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10811) );
  INV_X1 U8845 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10534) );
  INV_X1 U8846 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10296) );
  INV_X1 U8847 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10213) );
  INV_X1 U8848 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9764) );
  OR2_X1 U8849 ( .A1(n8748), .A2(n8747), .ZN(n11270) );
  INV_X1 U8850 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9566) );
  INV_X1 U8851 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9468) );
  INV_X1 U8852 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9382) );
  INV_X1 U8853 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9354) );
  INV_X1 U8854 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9349) );
  INV_X1 U8855 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9324) );
  INV_X1 U8856 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9311) );
  INV_X1 U8857 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9297) );
  INV_X1 U8858 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9287) );
  INV_X1 U8859 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9279) );
  INV_X1 U8860 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9313) );
  OAI211_X1 U8861 ( .C1(P2_IR_REG_31__SCAN_IN), .C2(P2_IR_REG_1__SCAN_IN), .A(
        n6903), .B(n8505), .ZN(n9453) );
  NAND2_X1 U8862 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6904), .ZN(n6903) );
  NOR2_X1 U8863 ( .A1(n8483), .A2(n8484), .ZN(n6904) );
  NAND2_X1 U8864 ( .A1(n14893), .A2(n12311), .ZN(n14894) );
  AND2_X1 U8865 ( .A1(n14895), .A2(n14892), .ZN(n12311) );
  NAND2_X1 U8866 ( .A1(n14105), .A2(n12369), .ZN(n14011) );
  OAI21_X1 U8867 ( .B1(n10038), .B2(n7579), .A(n7578), .ZN(n10123) );
  NAND2_X1 U8868 ( .A1(n7033), .A2(n12344), .ZN(n14019) );
  NAND2_X1 U8869 ( .A1(n7033), .A2(n7031), .ZN(n14020) );
  AND2_X1 U8870 ( .A1(n7572), .A2(n7569), .ZN(n7562) );
  NAND2_X1 U8871 ( .A1(n12408), .A2(n7566), .ZN(n7565) );
  INV_X1 U8872 ( .A(n7569), .ZN(n7566) );
  NAND2_X1 U8873 ( .A1(n7568), .A2(n12408), .ZN(n7567) );
  AND2_X1 U8874 ( .A1(n14318), .A2(n11916), .ZN(n14330) );
  NAND2_X1 U8875 ( .A1(n11058), .A2(n7588), .ZN(n11061) );
  INV_X1 U8876 ( .A(n9863), .ZN(n9864) );
  NAND2_X1 U8877 ( .A1(n14088), .A2(n12354), .ZN(n14028) );
  NAND2_X1 U8878 ( .A1(n7553), .A2(n7557), .ZN(n14038) );
  NAND2_X1 U8879 ( .A1(n14908), .A2(n7559), .ZN(n7553) );
  AOI21_X1 U8880 ( .B1(n7024), .B2(n7026), .A(n6510), .ZN(n7022) );
  NAND2_X1 U8881 ( .A1(n14135), .A2(n12321), .ZN(n14053) );
  AOI21_X1 U8882 ( .B1(n10633), .B2(n6631), .A(n6630), .ZN(n14064) );
  NAND2_X1 U8883 ( .A1(n6623), .A2(n6622), .ZN(n14073) );
  INV_X1 U8884 ( .A(n6624), .ZN(n6623) );
  OAI21_X1 U8885 ( .B1(n12321), .B2(n7583), .A(n12329), .ZN(n6624) );
  NAND2_X1 U8886 ( .A1(n7023), .A2(n7573), .ZN(n14081) );
  NAND2_X1 U8887 ( .A1(n14106), .A2(n7574), .ZN(n7023) );
  INV_X1 U8888 ( .A(n7552), .ZN(n7551) );
  AOI21_X1 U8889 ( .B1(n7031), .B2(n7029), .A(n6572), .ZN(n7028) );
  INV_X1 U8890 ( .A(n7031), .ZN(n7030) );
  NAND2_X1 U8891 ( .A1(n14036), .A2(n12298), .ZN(n14098) );
  NAND2_X1 U8892 ( .A1(n14906), .A2(n12286), .ZN(n14919) );
  INV_X1 U8893 ( .A(n10042), .ZN(n7580) );
  INV_X1 U8894 ( .A(n7581), .ZN(n10043) );
  NAND2_X1 U8895 ( .A1(n6632), .A2(n14060), .ZN(n10794) );
  NAND2_X1 U8896 ( .A1(n6629), .A2(n6626), .ZN(n6632) );
  INV_X1 U8897 ( .A(n6627), .ZN(n6626) );
  OR2_X1 U8898 ( .A1(n10633), .A2(n6630), .ZN(n6629) );
  INV_X1 U8899 ( .A(n14935), .ZN(n14113) );
  NAND2_X1 U8900 ( .A1(n12389), .A2(n12388), .ZN(n14125) );
  NAND2_X1 U8901 ( .A1(n11922), .A2(n11921), .ZN(n14583) );
  INV_X1 U8902 ( .A(n14133), .ZN(n14930) );
  NAND2_X1 U8903 ( .A1(n12240), .A2(n7042), .ZN(n12266) );
  NAND2_X1 U8904 ( .A1(n12239), .A2(n12238), .ZN(n7042) );
  OAI21_X1 U8905 ( .B1(n12239), .B2(n12238), .A(n12237), .ZN(n12240) );
  OR2_X1 U8906 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  NOR2_X1 U8907 ( .A1(n12243), .A2(n7088), .ZN(n12262) );
  NAND2_X1 U8908 ( .A1(n11974), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U8909 ( .A1(n12056), .A2(n12055), .ZN(n14389) );
  NAND2_X1 U8910 ( .A1(n6876), .A2(n7624), .ZN(n14377) );
  NAND2_X1 U8911 ( .A1(n14429), .A2(n6880), .ZN(n6876) );
  NAND2_X1 U8912 ( .A1(n14417), .A2(n7627), .ZN(n14392) );
  AND2_X1 U8913 ( .A1(n14417), .A2(n14277), .ZN(n14393) );
  NAND2_X1 U8914 ( .A1(n14412), .A2(n14416), .ZN(n14411) );
  NAND2_X1 U8915 ( .A1(n7129), .A2(n7130), .ZN(n14428) );
  NAND2_X1 U8916 ( .A1(n14458), .A2(n14272), .ZN(n14442) );
  NAND2_X1 U8917 ( .A1(n14453), .A2(n14298), .ZN(n14449) );
  NAND2_X1 U8918 ( .A1(n14270), .A2(n14269), .ZN(n14460) );
  NAND2_X1 U8919 ( .A1(n14295), .A2(n14294), .ZN(n14469) );
  NAND2_X1 U8920 ( .A1(n6871), .A2(n6873), .ZN(n14485) );
  NAND2_X1 U8921 ( .A1(n6872), .A2(n7600), .ZN(n6871) );
  INV_X1 U8922 ( .A(n14266), .ZN(n6872) );
  NAND2_X1 U8923 ( .A1(n7141), .A2(n14292), .ZN(n14505) );
  NAND2_X1 U8924 ( .A1(n14528), .A2(n14267), .ZN(n14502) );
  NAND2_X1 U8925 ( .A1(n14290), .A2(n14289), .ZN(n14522) );
  NAND2_X1 U8926 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  NAND2_X1 U8927 ( .A1(n11532), .A2(n11531), .ZN(n11530) );
  NAND2_X1 U8928 ( .A1(n11484), .A2(n11483), .ZN(n11532) );
  NAND2_X1 U8929 ( .A1(n10877), .A2(n10824), .ZN(n10835) );
  OAI21_X1 U8930 ( .B1(n10743), .B2(n6855), .A(n6439), .ZN(n10872) );
  NAND2_X1 U8931 ( .A1(n10838), .A2(n10837), .ZN(n10873) );
  NAND2_X1 U8932 ( .A1(n10460), .A2(n7607), .ZN(n7604) );
  NAND2_X1 U8933 ( .A1(n10231), .A2(n7607), .ZN(n7603) );
  NAND2_X1 U8934 ( .A1(n7609), .A2(n7607), .ZN(n10269) );
  NAND2_X1 U8935 ( .A1(n7610), .A2(n10459), .ZN(n7609) );
  NAND2_X1 U8936 ( .A1(n7406), .A2(n12118), .ZN(n10461) );
  AND2_X1 U8937 ( .A1(n10205), .A2(n10204), .ZN(n15018) );
  NAND2_X1 U8938 ( .A1(n10191), .A2(n10190), .ZN(n14544) );
  INV_X1 U8939 ( .A(n14520), .ZN(n14548) );
  INV_X2 U8940 ( .A(n14541), .ZN(n15022) );
  NAND2_X1 U8941 ( .A1(n11324), .A2(n11323), .ZN(n14547) );
  NAND2_X1 U8942 ( .A1(n10270), .A2(n6429), .ZN(n6866) );
  CLKBUF_X1 U8943 ( .A(n9971), .Z(n15123) );
  INV_X1 U8944 ( .A(n14251), .ZN(n14654) );
  INV_X1 U8945 ( .A(n14261), .ZN(n14659) );
  NAND2_X1 U8946 ( .A1(n14567), .A2(n15079), .ZN(n6845) );
  OAI21_X1 U8947 ( .B1(n14568), .B2(n15074), .A(n6844), .ZN(n6843) );
  INV_X1 U8948 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7395) );
  NAND2_X1 U8949 ( .A1(n7598), .A2(n7398), .ZN(n14661) );
  OR2_X1 U8950 ( .A1(n14574), .A2(n15074), .ZN(n7398) );
  AND2_X1 U8951 ( .A1(n14572), .A2(n14573), .ZN(n7598) );
  NOR2_X1 U8952 ( .A1(n14662), .A2(n14683), .ZN(n7396) );
  INV_X1 U8953 ( .A(n14389), .ZN(n14668) );
  AND2_X1 U8954 ( .A1(n11972), .A2(n11971), .ZN(n14679) );
  NOR2_X1 U8955 ( .A1(n10290), .A2(n10289), .ZN(n14655) );
  INV_X1 U8956 ( .A(n10045), .ZN(n10515) );
  OR2_X1 U8957 ( .A1(n9372), .A2(P1_U3086), .ZN(n9380) );
  NAND2_X1 U8958 ( .A1(n9124), .A2(n9088), .ZN(n14694) );
  NAND2_X1 U8959 ( .A1(n7491), .A2(n7489), .ZN(n9124) );
  NAND2_X1 U8960 ( .A1(n7491), .A2(n9084), .ZN(n9087) );
  NAND2_X1 U8961 ( .A1(n9725), .A2(n6469), .ZN(n6639) );
  NOR2_X1 U8962 ( .A1(n6642), .A2(n6641), .ZN(n6640) );
  AOI21_X1 U8963 ( .B1(n7041), .B2(n6468), .A(n7040), .ZN(n7039) );
  NOR2_X1 U8964 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n7040) );
  NAND2_X1 U8965 ( .A1(n7274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7590) );
  INV_X1 U8966 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12053) );
  XNOR2_X1 U8967 ( .A(n8996), .B(n8995), .ZN(n11941) );
  XNOR2_X1 U8968 ( .A(n9362), .B(P1_IR_REG_22__SCAN_IN), .ZN(n12072) );
  NAND2_X1 U8969 ( .A1(n9361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9362) );
  OR2_X1 U8970 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  INV_X1 U8971 ( .A(n9755), .ZN(n12075) );
  INV_X1 U8972 ( .A(n14433), .ZN(n14320) );
  INV_X1 U8973 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10814) );
  INV_X1 U8974 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n15443) );
  INV_X1 U8975 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10220) );
  INV_X1 U8976 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10063) );
  INV_X1 U8977 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9572) );
  INV_X1 U8978 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9465) );
  INV_X1 U8979 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9389) );
  INV_X1 U8980 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9351) );
  INV_X1 U8981 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9346) );
  INV_X1 U8982 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9329) );
  INV_X1 U8983 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9308) );
  INV_X1 U8984 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9300) );
  INV_X1 U8985 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10114) );
  INV_X1 U8986 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U8987 ( .A1(n7101), .A2(n14766), .ZN(n14811) );
  NAND2_X1 U8988 ( .A1(n15473), .A2(n15474), .ZN(n7101) );
  XNOR2_X1 U8989 ( .A(n14776), .B(n14775), .ZN(n15464) );
  XNOR2_X1 U8990 ( .A(n7107), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n14815) );
  XNOR2_X1 U8991 ( .A(n14782), .B(n7106), .ZN(n15467) );
  XNOR2_X1 U8992 ( .A(n14784), .B(n14785), .ZN(n14816) );
  XNOR2_X1 U8993 ( .A(n14788), .B(n7362), .ZN(n14817) );
  INV_X1 U8994 ( .A(n14789), .ZN(n7362) );
  INV_X1 U8995 ( .A(n7100), .ZN(n14947) );
  OAI21_X1 U8996 ( .B1(n14818), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6474), .ZN(
        n7100) );
  NAND2_X1 U8997 ( .A1(n6773), .A2(n7113), .ZN(n14958) );
  NAND2_X1 U8998 ( .A1(n14953), .A2(n7114), .ZN(n6773) );
  NOR2_X1 U8999 ( .A1(n14958), .A2(n14957), .ZN(n14956) );
  AOI21_X1 U9000 ( .B1(n14969), .B2(n14803), .A(n14966), .ZN(n14821) );
  OR2_X1 U9001 ( .A1(n10633), .A2(n10632), .ZN(n7550) );
  NAND2_X1 U9002 ( .A1(n10858), .A2(n10857), .ZN(n10865) );
  NAND2_X1 U9003 ( .A1(n7186), .A2(n10713), .ZN(n7228) );
  NAND2_X1 U9004 ( .A1(n6655), .A2(n6650), .ZN(P3_U3199) );
  NAND2_X1 U9005 ( .A1(n12834), .A2(n12835), .ZN(n6655) );
  INV_X1 U9006 ( .A(n6651), .ZN(n6650) );
  AOI21_X1 U9007 ( .B1(n7378), .B2(n12835), .A(n7376), .ZN(n12891) );
  OAI21_X1 U9008 ( .B1(n13239), .B2(n15295), .A(n6677), .ZN(P3_U3453) );
  INV_X1 U9009 ( .A(n6678), .ZN(n6677) );
  OAI22_X1 U9010 ( .A1(n13241), .A2(n13294), .B1(n15293), .B2(n13240), .ZN(
        n6678) );
  OAI21_X1 U9011 ( .B1(n11612), .B2(n11891), .A(n7184), .ZN(P3_U3268) );
  NOR2_X1 U9012 ( .A1(n11887), .A2(n11611), .ZN(n7185) );
  AND2_X1 U9013 ( .A1(n6829), .A2(n6464), .ZN(n14881) );
  NAND2_X1 U9014 ( .A1(n7636), .A2(n6587), .ZN(P2_U3528) );
  NAND2_X1 U9015 ( .A1(n13947), .A2(n15190), .ZN(n7636) );
  OAI21_X1 U9016 ( .B1(n13940), .B2(n15185), .A(n7115), .ZN(P2_U3498) );
  AOI21_X1 U9017 ( .B1(n9171), .B2(n13965), .A(n7116), .ZN(n7115) );
  NOR2_X1 U9018 ( .A1(n15187), .A2(n13941), .ZN(n7116) );
  NAND2_X1 U9019 ( .A1(n7003), .A2(n7314), .ZN(P2_U3496) );
  NAND2_X1 U9020 ( .A1(n15185), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U9021 ( .A1(n13947), .A2(n15187), .ZN(n7003) );
  XNOR2_X1 U9022 ( .A(n6647), .B(n7027), .ZN(n14010) );
  AOI211_X1 U9023 ( .C1(n14518), .C2(n14571), .A(n14342), .B(n14341), .ZN(
        n14343) );
  NAND2_X1 U9024 ( .A1(n7597), .A2(n7596), .ZN(P1_U3556) );
  AOI22_X1 U9025 ( .A1(n14335), .A2(n11847), .B1(P1_REG1_REG_28__SCAN_IN), 
        .B2(n15120), .ZN(n7596) );
  NAND2_X1 U9026 ( .A1(n14661), .A2(n15123), .ZN(n7597) );
  NAND2_X1 U9027 ( .A1(n7397), .A2(n7393), .ZN(P1_U3524) );
  NOR2_X1 U9028 ( .A1(n7396), .A2(n7394), .ZN(n7393) );
  NAND2_X1 U9029 ( .A1(n14661), .A2(n15111), .ZN(n7397) );
  NOR2_X1 U9030 ( .A1(n15111), .A2(n7395), .ZN(n7394) );
  NOR2_X1 U9031 ( .A1(n14953), .A2(n14952), .ZN(n14951) );
  INV_X1 U9032 ( .A(n7351), .ZN(n14962) );
  NAND2_X1 U9033 ( .A1(n6758), .A2(n6763), .ZN(n14964) );
  INV_X1 U9034 ( .A(n6769), .ZN(n14835) );
  OR2_X1 U9035 ( .A1(n12807), .A2(n12806), .ZN(n7259) );
  INV_X1 U9036 ( .A(n7259), .ZN(n6690) );
  OAI21_X1 U9037 ( .B1(n14529), .B2(n7602), .A(n14268), .ZN(n7601) );
  INV_X2 U9038 ( .A(n9680), .ZN(n10023) );
  NAND2_X1 U9039 ( .A1(n14961), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7104) );
  INV_X1 U9040 ( .A(n7104), .ZN(n6766) );
  INV_X1 U9041 ( .A(n6705), .ZN(n6704) );
  OAI21_X1 U9042 ( .B1(n12699), .B2(n12700), .A(n6707), .ZN(n6705) );
  INV_X1 U9043 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13982) );
  AND2_X2 U9044 ( .A1(n9665), .A2(n8466), .ZN(n8922) );
  INV_X2 U9045 ( .A(n9198), .ZN(n9196) );
  NOR2_X1 U9046 ( .A1(n13350), .A2(n7344), .ZN(n6436) );
  AND2_X1 U9047 ( .A1(n7281), .A2(n7280), .ZN(n6437) );
  AND2_X1 U9048 ( .A1(n14475), .A2(n14297), .ZN(n6438) );
  INV_X1 U9049 ( .A(n12018), .ZN(n7614) );
  AND2_X1 U9050 ( .A1(n6854), .A2(n12011), .ZN(n6439) );
  AND2_X1 U9051 ( .A1(n13705), .A2(n13629), .ZN(n6440) );
  INV_X1 U9052 ( .A(n12700), .ZN(n6706) );
  NAND4_X2 U9053 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .ZN(n12693)
         );
  XNOR2_X1 U9054 ( .A(n8458), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8466) );
  INV_X1 U9055 ( .A(n13148), .ZN(n6680) );
  NAND2_X1 U9056 ( .A1(n8625), .A2(SI_6_), .ZN(n6441) );
  AND2_X1 U9057 ( .A1(n14633), .A2(n14510), .ZN(n6442) );
  AND2_X1 U9058 ( .A1(n6841), .A2(n6840), .ZN(n6443) );
  AND2_X1 U9059 ( .A1(n13309), .A2(n13310), .ZN(n6444) );
  AND2_X1 U9060 ( .A1(n8207), .A2(n7217), .ZN(n6445) );
  INV_X1 U9061 ( .A(n14344), .ZN(n7620) );
  NAND2_X1 U9062 ( .A1(n7524), .A2(n7670), .ZN(n7739) );
  AND4_X1 U9063 ( .A1(n8230), .A2(n12905), .A3(n8229), .A4(n12921), .ZN(n6446)
         );
  NAND2_X1 U9064 ( .A1(n9154), .A2(n9153), .ZN(n13660) );
  NAND2_X1 U9065 ( .A1(n8353), .A2(n8356), .ZN(n12961) );
  NOR2_X1 U9066 ( .A1(n11062), .A2(n7589), .ZN(n7587) );
  INV_X1 U9067 ( .A(n7669), .ZN(n7518) );
  NAND2_X1 U9068 ( .A1(n10118), .A2(n10117), .ZN(n6447) );
  XOR2_X1 U9069 ( .A(n9171), .B(n13574), .Z(n6448) );
  AND2_X1 U9070 ( .A1(n12207), .A2(n7411), .ZN(n6449) );
  AND2_X1 U9071 ( .A1(n6799), .A2(n11160), .ZN(n6450) );
  AND2_X1 U9072 ( .A1(n6521), .A2(n10355), .ZN(n6451) );
  INV_X1 U9073 ( .A(n14961), .ZN(n7350) );
  INV_X1 U9074 ( .A(n8809), .ZN(n7477) );
  AND2_X1 U9075 ( .A1(n8681), .A2(n8680), .ZN(n6452) );
  OR2_X1 U9076 ( .A1(n7475), .A2(SI_14_), .ZN(n6453) );
  AND3_X1 U9077 ( .A1(n6441), .A2(n8597), .A3(n8577), .ZN(n6454) );
  AND2_X1 U9078 ( .A1(n7323), .A2(n13319), .ZN(n6455) );
  INV_X1 U9079 ( .A(n7601), .ZN(n7600) );
  INV_X1 U9080 ( .A(n14335), .ZN(n14662) );
  NAND2_X1 U9081 ( .A1(n11915), .A2(n11914), .ZN(n14335) );
  NAND2_X1 U9082 ( .A1(n9130), .A2(n9129), .ZN(n9171) );
  NOR2_X1 U9083 ( .A1(n7373), .A2(n12763), .ZN(n6456) );
  INV_X1 U9084 ( .A(n14501), .ZN(n7420) );
  INV_X1 U9085 ( .A(n12842), .ZN(n7368) );
  INV_X1 U9086 ( .A(n12827), .ZN(n7258) );
  INV_X2 U9087 ( .A(n8749), .ZN(n8907) );
  INV_X2 U9088 ( .A(n10786), .ZN(n12292) );
  CLKBUF_X3 U9089 ( .A(n10243), .Z(n12061) );
  AND2_X1 U9090 ( .A1(n14710), .A2(n9958), .ZN(n6457) );
  NAND2_X1 U9091 ( .A1(n8785), .A2(n9391), .ZN(n7478) );
  INV_X1 U9092 ( .A(n14448), .ZN(n7132) );
  NAND2_X1 U9093 ( .A1(n12446), .A2(n7501), .ZN(n7500) );
  INV_X1 U9094 ( .A(n8510), .ZN(n8560) );
  INV_X1 U9095 ( .A(n13636), .ZN(n7007) );
  NAND2_X2 U9096 ( .A1(n13986), .A2(n13988), .ZN(n8962) );
  INV_X2 U9097 ( .A(n8962), .ZN(n8511) );
  AND2_X1 U9098 ( .A1(n8104), .A2(n8352), .ZN(n6458) );
  OR2_X1 U9099 ( .A1(n11598), .A2(n6671), .ZN(n6459) );
  INV_X1 U9100 ( .A(n12408), .ZN(n7572) );
  OR2_X1 U9101 ( .A1(n13139), .A2(n12919), .ZN(n8214) );
  AND2_X1 U9102 ( .A1(n8662), .A2(n8661), .ZN(n6460) );
  AND2_X1 U9103 ( .A1(n6465), .A2(n7540), .ZN(n6461) );
  NOR2_X1 U9104 ( .A1(n11007), .A2(n7334), .ZN(n7333) );
  INV_X1 U9105 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9306) );
  OR2_X1 U9106 ( .A1(n6460), .A2(n7548), .ZN(n6462) );
  AND4_X1 U9107 ( .A1(n6702), .A2(n6700), .A3(n6699), .A4(n6697), .ZN(n6463)
         );
  NAND2_X1 U9108 ( .A1(n11816), .A2(n11817), .ZN(n6464) );
  INV_X1 U9109 ( .A(n7113), .ZN(n7112) );
  NAND2_X1 U9110 ( .A1(n14952), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7113) );
  AND2_X1 U9111 ( .A1(n8847), .A2(n8846), .ZN(n6465) );
  INV_X1 U9112 ( .A(n7503), .ZN(n7499) );
  NAND2_X1 U9113 ( .A1(n9736), .A2(n7038), .ZN(n10783) );
  OR2_X1 U9114 ( .A1(n14633), .A2(n14510), .ZN(n6466) );
  AND2_X1 U9115 ( .A1(n9491), .A2(n14173), .ZN(n6467) );
  AND2_X1 U9116 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n6468) );
  AND2_X1 U9117 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6469) );
  XNOR2_X1 U9118 ( .A(n14316), .B(n14261), .ZN(n6470) );
  AND2_X1 U9119 ( .A1(n12635), .A2(n15288), .ZN(n6471) );
  NOR2_X1 U9120 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9281) );
  INV_X1 U9121 ( .A(n14296), .ZN(n14473) );
  OAI21_X1 U9122 ( .B1(n12947), .B2(n7515), .A(n7514), .ZN(n12917) );
  AOI21_X1 U9123 ( .B1(n12456), .B2(n15218), .A(n12455), .ZN(n13138) );
  XNOR2_X1 U9124 ( .A(n12690), .B(n10918), .ZN(n11013) );
  AND2_X1 U9125 ( .A1(n13986), .A2(n8434), .ZN(n8536) );
  INV_X1 U9126 ( .A(n11688), .ZN(n11861) );
  AND2_X1 U9127 ( .A1(n13955), .A2(n13631), .ZN(n6472) );
  OR2_X1 U9128 ( .A1(n14785), .A2(n14784), .ZN(n6473) );
  OR2_X1 U9129 ( .A1(n14792), .A2(n14791), .ZN(n6474) );
  AND2_X1 U9130 ( .A1(n14429), .A2(n14276), .ZN(n6475) );
  NAND2_X1 U9131 ( .A1(n8774), .A2(n8773), .ZN(n11678) );
  OR2_X1 U9132 ( .A1(n12942), .A2(n12678), .ZN(n6476) );
  AND2_X1 U9133 ( .A1(n14600), .A2(n14304), .ZN(n6477) );
  AND2_X1 U9134 ( .A1(n9264), .A2(n9265), .ZN(n6478) );
  OR2_X1 U9135 ( .A1(n14776), .A2(n14775), .ZN(n6479) );
  INV_X1 U9136 ( .A(n11152), .ZN(n11142) );
  INV_X1 U9137 ( .A(n13334), .ZN(n7316) );
  OR2_X1 U9138 ( .A1(n14826), .A2(n14825), .ZN(n6480) );
  AND2_X1 U9139 ( .A1(n7190), .A2(n6598), .ZN(n6481) );
  AND2_X1 U9140 ( .A1(n13930), .A2(n13610), .ZN(n6482) );
  AND2_X1 U9141 ( .A1(n6680), .A2(n15289), .ZN(n6483) );
  AND2_X1 U9142 ( .A1(n8990), .A2(n8989), .ZN(n6484) );
  INV_X1 U9143 ( .A(n8704), .ZN(n7531) );
  AND2_X1 U9144 ( .A1(n13597), .A2(n13596), .ZN(n6485) );
  AND2_X1 U9145 ( .A1(n8780), .A2(n8779), .ZN(n6486) );
  AND2_X1 U9146 ( .A1(n14389), .A2(n14307), .ZN(n6487) );
  AND2_X1 U9147 ( .A1(n14283), .A2(n14282), .ZN(n6488) );
  AND2_X1 U9148 ( .A1(n11258), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6489) );
  AND2_X1 U9149 ( .A1(n11258), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6490) );
  AND2_X1 U9150 ( .A1(n10723), .A2(n13482), .ZN(n6491) );
  INV_X1 U9151 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13298) );
  AND2_X1 U9152 ( .A1(n12467), .A2(n7175), .ZN(n6492) );
  NOR2_X1 U9153 ( .A1(n12700), .A2(n11142), .ZN(n6493) );
  INV_X1 U9154 ( .A(n10546), .ZN(n7295) );
  NAND2_X1 U9155 ( .A1(n10827), .A2(n10826), .ZN(n14905) );
  OR2_X1 U9156 ( .A1(n13648), .A2(n13647), .ZN(n6494) );
  OR2_X1 U9157 ( .A1(n7232), .A2(n11196), .ZN(n6495) );
  AND2_X1 U9158 ( .A1(n6894), .A2(n9812), .ZN(n6496) );
  AND2_X1 U9159 ( .A1(n6804), .A2(n7663), .ZN(n6497) );
  NOR2_X1 U9160 ( .A1(n14289), .A2(n12228), .ZN(n6498) );
  NAND2_X1 U9161 ( .A1(n9710), .A2(n9709), .ZN(n10923) );
  OR2_X1 U9162 ( .A1(n8896), .A2(n8898), .ZN(n6499) );
  INV_X1 U9163 ( .A(n14535), .ZN(n14647) );
  NAND2_X1 U9164 ( .A1(n12025), .A2(n12024), .ZN(n14535) );
  AND2_X1 U9165 ( .A1(n13871), .A2(n13632), .ZN(n6500) );
  AND2_X1 U9166 ( .A1(n7350), .A2(n7349), .ZN(n6501) );
  OR2_X1 U9167 ( .A1(n7421), .A2(n6498), .ZN(n6502) );
  AND2_X1 U9168 ( .A1(n10238), .A2(n10240), .ZN(n6503) );
  INV_X1 U9169 ( .A(n7575), .ZN(n7574) );
  NAND2_X1 U9170 ( .A1(n7576), .A2(n14012), .ZN(n7575) );
  AND2_X1 U9171 ( .A1(n10484), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6504) );
  INV_X1 U9172 ( .A(n12164), .ZN(n7433) );
  INV_X1 U9173 ( .A(n12134), .ZN(n7431) );
  INV_X1 U9174 ( .A(n12150), .ZN(n7426) );
  INV_X1 U9175 ( .A(n7560), .ZN(n7559) );
  NAND2_X1 U9176 ( .A1(n12290), .A2(n14907), .ZN(n7560) );
  AND2_X1 U9177 ( .A1(n8446), .A2(n6745), .ZN(n6505) );
  INV_X1 U9178 ( .A(n12202), .ZN(n7428) );
  INV_X1 U9179 ( .A(n13565), .ZN(n13946) );
  NAND2_X1 U9180 ( .A1(n9091), .A2(n9090), .ZN(n13565) );
  OR2_X1 U9181 ( .A1(n8571), .A2(n8570), .ZN(n6506) );
  INV_X1 U9182 ( .A(n7589), .ZN(n7588) );
  AND2_X1 U9183 ( .A1(n10023), .A2(n10541), .ZN(n6507) );
  AND2_X1 U9184 ( .A1(n12308), .A2(n14148), .ZN(n6508) );
  AND2_X1 U9185 ( .A1(n12375), .A2(n12374), .ZN(n6509) );
  INV_X1 U9186 ( .A(n13622), .ZN(n6729) );
  AND2_X1 U9187 ( .A1(n12381), .A2(n12380), .ZN(n6510) );
  NAND2_X1 U9188 ( .A1(n7218), .A2(n8214), .ZN(n7217) );
  INV_X1 U9189 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7244) );
  AND2_X1 U9190 ( .A1(n12606), .A2(n7180), .ZN(n6511) );
  NOR2_X1 U9191 ( .A1(n6501), .A2(n14800), .ZN(n7103) );
  AND2_X1 U9192 ( .A1(n12403), .A2(n12402), .ZN(n6512) );
  AND2_X1 U9193 ( .A1(n11904), .A2(n11903), .ZN(n14564) );
  INV_X1 U9194 ( .A(n14564), .ZN(n14321) );
  NOR2_X1 U9195 ( .A1(n12291), .A2(n14924), .ZN(n6513) );
  NOR2_X1 U9196 ( .A1(n13089), .A2(n13100), .ZN(n6514) );
  NOR2_X1 U9197 ( .A1(n12148), .A2(n14909), .ZN(n6515) );
  NOR2_X1 U9198 ( .A1(n14637), .A2(n14488), .ZN(n6516) );
  NOR2_X1 U9199 ( .A1(n11863), .A2(n11854), .ZN(n6517) );
  NOR2_X1 U9200 ( .A1(n13753), .A2(n13620), .ZN(n6518) );
  NOR2_X1 U9201 ( .A1(n14443), .A2(n14300), .ZN(n6519) );
  OR2_X1 U9202 ( .A1(n7537), .A2(n6461), .ZN(n6520) );
  OR2_X1 U9203 ( .A1(n10552), .A2(n10551), .ZN(n6521) );
  INV_X1 U9204 ( .A(n7294), .ZN(n7293) );
  OAI21_X1 U9205 ( .B1(n7296), .B2(n7295), .A(n10554), .ZN(n7294) );
  NAND2_X1 U9206 ( .A1(n14697), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6522) );
  OR2_X1 U9207 ( .A1(n6828), .A2(n6444), .ZN(n6523) );
  AND2_X1 U9208 ( .A1(n11750), .A2(n11749), .ZN(n6524) );
  AND2_X1 U9209 ( .A1(n10334), .A2(n10333), .ZN(n6525) );
  NAND3_X1 U9210 ( .A1(n12173), .A2(n12172), .A3(n12171), .ZN(n6526) );
  NOR2_X1 U9211 ( .A1(n12133), .A2(n7431), .ZN(n6527) );
  AND2_X1 U9212 ( .A1(n6961), .A2(n6962), .ZN(n6528) );
  OR2_X1 U9213 ( .A1(n7679), .A2(n7522), .ZN(n6529) );
  INV_X1 U9214 ( .A(n12136), .ZN(n7069) );
  AND2_X1 U9215 ( .A1(n6952), .A2(n6955), .ZN(n6530) );
  AND2_X1 U9216 ( .A1(n7117), .A2(n13415), .ZN(n6531) );
  AND2_X1 U9217 ( .A1(n8691), .A2(SI_9_), .ZN(n6532) );
  OR2_X1 U9218 ( .A1(n8782), .A2(n6486), .ZN(n6533) );
  INV_X1 U9219 ( .A(n10632), .ZN(n7549) );
  INV_X1 U9220 ( .A(n7508), .ZN(n7507) );
  NAND2_X1 U9221 ( .A1(n7509), .A2(n15194), .ZN(n7508) );
  INV_X1 U9222 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9264) );
  AND2_X1 U9223 ( .A1(n9032), .A2(n9031), .ZN(n6534) );
  AND2_X1 U9224 ( .A1(n7169), .A2(n7171), .ZN(n6535) );
  NAND2_X1 U9225 ( .A1(n7657), .A2(n7523), .ZN(n7522) );
  AND2_X1 U9226 ( .A1(n8309), .A2(n8314), .ZN(n13087) );
  INV_X1 U9227 ( .A(n13087), .ZN(n7198) );
  OAI21_X1 U9228 ( .B1(n13225), .B2(n12895), .A(n8203), .ZN(n8383) );
  INV_X1 U9229 ( .A(n7181), .ZN(n7180) );
  OR2_X1 U9230 ( .A1(n12552), .A2(n7182), .ZN(n7181) );
  AND2_X1 U9231 ( .A1(n7428), .A2(n12201), .ZN(n6536) );
  INV_X1 U9232 ( .A(n7226), .ZN(n7225) );
  NAND2_X1 U9233 ( .A1(n8341), .A2(n7227), .ZN(n7226) );
  INV_X1 U9234 ( .A(n7221), .ZN(n7220) );
  NAND2_X1 U9235 ( .A1(n8214), .A2(n12921), .ZN(n7221) );
  NOR2_X1 U9236 ( .A1(n13241), .A2(n12948), .ZN(n6537) );
  AND2_X1 U9237 ( .A1(n8206), .A2(n8205), .ZN(n6538) );
  INV_X1 U9238 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8483) );
  INV_X1 U9239 ( .A(n8828), .ZN(n7475) );
  AND2_X1 U9240 ( .A1(n8830), .A2(n8813), .ZN(n8828) );
  INV_X1 U9241 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15313) );
  INV_X1 U9242 ( .A(n12217), .ZN(n7054) );
  INV_X1 U9243 ( .A(n12227), .ZN(n7059) );
  AND2_X1 U9244 ( .A1(n12004), .A2(n10250), .ZN(n6539) );
  OR2_X1 U9245 ( .A1(n12691), .A2(n10707), .ZN(n8251) );
  OR2_X1 U9246 ( .A1(n8947), .A2(n8949), .ZN(n6540) );
  AND3_X1 U9247 ( .A1(n8389), .A2(n8392), .A3(n7677), .ZN(n6541) );
  INV_X1 U9248 ( .A(n8590), .ZN(n6991) );
  AND2_X1 U9249 ( .A1(n8087), .A2(n8352), .ZN(n6542) );
  OR2_X1 U9250 ( .A1(n13628), .A2(n6440), .ZN(n6543) );
  NOR2_X1 U9251 ( .A1(n14337), .A2(n6856), .ZN(n6544) );
  AND2_X1 U9252 ( .A1(n8460), .A2(n7546), .ZN(n6545) );
  NOR2_X1 U9253 ( .A1(n13609), .A2(n7642), .ZN(n7641) );
  AND2_X1 U9254 ( .A1(n8329), .A2(n12436), .ZN(n6546) );
  INV_X1 U9255 ( .A(n14271), .ZN(n14461) );
  INV_X1 U9256 ( .A(n7236), .ZN(n7235) );
  OAI21_X1 U9257 ( .B1(n7848), .B2(n7237), .A(n7868), .ZN(n7236) );
  INV_X1 U9258 ( .A(n8597), .ZN(n7438) );
  AND2_X1 U9259 ( .A1(n7500), .A2(n7499), .ZN(n6547) );
  OR2_X1 U9260 ( .A1(n7428), .A2(n12201), .ZN(n6548) );
  AND2_X1 U9261 ( .A1(n9005), .A2(n9004), .ZN(n6549) );
  OR2_X1 U9262 ( .A1(n7433), .A2(n12163), .ZN(n6550) );
  AND3_X1 U9263 ( .A1(n9325), .A2(n9262), .A3(n9261), .ZN(n6551) );
  AOI21_X1 U9264 ( .B1(n6535), .B2(n7167), .A(n7166), .ZN(n7165) );
  OR2_X1 U9265 ( .A1(n7526), .A2(n8948), .ZN(n6552) );
  OR2_X1 U9266 ( .A1(n8704), .A2(n8705), .ZN(n6553) );
  OR2_X1 U9267 ( .A1(n7426), .A2(n12149), .ZN(n6554) );
  OR2_X1 U9268 ( .A1(n7064), .A2(n12129), .ZN(n6555) );
  NOR2_X1 U9269 ( .A1(n9363), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n6556) );
  OR2_X1 U9270 ( .A1(n7531), .A2(n7532), .ZN(n6557) );
  OR2_X1 U9271 ( .A1(n7535), .A2(n6484), .ZN(n6558) );
  AND2_X1 U9272 ( .A1(n6873), .A2(n6466), .ZN(n6870) );
  INV_X1 U9273 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6664) );
  INV_X1 U9274 ( .A(n6963), .ZN(n6962) );
  NAND2_X1 U9275 ( .A1(n6964), .A2(n7547), .ZN(n6963) );
  INV_X2 U9276 ( .A(n7733), .ZN(n8191) );
  NAND2_X1 U9277 ( .A1(n7853), .A2(n7511), .ZN(n7909) );
  INV_X1 U9278 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6931) );
  INV_X1 U9279 ( .A(n13635), .ZN(n7010) );
  INV_X1 U9280 ( .A(n11135), .ZN(n7384) );
  XNOR2_X1 U9281 ( .A(n14600), .B(n14398), .ZN(n14416) );
  INV_X1 U9282 ( .A(n14416), .ZN(n7628) );
  AND2_X1 U9283 ( .A1(n7672), .A2(n7756), .ZN(n7853) );
  NAND2_X1 U9284 ( .A1(n7853), .A2(n7673), .ZN(n7872) );
  INV_X1 U9285 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6848) );
  NOR2_X1 U9286 ( .A1(n14462), .A2(n14443), .ZN(n7285) );
  INV_X1 U9287 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9902) );
  INV_X1 U9288 ( .A(n11172), .ZN(n7232) );
  NAND2_X1 U9289 ( .A1(n14908), .A2(n14907), .ZN(n14906) );
  AND2_X1 U9290 ( .A1(n13533), .A2(n13538), .ZN(n13546) );
  INV_X1 U9291 ( .A(n13546), .ZN(n6887) );
  INV_X1 U9292 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U9293 ( .A1(n11933), .A2(n11932), .ZN(n14593) );
  INV_X1 U9294 ( .A(n14593), .ZN(n6832) );
  OR2_X1 U9295 ( .A1(n12772), .A2(n12771), .ZN(n6559) );
  AND2_X1 U9296 ( .A1(n12720), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6560) );
  AND2_X1 U9297 ( .A1(n12517), .A2(n13119), .ZN(n6561) );
  NAND2_X1 U9298 ( .A1(n7519), .A2(n12436), .ZN(n13044) );
  NAND2_X1 U9299 ( .A1(n9134), .A2(n9133), .ZN(n13864) );
  INV_X1 U9300 ( .A(n13864), .ZN(n7123) );
  AND2_X1 U9301 ( .A1(n9028), .A2(n9027), .ZN(n6562) );
  NAND2_X1 U9302 ( .A1(n6437), .A2(n6839), .ZN(n6563) );
  AND2_X1 U9303 ( .A1(n8332), .A2(n8322), .ZN(n6564) );
  AND2_X1 U9304 ( .A1(n12498), .A2(n13020), .ZN(n6565) );
  NOR2_X1 U9305 ( .A1(n13825), .A2(n13925), .ZN(n13797) );
  OR2_X1 U9306 ( .A1(n13098), .A2(n13097), .ZN(n13096) );
  AND2_X1 U9307 ( .A1(n7328), .A2(n7326), .ZN(n6566) );
  AND2_X1 U9308 ( .A1(n6768), .A2(n7103), .ZN(n6567) );
  AND2_X1 U9309 ( .A1(n11768), .A2(n7616), .ZN(n6568) );
  AND2_X1 U9310 ( .A1(n12356), .A2(n12354), .ZN(n6569) );
  AND2_X1 U9311 ( .A1(n7387), .A2(n7386), .ZN(n6570) );
  AND2_X1 U9312 ( .A1(n8069), .A2(n8068), .ZN(n13257) );
  NAND2_X1 U9313 ( .A1(n7853), .A2(n7512), .ZN(n7513) );
  NAND2_X1 U9314 ( .A1(n8390), .A2(n8389), .ZN(n6571) );
  AND2_X1 U9315 ( .A1(n12349), .A2(n12348), .ZN(n6572) );
  AND2_X1 U9316 ( .A1(n12720), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6573) );
  INV_X1 U9317 ( .A(n7947), .ZN(n6930) );
  AND2_X1 U9318 ( .A1(n7949), .A2(n7937), .ZN(n7947) );
  INV_X1 U9319 ( .A(n7650), .ZN(n8835) );
  OR2_X1 U9320 ( .A1(n7448), .A2(n7449), .ZN(n6574) );
  AND2_X1 U9321 ( .A1(n7351), .A2(n7350), .ZN(n6575) );
  OR2_X1 U9322 ( .A1(n12763), .A2(n7372), .ZN(n6576) );
  INV_X1 U9323 ( .A(n6688), .ZN(n12878) );
  NAND2_X1 U9324 ( .A1(n8029), .A2(n8028), .ZN(n6688) );
  NOR2_X1 U9325 ( .A1(n12004), .A2(n7608), .ZN(n7607) );
  INV_X1 U9326 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U9327 ( .A1(n11790), .A2(n11789), .ZN(n14264) );
  INV_X1 U9328 ( .A(n14264), .ZN(n7280) );
  INV_X1 U9329 ( .A(n10929), .ZN(n7646) );
  NOR2_X1 U9330 ( .A1(n10068), .A2(n10067), .ZN(n10072) );
  INV_X1 U9331 ( .A(n13435), .ZN(n7323) );
  INV_X2 U9332 ( .A(n15295), .ZN(n15293) );
  AND2_X1 U9333 ( .A1(n11360), .A2(n7117), .ZN(n6577) );
  NAND2_X1 U9334 ( .A1(n11983), .A2(n11982), .ZN(n14633) );
  INV_X1 U9335 ( .A(n14633), .ZN(n7286) );
  AND2_X1 U9336 ( .A1(n8452), .A2(n8446), .ZN(n6578) );
  INV_X1 U9337 ( .A(n11044), .ZN(n6670) );
  INV_X1 U9338 ( .A(n7550), .ZN(n10781) );
  INV_X1 U9339 ( .A(n7203), .ZN(n7202) );
  NOR2_X1 U9340 ( .A1(n13108), .A2(n8301), .ZN(n7203) );
  NOR2_X1 U9341 ( .A1(n12889), .A2(n7377), .ZN(n6579) );
  AND2_X1 U9342 ( .A1(n10350), .A2(n10349), .ZN(n6580) );
  AND2_X1 U9343 ( .A1(n7609), .A2(n10458), .ZN(n6581) );
  AND2_X1 U9344 ( .A1(n11058), .A2(n7587), .ZN(n6582) );
  INV_X1 U9345 ( .A(n7126), .ZN(n10361) );
  NOR2_X1 U9346 ( .A1(n10338), .A2(n15178), .ZN(n7126) );
  INV_X1 U9347 ( .A(n7283), .ZN(n11536) );
  AND2_X1 U9348 ( .A1(n6443), .A2(n10880), .ZN(n7283) );
  AND2_X1 U9349 ( .A1(n15351), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6583) );
  INV_X1 U9350 ( .A(n7256), .ZN(n7255) );
  OAI21_X1 U9351 ( .B1(n8065), .B2(n7257), .A(n8077), .ZN(n7256) );
  NOR2_X1 U9352 ( .A1(n10140), .A2(n10139), .ZN(n6584) );
  AND2_X1 U9353 ( .A1(n12748), .A2(n7374), .ZN(n6585) );
  OR2_X1 U9354 ( .A1(n10540), .A2(n9668), .ZN(n9680) );
  NAND2_X1 U9355 ( .A1(n11469), .A2(n11468), .ZN(n12291) );
  INV_X1 U9356 ( .A(n12291), .ZN(n6840) );
  NAND2_X1 U9357 ( .A1(n11475), .A2(n11474), .ZN(n12301) );
  INV_X1 U9358 ( .A(n12301), .ZN(n7282) );
  INV_X1 U9359 ( .A(n14067), .ZN(n6833) );
  NAND2_X1 U9360 ( .A1(n9624), .A2(n9623), .ZN(n13470) );
  INV_X1 U9361 ( .A(n13470), .ZN(n14883) );
  OR2_X1 U9362 ( .A1(n12811), .A2(n12830), .ZN(n6586) );
  INV_X1 U9363 ( .A(n12832), .ZN(n7369) );
  INV_X1 U9364 ( .A(n10552), .ZN(n7125) );
  NAND2_X1 U9365 ( .A1(n7315), .A2(n9628), .ZN(n9664) );
  OR2_X1 U9366 ( .A1(n15190), .A2(n15448), .ZN(n6587) );
  XNOR2_X1 U9367 ( .A(n8470), .B(n8469), .ZN(n9234) );
  AND2_X1 U9368 ( .A1(n7955), .A2(n7986), .ZN(n12809) );
  AND2_X1 U9369 ( .A1(n10768), .A2(n10767), .ZN(n15223) );
  INV_X1 U9370 ( .A(n15223), .ZN(n15201) );
  NAND2_X1 U9371 ( .A1(n12796), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6588) );
  AND2_X1 U9372 ( .A1(n12842), .A2(n7258), .ZN(n6589) );
  NAND2_X1 U9373 ( .A1(n6703), .A2(n6706), .ZN(n6590) );
  AND2_X1 U9374 ( .A1(n7581), .A2(n7580), .ZN(n6591) );
  OR2_X1 U9375 ( .A1(n13639), .A2(n13638), .ZN(n6592) );
  AND2_X1 U9376 ( .A1(n10242), .A2(n15064), .ZN(n15074) );
  INV_X1 U9377 ( .A(n15074), .ZN(n15108) );
  INV_X1 U9378 ( .A(n10268), .ZN(n7606) );
  AND2_X1 U9379 ( .A1(n8534), .A2(n8556), .ZN(n13505) );
  INV_X1 U9380 ( .A(n13505), .ZN(n6886) );
  XOR2_X1 U9381 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .Z(n6593) );
  XOR2_X1 U9382 ( .A(n12720), .B(P3_REG1_REG_8__SCAN_IN), .Z(n6594) );
  INV_X1 U9383 ( .A(n8434), .ZN(n13988) );
  AND2_X1 U9384 ( .A1(n15339), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6595) );
  INV_X1 U9385 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7349) );
  INV_X1 U9386 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7695) );
  INV_X1 U9387 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7001) );
  INV_X1 U9388 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7359) );
  INV_X1 U9389 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7360) );
  INV_X1 U9390 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7102) );
  INV_X1 U9391 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7106) );
  INV_X1 U9392 ( .A(n12771), .ZN(n7374) );
  NAND2_X1 U9393 ( .A1(n12749), .A2(n12771), .ZN(n6656) );
  OAI21_X2 U9394 ( .B1(n15192), .B2(n8288), .A(n8284), .ZN(n14851) );
  NAND2_X1 U9395 ( .A1(n11012), .A2(n11018), .ZN(n7785) );
  AOI21_X1 U9396 ( .B1(n10909), .B2(n8247), .A(n6602), .ZN(n6600) );
  NAND2_X1 U9397 ( .A1(n7743), .A2(n8251), .ZN(n10910) );
  INV_X1 U9398 ( .A(n8028), .ZN(n6603) );
  INV_X1 U9399 ( .A(n7702), .ZN(n6779) );
  NAND2_X1 U9400 ( .A1(n6605), .A2(n8250), .ZN(n10892) );
  XNOR2_X1 U9401 ( .A(n10576), .B(n10712), .ZN(n10762) );
  INV_X2 U9402 ( .A(n6608), .ZN(n11143) );
  NAND2_X2 U9403 ( .A1(n8404), .A2(n6608), .ZN(n11076) );
  MUX2_X1 U9404 ( .A(n11078), .B(n11079), .S(n11143), .Z(n11081) );
  MUX2_X1 U9405 ( .A(n11090), .B(n11091), .S(n11143), .Z(n11092) );
  MUX2_X1 U9406 ( .A(n15300), .B(n15230), .S(n11143), .Z(n11106) );
  MUX2_X1 U9407 ( .A(n11161), .B(n11162), .S(n11143), .Z(n11163) );
  MUX2_X1 U9408 ( .A(P3_REG1_REG_12__SCAN_IN), .B(P3_REG2_REG_12__SCAN_IN), 
        .S(n11143), .Z(n12740) );
  MUX2_X1 U9409 ( .A(P3_REG1_REG_18__SCAN_IN), .B(P3_REG2_REG_18__SCAN_IN), 
        .S(n11143), .Z(n12847) );
  NAND2_X1 U9410 ( .A1(n13329), .A2(n13330), .ZN(n6609) );
  NAND3_X1 U9411 ( .A1(n6616), .A2(n7458), .A3(n6615), .ZN(n6614) );
  NAND3_X1 U9412 ( .A1(n13416), .A2(n7324), .A3(n6455), .ZN(n6617) );
  NOR2_X2 U9413 ( .A1(n10024), .A2(n10319), .ZN(n10096) );
  NOR2_X4 U9414 ( .A1(n11415), .A2(n13847), .ZN(n11360) );
  OR2_X2 U9415 ( .A1(n10938), .A2(n11412), .ZN(n11415) );
  NAND2_X1 U9416 ( .A1(n6434), .A2(n10807), .ZN(n10938) );
  NAND2_X1 U9417 ( .A1(n13730), .A2(n13567), .ZN(n13731) );
  NOR2_X2 U9418 ( .A1(n13761), .A2(n13753), .ZN(n13730) );
  INV_X1 U9419 ( .A(n9644), .ZN(n10049) );
  NAND2_X2 U9420 ( .A1(n13996), .A2(n9247), .ZN(n9393) );
  XNOR2_X2 U9421 ( .A(n6619), .B(n8442), .ZN(n9247) );
  NAND3_X1 U9422 ( .A1(n7650), .A2(n7649), .A3(n8421), .ZN(n6620) );
  NAND2_X1 U9423 ( .A1(n14136), .A2(n7582), .ZN(n6622) );
  NAND2_X1 U9424 ( .A1(n6625), .A2(n12320), .ZN(n12321) );
  NAND3_X1 U9425 ( .A1(n7550), .A2(n7552), .A3(n10635), .ZN(n10782) );
  NAND2_X1 U9426 ( .A1(n9873), .A2(n6648), .ZN(n14155) );
  NOR2_X1 U9427 ( .A1(n6649), .A2(n6504), .ZN(n6648) );
  XNOR2_X1 U9428 ( .A(n11126), .B(n11152), .ZN(n11127) );
  INV_X1 U9429 ( .A(n6659), .ZN(n12795) );
  NAND2_X1 U9430 ( .A1(n6659), .A2(n6658), .ZN(n6657) );
  INV_X1 U9431 ( .A(n12794), .ZN(n6658) );
  NAND2_X1 U9432 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6663) );
  NAND3_X1 U9433 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6665) );
  OAI21_X2 U9434 ( .B1(n11601), .B2(n7508), .A(n7505), .ZN(n14853) );
  INV_X1 U9435 ( .A(n6667), .ZN(n6666) );
  OAI211_X1 U9436 ( .C1(n6676), .C2(n6675), .A(n11013), .B(n6673), .ZN(n11017)
         );
  NAND2_X1 U9437 ( .A1(n6674), .A2(n10772), .ZN(n6673) );
  AND2_X1 U9438 ( .A1(n10895), .A2(n10896), .ZN(n6676) );
  NAND2_X1 U9439 ( .A1(n10772), .A2(n10771), .ZN(n10897) );
  NAND2_X1 U9440 ( .A1(n10913), .A2(n10912), .ZN(n11014) );
  NAND2_X1 U9441 ( .A1(n6676), .A2(n10897), .ZN(n10913) );
  INV_X1 U9442 ( .A(n10912), .ZN(n6675) );
  NAND3_X1 U9443 ( .A1(n6704), .A2(n12701), .A3(n11142), .ZN(n6699) );
  NAND3_X1 U9444 ( .A1(n6712), .A2(P3_REG1_REG_15__SCAN_IN), .A3(n12787), .ZN(
        n7260) );
  NAND2_X1 U9445 ( .A1(n12788), .A2(n12797), .ZN(n12787) );
  INV_X1 U9446 ( .A(n12788), .ZN(n6711) );
  NAND2_X1 U9447 ( .A1(n6715), .A2(n6713), .ZN(n11237) );
  NAND3_X1 U9448 ( .A1(n11137), .A2(n6716), .A3(P3_REG1_REG_3__SCAN_IN), .ZN(
        n6715) );
  NAND2_X1 U9449 ( .A1(n11137), .A2(n11238), .ZN(n11582) );
  INV_X1 U9450 ( .A(n6719), .ZN(n6718) );
  NOR2_X1 U9451 ( .A1(n12755), .A2(n13208), .ZN(n12764) );
  NAND2_X1 U9452 ( .A1(n12754), .A2(n12771), .ZN(n6719) );
  NAND2_X1 U9453 ( .A1(n6721), .A2(n9842), .ZN(n9943) );
  NAND2_X1 U9454 ( .A1(n9841), .A2(n9840), .ZN(n6721) );
  NAND2_X1 U9455 ( .A1(n6724), .A2(n6722), .ZN(n9946) );
  INV_X1 U9456 ( .A(n6723), .ZN(n6722) );
  OAI21_X1 U9457 ( .B1(n9840), .B2(n6725), .A(n9942), .ZN(n6723) );
  NAND2_X1 U9458 ( .A1(n11697), .A2(n6739), .ZN(n6738) );
  OAI21_X4 U9459 ( .B1(n9247), .B2(n8598), .A(n6743), .ZN(n8786) );
  NAND3_X1 U9460 ( .A1(n6744), .A2(n8449), .A3(n11950), .ZN(n6743) );
  NAND2_X1 U9461 ( .A1(n6755), .A2(n6494), .ZN(n6751) );
  NAND2_X1 U9462 ( .A1(n13867), .A2(n6752), .ZN(n13948) );
  XNOR2_X1 U9463 ( .A(n14763), .B(n6756), .ZN(n14765) );
  NAND2_X1 U9464 ( .A1(n7351), .A2(n7104), .ZN(n6768) );
  INV_X1 U9465 ( .A(n14800), .ZN(n6767) );
  AND4_X2 U9466 ( .A1(n7511), .A2(n7672), .A3(n7756), .A4(n6774), .ZN(n8025)
         );
  NAND2_X1 U9467 ( .A1(n11618), .A2(n6780), .ZN(n6785) );
  NAND3_X1 U9468 ( .A1(n6786), .A2(n6791), .A3(n6785), .ZN(n6782) );
  XNOR2_X1 U9469 ( .A(n6811), .B(n12880), .ZN(n6810) );
  NOR2_X1 U9470 ( .A1(n12875), .A2(n6812), .ZN(n6811) );
  AND2_X1 U9471 ( .A1(n12877), .A2(n12876), .ZN(n6812) );
  OAI211_X1 U9472 ( .C1(n6435), .C2(P3_REG1_REG_0__SCAN_IN), .A(n6816), .B(
        n6813), .ZN(n11649) );
  NAND2_X1 U9473 ( .A1(n7704), .A2(n6814), .ZN(n6813) );
  INV_X1 U9474 ( .A(n6435), .ZN(n6815) );
  NAND2_X1 U9475 ( .A1(n13417), .A2(n13418), .ZN(n13416) );
  INV_X2 U9476 ( .A(n9958), .ZN(n12022) );
  NAND2_X1 U9477 ( .A1(n6845), .A2(n6842), .ZN(n14660) );
  AOI211_X1 U9478 ( .C1(n14329), .C2(n14321), .A(n14314), .B(n14640), .ZN(
        n14565) );
  NAND2_X1 U9479 ( .A1(n10743), .A2(n6439), .ZN(n6852) );
  NAND2_X1 U9480 ( .A1(n6852), .A2(n6853), .ZN(n10840) );
  NAND2_X1 U9481 ( .A1(n14345), .A2(n6544), .ZN(n14339) );
  NAND2_X1 U9482 ( .A1(n11484), .A2(n6860), .ZN(n6857) );
  NAND2_X1 U9483 ( .A1(n14266), .A2(n6870), .ZN(n6868) );
  MUX2_X1 U9484 ( .A(n10675), .B(P2_REG2_REG_1__SCAN_IN), .S(n9453), .Z(n9397)
         );
  NAND2_X1 U9485 ( .A1(n6905), .A2(n9796), .ZN(n9838) );
  OAI21_X1 U9486 ( .B1(n9796), .B2(n6905), .A(n9838), .ZN(n10572) );
  NAND2_X1 U9487 ( .A1(n13760), .A2(n13767), .ZN(n6906) );
  NAND2_X1 U9488 ( .A1(n13776), .A2(n13587), .ZN(n6907) );
  OAI21_X1 U9489 ( .B1(n10348), .B2(n7294), .A(n6908), .ZN(n10926) );
  NAND2_X1 U9490 ( .A1(n13597), .A2(n6919), .ZN(n13700) );
  NAND2_X1 U9491 ( .A1(n6912), .A2(n6913), .ZN(n13655) );
  NAND2_X1 U9492 ( .A1(n6924), .A2(n7983), .ZN(n7248) );
  XNOR2_X1 U9493 ( .A(n6924), .B(n7982), .ZN(n9654) );
  NAND2_X1 U9494 ( .A1(n7231), .A2(n7735), .ZN(n6925) );
  NAND2_X1 U9495 ( .A1(n7722), .A2(n7723), .ZN(n6926) );
  NAND2_X1 U9496 ( .A1(n8006), .A2(n6940), .ZN(n6939) );
  NAND2_X1 U9497 ( .A1(n8051), .A2(n8053), .ZN(n6944) );
  OAI21_X1 U9498 ( .B1(n7846), .B2(n7236), .A(n6946), .ZN(n7889) );
  NAND2_X1 U9499 ( .A1(n8093), .A2(n11748), .ZN(n6949) );
  NAND2_X1 U9500 ( .A1(n8121), .A2(n8120), .ZN(n6950) );
  OR2_X1 U9501 ( .A1(n9008), .A2(n6956), .ZN(n6952) );
  NAND2_X1 U9502 ( .A1(n9008), .A2(n6955), .ZN(n6954) );
  AOI21_X1 U9503 ( .B1(n8876), .B2(n8875), .A(n8874), .ZN(n8877) );
  NAND2_X1 U9504 ( .A1(n6958), .A2(n7536), .ZN(n8876) );
  NAND2_X1 U9505 ( .A1(n6959), .A2(n6520), .ZN(n6958) );
  NAND2_X1 U9506 ( .A1(n8639), .A2(n6966), .ZN(n6961) );
  OAI21_X1 U9507 ( .B1(n8639), .B2(n6963), .A(n6960), .ZN(n8685) );
  INV_X1 U9508 ( .A(n6967), .ZN(n6966) );
  NAND2_X1 U9509 ( .A1(n9033), .A2(n6974), .ZN(n6971) );
  OAI21_X1 U9510 ( .B1(n6971), .B2(n6534), .A(n6972), .ZN(n9071) );
  OAI21_X1 U9511 ( .B1(n6977), .B2(n6976), .A(n7529), .ZN(n8803) );
  NAND2_X1 U9512 ( .A1(n8617), .A2(n8618), .ZN(n8616) );
  OAI22_X1 U9513 ( .A1(n8592), .A2(n6978), .B1(n8590), .B2(n8591), .ZN(n8617)
         );
  NAND3_X1 U9514 ( .A1(n6984), .A2(n8926), .A3(n6540), .ZN(n7525) );
  NAND2_X1 U9515 ( .A1(n8572), .A2(n6506), .ZN(n8592) );
  OAI21_X1 U9516 ( .B1(n9204), .B2(n9203), .A(n9202), .ZN(n9252) );
  NAND2_X1 U9517 ( .A1(n8549), .A2(n7661), .ZN(n8571) );
  NAND2_X1 U9518 ( .A1(n10263), .A2(n10138), .ZN(n7339) );
  NAND3_X1 U9519 ( .A1(n6979), .A2(n13375), .A3(n14883), .ZN(n13356) );
  AOI21_X1 U9520 ( .B1(n9071), .B2(n9070), .A(n9069), .ZN(n9073) );
  AOI21_X1 U9521 ( .B1(n8571), .B2(n8570), .A(n8568), .ZN(n8569) );
  NAND2_X1 U9522 ( .A1(n8735), .A2(n8734), .ZN(n8763) );
  AND2_X1 U9523 ( .A1(n12810), .A2(n12809), .ZN(n6981) );
  NAND2_X1 U9524 ( .A1(n7375), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7373) );
  INV_X1 U9525 ( .A(n12747), .ZN(n12746) );
  NAND2_X1 U9526 ( .A1(n12747), .A2(n12748), .ZN(n12749) );
  NOR2_X1 U9527 ( .A1(n11181), .A2(n11182), .ZN(n11185) );
  NAND2_X1 U9528 ( .A1(n7525), .A2(n6552), .ZN(n8971) );
  NAND2_X1 U9529 ( .A1(n7533), .A2(n7534), .ZN(n9008) );
  NAND2_X1 U9530 ( .A1(n7530), .A2(n6553), .ZN(n8730) );
  NAND2_X1 U9531 ( .A1(n8622), .A2(n8621), .ZN(n8639) );
  NAND2_X1 U9532 ( .A1(n6986), .A2(n6985), .ZN(n8926) );
  INV_X1 U9533 ( .A(n8923), .ZN(n6985) );
  NAND2_X1 U9534 ( .A1(n8925), .A2(n8924), .ZN(n6986) );
  NAND3_X2 U9535 ( .A1(n8418), .A2(n8417), .A3(n8483), .ZN(n8579) );
  NAND3_X1 U9536 ( .A1(n8467), .A2(n9625), .A3(n8473), .ZN(n8475) );
  INV_X1 U9537 ( .A(n8881), .ZN(n8452) );
  NAND3_X1 U9538 ( .A1(n8423), .A2(n8424), .A3(n8422), .ZN(n8443) );
  NAND3_X1 U9539 ( .A1(n6987), .A2(n8521), .A3(n8520), .ZN(n6995) );
  NAND2_X1 U9540 ( .A1(n8494), .A2(n8493), .ZN(n6987) );
  NOR2_X2 U9541 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n8418) );
  NAND2_X1 U9542 ( .A1(n7650), .A2(n7345), .ZN(n8456) );
  NAND2_X1 U9543 ( .A1(n10053), .A2(n8922), .ZN(n8517) );
  NAND2_X1 U9544 ( .A1(n13460), .A2(n13347), .ZN(n13351) );
  NOR2_X1 U9545 ( .A1(n9073), .A2(n9072), .ZN(n9204) );
  OR2_X1 U9546 ( .A1(n8548), .A2(n8547), .ZN(n7661) );
  NAND2_X1 U9547 ( .A1(n6995), .A2(n8526), .ZN(n8548) );
  OAI22_X1 U9548 ( .A1(n7528), .A2(n8877), .B1(n8897), .B2(n7527), .ZN(n8925)
         );
  NOR2_X4 U9549 ( .A1(n8579), .A2(n8420), .ZN(n8421) );
  OAI21_X1 U9550 ( .B1(n8876), .B2(n8875), .A(n6499), .ZN(n7528) );
  MUX2_X1 U9551 ( .A(n9962), .B(n9279), .S(n11950), .Z(n8529) );
  NAND3_X1 U9552 ( .A1(n7695), .A2(n7694), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7002) );
  NAND2_X1 U9553 ( .A1(n7635), .A2(n7014), .ZN(n7012) );
  NAND2_X1 U9554 ( .A1(n14106), .A2(n7024), .ZN(n7021) );
  NAND2_X1 U9555 ( .A1(n7021), .A2(n7022), .ZN(n14045) );
  NAND2_X1 U9556 ( .A1(n9371), .A2(n9264), .ZN(n9711) );
  INV_X1 U9557 ( .A(n9361), .ZN(n9358) );
  NAND2_X1 U9558 ( .A1(n9269), .A2(n9265), .ZN(n7037) );
  NAND3_X1 U9559 ( .A1(n12162), .A2(n6550), .A3(n12161), .ZN(n7045) );
  INV_X1 U9560 ( .A(n7046), .ZN(n12206) );
  INV_X1 U9561 ( .A(n12203), .ZN(n7049) );
  NAND2_X1 U9562 ( .A1(n7050), .A2(n7053), .ZN(n12220) );
  NAND3_X1 U9563 ( .A1(n12215), .A2(n7051), .A3(n12214), .ZN(n7050) );
  NAND2_X1 U9564 ( .A1(n7055), .A2(n7058), .ZN(n12233) );
  NAND3_X1 U9565 ( .A1(n12225), .A2(n7056), .A3(n12224), .ZN(n7055) );
  NAND2_X1 U9566 ( .A1(n7061), .A2(n7060), .ZN(n7429) );
  NAND3_X1 U9567 ( .A1(n12128), .A2(n6555), .A3(n12127), .ZN(n7060) );
  OAI22_X1 U9568 ( .A1(n12137), .A2(n7067), .B1(n12138), .B2(n7069), .ZN(
        n12142) );
  NAND2_X1 U9569 ( .A1(n12152), .A2(n7073), .ZN(n7070) );
  OAI21_X1 U9570 ( .B1(n12152), .B2(n7074), .A(n7073), .ZN(n12157) );
  NAND2_X1 U9571 ( .A1(n7070), .A2(n7071), .ZN(n12156) );
  MUX2_X1 U9572 ( .A(n14164), .B(n14711), .S(n9958), .Z(n14999) );
  NAND2_X1 U9573 ( .A1(n8879), .A2(n7080), .ZN(n7076) );
  NAND2_X1 U9574 ( .A1(n7076), .A2(n7077), .ZN(n8953) );
  NAND2_X1 U9575 ( .A1(n8879), .A2(n8878), .ZN(n7079) );
  NAND2_X1 U9576 ( .A1(n8708), .A2(n8707), .ZN(n7083) );
  NAND2_X1 U9577 ( .A1(n8578), .A2(n6454), .ZN(n7097) );
  NAND2_X1 U9578 ( .A1(n8578), .A2(n8577), .ZN(n8595) );
  NAND3_X1 U9579 ( .A1(n7097), .A2(n8641), .A3(n7096), .ZN(n8645) );
  NAND4_X1 U9580 ( .A1(n14427), .A2(n14416), .A3(n7099), .A4(n12040), .ZN(
        n7098) );
  NAND2_X1 U9581 ( .A1(n14946), .A2(n7113), .ZN(n7108) );
  NAND3_X1 U9582 ( .A1(n7109), .A2(n7108), .A3(n7110), .ZN(n14797) );
  OR2_X2 U9583 ( .A1(n9940), .A2(n10644), .ZN(n10024) );
  NAND2_X1 U9584 ( .A1(n13670), .A2(n7120), .ZN(n13574) );
  NAND2_X1 U9585 ( .A1(n11336), .A2(n11335), .ZN(n11463) );
  NAND2_X1 U9586 ( .A1(n7129), .A2(n7127), .ZN(n14303) );
  NAND2_X1 U9587 ( .A1(n10248), .A2(n12116), .ZN(n7406) );
  NAND2_X1 U9588 ( .A1(n7133), .A2(n6539), .ZN(n10278) );
  NOR2_X1 U9589 ( .A1(n7399), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U9590 ( .A1(n14290), .A2(n7142), .ZN(n7141) );
  NAND2_X1 U9591 ( .A1(n7611), .A2(n9371), .ZN(n9725) );
  OAI21_X1 U9592 ( .B1(n12560), .B2(n7151), .A(n7148), .ZN(n12519) );
  NAND2_X1 U9593 ( .A1(n12560), .A2(n7148), .ZN(n7147) );
  OAI21_X1 U9594 ( .B1(n12560), .B2(n12474), .A(n7154), .ZN(n12616) );
  NAND2_X1 U9595 ( .A1(n12624), .A2(n13004), .ZN(n7168) );
  NAND2_X1 U9596 ( .A1(n12624), .A2(n7157), .ZN(n7156) );
  NAND3_X1 U9597 ( .A1(n7156), .A2(n7155), .A3(n7165), .ZN(n12542) );
  INV_X1 U9598 ( .A(n12502), .ZN(n7174) );
  NAND2_X1 U9599 ( .A1(n11566), .A2(n11565), .ZN(n12468) );
  NAND2_X1 U9600 ( .A1(n12468), .A2(n12467), .ZN(n12470) );
  INV_X1 U9601 ( .A(n10864), .ZN(n7177) );
  OAI21_X2 U9602 ( .B1(n12608), .B2(n7181), .A(n7178), .ZN(n12501) );
  OR2_X2 U9603 ( .A1(n8028), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U9604 ( .A1(n8390), .A2(n6541), .ZN(n8397) );
  NAND2_X1 U9605 ( .A1(n8390), .A2(n7183), .ZN(n8395) );
  NAND2_X1 U9606 ( .A1(n8397), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8393) );
  MUX2_X1 U9607 ( .A(n11130), .B(n11119), .S(n11143), .Z(n11087) );
  MUX2_X1 U9608 ( .A(n15297), .B(n15315), .S(n11143), .Z(n11097) );
  MUX2_X1 U9609 ( .A(n11101), .B(n11102), .S(n11143), .Z(n11103) );
  MUX2_X1 U9610 ( .A(n11110), .B(n11111), .S(n11143), .Z(n11112) );
  MUX2_X1 U9611 ( .A(n15303), .B(n11155), .S(n11143), .Z(n11157) );
  MUX2_X1 U9612 ( .A(n11186), .B(n15204), .S(n11143), .Z(n11187) );
  MUX2_X1 U9613 ( .A(P3_REG1_REG_11__SCAN_IN), .B(P3_REG2_REG_11__SCAN_IN), 
        .S(n11143), .Z(n11709) );
  MUX2_X1 U9614 ( .A(P3_REG1_REG_13__SCAN_IN), .B(P3_REG2_REG_13__SCAN_IN), 
        .S(n11143), .Z(n12772) );
  MUX2_X1 U9615 ( .A(P3_REG1_REG_14__SCAN_IN), .B(P3_REG2_REG_14__SCAN_IN), 
        .S(n11143), .Z(n12781) );
  MUX2_X1 U9616 ( .A(P3_REG1_REG_15__SCAN_IN), .B(P3_REG2_REG_15__SCAN_IN), 
        .S(n11143), .Z(n12782) );
  MUX2_X1 U9617 ( .A(n13195), .B(n13078), .S(n11143), .Z(n12811) );
  MUX2_X1 U9618 ( .A(P3_REG1_REG_17__SCAN_IN), .B(P3_REG2_REG_17__SCAN_IN), 
        .S(n11143), .Z(n12845) );
  MUX2_X1 U9619 ( .A(n12879), .B(n12884), .S(n11143), .Z(n12880) );
  MUX2_X1 U9620 ( .A(n12773), .B(n12794), .S(n11143), .Z(n12774) );
  AOI21_X1 U9621 ( .B1(n11143), .B2(P3_STATE_REG_SCAN_IN), .A(n7185), .ZN(
        n7184) );
  NAND2_X1 U9622 ( .A1(n11304), .A2(n7193), .ZN(n7189) );
  INV_X1 U9623 ( .A(n8302), .ZN(n7206) );
  INV_X1 U9624 ( .A(n12922), .ZN(n7213) );
  NAND2_X1 U9625 ( .A1(n12922), .A2(n7220), .ZN(n7214) );
  AOI21_X1 U9626 ( .B1(n12922), .B2(n12921), .A(n8370), .ZN(n12902) );
  OAI21_X1 U9627 ( .B1(n13016), .B2(n13017), .A(n8336), .ZN(n13012) );
  NAND2_X1 U9628 ( .A1(n7228), .A2(n8407), .ZN(P3_U3296) );
  NAND2_X1 U9629 ( .A1(n8233), .A2(n8232), .ZN(n7230) );
  NAND2_X1 U9630 ( .A1(n7752), .A2(n7751), .ZN(n7754) );
  INV_X1 U9631 ( .A(n7734), .ZN(n7231) );
  INV_X1 U9632 ( .A(n7260), .ZN(n12805) );
  INV_X1 U9633 ( .A(n7265), .ZN(n12765) );
  INV_X1 U9634 ( .A(n12785), .ZN(n12784) );
  NAND2_X1 U9635 ( .A1(n7265), .A2(n7264), .ZN(n12785) );
  OAI21_X1 U9636 ( .B1(n8177), .B2(n7268), .A(n7266), .ZN(n8180) );
  OAI21_X1 U9637 ( .B1(n8177), .B2(n8176), .A(n8178), .ZN(n8190) );
  AOI21_X1 U9638 ( .B1(n8176), .B2(n8178), .A(n6593), .ZN(n7269) );
  NAND3_X1 U9639 ( .A1(n8385), .A2(n6446), .A3(n8380), .ZN(n7270) );
  NAND2_X1 U9640 ( .A1(n9281), .A2(n7272), .ZN(n9284) );
  NOR2_X1 U9641 ( .A1(n10045), .A2(n15061), .ZN(n7273) );
  AND2_X1 U9642 ( .A1(n6551), .A2(n7278), .ZN(n7277) );
  NAND3_X1 U9643 ( .A1(n7275), .A2(n7276), .A3(n6556), .ZN(n7274) );
  AND2_X2 U9644 ( .A1(n7276), .A2(n7279), .ZN(n9371) );
  NOR2_X1 U9645 ( .A1(n9298), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9305) );
  INV_X1 U9646 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U9647 ( .A1(n7287), .A2(n7288), .ZN(n13776) );
  AND2_X4 U9648 ( .A1(n8416), .A2(n8415), .ZN(n7650) );
  OAI21_X1 U9649 ( .B1(n13749), .B2(n7311), .A(n7308), .ZN(n13713) );
  NAND2_X4 U9650 ( .A1(n9664), .A2(n9647), .ZN(n9828) );
  INV_X1 U9651 ( .A(n13332), .ZN(n13364) );
  INV_X1 U9652 ( .A(n7656), .ZN(n7318) );
  AOI21_X1 U9653 ( .B1(n7318), .B2(n13427), .A(n13337), .ZN(n7317) );
  NAND2_X1 U9654 ( .A1(n11003), .A2(n7335), .ZN(n11006) );
  NAND2_X1 U9655 ( .A1(n13462), .A2(n6436), .ZN(n7341) );
  NAND2_X1 U9656 ( .A1(n7341), .A2(n7342), .ZN(n13379) );
  AND2_X1 U9657 ( .A1(n8421), .A2(n8451), .ZN(n7345) );
  NAND2_X1 U9658 ( .A1(n7346), .A2(n7650), .ZN(n8464) );
  AND2_X1 U9659 ( .A1(n6545), .A2(n8451), .ZN(n7347) );
  NAND2_X1 U9660 ( .A1(n9688), .A2(n9689), .ZN(n9827) );
  AOI21_X1 U9661 ( .B1(n12818), .B2(n12832), .A(n7366), .ZN(n12850) );
  NAND2_X1 U9662 ( .A1(n12747), .A2(n6585), .ZN(n7375) );
  INV_X1 U9663 ( .A(n11123), .ZN(n7383) );
  NAND2_X1 U9664 ( .A1(n11760), .A2(n7614), .ZN(n11762) );
  NAND2_X1 U9665 ( .A1(n11533), .A2(n12015), .ZN(n7385) );
  NAND2_X1 U9666 ( .A1(n7390), .A2(n7389), .ZN(n14453) );
  OR2_X2 U9667 ( .A1(n14303), .A2(n7628), .ZN(n7401) );
  AND2_X2 U9668 ( .A1(n12098), .A2(n12079), .ZN(n12131) );
  NAND2_X1 U9669 ( .A1(n12210), .A2(n12211), .ZN(n12209) );
  MUX2_X1 U9670 ( .A(n12104), .B(n12107), .S(n12131), .Z(n7413) );
  INV_X1 U9671 ( .A(n12180), .ZN(n7418) );
  NAND2_X1 U9672 ( .A1(n7424), .A2(n7425), .ZN(n12152) );
  NAND3_X1 U9673 ( .A1(n12147), .A2(n6554), .A3(n12146), .ZN(n7424) );
  NAND3_X1 U9674 ( .A1(n12200), .A2(n12199), .A3(n6548), .ZN(n7427) );
  NAND2_X1 U9675 ( .A1(n7429), .A2(n7430), .ZN(n12137) );
  NAND2_X1 U9676 ( .A1(n9371), .A2(n7434), .ZN(n9709) );
  NAND2_X1 U9677 ( .A1(n9371), .A2(n6478), .ZN(n9707) );
  NAND2_X1 U9678 ( .A1(n9709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9356) );
  INV_X1 U9679 ( .A(n9057), .ZN(n7439) );
  NAND2_X1 U9680 ( .A1(n7439), .A2(n6574), .ZN(n7442) );
  NAND2_X1 U9681 ( .A1(n7442), .A2(n7440), .ZN(n9078) );
  NAND2_X1 U9682 ( .A1(n8666), .A2(n7455), .ZN(n7452) );
  OAI21_X1 U9683 ( .B1(n8738), .B2(n7463), .A(n7460), .ZN(n8783) );
  AOI21_X1 U9684 ( .B1(n7460), .B2(n7463), .A(n7459), .ZN(n7458) );
  OAI21_X1 U9685 ( .B1(n8527), .B2(n7465), .A(n8531), .ZN(n8552) );
  NAND2_X1 U9686 ( .A1(n7469), .A2(n7466), .ZN(n8555) );
  NAND2_X1 U9687 ( .A1(n8527), .A2(n8531), .ZN(n7469) );
  INV_X1 U9688 ( .A(n8785), .ZN(n7470) );
  NAND2_X1 U9689 ( .A1(n8979), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U9690 ( .A1(n9132), .A2(n9131), .ZN(n7491) );
  NAND2_X1 U9691 ( .A1(n12446), .A2(n12445), .ZN(n12976) );
  INV_X1 U9692 ( .A(n7500), .ZN(n12975) );
  INV_X1 U9693 ( .A(n12445), .ZN(n7502) );
  AND2_X1 U9694 ( .A1(n12974), .A2(n12988), .ZN(n7503) );
  NAND2_X1 U9695 ( .A1(n7519), .A2(n6546), .ZN(n13045) );
  NAND2_X1 U9696 ( .A1(n7521), .A2(n7520), .ZN(n13003) );
  NAND3_X1 U9697 ( .A1(n8687), .A2(n8686), .A3(n6557), .ZN(n7530) );
  INV_X1 U9698 ( .A(n8705), .ZN(n7532) );
  NAND3_X1 U9699 ( .A1(n8976), .A2(n8975), .A3(n6558), .ZN(n7533) );
  AOI22_X1 U9700 ( .A1(n7537), .A2(n7539), .B1(n6461), .B2(n7543), .ZN(n7536)
         );
  OR2_X1 U9701 ( .A1(n7543), .A2(n6465), .ZN(n7539) );
  NOR2_X1 U9702 ( .A1(n8456), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n8459) );
  INV_X1 U9703 ( .A(n8663), .ZN(n7548) );
  NOR2_X1 U9704 ( .A1(n7551), .A2(n10781), .ZN(n10634) );
  OAI211_X1 U9705 ( .C1(n14125), .C2(n7567), .A(n7563), .B(n7561), .ZN(n12415)
         );
  NAND2_X1 U9706 ( .A1(n14125), .A2(n7562), .ZN(n7561) );
  OAI21_X1 U9707 ( .B1(n7568), .B2(n7572), .A(n7564), .ZN(n7563) );
  NAND2_X1 U9708 ( .A1(n7568), .A2(n7565), .ZN(n7564) );
  NAND2_X1 U9709 ( .A1(n10042), .A2(n6447), .ZN(n7578) );
  NAND2_X1 U9710 ( .A1(n6447), .A2(n10036), .ZN(n7579) );
  NOR2_X1 U9711 ( .A1(n11059), .A2(n11060), .ZN(n7589) );
  NAND3_X2 U9712 ( .A1(n7594), .A2(n7593), .A3(n9728), .ZN(n15002) );
  AND2_X2 U9713 ( .A1(n9726), .A2(n14697), .ZN(n10484) );
  AND2_X2 U9714 ( .A1(n9726), .A2(n9727), .ZN(n11974) );
  INV_X1 U9715 ( .A(n10458), .ZN(n7608) );
  NAND3_X1 U9716 ( .A1(n7604), .A2(n7603), .A3(n10268), .ZN(n10272) );
  NAND2_X1 U9717 ( .A1(n14458), .A2(n7621), .ZN(n14274) );
  NAND2_X1 U9718 ( .A1(n7630), .A2(n7629), .ZN(n9672) );
  OR2_X1 U9719 ( .A1(n9667), .A2(n9666), .ZN(n7629) );
  NAND2_X1 U9720 ( .A1(n9667), .A2(n9666), .ZN(n7630) );
  NAND2_X1 U9721 ( .A1(n13697), .A2(n7634), .ZN(n7632) );
  NAND4_X1 U9722 ( .A1(n8421), .A2(n7649), .A3(n7650), .A4(n8442), .ZN(n8429)
         );
  NAND2_X1 U9723 ( .A1(n13213), .A2(n10660), .ZN(n13212) );
  NAND2_X1 U9724 ( .A1(n11453), .A2(n11452), .ZN(n11566) );
  INV_X1 U9725 ( .A(n11455), .ZN(n11453) );
  CLKBUF_X1 U9726 ( .A(n10415), .Z(n10610) );
  NAND2_X1 U9727 ( .A1(n9642), .A2(n9641), .ZN(n10415) );
  XNOR2_X1 U9728 ( .A(n12931), .B(n12933), .ZN(n13148) );
  XNOR2_X2 U9729 ( .A(n12501), .B(n12499), .ZN(n12624) );
  INV_X1 U9730 ( .A(n13222), .ZN(n7714) );
  NAND4_X2 U9731 ( .A1(n9732), .A2(n9731), .A3(n9730), .A4(n9729), .ZN(n15006)
         );
  AND2_X1 U9732 ( .A1(n12167), .A2(n12229), .ZN(n12181) );
  INV_X1 U9733 ( .A(n8803), .ZN(n8806) );
  AND4_X1 U9734 ( .A1(n8414), .A2(n8413), .A3(n8648), .A4(n8412), .ZN(n8415)
         );
  NAND2_X1 U9735 ( .A1(n8401), .A2(n8400), .ZN(n11301) );
  INV_X1 U9736 ( .A(n12113), .ZN(n12002) );
  AOI21_X1 U9737 ( .B1(n9252), .B2(n7653), .A(n9251), .ZN(n9253) );
  INV_X1 U9738 ( .A(n12693), .ZN(n7715) );
  NAND2_X1 U9739 ( .A1(n10036), .A2(n9866), .ZN(n9870) );
  OR2_X1 U9740 ( .A1(n12037), .A2(n9735), .ZN(n9731) );
  AND2_X1 U9741 ( .A1(n9233), .A2(n10304), .ZN(n7653) );
  OR2_X1 U9742 ( .A1(n14662), .A2(n14350), .ZN(n7654) );
  AND4_X1 U9743 ( .A1(n7678), .A2(n8209), .A3(n7677), .A4(n8392), .ZN(n7657)
         );
  AND4_X1 U9744 ( .A1(n8075), .A2(n8074), .A3(n8073), .A4(n8072), .ZN(n13004)
         );
  INV_X1 U9745 ( .A(n13004), .ZN(n12443) );
  XOR2_X1 U9746 ( .A(P2_IR_REG_27__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .Z(
        n7658) );
  AND2_X1 U9747 ( .A1(n8784), .A2(n8768), .ZN(n7659) );
  NAND2_X1 U9748 ( .A1(n8149), .A2(n8148), .ZN(n12677) );
  AND2_X1 U9749 ( .A1(n11191), .A2(n11165), .ZN(n7662) );
  INV_X1 U9750 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7838) );
  AND2_X1 U9751 ( .A1(n12716), .A2(n11114), .ZN(n7663) );
  OR2_X1 U9752 ( .A1(n9252), .A2(n9206), .ZN(n7664) );
  OR2_X1 U9753 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11658), .ZN(n7665) );
  AND2_X1 U9754 ( .A1(n8765), .A2(n8741), .ZN(n7666) );
  INV_X1 U9755 ( .A(n13011), .ZN(n12441) );
  NAND2_X2 U9756 ( .A1(n10303), .A2(n13841), .ZN(n13844) );
  NAND2_X1 U9757 ( .A1(n9768), .A2(n9767), .ZN(n15185) );
  AND2_X1 U9758 ( .A1(n8927), .A2(n8932), .ZN(n7668) );
  INV_X1 U9759 ( .A(n13920), .ZN(n13566) );
  INV_X1 U9760 ( .A(n12464), .ZN(n13238) );
  INV_X1 U9761 ( .A(n12961), .ZN(n8104) );
  INV_X1 U9762 ( .A(n13330), .ZN(n13328) );
  INV_X1 U9763 ( .A(n13257), .ZN(n12996) );
  AND2_X1 U9764 ( .A1(n12954), .A2(n12679), .ZN(n7669) );
  AND2_X2 U9765 ( .A1(n10659), .A2(n15234), .ZN(n15250) );
  OAI21_X1 U9766 ( .B1(n12111), .B2(n12131), .A(n12110), .ZN(n12112) );
  NAND2_X1 U9767 ( .A1(n12117), .A2(n12116), .ZN(n12121) );
  NAND2_X1 U9768 ( .A1(n8798), .A2(n8797), .ZN(n8804) );
  INV_X1 U9769 ( .A(n8804), .ZN(n8805) );
  OAI21_X1 U9770 ( .B1(n12179), .B2(n12178), .A(n12177), .ZN(n12180) );
  INV_X1 U9771 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U9772 ( .A1(n9232), .A2(n8481), .ZN(n9097) );
  INV_X1 U9773 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7675) );
  INV_X1 U9774 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8413) );
  INV_X1 U9775 ( .A(n12919), .ZN(n12449) );
  INV_X1 U9776 ( .A(n7792), .ZN(n7733) );
  INV_X1 U9777 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U9778 ( .A1(n8097), .A2(n8096), .ZN(n8112) );
  INV_X1 U9779 ( .A(n8035), .ZN(n8034) );
  NAND2_X1 U9780 ( .A1(n13139), .A2(n12449), .ZN(n12450) );
  OR2_X1 U9781 ( .A1(n7699), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9782 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  INV_X1 U9783 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U9784 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  INV_X1 U9785 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8604) );
  INV_X1 U9786 ( .A(n13730), .ZN(n13752) );
  INV_X1 U9787 ( .A(n10962), .ZN(n9668) );
  OR2_X1 U9788 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  INV_X1 U9789 ( .A(n8899), .ZN(n8929) );
  INV_X1 U9790 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9263) );
  INV_X1 U9791 ( .A(n11456), .ZN(n11452) );
  OR2_X1 U9792 ( .A1(n8126), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8142) );
  OR2_X1 U9793 ( .A1(n8081), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8098) );
  INV_X1 U9794 ( .A(n11222), .ZN(n11138) );
  AND2_X1 U9795 ( .A1(n8344), .A2(n8345), .ZN(n12986) );
  INV_X1 U9796 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11714) );
  OR2_X1 U9797 ( .A1(n10616), .A2(n10764), .ZN(n10652) );
  INV_X1 U9798 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U9799 ( .A1(n9170), .A2(n9187), .ZN(n9203) );
  AND2_X1 U9800 ( .A1(n8910), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8937) );
  INV_X1 U9801 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11555) );
  INV_X1 U9802 ( .A(n13964), .ZN(n13567) );
  INV_X1 U9803 ( .A(n11678), .ZN(n11359) );
  INV_X1 U9804 ( .A(n8786), .ZN(n9089) );
  INV_X1 U9805 ( .A(n9231), .ZN(n8481) );
  INV_X1 U9806 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8460) );
  INV_X1 U9807 ( .A(n10946), .ZN(n10947) );
  AND2_X1 U9808 ( .A1(n14320), .A2(n12072), .ZN(n9752) );
  AND2_X1 U9809 ( .A1(n10084), .A2(n10083), .ZN(n10087) );
  NAND2_X1 U9810 ( .A1(n10923), .A2(n9756), .ZN(n12068) );
  INV_X1 U9811 ( .A(n12072), .ZN(n9756) );
  INV_X1 U9812 ( .A(n14527), .ZN(n14509) );
  INV_X1 U9813 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14715) );
  NOR2_X1 U9814 ( .A1(n14787), .A2(n14786), .ZN(n14731) );
  INV_X1 U9815 ( .A(n12677), .ZN(n12934) );
  OR2_X1 U9816 ( .A1(n10589), .A2(n10411), .ZN(n12659) );
  OR2_X1 U9817 ( .A1(n8156), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8169) );
  INV_X1 U9818 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11736) );
  INV_X1 U9819 ( .A(n15191), .ZN(n12849) );
  INV_X1 U9820 ( .A(n12679), .ZN(n12964) );
  AND4_X1 U9821 ( .A1(n8064), .A2(n8063), .A3(n8062), .A4(n8061), .ZN(n13020)
         );
  INV_X1 U9822 ( .A(n13100), .ZN(n13074) );
  INV_X1 U9823 ( .A(n14857), .ZN(n15212) );
  NAND2_X1 U9824 ( .A1(n7839), .A2(n7838), .ZN(n7859) );
  INV_X1 U9825 ( .A(n13296), .ZN(n10620) );
  OR2_X1 U9826 ( .A1(n12895), .A2(n12894), .ZN(n13126) );
  INV_X1 U9827 ( .A(n11013), .ZN(n10909) );
  NOR2_X1 U9828 ( .A1(n10401), .A2(n10616), .ZN(n10592) );
  AND2_X1 U9829 ( .A1(n7795), .A2(n7776), .ZN(n7793) );
  NAND2_X1 U9830 ( .A1(n8818), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8865) );
  OR2_X1 U9831 ( .A1(n8865), .A2(n8864), .ZN(n8885) );
  NOR2_X1 U9832 ( .A1(n15379), .A2(n8984), .ZN(n8999) );
  INV_X1 U9833 ( .A(n14885), .ZN(n13447) );
  INV_X1 U9834 ( .A(n9250), .ZN(n9251) );
  AND2_X1 U9835 ( .A1(n8937), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8958) );
  NOR2_X1 U9836 ( .A1(n8775), .A2(n11555), .ZN(n8790) );
  OR2_X1 U9837 ( .A1(n13824), .A2(n13930), .ZN(n13825) );
  INV_X1 U9838 ( .A(n10548), .ZN(n10554) );
  XNOR2_X1 U9839 ( .A(n13489), .B(n9644), .ZN(n9666) );
  AND3_X1 U9840 ( .A1(n9658), .A2(n15176), .A3(n9657), .ZN(n10300) );
  OR2_X1 U9841 ( .A1(n10540), .A2(n9621), .ZN(n11874) );
  INV_X1 U9842 ( .A(n11360), .ZN(n11416) );
  INV_X1 U9843 ( .A(n11346), .ZN(n11420) );
  INV_X1 U9844 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U9845 ( .A1(n12105), .A2(n9752), .ZN(n10786) );
  OR2_X1 U9846 ( .A1(n10749), .A2(n10748), .ZN(n10828) );
  NAND2_X1 U9847 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  OR2_X1 U9848 ( .A1(n10188), .A2(n9724), .ZN(n14111) );
  AND2_X1 U9849 ( .A1(n12047), .A2(n12046), .ZN(n14355) );
  NOR2_X1 U9850 ( .A1(n11998), .A2(n15413), .ZN(n11984) );
  INV_X1 U9851 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14725) );
  OR2_X1 U9852 ( .A1(n10152), .A2(n10153), .ZN(n10979) );
  INV_X1 U9853 ( .A(n10923), .ZN(n12077) );
  INV_X1 U9854 ( .A(n12069), .ZN(n9871) );
  INV_X1 U9855 ( .A(n12012), .ZN(n10839) );
  INV_X1 U9856 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U9857 ( .A1(n8853), .A2(n8852), .ZN(n8879) );
  INV_X1 U9858 ( .A(n12988), .ZN(n12965) );
  INV_X1 U9859 ( .A(n12674), .ZN(n12644) );
  INV_X1 U9860 ( .A(n7744), .ZN(n8170) );
  AND4_X1 U9861 ( .A1(n8050), .A2(n8049), .A3(n8048), .A4(n8047), .ZN(n13028)
         );
  INV_X1 U9862 ( .A(n12888), .ZN(n12835) );
  INV_X1 U9863 ( .A(n12892), .ZN(n12864) );
  AND2_X1 U9864 ( .A1(P3_U3897), .A2(n8404), .ZN(n12890) );
  INV_X1 U9865 ( .A(n8362), .ZN(n12933) );
  INV_X1 U9866 ( .A(n13125), .ZN(n14847) );
  AND2_X1 U9867 ( .A1(n11070), .A2(n15287), .ZN(n10658) );
  INV_X1 U9868 ( .A(n10917), .ZN(n15228) );
  AND2_X1 U9869 ( .A1(n15248), .A2(n15238), .ZN(n15246) );
  AND2_X1 U9870 ( .A1(n10613), .A2(n10612), .ZN(n10657) );
  AND2_X1 U9871 ( .A1(n13203), .A2(n13202), .ZN(n13287) );
  INV_X1 U9872 ( .A(n13152), .ZN(n14874) );
  INV_X1 U9873 ( .A(n13143), .ZN(n15289) );
  NAND2_X1 U9874 ( .A1(n10777), .A2(n10416), .ZN(n15281) );
  INV_X1 U9875 ( .A(n14891), .ZN(n13449) );
  AND2_X1 U9876 ( .A1(n9410), .A2(n9409), .ZN(n15155) );
  AND2_X1 U9877 ( .A1(n9404), .A2(n9425), .ZN(n15158) );
  AND2_X1 U9878 ( .A1(n9159), .A2(n9158), .ZN(n13653) );
  AND2_X1 U9879 ( .A1(n13586), .A2(n13585), .ZN(n13793) );
  INV_X1 U9880 ( .A(n13816), .ZN(n13846) );
  AND2_X1 U9881 ( .A1(n13844), .A2(n9628), .ZN(n13850) );
  AND2_X1 U9882 ( .A1(n15170), .A2(n10300), .ZN(n9660) );
  INV_X1 U9883 ( .A(n11874), .ZN(n15179) );
  AND2_X1 U9884 ( .A1(n9664), .A2(n13891), .ZN(n15182) );
  INV_X1 U9885 ( .A(n15182), .ZN(n13905) );
  AND2_X1 U9886 ( .A1(n8671), .A2(n8714), .ZN(n9912) );
  OR2_X1 U9887 ( .A1(n11488), .A2(n11487), .ZN(n11773) );
  INV_X1 U9888 ( .A(n14927), .ZN(n14131) );
  INV_X1 U9889 ( .A(n10484), .ZN(n11900) );
  AND2_X1 U9890 ( .A1(n11979), .A2(n11978), .ZN(n14471) );
  INV_X1 U9891 ( .A(n11974), .ZN(n11779) );
  INV_X1 U9892 ( .A(n14987), .ZN(n14245) );
  INV_X1 U9893 ( .A(n14992), .ZN(n14219) );
  INV_X1 U9894 ( .A(n14983), .ZN(n14243) );
  INV_X1 U9895 ( .A(n14640), .ZN(n15016) );
  NAND2_X1 U9896 ( .A1(n14339), .A2(n7654), .ZN(n14286) );
  NAND2_X1 U9897 ( .A1(n10192), .A2(n14544), .ZN(n14541) );
  INV_X1 U9898 ( .A(n14630), .ZN(n11847) );
  NAND2_X1 U9899 ( .A1(n12076), .A2(n12074), .ZN(n15079) );
  NAND2_X1 U9900 ( .A1(n9377), .A2(n9378), .ZN(n9705) );
  AND2_X1 U9901 ( .A1(n10531), .A2(n10812), .ZN(n11992) );
  AND2_X1 U9902 ( .A1(n9463), .A2(n9388), .ZN(n10821) );
  AND2_X1 U9903 ( .A1(n11129), .A2(n11128), .ZN(n15191) );
  NAND2_X1 U9904 ( .A1(n10400), .A2(n10658), .ZN(n12652) );
  AND2_X1 U9905 ( .A1(n8202), .A2(n8201), .ZN(n12454) );
  INV_X1 U9906 ( .A(n12692), .ZN(n12680) );
  INV_X1 U9907 ( .A(n13119), .ZN(n12686) );
  NOR2_X2 U9908 ( .A1(n10394), .A2(n11882), .ZN(n12692) );
  OR2_X1 U9909 ( .A1(n11144), .A2(n11118), .ZN(n12888) );
  INV_X1 U9910 ( .A(n12890), .ZN(n12868) );
  AND2_X1 U9911 ( .A1(n13102), .A2(n13101), .ZN(n13202) );
  NAND2_X1 U9912 ( .A1(n10658), .A2(n15232), .ZN(n15234) );
  INV_X1 U9913 ( .A(n15246), .ZN(n12945) );
  INV_X1 U9914 ( .A(n15308), .ZN(n15306) );
  AND2_X1 U9915 ( .A1(n15274), .A2(n15273), .ZN(n15302) );
  AND2_X1 U9916 ( .A1(n10595), .A2(n10594), .ZN(n15295) );
  OR2_X1 U9917 ( .A1(n11883), .A2(n11882), .ZN(n15425) );
  INV_X1 U9918 ( .A(SI_14_), .ZN(n9391) );
  INV_X1 U9919 ( .A(SI_10_), .ZN(n9294) );
  INV_X1 U9920 ( .A(n10606), .ZN(n11891) );
  INV_X1 U9921 ( .A(n9631), .ZN(n13452) );
  OR2_X1 U9922 ( .A1(n9426), .A2(n9425), .ZN(n13556) );
  INV_X1 U9923 ( .A(n15155), .ZN(n15143) );
  INV_X1 U9924 ( .A(n15158), .ZN(n15129) );
  NAND2_X1 U9925 ( .A1(n13844), .A2(n10306), .ZN(n13835) );
  INV_X1 U9926 ( .A(n15190), .ZN(n15188) );
  INV_X1 U9927 ( .A(n13705), .ZN(n13960) );
  INV_X1 U9928 ( .A(n13763), .ZN(n13975) );
  NOR2_X1 U9929 ( .A1(n15173), .A2(n15167), .ZN(n15168) );
  AND2_X1 U9930 ( .A1(n9634), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15176) );
  XNOR2_X1 U9931 ( .A(n9237), .B(n9236), .ZN(n14002) );
  AND2_X1 U9932 ( .A1(n9373), .A2(n9490), .ZN(n14977) );
  OR2_X1 U9933 ( .A1(n14913), .A2(n15072), .ZN(n14927) );
  INV_X1 U9934 ( .A(n14297), .ZN(n14489) );
  OR2_X1 U9935 ( .A1(n14980), .A2(n12253), .ZN(n14987) );
  OR2_X1 U9936 ( .A1(n14980), .A2(n9895), .ZN(n14992) );
  OR3_X1 U9937 ( .A1(n15022), .A2(n12072), .A3(n12091), .ZN(n15012) );
  OR2_X1 U9938 ( .A1(n15022), .A2(n10194), .ZN(n14520) );
  INV_X1 U9939 ( .A(n15123), .ZN(n15120) );
  INV_X1 U9940 ( .A(n14655), .ZN(n15109) );
  INV_X2 U9941 ( .A(n15109), .ZN(n15111) );
  INV_X1 U9942 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10532) );
  INV_X1 U9943 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9763) );
  INV_X1 U9944 ( .A(n12680), .ZN(P3_U3897) );
  NOR2_X1 U9945 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7678) );
  INV_X1 U9946 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U9947 ( .A1(n7683), .A2(n7680), .ZN(n13299) );
  INV_X1 U9948 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7681) );
  XNOR2_X2 U9949 ( .A(n7682), .B(n7681), .ZN(n7685) );
  NAND2_X1 U9950 ( .A1(n8194), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7691) );
  INV_X1 U9951 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10407) );
  OR2_X1 U9952 ( .A1(n7744), .A2(n10407), .ZN(n7690) );
  INV_X1 U9953 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11084) );
  NAND2_X4 U9954 ( .A1(n7687), .A2(n12417), .ZN(n8199) );
  INV_X1 U9955 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11085) );
  OR2_X1 U9956 ( .A1(n8199), .A2(n11085), .ZN(n7688) );
  INV_X1 U9957 ( .A(n7722), .ZN(n7693) );
  INV_X1 U9958 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U9959 ( .A1(n9714), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9960 ( .A1(n7693), .A2(n7692), .ZN(n7698) );
  MUX2_X1 U9961 ( .A(n7698), .B(SI_0_), .S(n11950), .Z(n13305) );
  XNOR2_X2 U9962 ( .A(n7701), .B(n7700), .ZN(n8404) );
  MUX2_X1 U9963 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13305), .S(n11076), .Z(n10660)
         );
  INV_X1 U9964 ( .A(n10660), .ZN(n10626) );
  INV_X1 U9965 ( .A(n13219), .ZN(n7713) );
  NAND2_X1 U9966 ( .A1(n8195), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7709) );
  INV_X1 U9967 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11079) );
  INV_X1 U9968 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7705) );
  INV_X1 U9969 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11624) );
  OR2_X1 U9970 ( .A1(n7744), .A2(n11624), .ZN(n7706) );
  NAND2_X1 U9971 ( .A1(n7721), .A2(SI_1_), .ZN(n7712) );
  XNOR2_X1 U9972 ( .A(n7723), .B(n7722), .ZN(n9330) );
  NAND2_X1 U9973 ( .A1(n7792), .A2(n9330), .ZN(n7711) );
  INV_X1 U9974 ( .A(n11629), .ZN(n11080) );
  NAND2_X1 U9975 ( .A1(n8030), .A2(n11080), .ZN(n7710) );
  NAND2_X1 U9976 ( .A1(n12693), .A2(n13222), .ZN(n8237) );
  NAND2_X1 U9977 ( .A1(n7713), .A2(n8237), .ZN(n10424) );
  NAND2_X1 U9978 ( .A1(n10424), .A2(n8216), .ZN(n10763) );
  NAND2_X1 U9979 ( .A1(n8195), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7720) );
  INV_X1 U9980 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7716) );
  OR2_X1 U9981 ( .A1(n8184), .A2(n7716), .ZN(n7719) );
  INV_X1 U9982 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11119) );
  OR2_X1 U9983 ( .A1(n8199), .A2(n11119), .ZN(n7718) );
  INV_X1 U9984 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10585) );
  OR2_X1 U9985 ( .A1(n7744), .A2(n10585), .ZN(n7717) );
  NAND4_X2 U9986 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n13214)
         );
  NAND2_X1 U9987 ( .A1(n9313), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U9988 ( .A1(n9279), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U9989 ( .A1(n9962), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U9990 ( .A1(n7736), .A2(n7725), .ZN(n7734) );
  XNOR2_X1 U9991 ( .A(n7735), .B(n7734), .ZN(n9340) );
  NAND2_X1 U9992 ( .A1(n7792), .A2(n9340), .ZN(n7728) );
  NAND2_X1 U9993 ( .A1(n6432), .A2(n11299), .ZN(n7727) );
  OR2_X1 U9994 ( .A1(n13214), .A2(n10576), .ZN(n8250) );
  NAND2_X1 U9995 ( .A1(n6428), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7732) );
  OR2_X1 U9996 ( .A1(n7744), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n7731) );
  INV_X1 U9997 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11090) );
  INV_X1 U9998 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11091) );
  OR2_X1 U9999 ( .A1(n8199), .A2(n11091), .ZN(n7729) );
  NAND2_X1 U10000 ( .A1(n9287), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10001 ( .A1(n10114), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10002 ( .A1(n7753), .A2(n7737), .ZN(n7750) );
  XNOR2_X1 U10003 ( .A(n7752), .B(n7750), .ZN(n9338) );
  NAND2_X1 U10004 ( .A1(n7792), .A2(n9338), .ZN(n7742) );
  NAND2_X1 U10005 ( .A1(n7726), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7738) );
  MUX2_X1 U10006 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7738), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n7740) );
  NAND2_X1 U10007 ( .A1(n7740), .A2(n7739), .ZN(n11135) );
  NAND2_X1 U10008 ( .A1(n6432), .A2(n11135), .ZN(n7741) );
  OAI211_X1 U10009 ( .C1(n7770), .C2(SI_3_), .A(n7742), .B(n7741), .ZN(n10707)
         );
  NAND2_X1 U10010 ( .A1(n12691), .A2(n10707), .ZN(n8252) );
  INV_X1 U10011 ( .A(n10895), .ZN(n10891) );
  NAND2_X1 U10012 ( .A1(n10892), .A2(n10891), .ZN(n7743) );
  NAND2_X1 U10013 ( .A1(n6428), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7749) );
  INV_X1 U10014 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15297) );
  OR2_X1 U10015 ( .A1(n8060), .A2(n15297), .ZN(n7748) );
  INV_X1 U10016 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15315) );
  OR2_X1 U10017 ( .A1(n8199), .A2(n15315), .ZN(n7747) );
  AND2_X1 U10018 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7745) );
  NOR2_X1 U10019 ( .A1(n7764), .A2(n7745), .ZN(n10866) );
  OR2_X1 U10020 ( .A1(n7744), .A2(n10866), .ZN(n7746) );
  NAND4_X1 U10021 ( .A1(n7749), .A2(n7748), .A3(n7747), .A4(n7746), .ZN(n12690) );
  INV_X1 U10022 ( .A(n7750), .ZN(n7751) );
  NAND2_X1 U10023 ( .A1(n7754), .A2(n7753), .ZN(n7773) );
  NAND2_X1 U10024 ( .A1(n9297), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10025 ( .A1(n9300), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U10026 ( .A1(n7774), .A2(n7755), .ZN(n7771) );
  XNOR2_X1 U10027 ( .A(n7773), .B(n7771), .ZN(n9316) );
  NAND2_X1 U10028 ( .A1(n7792), .A2(n9316), .ZN(n7762) );
  INV_X1 U10029 ( .A(n7757), .ZN(n7760) );
  NAND2_X1 U10030 ( .A1(n7739), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7758) );
  MUX2_X1 U10031 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7758), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7759) );
  NAND2_X1 U10032 ( .A1(n6433), .A2(n11258), .ZN(n7761) );
  OAI211_X1 U10033 ( .C1(n7770), .C2(SI_4_), .A(n7762), .B(n7761), .ZN(n10918)
         );
  OR2_X1 U10034 ( .A1(n12690), .A2(n10918), .ZN(n8259) );
  NAND2_X1 U10035 ( .A1(n6428), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7769) );
  INV_X1 U10036 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11102) );
  OR2_X1 U10037 ( .A1(n8199), .A2(n11102), .ZN(n7768) );
  INV_X1 U10038 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11101) );
  OR2_X1 U10039 ( .A1(n8060), .A2(n11101), .ZN(n7767) );
  NAND2_X1 U10040 ( .A1(n7764), .A2(n7763), .ZN(n7786) );
  OR2_X1 U10041 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  AND2_X1 U10042 ( .A1(n7786), .A2(n7765), .ZN(n11025) );
  OR2_X1 U10043 ( .A1(n7744), .A2(n11025), .ZN(n7766) );
  NAND4_X1 U10044 ( .A1(n7769), .A2(n7768), .A3(n7767), .A4(n7766), .ZN(n15213) );
  INV_X1 U10045 ( .A(SI_5_), .ZN(n9315) );
  NAND2_X1 U10046 ( .A1(n8166), .A2(n9315), .ZN(n7784) );
  INV_X1 U10047 ( .A(n7771), .ZN(n7772) );
  NAND2_X1 U10048 ( .A1(n7773), .A2(n7772), .ZN(n7775) );
  NAND2_X1 U10049 ( .A1(n9311), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10050 ( .A1(n9308), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7776) );
  INV_X1 U10051 ( .A(n7793), .ZN(n7777) );
  XNOR2_X1 U10052 ( .A(n7794), .B(n7777), .ZN(n9314) );
  NAND2_X1 U10053 ( .A1(n7792), .A2(n9314), .ZN(n7783) );
  NOR2_X1 U10054 ( .A1(n7757), .A2(n13298), .ZN(n7778) );
  MUX2_X1 U10055 ( .A(n13298), .B(n7778), .S(P3_IR_REG_5__SCAN_IN), .Z(n7781)
         );
  NAND2_X1 U10056 ( .A1(n7757), .A2(n7779), .ZN(n7813) );
  INV_X1 U10057 ( .A(n7813), .ZN(n7780) );
  NAND2_X1 U10058 ( .A1(n6432), .A2(n11222), .ZN(n7782) );
  NAND2_X1 U10059 ( .A1(n15213), .A2(n11024), .ZN(n8258) );
  NAND2_X1 U10060 ( .A1(n8266), .A2(n8258), .ZN(n11039) );
  INV_X1 U10061 ( .A(n11039), .ZN(n11018) );
  NAND2_X1 U10062 ( .A1(n7785), .A2(n8266), .ZN(n15211) );
  NAND2_X1 U10063 ( .A1(n6428), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7791) );
  INV_X1 U10064 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15300) );
  OR2_X1 U10065 ( .A1(n8060), .A2(n15300), .ZN(n7790) );
  INV_X1 U10066 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15230) );
  OR2_X1 U10067 ( .A1(n8199), .A2(n15230), .ZN(n7789) );
  NAND2_X1 U10068 ( .A1(n7786), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7787) );
  AND2_X1 U10069 ( .A1(n7803), .A2(n7787), .ZN(n15226) );
  OR2_X1 U10070 ( .A1(n7744), .A2(n15226), .ZN(n7788) );
  NAND4_X1 U10071 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7788), .ZN(n12689) );
  NAND2_X1 U10072 ( .A1(n8166), .A2(SI_6_), .ZN(n7801) );
  NAND2_X1 U10073 ( .A1(n7794), .A2(n7793), .ZN(n7796) );
  XNOR2_X1 U10074 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7797) );
  XNOR2_X1 U10075 ( .A(n7806), .B(n7797), .ZN(n9335) );
  NAND2_X1 U10076 ( .A1(n7792), .A2(n9335), .ZN(n7800) );
  NAND2_X1 U10077 ( .A1(n7813), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7798) );
  XNOR2_X1 U10078 ( .A(n7798), .B(P3_IR_REG_6__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U10079 ( .A1(n6433), .A2(n12705), .ZN(n7799) );
  AND3_X2 U10080 ( .A1(n7801), .A2(n7800), .A3(n7799), .ZN(n15225) );
  OR2_X2 U10081 ( .A1(n12689), .A2(n15225), .ZN(n8268) );
  NAND2_X1 U10082 ( .A1(n12689), .A2(n15225), .ZN(n8267) );
  NAND2_X1 U10083 ( .A1(n8268), .A2(n8267), .ZN(n11041) );
  INV_X1 U10084 ( .A(n11041), .ZN(n8220) );
  NAND2_X1 U10085 ( .A1(n15211), .A2(n8220), .ZN(n7802) );
  NAND2_X1 U10086 ( .A1(n7802), .A2(n8268), .ZN(n11304) );
  NAND2_X1 U10087 ( .A1(n6428), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n11230) );
  INV_X1 U10088 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11110) );
  OR2_X1 U10089 ( .A1(n8060), .A2(n11110), .ZN(n11229) );
  INV_X1 U10090 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11111) );
  OR2_X1 U10091 ( .A1(n8199), .A2(n11111), .ZN(n11228) );
  AND2_X1 U10092 ( .A1(n7803), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7804) );
  NOR2_X1 U10093 ( .A1(n7818), .A2(n7804), .ZN(n11529) );
  OR2_X1 U10094 ( .A1(n7744), .A2(n11529), .ZN(n11227) );
  NAND4_X1 U10095 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(
        n15214) );
  NAND2_X1 U10096 ( .A1(n9329), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10097 ( .A1(n7806), .A2(n7805), .ZN(n7808) );
  NAND2_X1 U10098 ( .A1(n9324), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10099 ( .A1(n9346), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10100 ( .A1(n9349), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10101 ( .A1(n7825), .A2(n7809), .ZN(n7810) );
  NAND2_X1 U10102 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  NAND2_X1 U10103 ( .A1(n7826), .A2(n7812), .ZN(n9318) );
  NAND2_X1 U10104 ( .A1(n7792), .A2(n9318), .ZN(n7817) );
  NAND2_X1 U10105 ( .A1(n7831), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7815) );
  INV_X1 U10106 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7814) );
  XNOR2_X1 U10107 ( .A(n7815), .B(n7814), .ZN(n11152) );
  NAND2_X1 U10108 ( .A1(n6432), .A2(n11152), .ZN(n7816) );
  OAI211_X1 U10109 ( .C1(n7770), .C2(SI_7_), .A(n7817), .B(n7816), .ZN(n11522)
         );
  OR2_X1 U10110 ( .A1(n15214), .A2(n11522), .ZN(n8273) );
  NAND2_X1 U10111 ( .A1(n15214), .A2(n11522), .ZN(n8272) );
  NAND2_X1 U10112 ( .A1(n8100), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7824) );
  INV_X1 U10113 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15303) );
  OR2_X1 U10114 ( .A1(n8060), .A2(n15303), .ZN(n7823) );
  NOR2_X1 U10115 ( .A1(n7818), .A2(n11736), .ZN(n7819) );
  OR2_X1 U10116 ( .A1(n7839), .A2(n7819), .ZN(n11052) );
  INV_X1 U10117 ( .A(n11052), .ZN(n11743) );
  OR2_X1 U10118 ( .A1(n7744), .A2(n11743), .ZN(n7822) );
  INV_X1 U10119 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n7820) );
  OR2_X1 U10120 ( .A1(n8184), .A2(n7820), .ZN(n7821) );
  NAND4_X1 U10121 ( .A1(n7824), .A2(n7823), .A3(n7822), .A4(n7821), .ZN(n12688) );
  NAND2_X1 U10122 ( .A1(n9351), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10123 ( .A1(n9354), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7827) );
  OR2_X1 U10124 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U10125 ( .A1(n7846), .A2(n7830), .ZN(n9334) );
  INV_X4 U10126 ( .A(n7770), .ZN(n8166) );
  NAND2_X1 U10127 ( .A1(n8166), .A2(SI_8_), .ZN(n7837) );
  NOR2_X1 U10128 ( .A1(n7831), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7834) );
  OR2_X1 U10129 ( .A1(n7834), .A2(n13298), .ZN(n7832) );
  MUX2_X1 U10130 ( .A(n7832), .B(P3_IR_REG_31__SCAN_IN), .S(n7833), .Z(n7835)
         );
  NAND2_X1 U10131 ( .A1(n7834), .A2(n7833), .ZN(n7851) );
  NAND2_X1 U10132 ( .A1(n7835), .A2(n7851), .ZN(n12720) );
  INV_X1 U10133 ( .A(n12720), .ZN(n11156) );
  NAND2_X1 U10134 ( .A1(n6433), .A2(n11156), .ZN(n7836) );
  OAI211_X1 U10135 ( .C1(n7733), .C2(n9334), .A(n7837), .B(n7836), .ZN(n11596)
         );
  XNOR2_X1 U10136 ( .A(n12688), .B(n11596), .ZN(n11047) );
  INV_X1 U10137 ( .A(n11596), .ZN(n11735) );
  OR2_X1 U10138 ( .A1(n12688), .A2(n11735), .ZN(n8277) );
  NAND2_X1 U10139 ( .A1(n6428), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7844) );
  INV_X1 U10140 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11162) );
  OR2_X1 U10141 ( .A1(n8199), .A2(n11162), .ZN(n7843) );
  INV_X1 U10142 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11161) );
  OR2_X1 U10143 ( .A1(n8060), .A2(n11161), .ZN(n7842) );
  OR2_X1 U10144 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  AND2_X1 U10145 ( .A1(n7859), .A2(n7840), .ZN(n11606) );
  OR2_X1 U10146 ( .A1(n7744), .A2(n11606), .ZN(n7841) );
  NAND4_X1 U10147 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n15196) );
  INV_X1 U10148 ( .A(SI_9_), .ZN(n9296) );
  NAND2_X1 U10149 ( .A1(n8166), .A2(n9296), .ZN(n7858) );
  NAND2_X1 U10150 ( .A1(n9389), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10151 ( .A1(n9382), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7847) );
  OR2_X1 U10152 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  NAND2_X1 U10153 ( .A1(n7866), .A2(n7850), .ZN(n9295) );
  NAND2_X1 U10154 ( .A1(n8191), .A2(n9295), .ZN(n7857) );
  NAND2_X1 U10155 ( .A1(n7851), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7852) );
  MUX2_X1 U10156 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7852), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7855) );
  INV_X1 U10157 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U10158 ( .A1(n7855), .A2(n7854), .ZN(n11172) );
  NAND2_X1 U10159 ( .A1(n6433), .A2(n11172), .ZN(n7856) );
  NOR2_X1 U10160 ( .A1(n15196), .A2(n15282), .ZN(n8282) );
  NAND2_X1 U10161 ( .A1(n15196), .A2(n15282), .ZN(n8280) );
  NAND2_X1 U10162 ( .A1(n6428), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7864) );
  INV_X1 U10163 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11186) );
  OR2_X1 U10164 ( .A1(n8060), .A2(n11186), .ZN(n7863) );
  INV_X1 U10165 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15204) );
  OR2_X1 U10166 ( .A1(n8199), .A2(n15204), .ZN(n7862) );
  NAND2_X1 U10167 ( .A1(n7859), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7860) );
  AND2_X1 U10168 ( .A1(n7877), .A2(n7860), .ZN(n15210) );
  OR2_X1 U10169 ( .A1(n7744), .A2(n15210), .ZN(n7861) );
  NAND4_X1 U10170 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n12635) );
  NAND2_X1 U10171 ( .A1(n9465), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10172 ( .A1(n9468), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7867) );
  OR2_X1 U10173 ( .A1(n7869), .A2(n7868), .ZN(n7870) );
  NAND2_X1 U10174 ( .A1(n7886), .A2(n7870), .ZN(n9293) );
  NAND2_X1 U10175 ( .A1(n8191), .A2(n9293), .ZN(n7876) );
  NOR2_X1 U10176 ( .A1(n7853), .A2(n13298), .ZN(n7871) );
  MUX2_X1 U10177 ( .A(n13298), .B(n7871), .S(P3_IR_REG_10__SCAN_IN), .Z(n7874)
         );
  INV_X1 U10178 ( .A(n7872), .ZN(n7873) );
  NAND2_X1 U10179 ( .A1(n6432), .A2(n11393), .ZN(n7875) );
  OAI211_X1 U10180 ( .C1(n7770), .C2(SI_10_), .A(n7876), .B(n7875), .ZN(n15205) );
  NAND2_X1 U10181 ( .A1(n12635), .A2(n15205), .ZN(n8219) );
  INV_X1 U10182 ( .A(n8219), .ZN(n8288) );
  OR2_X1 U10183 ( .A1(n12635), .A2(n15205), .ZN(n8284) );
  NAND2_X1 U10184 ( .A1(n6428), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7884) );
  AND2_X1 U10185 ( .A1(n7877), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7878) );
  NOR2_X1 U10186 ( .A1(n7895), .A2(n7878), .ZN(n14862) );
  OR2_X1 U10187 ( .A1(n7744), .A2(n14862), .ZN(n7883) );
  INV_X1 U10188 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7879) );
  OR2_X1 U10189 ( .A1(n8060), .A2(n7879), .ZN(n7882) );
  INV_X1 U10190 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7880) );
  OR2_X1 U10191 ( .A1(n8199), .A2(n7880), .ZN(n7881) );
  NAND4_X1 U10192 ( .A1(n7884), .A2(n7883), .A3(n7882), .A4(n7881), .ZN(n15197) );
  NAND2_X1 U10193 ( .A1(n9572), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10194 ( .A1(n9566), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7887) );
  OR2_X1 U10195 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  NAND2_X1 U10196 ( .A1(n7903), .A2(n7890), .ZN(n9303) );
  NAND2_X1 U10197 ( .A1(n8191), .A2(n9303), .ZN(n7894) );
  NAND2_X1 U10198 ( .A1(n8166), .A2(n9304), .ZN(n7893) );
  NAND2_X1 U10199 ( .A1(n7872), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7891) );
  INV_X1 U10200 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n15451) );
  XNOR2_X1 U10201 ( .A(n7891), .B(n15451), .ZN(n11394) );
  NAND2_X1 U10202 ( .A1(n6432), .A2(n11394), .ZN(n7892) );
  NAND2_X1 U10203 ( .A1(n15197), .A2(n12636), .ZN(n8290) );
  NAND2_X1 U10204 ( .A1(n6428), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10205 ( .A1(n7895), .A2(n11714), .ZN(n7930) );
  INV_X1 U10206 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U10207 ( .A1(n7896), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10208 ( .A1(n7930), .A2(n7897), .ZN(n14841) );
  INV_X1 U10209 ( .A(n14841), .ZN(n12568) );
  OR2_X1 U10210 ( .A1(n7744), .A2(n12568), .ZN(n7900) );
  INV_X1 U10211 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14871) );
  OR2_X1 U10212 ( .A1(n8060), .A2(n14871), .ZN(n7899) );
  INV_X1 U10213 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n15329) );
  OR2_X1 U10214 ( .A1(n8199), .A2(n15329), .ZN(n7898) );
  NAND4_X1 U10215 ( .A1(n7901), .A2(n7900), .A3(n7899), .A4(n7898), .ZN(n12687) );
  NAND2_X1 U10216 ( .A1(n9763), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10217 ( .A1(n9764), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7904) );
  OR2_X1 U10218 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  AND2_X1 U10219 ( .A1(n7922), .A2(n7907), .ZN(n9320) );
  NAND2_X1 U10220 ( .A1(n8191), .A2(n9320), .ZN(n7913) );
  NAND2_X1 U10221 ( .A1(n8166), .A2(SI_12_), .ZN(n7912) );
  NAND2_X1 U10222 ( .A1(n7513), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7908) );
  MUX2_X1 U10223 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7908), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7910) );
  NAND2_X1 U10224 ( .A1(n7910), .A2(n7909), .ZN(n12739) );
  INV_X1 U10225 ( .A(n12739), .ZN(n11725) );
  NAND2_X1 U10226 ( .A1(n6432), .A2(n11725), .ZN(n7911) );
  INV_X1 U10227 ( .A(n8296), .ZN(n7914) );
  NAND2_X1 U10228 ( .A1(n12687), .A2(n14846), .ZN(n8289) );
  NAND2_X1 U10229 ( .A1(n8296), .A2(n8289), .ZN(n12426) );
  AND2_X1 U10230 ( .A1(n14850), .A2(n7916), .ZN(n7915) );
  INV_X1 U10231 ( .A(n7916), .ZN(n7918) );
  AND2_X1 U10232 ( .A1(n14842), .A2(n8296), .ZN(n7917) );
  NAND2_X1 U10233 ( .A1(n7920), .A2(n7919), .ZN(n13115) );
  XNOR2_X1 U10234 ( .A(n7936), .B(n6931), .ZN(n9374) );
  NAND2_X1 U10235 ( .A1(n9374), .A2(n8191), .ZN(n7927) );
  NAND2_X1 U10236 ( .A1(n7909), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7925) );
  AOI22_X1 U10237 ( .A1(n8166), .A2(n9375), .B1(n6433), .B2(n12771), .ZN(n7926) );
  NAND2_X1 U10238 ( .A1(n6428), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7935) );
  INV_X1 U10239 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15428) );
  OR2_X1 U10240 ( .A1(n8199), .A2(n15428), .ZN(n7934) );
  INV_X1 U10241 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13208) );
  OR2_X1 U10242 ( .A1(n8060), .A2(n13208), .ZN(n7933) );
  INV_X1 U10243 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U10244 ( .A1(n7930), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7931) );
  AND2_X1 U10245 ( .A1(n7941), .A2(n7931), .ZN(n13120) );
  OR2_X1 U10246 ( .A1(n7744), .A2(n13120), .ZN(n7932) );
  NAND4_X1 U10247 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n14838) );
  NOR2_X1 U10248 ( .A1(n13293), .A2(n14838), .ZN(n8302) );
  NAND2_X1 U10249 ( .A1(n13293), .A2(n14838), .ZN(n8215) );
  NAND2_X1 U10250 ( .A1(n10063), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7949) );
  INV_X1 U10251 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10065) );
  NAND2_X1 U10252 ( .A1(n10065), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7937) );
  XNOR2_X1 U10253 ( .A(n7948), .B(n7947), .ZN(n9392) );
  NAND2_X1 U10254 ( .A1(n9392), .A2(n8191), .ZN(n7940) );
  NOR2_X1 U10255 ( .A1(n7909), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7952) );
  OR2_X1 U10256 ( .A1(n7952), .A2(n13298), .ZN(n7938) );
  INV_X1 U10257 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7951) );
  XNOR2_X1 U10258 ( .A(n7938), .B(n7951), .ZN(n12796) );
  AOI22_X1 U10259 ( .A1(n8166), .A2(n9391), .B1(n6433), .B2(n12796), .ZN(n7939) );
  NAND2_X1 U10260 ( .A1(n6428), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7946) );
  INV_X1 U10261 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13104) );
  OR2_X1 U10262 ( .A1(n8199), .A2(n13104), .ZN(n7945) );
  INV_X1 U10263 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13204) );
  OR2_X1 U10264 ( .A1(n8060), .A2(n13204), .ZN(n7944) );
  NAND2_X1 U10265 ( .A1(n7941), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7942) );
  AND2_X1 U10266 ( .A1(n7960), .A2(n7942), .ZN(n13103) );
  OR2_X1 U10267 ( .A1(n7744), .A2(n13103), .ZN(n7943) );
  XNOR2_X1 U10268 ( .A(n13289), .B(n13119), .ZN(n13097) );
  INV_X1 U10269 ( .A(n13097), .ZN(n13108) );
  OR2_X1 U10270 ( .A1(n13289), .A2(n12686), .ZN(n8305) );
  NAND2_X1 U10271 ( .A1(n10220), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10272 ( .A1(n10213), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10273 ( .A1(n7969), .A2(n7950), .ZN(n7966) );
  XNOR2_X1 U10274 ( .A(n7968), .B(n7966), .ZN(n9603) );
  NAND2_X1 U10275 ( .A1(n9603), .A2(n8191), .ZN(n7957) );
  NAND2_X1 U10276 ( .A1(n7952), .A2(n7951), .ZN(n7954) );
  NAND2_X1 U10277 ( .A1(n7954), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7953) );
  MUX2_X1 U10278 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7953), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n7955) );
  AOI22_X1 U10279 ( .A1(n8166), .A2(SI_15_), .B1(n6432), .B2(n12809), .ZN(
        n7956) );
  NAND2_X1 U10280 ( .A1(n7957), .A2(n7956), .ZN(n13089) );
  NAND2_X1 U10281 ( .A1(n6428), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7965) );
  INV_X1 U10282 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13091) );
  OR2_X1 U10283 ( .A1(n8199), .A2(n13091), .ZN(n7964) );
  INV_X1 U10284 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13199) );
  OR2_X1 U10285 ( .A1(n8060), .A2(n13199), .ZN(n7963) );
  INV_X1 U10286 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10287 ( .A1(n7960), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7961) );
  AND2_X1 U10288 ( .A1(n7975), .A2(n7961), .ZN(n13090) );
  OR2_X1 U10289 ( .A1(n7744), .A2(n13090), .ZN(n7962) );
  NAND4_X1 U10290 ( .A1(n7965), .A2(n7964), .A3(n7963), .A4(n7962), .ZN(n13100) );
  OR2_X1 U10291 ( .A1(n13089), .A2(n13074), .ZN(n8309) );
  NAND2_X1 U10292 ( .A1(n13089), .A2(n13074), .ZN(n8314) );
  NAND2_X1 U10293 ( .A1(n13086), .A2(n8314), .ZN(n13070) );
  INV_X1 U10294 ( .A(n7966), .ZN(n7967) );
  NAND2_X1 U10295 ( .A1(n15443), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10296 ( .A1(n10296), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10297 ( .A1(n7984), .A2(n7971), .ZN(n7982) );
  NAND2_X1 U10298 ( .A1(n9654), .A2(n8191), .ZN(n7974) );
  NAND2_X1 U10299 ( .A1(n7986), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7972) );
  XNOR2_X1 U10300 ( .A(n7972), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U10301 ( .A1(n8166), .A2(SI_16_), .B1(n6433), .B2(n12830), .ZN(
        n7973) );
  NAND2_X1 U10302 ( .A1(n7974), .A2(n7973), .ZN(n13076) );
  NAND2_X1 U10303 ( .A1(n6428), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7980) );
  INV_X1 U10304 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13078) );
  OR2_X1 U10305 ( .A1(n8199), .A2(n13078), .ZN(n7979) );
  INV_X1 U10306 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13195) );
  OR2_X1 U10307 ( .A1(n8060), .A2(n13195), .ZN(n7978) );
  OR2_X2 U10308 ( .A1(n7975), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10309 ( .A1(n7975), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7976) );
  AND2_X1 U10310 ( .A1(n7994), .A2(n7976), .ZN(n13077) );
  OR2_X1 U10311 ( .A1(n7744), .A2(n13077), .ZN(n7977) );
  OR2_X1 U10312 ( .A1(n13076), .A2(n13085), .ZN(n8316) );
  NAND2_X1 U10313 ( .A1(n13076), .A2(n13085), .ZN(n8315) );
  NAND2_X1 U10314 ( .A1(n8316), .A2(n8315), .ZN(n13072) );
  INV_X1 U10315 ( .A(n13072), .ZN(n13069) );
  NAND2_X1 U10316 ( .A1(n13070), .A2(n13069), .ZN(n7981) );
  NAND2_X1 U10317 ( .A1(n7981), .A2(n8315), .ZN(n13062) );
  INV_X1 U10318 ( .A(n7982), .ZN(n7983) );
  NAND2_X1 U10319 ( .A1(n10532), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10320 ( .A1(n10534), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10321 ( .A1(n8003), .A2(n7985), .ZN(n8000) );
  XNOR2_X1 U10322 ( .A(n8002), .B(n8000), .ZN(n9834) );
  NAND2_X1 U10323 ( .A1(n9834), .A2(n8191), .ZN(n7991) );
  INV_X1 U10324 ( .A(n7986), .ZN(n7988) );
  INV_X1 U10325 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U10326 ( .A1(n7988), .A2(n7987), .ZN(n8008) );
  NAND2_X1 U10327 ( .A1(n8008), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7989) );
  XNOR2_X1 U10328 ( .A(n7989), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U10329 ( .A1(n8166), .A2(SI_17_), .B1(n6432), .B2(n12842), .ZN(
        n7990) );
  NAND2_X1 U10330 ( .A1(n7991), .A2(n7990), .ZN(n12584) );
  NAND2_X1 U10331 ( .A1(n8100), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7999) );
  INV_X1 U10332 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13191) );
  OR2_X1 U10333 ( .A1(n8060), .A2(n13191), .ZN(n7998) );
  INV_X1 U10334 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10335 ( .A1(n7994), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7995) );
  AND2_X1 U10336 ( .A1(n8012), .A2(n7995), .ZN(n13063) );
  OR2_X1 U10337 ( .A1(n7744), .A2(n13063), .ZN(n7997) );
  INV_X1 U10338 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13275) );
  OR2_X1 U10339 ( .A1(n8184), .A2(n13275), .ZN(n7996) );
  OR2_X1 U10340 ( .A1(n12584), .A2(n13075), .ZN(n8319) );
  NAND2_X1 U10341 ( .A1(n12584), .A2(n13075), .ZN(n13041) );
  INV_X1 U10342 ( .A(n13057), .ZN(n13061) );
  NAND2_X1 U10343 ( .A1(n13062), .A2(n13061), .ZN(n13060) );
  INV_X1 U10344 ( .A(n8000), .ZN(n8001) );
  NAND2_X1 U10345 ( .A1(n10814), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10346 ( .A1(n10811), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8004) );
  OR2_X1 U10347 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  NAND2_X1 U10348 ( .A1(n8020), .A2(n8007), .ZN(n9904) );
  OR2_X1 U10349 ( .A1(n9904), .A2(n7733), .ZN(n8011) );
  OAI21_X1 U10350 ( .B1(n8008), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8009) );
  XNOR2_X1 U10351 ( .A(n8009), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U10352 ( .A1(n8166), .A2(SI_18_), .B1(n6433), .B2(n12876), .ZN(
        n8010) );
  NAND2_X1 U10353 ( .A1(n8011), .A2(n8010), .ZN(n12643) );
  NAND2_X1 U10354 ( .A1(n8195), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8017) );
  INV_X1 U10355 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13271) );
  OR2_X1 U10356 ( .A1(n8184), .A2(n13271), .ZN(n8016) );
  OR2_X2 U10357 ( .A1(n8012), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10358 ( .A1(n8012), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8013) );
  AND2_X1 U10359 ( .A1(n8035), .A2(n8013), .ZN(n13050) );
  OR2_X1 U10360 ( .A1(n7744), .A2(n13050), .ZN(n8015) );
  INV_X1 U10361 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13051) );
  OR2_X1 U10362 ( .A1(n8199), .A2(n13051), .ZN(n8014) );
  NAND2_X1 U10363 ( .A1(n12643), .A2(n13059), .ZN(n8325) );
  INV_X1 U10364 ( .A(n13047), .ZN(n8329) );
  INV_X1 U10365 ( .A(n13041), .ZN(n8323) );
  NOR2_X1 U10366 ( .A1(n8329), .A2(n8323), .ZN(n8018) );
  INV_X1 U10367 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U10368 ( .A1(n10888), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8041) );
  INV_X1 U10369 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10890) );
  NAND2_X1 U10370 ( .A1(n10890), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8021) );
  OR2_X1 U10371 ( .A1(n8023), .A2(n8022), .ZN(n8024) );
  NAND2_X1 U10372 ( .A1(n8042), .A2(n8024), .ZN(n9992) );
  NAND2_X1 U10373 ( .A1(n9992), .A2(n8191), .ZN(n8032) );
  INV_X1 U10374 ( .A(SI_19_), .ZN(n9991) );
  INV_X1 U10375 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U10376 ( .A1(n8026), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8027) );
  MUX2_X1 U10377 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8027), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8029) );
  AOI22_X1 U10378 ( .A1(n8166), .A2(n9991), .B1(n6432), .B2(n6688), .ZN(n8031)
         );
  NAND2_X1 U10379 ( .A1(n6428), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8040) );
  INV_X1 U10380 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13033) );
  OR2_X1 U10381 ( .A1(n8199), .A2(n13033), .ZN(n8039) );
  INV_X1 U10382 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13183) );
  OR2_X1 U10383 ( .A1(n8060), .A2(n13183), .ZN(n8038) );
  INV_X1 U10384 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10385 ( .A1(n8035), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8036) );
  AND2_X1 U10386 ( .A1(n8045), .A2(n8036), .ZN(n13032) );
  OR2_X1 U10387 ( .A1(n7744), .A2(n13032), .ZN(n8037) );
  NAND4_X1 U10388 ( .A1(n8040), .A2(n8039), .A3(n8038), .A4(n8037), .ZN(n12682) );
  NAND2_X1 U10389 ( .A1(n13269), .A2(n12682), .ZN(n8332) );
  XNOR2_X1 U10390 ( .A(n8051), .B(n6945), .ZN(n10184) );
  NAND2_X1 U10391 ( .A1(n10184), .A2(n8191), .ZN(n8044) );
  NAND2_X1 U10392 ( .A1(n8166), .A2(SI_20_), .ZN(n8043) );
  NAND2_X1 U10393 ( .A1(n8100), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8050) );
  INV_X1 U10394 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13178) );
  OR2_X1 U10395 ( .A1(n8060), .A2(n13178), .ZN(n8049) );
  OR2_X2 U10396 ( .A1(n8045), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10397 ( .A1(n8045), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8046) );
  AND2_X1 U10398 ( .A1(n8058), .A2(n8046), .ZN(n12609) );
  OR2_X1 U10399 ( .A1(n7744), .A2(n12609), .ZN(n8048) );
  INV_X1 U10400 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13263) );
  OR2_X1 U10401 ( .A1(n8184), .A2(n13263), .ZN(n8047) );
  NAND2_X1 U10402 ( .A1(n12605), .A2(n13028), .ZN(n8337) );
  XNOR2_X1 U10403 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n8065) );
  XNOR2_X1 U10404 ( .A(n8066), .B(n8065), .ZN(n10345) );
  NAND2_X1 U10405 ( .A1(n10345), .A2(n8191), .ZN(n8055) );
  NAND2_X1 U10406 ( .A1(n8166), .A2(SI_21_), .ZN(n8054) );
  INV_X1 U10407 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U10408 ( .A1(n8058), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10409 ( .A1(n8070), .A2(n8059), .ZN(n13007) );
  NAND2_X1 U10410 ( .A1(n8170), .A2(n13007), .ZN(n8064) );
  INV_X1 U10411 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13009) );
  OR2_X1 U10412 ( .A1(n8199), .A2(n13009), .ZN(n8063) );
  INV_X1 U10413 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13174) );
  OR2_X1 U10414 ( .A1(n8060), .A2(n13174), .ZN(n8062) );
  INV_X1 U10415 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13259) );
  OR2_X1 U10416 ( .A1(n8184), .A2(n13259), .ZN(n8061) );
  NAND2_X1 U10417 ( .A1(n13170), .A2(n13020), .ZN(n8341) );
  INV_X1 U10418 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U10419 ( .A1(n11036), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8067) );
  XNOR2_X1 U10420 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n8077) );
  XNOR2_X1 U10421 ( .A(n8078), .B(n8077), .ZN(n10446) );
  NAND2_X1 U10422 ( .A1(n10446), .A2(n8191), .ZN(n8069) );
  NAND2_X1 U10423 ( .A1(n8166), .A2(SI_22_), .ZN(n8068) );
  NAND2_X1 U10424 ( .A1(n8070), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10425 ( .A1(n8081), .A2(n8071), .ZN(n12992) );
  NAND2_X1 U10426 ( .A1(n12992), .A2(n8170), .ZN(n8075) );
  NAND2_X1 U10427 ( .A1(n8100), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10428 ( .A1(n8195), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8073) );
  INV_X1 U10429 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13255) );
  OR2_X1 U10430 ( .A1(n8184), .A2(n13255), .ZN(n8072) );
  NAND2_X1 U10431 ( .A1(n12996), .A2(n13004), .ZN(n8345) );
  NAND2_X1 U10432 ( .A1(n12998), .A2(n8345), .ZN(n8076) );
  NAND2_X1 U10433 ( .A1(n8076), .A2(n8344), .ZN(n12973) );
  INV_X1 U10434 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15351) );
  XNOR2_X1 U10435 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8088) );
  XNOR2_X1 U10436 ( .A(n8089), .B(n8088), .ZN(n10607) );
  NAND2_X1 U10437 ( .A1(n10607), .A2(n8191), .ZN(n8080) );
  NAND2_X1 U10438 ( .A1(n8166), .A2(SI_23_), .ZN(n8079) );
  INV_X1 U10439 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U10440 ( .A1(n8081), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10441 ( .A1(n8098), .A2(n8082), .ZN(n12981) );
  NAND2_X1 U10442 ( .A1(n12981), .A2(n8170), .ZN(n8086) );
  NAND2_X1 U10443 ( .A1(n8100), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U10444 ( .A1(n8195), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8083) );
  AND2_X1 U10445 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U10446 ( .A1(n12973), .A2(n12977), .ZN(n8087) );
  INV_X1 U10447 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U10448 ( .A1(n11666), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8090) );
  INV_X1 U10449 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U10450 ( .A1(n8092), .A2(n11745), .ZN(n8093) );
  INV_X1 U10451 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11748) );
  XNOR2_X1 U10452 ( .A(n8105), .B(n11748), .ZN(n10905) );
  NAND2_X1 U10453 ( .A1(n10905), .A2(n8191), .ZN(n8095) );
  NAND2_X1 U10454 ( .A1(n8166), .A2(SI_24_), .ZN(n8094) );
  INV_X1 U10455 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10456 ( .A1(n8098), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10457 ( .A1(n8112), .A2(n8099), .ZN(n12968) );
  NAND2_X1 U10458 ( .A1(n12968), .A2(n8170), .ZN(n8103) );
  AOI22_X1 U10459 ( .A1(n8100), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n8195), .B2(
        P3_REG1_REG_24__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10460 ( .A1(n6428), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10461 ( .A1(n12967), .A2(n12978), .ZN(n8356) );
  XNOR2_X1 U10462 ( .A(n12053), .B(P1_DATAO_REG_25__SCAN_IN), .ZN(n8107) );
  XNOR2_X1 U10463 ( .A(n8121), .B(n8107), .ZN(n11031) );
  NAND2_X1 U10464 ( .A1(n11031), .A2(n8191), .ZN(n8109) );
  NAND2_X1 U10465 ( .A1(n8166), .A2(SI_25_), .ZN(n8108) );
  INV_X1 U10466 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U10467 ( .A1(n8112), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10468 ( .A1(n8126), .A2(n8113), .ZN(n12955) );
  NAND2_X1 U10469 ( .A1(n12955), .A2(n8170), .ZN(n8119) );
  INV_X1 U10470 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U10471 ( .A1(n6428), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10472 ( .A1(n8195), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8114) );
  OAI211_X1 U10473 ( .C1(n8199), .C2(n8116), .A(n8115), .B(n8114), .ZN(n8117)
         );
  INV_X1 U10474 ( .A(n8117), .ZN(n8118) );
  NAND2_X1 U10475 ( .A1(n12954), .A2(n12964), .ZN(n8359) );
  NAND2_X1 U10476 ( .A1(n12951), .A2(n8359), .ZN(n12931) );
  NAND2_X1 U10477 ( .A1(n15327), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10478 ( .A1(n12053), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8122) );
  INV_X1 U10479 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14000) );
  XNOR2_X1 U10480 ( .A(n14000), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8123) );
  XNOR2_X1 U10481 ( .A(n8134), .B(n8123), .ZN(n11300) );
  NAND2_X1 U10482 ( .A1(n11300), .A2(n8191), .ZN(n8125) );
  NAND2_X1 U10483 ( .A1(n8166), .A2(SI_26_), .ZN(n8124) );
  NAND2_X1 U10484 ( .A1(n8126), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10485 ( .A1(n8142), .A2(n8127), .ZN(n12938) );
  NAND2_X1 U10486 ( .A1(n12938), .A2(n8170), .ZN(n8132) );
  INV_X1 U10487 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U10488 ( .A1(n8195), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U10489 ( .A1(n6428), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8128) );
  OAI211_X1 U10490 ( .C1(n12940), .C2(n8199), .A(n8129), .B(n8128), .ZN(n8130)
         );
  INV_X1 U10491 ( .A(n8130), .ZN(n8131) );
  NAND2_X1 U10492 ( .A1(n12942), .A2(n12948), .ZN(n8365) );
  INV_X1 U10493 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14708) );
  AND2_X1 U10494 ( .A1(n14708), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10495 ( .A1(n14000), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8135) );
  XNOR2_X1 U10496 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8137) );
  XNOR2_X1 U10497 ( .A(n8151), .B(n8137), .ZN(n11610) );
  NAND2_X1 U10498 ( .A1(n11610), .A2(n8191), .ZN(n8139) );
  NAND2_X1 U10499 ( .A1(n8166), .A2(SI_27_), .ZN(n8138) );
  INV_X1 U10500 ( .A(n8142), .ZN(n8141) );
  INV_X1 U10501 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10502 ( .A1(n8141), .A2(n8140), .ZN(n8156) );
  NAND2_X1 U10503 ( .A1(n8142), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10504 ( .A1(n8156), .A2(n8143), .ZN(n12926) );
  NAND2_X1 U10505 ( .A1(n12926), .A2(n8170), .ZN(n8149) );
  INV_X1 U10506 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U10507 ( .A1(n6428), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10508 ( .A1(n8195), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8144) );
  OAI211_X1 U10509 ( .C1(n8199), .C2(n8146), .A(n8145), .B(n8144), .ZN(n8147)
         );
  INV_X1 U10510 ( .A(n8147), .ZN(n8148) );
  NOR2_X1 U10511 ( .A1(n13238), .A2(n12677), .ZN(n8370) );
  INV_X1 U10512 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13997) );
  AND2_X1 U10513 ( .A1(n13997), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8150) );
  INV_X1 U10514 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14702) );
  NAND2_X1 U10515 ( .A1(n14702), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8152) );
  INV_X1 U10516 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9151) );
  XNOR2_X1 U10517 ( .A(n9151), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8153) );
  XNOR2_X1 U10518 ( .A(n8163), .B(n8153), .ZN(n11888) );
  NAND2_X1 U10519 ( .A1(n11888), .A2(n8191), .ZN(n8155) );
  NAND2_X1 U10520 ( .A1(n7721), .A2(SI_28_), .ZN(n8154) );
  NAND2_X1 U10521 ( .A1(n8156), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10522 ( .A1(n8169), .A2(n8157), .ZN(n12911) );
  INV_X1 U10523 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U10524 ( .A1(n6428), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10525 ( .A1(n8195), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8158) );
  OAI211_X1 U10526 ( .C1(n8199), .C2(n8160), .A(n8159), .B(n8158), .ZN(n8161)
         );
  NAND2_X1 U10527 ( .A1(n13139), .A2(n12919), .ZN(n8371) );
  INV_X1 U10528 ( .A(n8214), .ZN(n8377) );
  INV_X1 U10529 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14698) );
  AND2_X1 U10530 ( .A1(n14698), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10531 ( .A1(n9151), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8164) );
  XNOR2_X1 U10532 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8175) );
  XNOR2_X1 U10533 ( .A(n8177), .B(n8175), .ZN(n12416) );
  NAND2_X1 U10534 ( .A1(n12416), .A2(n8191), .ZN(n8168) );
  NAND2_X1 U10535 ( .A1(n8166), .A2(SI_29_), .ZN(n8167) );
  NAND2_X1 U10536 ( .A1(n12457), .A2(n8170), .ZN(n8202) );
  INV_X1 U10537 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U10538 ( .A1(n6428), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U10539 ( .A1(n8195), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8171) );
  OAI211_X1 U10540 ( .C1(n8199), .C2(n12458), .A(n8172), .B(n8171), .ZN(n8173)
         );
  INV_X1 U10541 ( .A(n8173), .ZN(n8174) );
  INV_X1 U10542 ( .A(n8175), .ZN(n8176) );
  INV_X1 U10543 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14695) );
  NAND2_X1 U10544 ( .A1(n14695), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8178) );
  INV_X1 U10545 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15339) );
  INV_X1 U10546 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9128) );
  XNOR2_X1 U10547 ( .A(n9128), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n8179) );
  XNOR2_X1 U10548 ( .A(n8180), .B(n8179), .ZN(n13297) );
  NAND2_X1 U10549 ( .A1(n13297), .A2(n8191), .ZN(n8182) );
  NAND2_X1 U10550 ( .A1(n7721), .A2(SI_31_), .ZN(n8181) );
  INV_X1 U10551 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10552 ( .A1(n8195), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8186) );
  INV_X1 U10553 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n8183) );
  OR2_X1 U10554 ( .A1(n8184), .A2(n8183), .ZN(n8185) );
  OAI211_X1 U10555 ( .C1(n8199), .C2(n8187), .A(n8186), .B(n8185), .ZN(n8188)
         );
  INV_X1 U10556 ( .A(n8188), .ZN(n8189) );
  XNOR2_X1 U10557 ( .A(n8190), .B(n6593), .ZN(n11884) );
  NAND2_X1 U10558 ( .A1(n11884), .A2(n8191), .ZN(n8193) );
  NAND2_X1 U10559 ( .A1(n7721), .A2(SI_30_), .ZN(n8192) );
  INV_X1 U10560 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10561 ( .A1(n6428), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10562 ( .A1(n8195), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U10563 ( .C1(n8199), .C2(n8198), .A(n8197), .B(n8196), .ZN(n8200)
         );
  INV_X1 U10564 ( .A(n8200), .ZN(n8201) );
  NAND2_X1 U10565 ( .A1(n13229), .A2(n12454), .ZN(n8203) );
  INV_X1 U10566 ( .A(n13229), .ZN(n12901) );
  INV_X1 U10567 ( .A(n12895), .ZN(n12676) );
  NAND2_X1 U10568 ( .A1(n13133), .A2(n12907), .ZN(n8376) );
  OAI21_X1 U10569 ( .B1(n12901), .B2(n12676), .A(n8376), .ZN(n8204) );
  NOR2_X1 U10570 ( .A1(n8383), .A2(n8204), .ZN(n8207) );
  INV_X1 U10571 ( .A(n8384), .ZN(n8206) );
  NOR2_X1 U10572 ( .A1(n13229), .A2(n12454), .ZN(n8379) );
  NAND2_X1 U10573 ( .A1(n8379), .A2(n13225), .ZN(n8205) );
  XNOR2_X1 U10574 ( .A(n8208), .B(n6688), .ZN(n8213) );
  NAND2_X1 U10575 ( .A1(n8234), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U10576 ( .A1(n10893), .A2(n10617), .ZN(n10596) );
  INV_X1 U10577 ( .A(n10596), .ZN(n8212) );
  NAND2_X1 U10578 ( .A1(n8381), .A2(n8376), .ZN(n12459) );
  INV_X1 U10579 ( .A(n12459), .ZN(n8230) );
  NAND2_X1 U10580 ( .A1(n8214), .A2(n8371), .ZN(n12903) );
  INV_X1 U10581 ( .A(n12903), .ZN(n12905) );
  INV_X1 U10582 ( .A(n12952), .ZN(n8228) );
  INV_X1 U10583 ( .A(n8215), .ZN(n8301) );
  OR2_X1 U10584 ( .A1(n8302), .A2(n8301), .ZN(n13116) );
  INV_X1 U10585 ( .A(n11441), .ZN(n8217) );
  NOR3_X1 U10586 ( .A1(n8217), .A2(n11039), .A3(n10769), .ZN(n8218) );
  XNOR2_X1 U10587 ( .A(n15196), .B(n12421), .ZN(n11600) );
  NAND4_X1 U10588 ( .A1(n8218), .A2(n14850), .A3(n14844), .A4(n11600), .ZN(
        n8223) );
  NAND2_X1 U10589 ( .A1(n8284), .A2(n8219), .ZN(n15194) );
  NAND2_X1 U10590 ( .A1(n13213), .A2(n10626), .ZN(n8238) );
  NAND2_X1 U10591 ( .A1(n13219), .A2(n8238), .ZN(n10600) );
  NOR4_X1 U10592 ( .A1(n10895), .A2(n15194), .A3(n11041), .A4(n10600), .ZN(
        n8221) );
  NAND4_X1 U10593 ( .A1(n8221), .A2(n10762), .A3(n10909), .A4(n11047), .ZN(
        n8222) );
  NOR4_X1 U10594 ( .A1(n7198), .A2(n13116), .A3(n8223), .A4(n8222), .ZN(n8224)
         );
  NAND4_X1 U10595 ( .A1(n13047), .A2(n13097), .A3(n13069), .A4(n8224), .ZN(
        n8225) );
  INV_X1 U10596 ( .A(n13026), .ZN(n13036) );
  NOR4_X1 U10597 ( .A1(n13057), .A2(n13017), .A3(n8225), .A4(n13036), .ZN(
        n8226) );
  NAND4_X1 U10598 ( .A1(n12986), .A2(n13011), .A3(n8226), .A4(n12977), .ZN(
        n8227) );
  NOR4_X1 U10599 ( .A1(n12933), .A2(n8228), .A3(n12961), .A4(n8227), .ZN(n8229) );
  XNOR2_X1 U10600 ( .A(n8231), .B(n6688), .ZN(n8233) );
  NAND2_X1 U10601 ( .A1(n10416), .A2(n10617), .ZN(n10414) );
  INV_X1 U10602 ( .A(n10414), .ZN(n8232) );
  NAND2_X1 U10603 ( .A1(n10417), .A2(n6688), .ZN(n10618) );
  INV_X1 U10604 ( .A(n10618), .ZN(n10764) );
  INV_X1 U10605 ( .A(n8390), .ZN(n8235) );
  NAND2_X1 U10606 ( .A1(n8235), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8236) );
  MUX2_X1 U10607 ( .A(n8216), .B(n8237), .S(n10616), .Z(n8244) );
  NAND2_X1 U10608 ( .A1(n8238), .A2(n10615), .ZN(n8241) );
  NAND2_X1 U10609 ( .A1(n8238), .A2(n10893), .ZN(n8239) );
  NAND3_X1 U10610 ( .A1(n8239), .A2(n10616), .A3(n8216), .ZN(n8240) );
  OAI21_X1 U10611 ( .B1(n10769), .B2(n8241), .A(n8240), .ZN(n8242) );
  OAI21_X1 U10612 ( .B1(n10893), .B2(n13219), .A(n8242), .ZN(n8243) );
  NAND3_X1 U10613 ( .A1(n8244), .A2(n10762), .A3(n8243), .ZN(n8249) );
  NAND2_X1 U10614 ( .A1(n13214), .A2(n10576), .ZN(n8245) );
  NAND2_X1 U10615 ( .A1(n8252), .A2(n8245), .ZN(n8246) );
  NAND2_X1 U10616 ( .A1(n8246), .A2(n11074), .ZN(n8248) );
  INV_X1 U10617 ( .A(n8251), .ZN(n8247) );
  AOI21_X1 U10618 ( .B1(n8249), .B2(n8248), .A(n8247), .ZN(n8256) );
  AOI21_X1 U10619 ( .B1(n8251), .B2(n8250), .A(n11074), .ZN(n8255) );
  NOR2_X1 U10620 ( .A1(n8252), .A2(n11074), .ZN(n8253) );
  NOR2_X1 U10621 ( .A1(n11013), .A2(n8253), .ZN(n8254) );
  OAI21_X1 U10622 ( .B1(n8256), .B2(n8255), .A(n8254), .ZN(n8257) );
  NAND2_X1 U10623 ( .A1(n8257), .A2(n11018), .ZN(n8265) );
  NAND2_X1 U10624 ( .A1(n8267), .A2(n8258), .ZN(n8260) );
  NAND2_X1 U10625 ( .A1(n8260), .A2(n10616), .ZN(n8264) );
  NOR2_X1 U10626 ( .A1(n8260), .A2(n8259), .ZN(n8262) );
  AND2_X1 U10627 ( .A1(n12690), .A2(n10918), .ZN(n8261) );
  MUX2_X1 U10628 ( .A(n8262), .B(n8261), .S(n11074), .Z(n8263) );
  AOI21_X1 U10629 ( .B1(n8265), .B2(n8264), .A(n8263), .ZN(n8271) );
  AOI21_X1 U10630 ( .B1(n8268), .B2(n8266), .A(n10616), .ZN(n8270) );
  MUX2_X1 U10631 ( .A(n8268), .B(n8267), .S(n11074), .Z(n8269) );
  OAI211_X1 U10632 ( .C1(n8271), .C2(n8270), .A(n11441), .B(n8269), .ZN(n8275)
         );
  MUX2_X1 U10633 ( .A(n8273), .B(n8272), .S(n10616), .Z(n8274) );
  NAND3_X1 U10634 ( .A1(n8275), .A2(n11047), .A3(n8274), .ZN(n8279) );
  NAND2_X1 U10635 ( .A1(n12688), .A2(n11735), .ZN(n8276) );
  MUX2_X1 U10636 ( .A(n8277), .B(n8276), .S(n11074), .Z(n8278) );
  NAND3_X1 U10637 ( .A1(n8279), .A2(n11600), .A3(n8278), .ZN(n8287) );
  INV_X1 U10638 ( .A(n8280), .ZN(n8281) );
  MUX2_X1 U10639 ( .A(n8282), .B(n8281), .S(n10616), .Z(n8283) );
  NOR2_X1 U10640 ( .A1(n8283), .A2(n15194), .ZN(n8286) );
  NOR2_X1 U10641 ( .A1(n8284), .A2(n11074), .ZN(n8285) );
  AOI21_X1 U10642 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8294) );
  INV_X1 U10643 ( .A(n14850), .ZN(n14852) );
  NAND2_X1 U10644 ( .A1(n14850), .A2(n8288), .ZN(n8291) );
  NAND3_X1 U10645 ( .A1(n8291), .A2(n8290), .A3(n8289), .ZN(n8292) );
  NAND2_X1 U10646 ( .A1(n8292), .A2(n11074), .ZN(n8293) );
  OAI21_X1 U10647 ( .B1(n8294), .B2(n14852), .A(n8293), .ZN(n8297) );
  AOI21_X1 U10648 ( .B1(n8296), .B2(n14842), .A(n11074), .ZN(n8295) );
  AOI21_X1 U10649 ( .B1(n8297), .B2(n8296), .A(n8295), .ZN(n8300) );
  INV_X1 U10650 ( .A(n13116), .ZN(n13114) );
  NAND3_X1 U10651 ( .A1(n12687), .A2(n14846), .A3(n10616), .ZN(n8298) );
  NAND3_X1 U10652 ( .A1(n13097), .A2(n13114), .A3(n8298), .ZN(n8299) );
  OR2_X1 U10653 ( .A1(n8300), .A2(n8299), .ZN(n8308) );
  MUX2_X1 U10654 ( .A(n8302), .B(n8301), .S(n11074), .Z(n8303) );
  NAND2_X1 U10655 ( .A1(n13097), .A2(n8303), .ZN(n8307) );
  NAND2_X1 U10656 ( .A1(n13289), .A2(n12686), .ZN(n8304) );
  MUX2_X1 U10657 ( .A(n8305), .B(n8304), .S(n11074), .Z(n8306) );
  NAND4_X1 U10658 ( .A1(n8308), .A2(n13087), .A3(n8307), .A4(n8306), .ZN(n8313) );
  NAND2_X1 U10659 ( .A1(n8316), .A2(n8309), .ZN(n8310) );
  NAND2_X1 U10660 ( .A1(n8310), .A2(n10616), .ZN(n8312) );
  INV_X1 U10661 ( .A(n8315), .ZN(n8311) );
  AOI21_X1 U10662 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(n8318) );
  AOI21_X1 U10663 ( .B1(n8315), .B2(n8314), .A(n10616), .ZN(n8317) );
  OAI22_X1 U10664 ( .A1(n8318), .A2(n8317), .B1(n10616), .B2(n8316), .ZN(n8324) );
  INV_X1 U10665 ( .A(n8319), .ZN(n8320) );
  NAND2_X1 U10666 ( .A1(n8325), .A2(n8320), .ZN(n8321) );
  NAND4_X1 U10667 ( .A1(n8332), .A2(n11074), .A3(n8322), .A4(n8321), .ZN(n8327) );
  AOI22_X1 U10668 ( .A1(n8324), .A2(n13061), .B1(n8323), .B2(n8327), .ZN(n8330) );
  NAND3_X1 U10669 ( .A1(n8331), .A2(n10616), .A3(n8325), .ZN(n8326) );
  NAND2_X1 U10670 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  OAI21_X1 U10671 ( .B1(n8330), .B2(n8329), .A(n8328), .ZN(n8334) );
  MUX2_X1 U10672 ( .A(n8332), .B(n8331), .S(n11074), .Z(n8333) );
  NAND2_X1 U10673 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  INV_X1 U10674 ( .A(n13017), .ZN(n13015) );
  NAND2_X1 U10675 ( .A1(n8335), .A2(n13015), .ZN(n8339) );
  MUX2_X1 U10676 ( .A(n8337), .B(n8336), .S(n10616), .Z(n8338) );
  NAND3_X1 U10677 ( .A1(n8339), .A2(n13011), .A3(n8338), .ZN(n8343) );
  MUX2_X1 U10678 ( .A(n8341), .B(n8340), .S(n11074), .Z(n8342) );
  NAND3_X1 U10679 ( .A1(n8343), .A2(n12986), .A3(n8342), .ZN(n8347) );
  MUX2_X1 U10680 ( .A(n8345), .B(n8344), .S(n10616), .Z(n8346) );
  NAND2_X1 U10681 ( .A1(n8347), .A2(n8346), .ZN(n8348) );
  NAND2_X1 U10682 ( .A1(n8348), .A2(n12977), .ZN(n8350) );
  NAND3_X1 U10683 ( .A1(n12974), .A2(n12965), .A3(n11074), .ZN(n8349) );
  NAND2_X1 U10684 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  NAND2_X1 U10685 ( .A1(n8351), .A2(n8104), .ZN(n8358) );
  NAND2_X1 U10686 ( .A1(n8353), .A2(n8352), .ZN(n8354) );
  NAND2_X1 U10687 ( .A1(n8354), .A2(n8356), .ZN(n8355) );
  MUX2_X1 U10688 ( .A(n8356), .B(n8355), .S(n10616), .Z(n8357) );
  NAND3_X1 U10689 ( .A1(n8358), .A2(n12952), .A3(n8357), .ZN(n8363) );
  OR2_X1 U10690 ( .A1(n12954), .A2(n12964), .ZN(n8360) );
  MUX2_X1 U10691 ( .A(n8360), .B(n8359), .S(n10616), .Z(n8361) );
  NAND3_X1 U10692 ( .A1(n8363), .A2(n8362), .A3(n8361), .ZN(n8367) );
  MUX2_X1 U10693 ( .A(n8365), .B(n8364), .S(n10616), .Z(n8366) );
  NAND2_X1 U10694 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND2_X1 U10695 ( .A1(n8368), .A2(n12921), .ZN(n8369) );
  INV_X1 U10696 ( .A(n8369), .ZN(n8375) );
  OAI21_X1 U10697 ( .B1(n12934), .B2(n12464), .A(n8369), .ZN(n8373) );
  NOR2_X1 U10698 ( .A1(n8370), .A2(n10616), .ZN(n8372) );
  AOI22_X1 U10699 ( .A1(n8373), .A2(n12905), .B1(n8372), .B2(n8371), .ZN(n8374) );
  AOI21_X1 U10700 ( .B1(n8375), .B2(n11074), .A(n8374), .ZN(n8378) );
  OAI21_X1 U10701 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8382) );
  INV_X1 U10702 ( .A(n8379), .ZN(n8380) );
  NAND3_X1 U10703 ( .A1(n8382), .A2(n8381), .A3(n8380), .ZN(n8386) );
  INV_X1 U10704 ( .A(n8383), .ZN(n8385) );
  AOI21_X1 U10705 ( .B1(n8386), .B2(n8385), .A(n8384), .ZN(n8387) );
  MUX2_X1 U10706 ( .A(n15232), .B(n10764), .S(n8387), .Z(n8388) );
  NAND2_X1 U10707 ( .A1(n6571), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8391) );
  NOR2_X1 U10708 ( .A1(n11073), .A2(P3_U3151), .ZN(n10713) );
  INV_X1 U10709 ( .A(n10713), .ZN(n11071) );
  NAND2_X1 U10710 ( .A1(n8394), .A2(n7702), .ZN(n11032) );
  INV_X1 U10711 ( .A(n11032), .ZN(n8403) );
  NAND2_X1 U10712 ( .A1(n8395), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8396) );
  MUX2_X1 U10713 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8396), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8398) );
  NAND2_X1 U10714 ( .A1(n7702), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8399) );
  MUX2_X1 U10715 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8399), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8401) );
  NOR2_X1 U10716 ( .A1(n10908), .A2(n11301), .ZN(n8402) );
  INV_X1 U10717 ( .A(n8404), .ZN(n12452) );
  NAND2_X1 U10718 ( .A1(n12452), .A2(n11143), .ZN(n11118) );
  NOR2_X1 U10719 ( .A1(n14857), .A2(n10618), .ZN(n8405) );
  NAND2_X1 U10720 ( .A1(n11070), .A2(n8405), .ZN(n10411) );
  NAND2_X1 U10721 ( .A1(n10713), .A2(n10777), .ZN(n8406) );
  OAI211_X1 U10722 ( .C1(n10411), .C2(n8404), .A(P3_B_REG_SCAN_IN), .B(n8406), 
        .ZN(n8407) );
  NOR2_X2 U10723 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n8411) );
  NOR2_X2 U10724 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8410) );
  AND4_X2 U10725 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n8416)
         );
  INV_X1 U10726 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8412) );
  NOR2_X2 U10727 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8417) );
  NAND3_X1 U10728 ( .A1(n8837), .A2(n8599), .A3(n8419), .ZN(n8420) );
  NOR2_X1 U10729 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8424) );
  NOR2_X1 U10730 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8423) );
  NOR2_X1 U10731 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8422) );
  INV_X1 U10732 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8425) );
  INV_X1 U10733 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8444) );
  NAND4_X1 U10734 ( .A1(n8425), .A2(n8444), .A3(n9235), .A4(n9236), .ZN(n8450)
         );
  INV_X1 U10735 ( .A(n8429), .ZN(n8427) );
  NAND2_X1 U10736 ( .A1(n8427), .A2(n8426), .ZN(n13981) );
  NAND2_X1 U10737 ( .A1(n8536), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U10738 ( .A1(n8510), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10739 ( .A1(n8511), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10740 ( .A1(n9160), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8435) );
  INV_X1 U10741 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10742 ( .A1(n9716), .A2(SI_0_), .ZN(n8439) );
  NAND2_X1 U10743 ( .A1(n8439), .A2(n8438), .ZN(n8441) );
  INV_X4 U10744 ( .A(n8598), .ZN(n9716) );
  AND2_X1 U10745 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10746 ( .A1(n9716), .A2(n8440), .ZN(n8486) );
  NAND2_X1 U10747 ( .A1(n8441), .A2(n8486), .ZN(n14003) );
  AND2_X1 U10748 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n8448) );
  AND3_X1 U10749 ( .A1(n8444), .A2(n9235), .A3(n9236), .ZN(n8445) );
  NAND2_X1 U10750 ( .A1(n9211), .A2(n9673), .ZN(n9625) );
  INV_X1 U10751 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8451) );
  INV_X1 U10752 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8453) );
  INV_X1 U10753 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10754 ( .A1(n8456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8457) );
  XNOR2_X2 U10755 ( .A(n8457), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U10756 ( .A1(n8482), .A2(n10304), .ZN(n8465) );
  OAI21_X1 U10757 ( .B1(n8459), .B2(n13982), .A(P2_IR_REG_20__SCAN_IN), .ZN(
        n8462) );
  NAND2_X1 U10758 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8460), .ZN(n8461) );
  NAND2_X1 U10759 ( .A1(n8462), .A2(n8461), .ZN(n8463) );
  NAND2_X1 U10760 ( .A1(n8465), .A2(n10305), .ZN(n8473) );
  NAND2_X1 U10761 ( .A1(n8471), .A2(n8466), .ZN(n9095) );
  OAI21_X1 U10762 ( .B1(n9095), .B2(n9231), .A(n10541), .ZN(n8467) );
  INV_X1 U10763 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8469) );
  INV_X1 U10764 ( .A(n9234), .ZN(n9141) );
  INV_X1 U10765 ( .A(n8471), .ZN(n9621) );
  INV_X1 U10766 ( .A(n8482), .ZN(n9232) );
  NAND3_X2 U10767 ( .A1(n8472), .A2(n10305), .A3(n9097), .ZN(n8544) );
  OAI211_X1 U10768 ( .C1(n9673), .C2(n8473), .A(n8544), .B(n9211), .ZN(n8474)
         );
  NAND2_X1 U10769 ( .A1(n8475), .A2(n8474), .ZN(n8495) );
  NAND2_X1 U10770 ( .A1(n8510), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8480) );
  INV_X1 U10771 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10772 ( .A1(n9160), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10773 ( .A1(n8536), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U10774 ( .A1(n8544), .A2(n13489), .ZN(n8490) );
  NAND2_X1 U10775 ( .A1(n8484), .A2(n8483), .ZN(n8505) );
  AND2_X1 U10776 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8485) );
  NAND2_X1 U10777 ( .A1(n8598), .A2(n8485), .ZN(n9718) );
  NAND2_X1 U10778 ( .A1(n9718), .A2(n8486), .ZN(n8503) );
  XNOR2_X1 U10779 ( .A(n8499), .B(n8503), .ZN(n9855) );
  NAND2_X1 U10780 ( .A1(n9855), .A2(n8786), .ZN(n8488) );
  NAND2_X1 U10781 ( .A1(n8922), .A2(n9644), .ZN(n8489) );
  NAND2_X1 U10782 ( .A1(n8490), .A2(n8489), .ZN(n8496) );
  NAND2_X1 U10783 ( .A1(n8495), .A2(n8496), .ZN(n8494) );
  NAND2_X1 U10784 ( .A1(n8922), .A2(n13489), .ZN(n8492) );
  NAND2_X1 U10785 ( .A1(n8544), .A2(n9644), .ZN(n8491) );
  NAND2_X1 U10786 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  INV_X1 U10787 ( .A(n8495), .ZN(n8498) );
  INV_X1 U10788 ( .A(n8496), .ZN(n8497) );
  NAND2_X1 U10789 ( .A1(n8498), .A2(n8497), .ZN(n8521) );
  INV_X1 U10790 ( .A(n8500), .ZN(n8501) );
  INV_X1 U10791 ( .A(SI_1_), .ZN(n9331) );
  NOR2_X1 U10792 ( .A1(n8501), .A2(n9331), .ZN(n8502) );
  XNOR2_X1 U10793 ( .A(n8527), .B(n8528), .ZN(n9959) );
  NAND2_X1 U10794 ( .A1(n9959), .A2(n8786), .ZN(n8509) );
  NAND2_X1 U10795 ( .A1(n8505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8504) );
  MUX2_X1 U10796 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8504), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8508) );
  INV_X1 U10797 ( .A(n8505), .ZN(n8507) );
  INV_X1 U10798 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U10799 ( .A1(n8507), .A2(n8506), .ZN(n8533) );
  NAND2_X1 U10800 ( .A1(n8508), .A2(n8533), .ZN(n13496) );
  INV_X1 U10801 ( .A(n13496), .ZN(n9415) );
  NAND2_X1 U10802 ( .A1(n8510), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10803 ( .A1(n9160), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10804 ( .A1(n8536), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U10805 ( .A1(n8511), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8512) );
  NAND4_X2 U10806 ( .A1(n8515), .A2(n8514), .A3(n8513), .A4(n8512), .ZN(n9210)
         );
  NAND2_X1 U10807 ( .A1(n8544), .A2(n9210), .ZN(n8516) );
  NAND2_X1 U10808 ( .A1(n8544), .A2(n10053), .ZN(n8519) );
  NAND2_X1 U10809 ( .A1(n8922), .A2(n9210), .ZN(n8518) );
  NAND2_X1 U10810 ( .A1(n8519), .A2(n8518), .ZN(n8522) );
  NAND2_X1 U10811 ( .A1(n8523), .A2(n8522), .ZN(n8520) );
  INV_X1 U10812 ( .A(n8522), .ZN(n8525) );
  INV_X1 U10813 ( .A(n8523), .ZN(n8524) );
  NAND2_X1 U10814 ( .A1(n8525), .A2(n8524), .ZN(n8526) );
  INV_X1 U10815 ( .A(n8529), .ZN(n8530) );
  NAND2_X1 U10816 ( .A1(n8530), .A2(SI_2_), .ZN(n8531) );
  MUX2_X1 U10817 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n11950), .Z(n8553) );
  XNOR2_X1 U10818 ( .A(n8553), .B(SI_3_), .ZN(n8550) );
  NAND2_X1 U10819 ( .A1(n8533), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10820 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8532), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8534) );
  OR2_X1 U10821 ( .A1(n8533), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10822 ( .A1(n10684), .A2(n8922), .ZN(n8543) );
  NAND2_X1 U10823 ( .A1(n8510), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8541) );
  INV_X1 U10824 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10825 ( .A1(n9160), .A2(n8535), .ZN(n8540) );
  INV_X1 U10826 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10827 ( .A1(n8511), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10828 ( .A1(n8544), .A2(n13488), .ZN(n8542) );
  NAND2_X1 U10829 ( .A1(n8543), .A2(n8542), .ZN(n8547) );
  AOI22_X1 U10830 ( .A1(n8544), .A2(n10684), .B1(n13488), .B2(n8922), .ZN(
        n8545) );
  AOI21_X1 U10831 ( .B1(n8548), .B2(n8547), .A(n8545), .ZN(n8546) );
  INV_X1 U10832 ( .A(n8546), .ZN(n8549) );
  INV_X1 U10833 ( .A(n8550), .ZN(n8551) );
  NAND2_X1 U10834 ( .A1(n8553), .A2(SI_3_), .ZN(n8554) );
  NAND2_X1 U10835 ( .A1(n8555), .A2(n8554), .ZN(n8575) );
  MUX2_X1 U10836 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n11950), .Z(n8576) );
  XNOR2_X1 U10837 ( .A(n8576), .B(SI_4_), .ZN(n8573) );
  XNOR2_X1 U10838 ( .A(n8575), .B(n8573), .ZN(n10227) );
  NAND2_X1 U10839 ( .A1(n10227), .A2(n8786), .ZN(n8559) );
  NAND2_X1 U10840 ( .A1(n8556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8557) );
  XNOR2_X1 U10841 ( .A(n8557), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U10842 ( .A1(n8907), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8906), .B2(
        n9599), .ZN(n8558) );
  NAND2_X1 U10843 ( .A1(n8559), .A2(n8558), .ZN(n10644) );
  NAND2_X1 U10844 ( .A1(n10644), .A2(n9165), .ZN(n8567) );
  INV_X1 U10845 ( .A(n8922), .ZN(n9198) );
  NAND2_X1 U10846 ( .A1(n8511), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10847 ( .A1(n8510), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8564) );
  NOR2_X1 U10848 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8561) );
  NOR2_X1 U10849 ( .A1(n8583), .A2(n8561), .ZN(n10643) );
  NAND2_X1 U10850 ( .A1(n9160), .A2(n10643), .ZN(n8563) );
  INV_X2 U10851 ( .A(n9094), .ZN(n9136) );
  NAND2_X1 U10852 ( .A1(n9136), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8562) );
  NAND4_X1 U10853 ( .A1(n8565), .A2(n8564), .A3(n8563), .A4(n8562), .ZN(n13487) );
  NAND2_X1 U10854 ( .A1(n9196), .A2(n13487), .ZN(n8566) );
  NAND2_X1 U10855 ( .A1(n8567), .A2(n8566), .ZN(n8570) );
  AOI22_X1 U10856 ( .A1(n10644), .A2(n9172), .B1(n13487), .B2(n9165), .ZN(
        n8568) );
  INV_X1 U10857 ( .A(n8569), .ZN(n8572) );
  INV_X1 U10858 ( .A(n8573), .ZN(n8574) );
  NAND2_X1 U10859 ( .A1(n8575), .A2(n8574), .ZN(n8578) );
  NAND2_X1 U10860 ( .A1(n8576), .A2(SI_4_), .ZN(n8577) );
  MUX2_X1 U10861 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9716), .Z(n8596) );
  XNOR2_X1 U10862 ( .A(n8596), .B(SI_5_), .ZN(n8593) );
  XNOR2_X1 U10863 ( .A(n8595), .B(n8593), .ZN(n10232) );
  NAND2_X1 U10864 ( .A1(n10232), .A2(n8786), .ZN(n8582) );
  INV_X1 U10865 ( .A(n8579), .ZN(n8600) );
  OR2_X1 U10866 ( .A1(n8600), .A2(n13982), .ZN(n8580) );
  XNOR2_X1 U10867 ( .A(n8580), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9443) );
  AOI22_X1 U10868 ( .A1(n8907), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8906), .B2(
        n9443), .ZN(n8581) );
  NAND2_X1 U10869 ( .A1(n8582), .A2(n8581), .ZN(n10319) );
  NAND2_X1 U10870 ( .A1(n10319), .A2(n9172), .ZN(n8589) );
  NAND2_X1 U10871 ( .A1(n8583), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8605) );
  OAI21_X1 U10872 ( .B1(n8583), .B2(P2_REG3_REG_5__SCAN_IN), .A(n8605), .ZN(
        n10320) );
  OR2_X1 U10873 ( .A1(n9114), .A2(n10320), .ZN(n8587) );
  NAND2_X1 U10874 ( .A1(n8510), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U10875 ( .A1(n8511), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U10876 ( .A1(n9136), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8584) );
  NAND4_X1 U10877 ( .A1(n8587), .A2(n8586), .A3(n8585), .A4(n8584), .ZN(n13486) );
  NAND2_X1 U10878 ( .A1(n9165), .A2(n13486), .ZN(n8588) );
  NAND2_X1 U10879 ( .A1(n8589), .A2(n8588), .ZN(n8591) );
  INV_X1 U10880 ( .A(n9198), .ZN(n9172) );
  AOI22_X1 U10881 ( .A1(n10319), .A2(n9165), .B1(n9172), .B2(n13486), .ZN(
        n8590) );
  INV_X1 U10882 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U10883 ( .A1(n8596), .A2(SI_5_), .ZN(n8597) );
  MUX2_X1 U10884 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9040), .Z(n8625) );
  XNOR2_X1 U10885 ( .A(n8625), .B(SI_6_), .ZN(n8623) );
  NAND2_X1 U10886 ( .A1(n10270), .A2(n8786), .ZN(n8603) );
  NAND2_X1 U10887 ( .A1(n8600), .A2(n8599), .ZN(n8836) );
  NAND2_X1 U10888 ( .A1(n8836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U10889 ( .A(n8601), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9544) );
  AOI22_X1 U10890 ( .A1(n8907), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8906), .B2(
        n9544), .ZN(n8602) );
  NAND2_X1 U10891 ( .A1(n10334), .A2(n9165), .ZN(n8612) );
  NAND2_X1 U10892 ( .A1(n8510), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10893 ( .A1(n9136), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8609) );
  AND2_X1 U10894 ( .A1(n8605), .A2(n8604), .ZN(n8606) );
  NOR2_X1 U10895 ( .A1(n8629), .A2(n8606), .ZN(n10141) );
  NAND2_X1 U10896 ( .A1(n9160), .A2(n10141), .ZN(n8608) );
  NAND2_X1 U10897 ( .A1(n8511), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8607) );
  NAND4_X1 U10898 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), .ZN(n13485) );
  NAND2_X1 U10899 ( .A1(n9172), .A2(n13485), .ZN(n8611) );
  NAND2_X1 U10900 ( .A1(n8612), .A2(n8611), .ZN(n8618) );
  INV_X1 U10901 ( .A(n13485), .ZN(n10333) );
  NAND2_X1 U10902 ( .A1(n10334), .A2(n9196), .ZN(n8613) );
  OAI21_X1 U10903 ( .B1(n10333), .B2(n8614), .A(n8613), .ZN(n8615) );
  NAND2_X1 U10904 ( .A1(n8616), .A2(n8615), .ZN(n8622) );
  INV_X1 U10905 ( .A(n8617), .ZN(n8620) );
  INV_X1 U10906 ( .A(n8618), .ZN(n8619) );
  NAND2_X1 U10907 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  INV_X1 U10908 ( .A(n8623), .ZN(n8624) );
  MUX2_X1 U10909 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9040), .Z(n8643) );
  XNOR2_X1 U10910 ( .A(n8643), .B(SI_7_), .ZN(n8640) );
  XNOR2_X1 U10911 ( .A(n8642), .B(n8640), .ZN(n10476) );
  NAND2_X1 U10912 ( .A1(n10476), .A2(n8786), .ZN(n8628) );
  NAND2_X1 U10913 ( .A1(n8646), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8626) );
  XNOR2_X1 U10914 ( .A(n8626), .B(P2_IR_REG_7__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U10915 ( .A1(n8907), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8906), .B2(
        n15124), .ZN(n8627) );
  NAND2_X1 U10916 ( .A1(n8628), .A2(n8627), .ZN(n15178) );
  NAND2_X1 U10917 ( .A1(n15178), .A2(n9196), .ZN(n8636) );
  NAND2_X1 U10918 ( .A1(n9155), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U10919 ( .A1(n8510), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U10920 ( .A1(n8629), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8655) );
  OR2_X1 U10921 ( .A1(n8629), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8630) );
  AND2_X1 U10922 ( .A1(n8655), .A2(n8630), .ZN(n10339) );
  NAND2_X1 U10923 ( .A1(n9160), .A2(n10339), .ZN(n8632) );
  NAND2_X1 U10924 ( .A1(n9136), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8631) );
  NAND4_X1 U10925 ( .A1(n8634), .A2(n8633), .A3(n8632), .A4(n8631), .ZN(n13484) );
  NAND2_X1 U10926 ( .A1(n9165), .A2(n13484), .ZN(n8635) );
  NAND2_X1 U10927 ( .A1(n8636), .A2(n8635), .ZN(n8638) );
  AOI22_X1 U10928 ( .A1(n15178), .A2(n9165), .B1(n9172), .B2(n13484), .ZN(
        n8637) );
  INV_X1 U10929 ( .A(n8640), .ZN(n8641) );
  NAND2_X1 U10930 ( .A1(n8643), .A2(SI_7_), .ZN(n8644) );
  NAND2_X1 U10931 ( .A1(n8645), .A2(n8644), .ZN(n8666) );
  MUX2_X1 U10932 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9040), .Z(n8667) );
  XNOR2_X1 U10933 ( .A(n8667), .B(SI_8_), .ZN(n8664) );
  XNOR2_X1 U10934 ( .A(n8666), .B(n8664), .ZN(n10739) );
  NAND2_X1 U10935 ( .A1(n10739), .A2(n8786), .ZN(n8653) );
  NOR2_X1 U10936 ( .A1(n8649), .A2(n13982), .ZN(n8647) );
  MUX2_X1 U10937 ( .A(n13982), .B(n8647), .S(P2_IR_REG_8__SCAN_IN), .Z(n8651)
         );
  NAND2_X1 U10938 ( .A1(n8649), .A2(n8648), .ZN(n8670) );
  INV_X1 U10939 ( .A(n8670), .ZN(n8650) );
  NOR2_X1 U10940 ( .A1(n8651), .A2(n8650), .ZN(n9807) );
  AOI22_X1 U10941 ( .A1(n8906), .A2(n9807), .B1(n8907), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U10942 ( .A1(n10552), .A2(n9165), .ZN(n8662) );
  NAND2_X1 U10943 ( .A1(n9155), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U10944 ( .A1(n8510), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8659) );
  INV_X1 U10945 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10946 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  AND2_X1 U10947 ( .A1(n8674), .A2(n8656), .ZN(n10439) );
  NAND2_X1 U10948 ( .A1(n9160), .A2(n10439), .ZN(n8658) );
  NAND2_X1 U10949 ( .A1(n9136), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8657) );
  NAND4_X1 U10950 ( .A1(n8660), .A2(n8659), .A3(n8658), .A4(n8657), .ZN(n13483) );
  NAND2_X1 U10951 ( .A1(n9172), .A2(n13483), .ZN(n8661) );
  AOI22_X1 U10952 ( .A1(n10552), .A2(n9196), .B1(n13483), .B2(n9165), .ZN(
        n8663) );
  INV_X1 U10953 ( .A(n8664), .ZN(n8665) );
  NAND2_X1 U10954 ( .A1(n8667), .A2(SI_8_), .ZN(n8668) );
  MUX2_X1 U10955 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9040), .Z(n8691) );
  XNOR2_X1 U10956 ( .A(n8691), .B(SI_9_), .ZN(n8688) );
  XNOR2_X1 U10957 ( .A(n8690), .B(n8688), .ZN(n10820) );
  NAND2_X1 U10958 ( .A1(n10820), .A2(n8786), .ZN(n8673) );
  NAND2_X1 U10959 ( .A1(n8670), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8669) );
  MUX2_X1 U10960 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8669), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8671) );
  AOI22_X1 U10961 ( .A1(n8906), .A2(n9912), .B1(n8907), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U10962 ( .A1(n10723), .A2(n9196), .ZN(n8681) );
  NAND2_X1 U10963 ( .A1(n9155), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U10964 ( .A1(n8510), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8678) );
  AND2_X1 U10965 ( .A1(n8674), .A2(n10729), .ZN(n8675) );
  NOR2_X1 U10966 ( .A1(n8696), .A2(n8675), .ZN(n10731) );
  NAND2_X1 U10967 ( .A1(n9160), .A2(n10731), .ZN(n8677) );
  NAND2_X1 U10968 ( .A1(n9136), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8676) );
  NAND4_X1 U10969 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n13482) );
  NAND2_X1 U10970 ( .A1(n9165), .A2(n13482), .ZN(n8680) );
  NAND2_X1 U10971 ( .A1(n10723), .A2(n9165), .ZN(n8683) );
  NAND2_X1 U10972 ( .A1(n8922), .A2(n13482), .ZN(n8682) );
  NAND2_X1 U10973 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  NAND2_X1 U10974 ( .A1(n8685), .A2(n8684), .ZN(n8687) );
  NAND2_X1 U10975 ( .A1(n6528), .A2(n6452), .ZN(n8686) );
  INV_X1 U10976 ( .A(n8688), .ZN(n8689) );
  MUX2_X1 U10977 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9040), .Z(n8709) );
  XNOR2_X1 U10978 ( .A(n8709), .B(SI_10_), .ZN(n8692) );
  XNOR2_X1 U10979 ( .A(n8708), .B(n8692), .ZN(n10825) );
  NAND2_X1 U10980 ( .A1(n10825), .A2(n8786), .ZN(n8695) );
  NAND2_X1 U10981 ( .A1(n8714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8693) );
  XNOR2_X1 U10982 ( .A(n8693), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U10983 ( .A1(n9994), .A2(n8906), .B1(n8907), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U10984 ( .A1(n11010), .A2(n9165), .ZN(n8703) );
  NOR2_X1 U10985 ( .A1(n8696), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8697) );
  OR2_X1 U10986 ( .A1(n8718), .A2(n8697), .ZN(n10999) );
  OR2_X1 U10987 ( .A1(n9114), .A2(n10999), .ZN(n8701) );
  NAND2_X1 U10988 ( .A1(n8510), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U10989 ( .A1(n8511), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U10990 ( .A1(n9136), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8698) );
  NAND4_X1 U10991 ( .A1(n8701), .A2(n8700), .A3(n8699), .A4(n8698), .ZN(n13481) );
  NAND2_X1 U10992 ( .A1(n9196), .A2(n13481), .ZN(n8702) );
  NAND2_X1 U10993 ( .A1(n8703), .A2(n8702), .ZN(n8705) );
  AOI22_X1 U10994 ( .A1(n11010), .A2(n9196), .B1(n13481), .B2(n9165), .ZN(
        n8704) );
  INV_X1 U10995 ( .A(n8709), .ZN(n8706) );
  NAND2_X1 U10996 ( .A1(n8706), .A2(n9294), .ZN(n8707) );
  NAND2_X1 U10997 ( .A1(n8709), .A2(SI_10_), .ZN(n8710) );
  MUX2_X1 U10998 ( .A(n9572), .B(n9566), .S(n9040), .Z(n8711) );
  INV_X1 U10999 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U11000 ( .A1(n8712), .A2(SI_11_), .ZN(n8713) );
  XNOR2_X1 U11001 ( .A(n8738), .B(n8737), .ZN(n11321) );
  NAND2_X1 U11002 ( .A1(n11321), .A2(n8786), .ZN(n8717) );
  OR2_X1 U11003 ( .A1(n8743), .A2(n13982), .ZN(n8715) );
  XNOR2_X1 U11004 ( .A(n8715), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U11005 ( .A1(n10006), .A2(n8906), .B1(n8907), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11006 ( .A1(n11412), .A2(n9196), .ZN(n8725) );
  NAND2_X1 U11007 ( .A1(n8510), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11008 ( .A1(n8511), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8722) );
  OR2_X1 U11009 ( .A1(n8718), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8719) );
  AND2_X1 U11010 ( .A1(n8753), .A2(n8719), .ZN(n11401) );
  NAND2_X1 U11011 ( .A1(n9160), .A2(n11401), .ZN(n8721) );
  NAND2_X1 U11012 ( .A1(n9136), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8720) );
  NAND4_X1 U11013 ( .A1(n8723), .A2(n8722), .A3(n8721), .A4(n8720), .ZN(n13480) );
  NAND2_X1 U11014 ( .A1(n9165), .A2(n13480), .ZN(n8724) );
  NAND2_X1 U11015 ( .A1(n8725), .A2(n8724), .ZN(n8731) );
  NAND2_X1 U11016 ( .A1(n8730), .A2(n8731), .ZN(n8729) );
  NAND2_X1 U11017 ( .A1(n11412), .A2(n9165), .ZN(n8727) );
  NAND2_X1 U11018 ( .A1(n8922), .A2(n13480), .ZN(n8726) );
  NAND2_X1 U11019 ( .A1(n8727), .A2(n8726), .ZN(n8728) );
  NAND2_X1 U11020 ( .A1(n8729), .A2(n8728), .ZN(n8735) );
  INV_X1 U11021 ( .A(n8730), .ZN(n8733) );
  INV_X1 U11022 ( .A(n8731), .ZN(n8732) );
  NAND2_X1 U11023 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  MUX2_X1 U11024 ( .A(n9763), .B(n9764), .S(n9040), .Z(n8739) );
  INV_X1 U11025 ( .A(n8739), .ZN(n8740) );
  NAND2_X1 U11026 ( .A1(n8740), .A2(SI_12_), .ZN(n8741) );
  XNOR2_X1 U11027 ( .A(n8764), .B(n7666), .ZN(n11466) );
  NAND2_X1 U11028 ( .A1(n11466), .A2(n8786), .ZN(n8752) );
  INV_X1 U11029 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8742) );
  NOR2_X1 U11030 ( .A1(n8746), .A2(n13982), .ZN(n8744) );
  MUX2_X1 U11031 ( .A(n13982), .B(n8744), .S(P2_IR_REG_12__SCAN_IN), .Z(n8748)
         );
  INV_X1 U11032 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11033 ( .A1(n8746), .A2(n8745), .ZN(n8770) );
  INV_X1 U11034 ( .A(n8770), .ZN(n8747) );
  OAI22_X1 U11035 ( .A1(n11270), .A2(n9393), .B1(n9152), .B2(n9764), .ZN(n8750) );
  INV_X1 U11036 ( .A(n8750), .ZN(n8751) );
  NAND2_X1 U11037 ( .A1(n13847), .A2(n9165), .ZN(n8760) );
  NAND2_X1 U11038 ( .A1(n9155), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11039 ( .A1(n8510), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11040 ( .A1(n8753), .A2(n11435), .ZN(n8754) );
  AND2_X1 U11041 ( .A1(n8775), .A2(n8754), .ZN(n13840) );
  NAND2_X1 U11042 ( .A1(n9160), .A2(n13840), .ZN(n8756) );
  NAND2_X1 U11043 ( .A1(n9136), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8755) );
  NAND4_X1 U11044 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n13479) );
  NAND2_X1 U11045 ( .A1(n9172), .A2(n13479), .ZN(n8759) );
  NAND2_X1 U11046 ( .A1(n8760), .A2(n8759), .ZN(n8762) );
  AOI22_X1 U11047 ( .A1(n13847), .A2(n9196), .B1(n13479), .B2(n9165), .ZN(
        n8761) );
  MUX2_X1 U11048 ( .A(n9902), .B(n6931), .S(n9040), .Z(n8766) );
  NAND2_X1 U11049 ( .A1(n8766), .A2(n9375), .ZN(n8784) );
  INV_X1 U11050 ( .A(n8766), .ZN(n8767) );
  NAND2_X1 U11051 ( .A1(n8767), .A2(SI_13_), .ZN(n8768) );
  XNOR2_X1 U11052 ( .A(n8783), .B(n7659), .ZN(n11472) );
  NAND2_X1 U11053 ( .A1(n11472), .A2(n8786), .ZN(n8774) );
  NAND2_X1 U11054 ( .A1(n8770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8769) );
  MUX2_X1 U11055 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8769), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8771) );
  NAND2_X1 U11056 ( .A1(n8771), .A2(n8814), .ZN(n15142) );
  OAI22_X1 U11057 ( .A1(n15142), .A2(n9393), .B1(n9152), .B2(n6931), .ZN(n8772) );
  INV_X1 U11058 ( .A(n8772), .ZN(n8773) );
  NAND2_X1 U11059 ( .A1(n11678), .A2(n9196), .ZN(n8780) );
  AND2_X1 U11060 ( .A1(n8775), .A2(n11555), .ZN(n8776) );
  OR2_X1 U11061 ( .A1(n8790), .A2(n8776), .ZN(n11558) );
  AOI22_X1 U11062 ( .A1(n9155), .A2(P2_REG0_REG_13__SCAN_IN), .B1(n9136), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11063 ( .A1(n8510), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8777) );
  OAI211_X1 U11064 ( .C1(n11558), .C2(n9114), .A(n8778), .B(n8777), .ZN(n13478) );
  NAND2_X1 U11065 ( .A1(n13478), .A2(n9165), .ZN(n8779) );
  AOI22_X1 U11066 ( .A1(n11678), .A2(n9165), .B1(n9172), .B2(n13478), .ZN(
        n8781) );
  INV_X1 U11067 ( .A(n8781), .ZN(n8782) );
  MUX2_X1 U11068 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9040), .Z(n8809) );
  XNOR2_X1 U11069 ( .A(n8810), .B(n8809), .ZN(n11763) );
  NAND2_X1 U11070 ( .A1(n11763), .A2(n8786), .ZN(n8789) );
  NAND2_X1 U11071 ( .A1(n8814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8787) );
  XNOR2_X1 U11072 ( .A(n8787), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U11073 ( .A1(n13524), .A2(n8906), .B1(n8907), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U11074 ( .A1(n14887), .A2(n9165), .ZN(n8798) );
  INV_X1 U11075 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8796) );
  INV_X1 U11076 ( .A(n8790), .ZN(n8792) );
  INV_X1 U11077 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11078 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  NAND2_X1 U11079 ( .A1(n8819), .A2(n8793), .ZN(n14890) );
  OR2_X1 U11080 ( .A1(n14890), .A2(n9114), .ZN(n8795) );
  AOI22_X1 U11081 ( .A1(n8510), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9136), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n8794) );
  OAI211_X1 U11082 ( .C1(n8962), .C2(n8796), .A(n8795), .B(n8794), .ZN(n13477)
         );
  NAND2_X1 U11083 ( .A1(n13477), .A2(n9196), .ZN(n8797) );
  NAND2_X1 U11084 ( .A1(n14887), .A2(n9196), .ZN(n8800) );
  NAND2_X1 U11085 ( .A1(n13477), .A2(n9165), .ZN(n8799) );
  NAND2_X1 U11086 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  NAND2_X1 U11087 ( .A1(n8802), .A2(n8801), .ZN(n8808) );
  NAND2_X1 U11088 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  MUX2_X1 U11089 ( .A(n10220), .B(n10213), .S(n9040), .Z(n8811) );
  NAND2_X1 U11090 ( .A1(n8811), .A2(n9604), .ZN(n8830) );
  INV_X1 U11091 ( .A(n8811), .ZN(n8812) );
  NAND2_X1 U11092 ( .A1(n8812), .A2(SI_15_), .ZN(n8813) );
  XNOR2_X1 U11093 ( .A(n8829), .B(n8828), .ZN(n11787) );
  NAND2_X1 U11094 ( .A1(n11787), .A2(n8786), .ZN(n8817) );
  OAI21_X1 U11095 ( .B1(n8814), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U11096 ( .A(n8815), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15156) );
  AOI22_X1 U11097 ( .A1(n15156), .A2(n8906), .B1(n8907), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11098 ( .A1(n11863), .A2(n9196), .ZN(n8825) );
  INV_X1 U11099 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8823) );
  INV_X1 U11100 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n15406) );
  NAND2_X1 U11101 ( .A1(n8819), .A2(n15406), .ZN(n8820) );
  NAND2_X1 U11102 ( .A1(n8865), .A2(n8820), .ZN(n11829) );
  OR2_X1 U11103 ( .A1(n11829), .A2(n9114), .ZN(n8822) );
  AOI22_X1 U11104 ( .A1(n8511), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n8510), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U11105 ( .C1(n9094), .C2(n8823), .A(n8822), .B(n8821), .ZN(n13476)
         );
  NAND2_X1 U11106 ( .A1(n13476), .A2(n9165), .ZN(n8824) );
  NAND2_X1 U11107 ( .A1(n8825), .A2(n8824), .ZN(n8827) );
  AOI22_X1 U11108 ( .A1(n11863), .A2(n9165), .B1(n9172), .B2(n13476), .ZN(
        n8826) );
  MUX2_X1 U11109 ( .A(n15443), .B(n10296), .S(n9040), .Z(n8832) );
  NAND2_X1 U11110 ( .A1(n8832), .A2(n9655), .ZN(n8852) );
  INV_X1 U11111 ( .A(n8832), .ZN(n8833) );
  NAND2_X1 U11112 ( .A1(n8833), .A2(SI_16_), .ZN(n8834) );
  XNOR2_X1 U11113 ( .A(n8851), .B(n8850), .ZN(n12020) );
  NAND2_X1 U11114 ( .A1(n12020), .A2(n8786), .ZN(n8840) );
  OR2_X1 U11115 ( .A1(n8836), .A2(n8835), .ZN(n8857) );
  NAND2_X1 U11116 ( .A1(n8857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8838) );
  XNOR2_X1 U11117 ( .A(n8838), .B(n8837), .ZN(n11511) );
  INV_X1 U11118 ( .A(n11511), .ZN(n11277) );
  AOI22_X1 U11119 ( .A1(n8907), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8906), 
        .B2(n11277), .ZN(n8839) );
  NAND2_X1 U11120 ( .A1(n13607), .A2(n9165), .ZN(n8847) );
  XNOR2_X1 U11121 ( .A(n8865), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U11122 ( .A1(n13412), .A2(n9160), .ZN(n8845) );
  INV_X1 U11123 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11858) );
  NAND2_X1 U11124 ( .A1(n9155), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11125 ( .A1(n9136), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8841) );
  OAI211_X1 U11126 ( .C1(n8560), .C2(n11858), .A(n8842), .B(n8841), .ZN(n8843)
         );
  INV_X1 U11127 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U11128 ( .A1(n8845), .A2(n8844), .ZN(n13578) );
  NAND2_X1 U11129 ( .A1(n13578), .A2(n9196), .ZN(n8846) );
  INV_X1 U11130 ( .A(n13578), .ZN(n13606) );
  NAND2_X1 U11131 ( .A1(n13607), .A2(n9196), .ZN(n8848) );
  OAI21_X1 U11132 ( .B1(n13606), .B2(n8614), .A(n8848), .ZN(n8849) );
  NAND2_X1 U11133 ( .A1(n8851), .A2(n8850), .ZN(n8853) );
  MUX2_X1 U11134 ( .A(n10532), .B(n10534), .S(n9040), .Z(n8854) );
  INV_X1 U11135 ( .A(SI_17_), .ZN(n9835) );
  NAND2_X1 U11136 ( .A1(n8854), .A2(n9835), .ZN(n8880) );
  INV_X1 U11137 ( .A(n8854), .ZN(n8855) );
  NAND2_X1 U11138 ( .A1(n8855), .A2(SI_17_), .ZN(n8856) );
  XNOR2_X1 U11139 ( .A(n8879), .B(n8878), .ZN(n11991) );
  NAND2_X1 U11140 ( .A1(n11991), .A2(n8786), .ZN(n8861) );
  OAI21_X1 U11141 ( .B1(n8857), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8858) );
  MUX2_X1 U11142 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8858), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8859) );
  NAND2_X1 U11143 ( .A1(n8859), .A2(n8881), .ZN(n13537) );
  INV_X1 U11144 ( .A(n13537), .ZN(n13530) );
  AOI22_X1 U11145 ( .A1(n8907), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8906), 
        .B2(n13530), .ZN(n8860) );
  NAND2_X1 U11146 ( .A1(n13930), .A2(n9196), .ZN(n8873) );
  INV_X1 U11147 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8863) );
  INV_X1 U11148 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8862) );
  OAI21_X1 U11149 ( .B1(n8865), .B2(n8863), .A(n8862), .ZN(n8866) );
  NAND2_X1 U11150 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8864) );
  AND2_X1 U11151 ( .A1(n8866), .A2(n8885), .ZN(n13827) );
  NAND2_X1 U11152 ( .A1(n13827), .A2(n9160), .ZN(n8871) );
  INV_X1 U11153 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13831) );
  NAND2_X1 U11154 ( .A1(n8511), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U11155 ( .A1(n9136), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8867) );
  OAI211_X1 U11156 ( .C1(n8560), .C2(n13831), .A(n8868), .B(n8867), .ZN(n8869)
         );
  INV_X1 U11157 ( .A(n8869), .ZN(n8870) );
  NAND2_X1 U11158 ( .A1(n8871), .A2(n8870), .ZN(n13581) );
  NAND2_X1 U11159 ( .A1(n13581), .A2(n9165), .ZN(n8872) );
  NAND2_X1 U11160 ( .A1(n8873), .A2(n8872), .ZN(n8875) );
  AOI22_X1 U11161 ( .A1(n13930), .A2(n9165), .B1(n9172), .B2(n13581), .ZN(
        n8874) );
  MUX2_X1 U11162 ( .A(n10814), .B(n10811), .S(n9716), .Z(n8899) );
  XNOR2_X1 U11163 ( .A(n8900), .B(n8899), .ZN(n11981) );
  NAND2_X1 U11164 ( .A1(n11981), .A2(n8786), .ZN(n8884) );
  NAND2_X1 U11165 ( .A1(n8881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8882) );
  XNOR2_X1 U11166 ( .A(n8882), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U11167 ( .A1(n8907), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8906), 
        .B2(n13550), .ZN(n8883) );
  NAND2_X1 U11168 ( .A1(n13925), .A2(n9165), .ZN(n8894) );
  INV_X1 U11169 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n15444) );
  INV_X1 U11170 ( .A(n8910), .ZN(n8912) );
  NAND2_X1 U11171 ( .A1(n8885), .A2(n15444), .ZN(n8886) );
  NAND2_X1 U11172 ( .A1(n8912), .A2(n8886), .ZN(n13812) );
  OR2_X1 U11173 ( .A1(n13812), .A2(n9114), .ZN(n8892) );
  INV_X1 U11174 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11175 ( .A1(n9136), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11176 ( .A1(n8510), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8887) );
  OAI211_X1 U11177 ( .C1(n8962), .C2(n8889), .A(n8888), .B(n8887), .ZN(n8890)
         );
  INV_X1 U11178 ( .A(n8890), .ZN(n8891) );
  NAND2_X1 U11179 ( .A1(n8892), .A2(n8891), .ZN(n13583) );
  NAND2_X1 U11180 ( .A1(n13583), .A2(n9196), .ZN(n8893) );
  NAND2_X1 U11181 ( .A1(n8894), .A2(n8893), .ZN(n8897) );
  INV_X1 U11182 ( .A(n13583), .ZN(n13611) );
  NAND2_X1 U11183 ( .A1(n13925), .A2(n9196), .ZN(n8895) );
  OAI21_X1 U11184 ( .B1(n13611), .B2(n8614), .A(n8895), .ZN(n8896) );
  INV_X1 U11185 ( .A(n8897), .ZN(n8898) );
  INV_X1 U11186 ( .A(n8928), .ZN(n8901) );
  NAND2_X1 U11187 ( .A1(n8901), .A2(SI_18_), .ZN(n8902) );
  MUX2_X1 U11188 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9716), .Z(n8903) );
  NAND2_X1 U11189 ( .A1(n8903), .A2(SI_19_), .ZN(n8932) );
  INV_X1 U11190 ( .A(n8903), .ZN(n8904) );
  NAND2_X1 U11191 ( .A1(n8904), .A2(n9991), .ZN(n8930) );
  NAND2_X1 U11192 ( .A1(n8932), .A2(n8930), .ZN(n8905) );
  NAND2_X1 U11193 ( .A1(n11961), .A2(n8786), .ZN(n8909) );
  AOI22_X1 U11194 ( .A1(n8907), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8906), 
        .B2(n10304), .ZN(n8908) );
  NAND2_X1 U11195 ( .A1(n13920), .A2(n9196), .ZN(n8921) );
  INV_X1 U11196 ( .A(n8937), .ZN(n8914) );
  INV_X1 U11197 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11198 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  AND2_X1 U11199 ( .A1(n8914), .A2(n8913), .ZN(n13800) );
  NAND2_X1 U11200 ( .A1(n13800), .A2(n9160), .ZN(n8919) );
  INV_X1 U11201 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15348) );
  NAND2_X1 U11202 ( .A1(n9136), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11203 ( .A1(n8510), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8915) );
  OAI211_X1 U11204 ( .C1(n8962), .C2(n15348), .A(n8916), .B(n8915), .ZN(n8917)
         );
  INV_X1 U11205 ( .A(n8917), .ZN(n8918) );
  NAND2_X1 U11206 ( .A1(n8919), .A2(n8918), .ZN(n13475) );
  NAND2_X1 U11207 ( .A1(n13475), .A2(n9165), .ZN(n8920) );
  NAND2_X1 U11208 ( .A1(n8921), .A2(n8920), .ZN(n8924) );
  AOI22_X1 U11209 ( .A1(n13920), .A2(n9165), .B1(n8922), .B2(n13475), .ZN(
        n8923) );
  NAND2_X1 U11210 ( .A1(n8929), .A2(SI_18_), .ZN(n8927) );
  NOR2_X1 U11211 ( .A1(n8929), .A2(SI_18_), .ZN(n8933) );
  INV_X1 U11212 ( .A(n8930), .ZN(n8931) );
  AOI21_X1 U11213 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8934) );
  INV_X1 U11214 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n15429) );
  MUX2_X1 U11215 ( .A(n6945), .B(n15429), .S(n9716), .Z(n8950) );
  XNOR2_X1 U11216 ( .A(n8952), .B(n8950), .ZN(n11970) );
  NAND2_X1 U11217 ( .A1(n11970), .A2(n8786), .ZN(n8936) );
  OR2_X1 U11218 ( .A1(n9152), .A2(n15429), .ZN(n8935) );
  NAND2_X1 U11219 ( .A1(n13915), .A2(n9165), .ZN(n8945) );
  NOR2_X1 U11220 ( .A1(n8937), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8938) );
  OR2_X1 U11221 ( .A1(n8958), .A2(n8938), .ZN(n13784) );
  INV_X1 U11222 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11223 ( .A1(n9136), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11224 ( .A1(n8510), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8939) );
  OAI211_X1 U11225 ( .C1(n8962), .C2(n8941), .A(n8940), .B(n8939), .ZN(n8942)
         );
  INV_X1 U11226 ( .A(n8942), .ZN(n8943) );
  OAI21_X1 U11227 ( .B1(n13784), .B2(n9114), .A(n8943), .ZN(n13588) );
  NAND2_X1 U11228 ( .A1(n13588), .A2(n9196), .ZN(n8944) );
  NAND2_X1 U11229 ( .A1(n8945), .A2(n8944), .ZN(n8948) );
  INV_X1 U11230 ( .A(n13588), .ZN(n13616) );
  NAND2_X1 U11231 ( .A1(n13915), .A2(n9196), .ZN(n8946) );
  OAI21_X1 U11232 ( .B1(n13616), .B2(n8614), .A(n8946), .ZN(n8947) );
  INV_X1 U11233 ( .A(n8950), .ZN(n8951) );
  INV_X1 U11234 ( .A(SI_20_), .ZN(n10185) );
  MUX2_X1 U11235 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9716), .Z(n8980) );
  XNOR2_X1 U11236 ( .A(n8980), .B(SI_21_), .ZN(n8977) );
  XNOR2_X1 U11237 ( .A(n8979), .B(n8977), .ZN(n12028) );
  NAND2_X1 U11238 ( .A1(n12028), .A2(n8786), .ZN(n8957) );
  OR2_X1 U11239 ( .A1(n9152), .A2(n11036), .ZN(n8956) );
  NAND2_X1 U11240 ( .A1(n13763), .A2(n9196), .ZN(n8967) );
  OR2_X1 U11241 ( .A1(n8958), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8959) );
  AND2_X1 U11242 ( .A1(n8959), .A2(n8984), .ZN(n13762) );
  NAND2_X1 U11243 ( .A1(n13762), .A2(n9160), .ZN(n8965) );
  INV_X1 U11244 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U11245 ( .A1(n9136), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U11246 ( .A1(n8510), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8960) );
  OAI211_X1 U11247 ( .C1(n8962), .C2(n13972), .A(n8961), .B(n8960), .ZN(n8963)
         );
  INV_X1 U11248 ( .A(n8963), .ZN(n8964) );
  NAND2_X1 U11249 ( .A1(n8965), .A2(n8964), .ZN(n13590) );
  NAND2_X1 U11250 ( .A1(n13590), .A2(n9165), .ZN(n8966) );
  NAND2_X1 U11251 ( .A1(n8967), .A2(n8966), .ZN(n8972) );
  NAND2_X1 U11252 ( .A1(n8971), .A2(n8972), .ZN(n8970) );
  INV_X1 U11253 ( .A(n13590), .ZN(n13618) );
  NAND2_X1 U11254 ( .A1(n13763), .A2(n9165), .ZN(n8968) );
  OAI21_X1 U11255 ( .B1(n13618), .B2(n9198), .A(n8968), .ZN(n8969) );
  NAND2_X1 U11256 ( .A1(n8970), .A2(n8969), .ZN(n8976) );
  INV_X1 U11257 ( .A(n8971), .ZN(n8974) );
  INV_X1 U11258 ( .A(n8972), .ZN(n8973) );
  NAND2_X1 U11259 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  INV_X1 U11260 ( .A(n8977), .ZN(n8978) );
  NAND2_X1 U11261 ( .A1(n8980), .A2(SI_21_), .ZN(n8981) );
  MUX2_X1 U11262 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9716), .Z(n9013) );
  XNOR2_X1 U11263 ( .A(n11951), .B(n9013), .ZN(n11574) );
  NAND2_X1 U11264 ( .A1(n11574), .A2(n8786), .ZN(n8983) );
  OR2_X1 U11265 ( .A1(n9152), .A2(n15351), .ZN(n8982) );
  NAND2_X1 U11266 ( .A1(n13753), .A2(n9165), .ZN(n8990) );
  NAND2_X1 U11267 ( .A1(n9155), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11268 ( .A1(n8510), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8987) );
  INV_X1 U11269 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n15379) );
  AOI21_X1 U11270 ( .B1(n15379), .B2(n8984), .A(n8999), .ZN(n13754) );
  NAND2_X1 U11271 ( .A1(n9160), .A2(n13754), .ZN(n8986) );
  NAND2_X1 U11272 ( .A1(n9136), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8985) );
  NAND4_X1 U11273 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n13592) );
  NAND2_X1 U11274 ( .A1(n8922), .A2(n13592), .ZN(n8989) );
  AOI22_X1 U11275 ( .A1(n13753), .A2(n8922), .B1(n13592), .B2(n9165), .ZN(
        n8991) );
  NAND2_X1 U11276 ( .A1(n8992), .A2(n9013), .ZN(n8994) );
  NAND2_X1 U11277 ( .A1(n9012), .A2(SI_22_), .ZN(n8993) );
  NAND2_X1 U11278 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  MUX2_X1 U11279 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9716), .Z(n9016) );
  XNOR2_X1 U11280 ( .A(n9016), .B(SI_23_), .ZN(n8995) );
  NAND2_X1 U11281 ( .A1(n11941), .A2(n8786), .ZN(n8998) );
  OR2_X1 U11282 ( .A1(n9152), .A2(n11666), .ZN(n8997) );
  NAND2_X1 U11283 ( .A1(n13964), .A2(n9196), .ZN(n9005) );
  NAND2_X1 U11284 ( .A1(n8999), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9022) );
  OAI21_X1 U11285 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8999), .A(n9022), .ZN(
        n13733) );
  OR2_X1 U11286 ( .A1(n9114), .A2(n13733), .ZN(n9003) );
  NAND2_X1 U11287 ( .A1(n9155), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11288 ( .A1(n8510), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U11289 ( .A1(n9136), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9000) );
  NAND4_X1 U11290 ( .A1(n9003), .A2(n9002), .A3(n9001), .A4(n9000), .ZN(n13621) );
  NAND2_X1 U11291 ( .A1(n9165), .A2(n13621), .ZN(n9004) );
  AOI22_X1 U11292 ( .A1(n13964), .A2(n9165), .B1(n8922), .B2(n13621), .ZN(
        n9006) );
  INV_X1 U11293 ( .A(n9006), .ZN(n9007) );
  INV_X1 U11294 ( .A(n9016), .ZN(n9009) );
  INV_X1 U11295 ( .A(SI_23_), .ZN(n10609) );
  NAND2_X1 U11296 ( .A1(n9009), .A2(n10609), .ZN(n9017) );
  OAI21_X1 U11297 ( .B1(SI_22_), .B2(n9013), .A(n9017), .ZN(n9010) );
  INV_X1 U11298 ( .A(n9010), .ZN(n9011) );
  INV_X1 U11299 ( .A(n9013), .ZN(n9015) );
  INV_X1 U11300 ( .A(SI_22_), .ZN(n9014) );
  NOR2_X1 U11301 ( .A1(n9015), .A2(n9014), .ZN(n9018) );
  AOI22_X1 U11302 ( .A1(n9018), .A2(n9017), .B1(n9016), .B2(SI_23_), .ZN(n9019) );
  MUX2_X1 U11303 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9040), .Z(n9035) );
  XNOR2_X1 U11304 ( .A(n9034), .B(n9035), .ZN(n11931) );
  NAND2_X1 U11305 ( .A1(n11931), .A2(n8786), .ZN(n9021) );
  OR2_X1 U11306 ( .A1(n9152), .A2(n11745), .ZN(n9020) );
  NAND2_X1 U11307 ( .A1(n13888), .A2(n9165), .ZN(n9028) );
  NAND2_X1 U11308 ( .A1(n8511), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U11309 ( .A1(n8510), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9025) );
  INV_X1 U11310 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13431) );
  AOI21_X1 U11311 ( .B1(n13431), .B2(n9022), .A(n9046), .ZN(n13721) );
  NAND2_X1 U11312 ( .A1(n9160), .A2(n13721), .ZN(n9024) );
  NAND2_X1 U11313 ( .A1(n9136), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9023) );
  NAND4_X1 U11314 ( .A1(n9026), .A2(n9025), .A3(n9024), .A4(n9023), .ZN(n13625) );
  NAND2_X1 U11315 ( .A1(n9172), .A2(n13625), .ZN(n9027) );
  NAND2_X1 U11316 ( .A1(n13888), .A2(n9196), .ZN(n9030) );
  NAND2_X1 U11317 ( .A1(n9165), .A2(n13625), .ZN(n9029) );
  NAND2_X1 U11318 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  NAND2_X1 U11319 ( .A1(n6530), .A2(n6562), .ZN(n9033) );
  INV_X1 U11320 ( .A(n9034), .ZN(n9036) );
  NAND2_X1 U11321 ( .A1(n9036), .A2(n9035), .ZN(n9039) );
  NAND2_X1 U11322 ( .A1(n9037), .A2(SI_24_), .ZN(n9038) );
  NAND2_X1 U11323 ( .A1(n9039), .A2(n9038), .ZN(n9057) );
  MUX2_X1 U11324 ( .A(n12053), .B(n15327), .S(n9040), .Z(n9041) );
  INV_X1 U11325 ( .A(SI_25_), .ZN(n11033) );
  NAND2_X1 U11326 ( .A1(n9041), .A2(n11033), .ZN(n9055) );
  INV_X1 U11327 ( .A(n9041), .ZN(n9042) );
  NAND2_X1 U11328 ( .A1(n9042), .A2(SI_25_), .ZN(n9043) );
  NAND2_X1 U11329 ( .A1(n9055), .A2(n9043), .ZN(n9056) );
  XNOR2_X1 U11330 ( .A(n9057), .B(n9056), .ZN(n12052) );
  NAND2_X1 U11331 ( .A1(n12052), .A2(n8786), .ZN(n9045) );
  OR2_X1 U11332 ( .A1(n9152), .A2(n15327), .ZN(n9044) );
  NAND2_X1 U11333 ( .A1(n13705), .A2(n9196), .ZN(n9052) );
  NAND2_X1 U11334 ( .A1(n9046), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9061) );
  OAI21_X1 U11335 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n9046), .A(n9061), .ZN(
        n13400) );
  OR2_X1 U11336 ( .A1(n9114), .A2(n13400), .ZN(n9050) );
  NAND2_X1 U11337 ( .A1(n9155), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11338 ( .A1(n8510), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11339 ( .A1(n9136), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9047) );
  NAND4_X1 U11340 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n13598) );
  NAND2_X1 U11341 ( .A1(n9165), .A2(n13598), .ZN(n9051) );
  NAND2_X1 U11342 ( .A1(n9052), .A2(n9051), .ZN(n9054) );
  AOI22_X1 U11343 ( .A1(n13705), .A2(n9165), .B1(n9172), .B2(n13598), .ZN(
        n9053) );
  MUX2_X1 U11344 ( .A(n14708), .B(n14000), .S(n9716), .Z(n9074) );
  XNOR2_X1 U11345 ( .A(n9074), .B(SI_26_), .ZN(n9058) );
  XNOR2_X1 U11346 ( .A(n9075), .B(n9058), .ZN(n13998) );
  NAND2_X1 U11347 ( .A1(n13998), .A2(n8786), .ZN(n9060) );
  OR2_X1 U11348 ( .A1(n9152), .A2(n14000), .ZN(n9059) );
  NAND2_X1 U11349 ( .A1(n13955), .A2(n8544), .ZN(n9068) );
  INV_X1 U11350 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U11351 ( .A1(n9062), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9112) );
  OAI21_X1 U11352 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n9062), .A(n9112), .ZN(
        n13690) );
  OR2_X1 U11353 ( .A1(n9114), .A2(n13690), .ZN(n9066) );
  NAND2_X1 U11354 ( .A1(n8510), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11355 ( .A1(n9136), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11356 ( .A1(n9155), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9063) );
  NAND4_X1 U11357 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n13630) );
  NAND2_X1 U11358 ( .A1(n9172), .A2(n13630), .ZN(n9067) );
  NAND2_X1 U11359 ( .A1(n9068), .A2(n9067), .ZN(n9070) );
  AOI22_X1 U11360 ( .A1(n13955), .A2(n8922), .B1(n13630), .B2(n9165), .ZN(
        n9069) );
  NOR2_X1 U11361 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  INV_X1 U11362 ( .A(SI_26_), .ZN(n11302) );
  MUX2_X1 U11363 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9716), .Z(n9106) );
  NOR2_X1 U11364 ( .A1(n9106), .A2(SI_27_), .ZN(n9076) );
  NAND2_X1 U11365 ( .A1(n9106), .A2(SI_27_), .ZN(n9077) );
  NAND2_X1 U11366 ( .A1(n9078), .A2(n9077), .ZN(n9148) );
  MUX2_X1 U11367 ( .A(n14698), .B(n9151), .S(n9716), .Z(n9079) );
  INV_X1 U11368 ( .A(SI_28_), .ZN(n11889) );
  NAND2_X1 U11369 ( .A1(n9079), .A2(n11889), .ZN(n9082) );
  INV_X1 U11370 ( .A(n9079), .ZN(n9080) );
  NAND2_X1 U11371 ( .A1(n9080), .A2(SI_28_), .ZN(n9081) );
  NAND2_X1 U11372 ( .A1(n9082), .A2(n9081), .ZN(n9147) );
  INV_X1 U11373 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13989) );
  MUX2_X1 U11374 ( .A(n14695), .B(n13989), .S(n9716), .Z(n9083) );
  XNOR2_X1 U11375 ( .A(n9083), .B(SI_29_), .ZN(n9131) );
  INV_X1 U11376 ( .A(SI_29_), .ZN(n12419) );
  NAND2_X1 U11377 ( .A1(n9083), .A2(n12419), .ZN(n9084) );
  MUX2_X1 U11378 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9716), .Z(n9085) );
  NAND2_X1 U11379 ( .A1(n9085), .A2(SI_30_), .ZN(n9123) );
  OAI21_X1 U11380 ( .B1(SI_30_), .B2(n9085), .A(n9123), .ZN(n9086) );
  NAND2_X1 U11381 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  INV_X1 U11382 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13985) );
  OR2_X1 U11383 ( .A1(n9152), .A2(n13985), .ZN(n9090) );
  INV_X1 U11384 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U11385 ( .A1(n8510), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11386 ( .A1(n8511), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9092) );
  OAI211_X1 U11387 ( .C1(n9094), .C2(n15445), .A(n9093), .B(n9092), .ZN(n13472) );
  NAND2_X1 U11388 ( .A1(n9165), .A2(n13472), .ZN(n9102) );
  INV_X1 U11389 ( .A(n9095), .ZN(n9096) );
  AND2_X1 U11390 ( .A1(n9097), .A2(n9096), .ZN(n9101) );
  NAND2_X1 U11391 ( .A1(n9136), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11392 ( .A1(n8510), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9099) );
  NAND2_X1 U11393 ( .A1(n9155), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9098) );
  AND3_X1 U11394 ( .A1(n9100), .A2(n9099), .A3(n9098), .ZN(n13638) );
  AOI21_X1 U11395 ( .B1(n9102), .B2(n9101), .A(n13638), .ZN(n9103) );
  AOI21_X1 U11396 ( .B1(n13565), .B2(n8922), .A(n9103), .ZN(n9176) );
  NAND2_X1 U11397 ( .A1(n13565), .A2(n9165), .ZN(n9105) );
  INV_X1 U11398 ( .A(n13638), .ZN(n13473) );
  NAND2_X1 U11399 ( .A1(n9172), .A2(n13473), .ZN(n9104) );
  NAND2_X1 U11400 ( .A1(n9105), .A2(n9104), .ZN(n9175) );
  NAND2_X1 U11401 ( .A1(n9176), .A2(n9175), .ZN(n9195) );
  INV_X1 U11402 ( .A(n9106), .ZN(n9107) );
  XNOR2_X1 U11403 ( .A(n9107), .B(SI_27_), .ZN(n9108) );
  XNOR2_X1 U11404 ( .A(n9109), .B(n9108), .ZN(n13995) );
  NAND2_X1 U11405 ( .A1(n13995), .A2(n8786), .ZN(n9111) );
  OR2_X1 U11406 ( .A1(n9152), .A2(n13997), .ZN(n9110) );
  INV_X1 U11407 ( .A(n9112), .ZN(n9113) );
  INV_X1 U11408 ( .A(n9135), .ZN(n9157) );
  OAI21_X1 U11409 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n9113), .A(n9157), .ZN(
        n13673) );
  OR2_X1 U11410 ( .A1(n9114), .A2(n13673), .ZN(n9118) );
  NAND2_X1 U11411 ( .A1(n8511), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11412 ( .A1(n8510), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U11413 ( .A1(n9136), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9115) );
  NAND4_X1 U11414 ( .A1(n9118), .A2(n9117), .A3(n9116), .A4(n9115), .ZN(n13632) );
  AND2_X1 U11415 ( .A1(n9165), .A2(n13632), .ZN(n9119) );
  AOI21_X1 U11416 ( .B1(n13871), .B2(n8922), .A(n9119), .ZN(n9183) );
  NAND2_X1 U11417 ( .A1(n13871), .A2(n8544), .ZN(n9121) );
  NAND2_X1 U11418 ( .A1(n9172), .A2(n13632), .ZN(n9120) );
  NAND2_X1 U11419 ( .A1(n9121), .A2(n9120), .ZN(n9184) );
  NAND2_X1 U11420 ( .A1(n9183), .A2(n9184), .ZN(n9122) );
  AND2_X1 U11421 ( .A1(n9195), .A2(n9122), .ZN(n9170) );
  MUX2_X1 U11422 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9716), .Z(n9125) );
  XNOR2_X1 U11423 ( .A(n9125), .B(SI_31_), .ZN(n9126) );
  NAND2_X1 U11424 ( .A1(n11892), .A2(n8786), .ZN(n9130) );
  OR2_X1 U11425 ( .A1(n9152), .A2(n9128), .ZN(n9129) );
  XNOR2_X1 U11426 ( .A(n9171), .B(n13472), .ZN(n9228) );
  NAND2_X1 U11427 ( .A1(n13987), .A2(n8786), .ZN(n9134) );
  OR2_X1 U11428 ( .A1(n9152), .A2(n13989), .ZN(n9133) );
  NAND2_X1 U11429 ( .A1(n9155), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U11430 ( .A1(n8510), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U11431 ( .A1(n9160), .A2(n13642), .ZN(n9138) );
  NAND2_X1 U11432 ( .A1(n9136), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9137) );
  NAND4_X1 U11433 ( .A1(n9140), .A2(n9139), .A3(n9138), .A4(n9137), .ZN(n13474) );
  NAND2_X1 U11434 ( .A1(n9165), .A2(n13474), .ZN(n9142) );
  NAND2_X1 U11435 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  AOI21_X1 U11436 ( .B1(n13864), .B2(n8922), .A(n9143), .ZN(n9178) );
  NAND2_X1 U11437 ( .A1(n13864), .A2(n9165), .ZN(n9145) );
  NAND2_X1 U11438 ( .A1(n9172), .A2(n13474), .ZN(n9144) );
  NAND2_X1 U11439 ( .A1(n9145), .A2(n9144), .ZN(n9177) );
  NAND2_X1 U11440 ( .A1(n9178), .A2(n9177), .ZN(n9146) );
  AND2_X1 U11441 ( .A1(n9228), .A2(n9146), .ZN(n9188) );
  NAND2_X1 U11442 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  NAND2_X1 U11443 ( .A1(n9150), .A2(n9149), .ZN(n13990) );
  NAND2_X1 U11444 ( .A1(n13990), .A2(n8786), .ZN(n9154) );
  OR2_X1 U11445 ( .A1(n9152), .A2(n9151), .ZN(n9153) );
  NAND2_X1 U11446 ( .A1(n9155), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U11447 ( .A1(n8510), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9163) );
  INV_X1 U11448 ( .A(n13642), .ZN(n9159) );
  INV_X1 U11449 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11450 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  NAND2_X1 U11451 ( .A1(n9160), .A2(n13653), .ZN(n9162) );
  NAND2_X1 U11452 ( .A1(n9136), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9161) );
  NAND4_X1 U11453 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), .ZN(n13635) );
  AND2_X1 U11454 ( .A1(n9165), .A2(n13635), .ZN(n9166) );
  AOI21_X1 U11455 ( .B1(n13660), .B2(n8922), .A(n9166), .ZN(n9190) );
  NAND2_X1 U11456 ( .A1(n13660), .A2(n9165), .ZN(n9168) );
  NAND2_X1 U11457 ( .A1(n8922), .A2(n13635), .ZN(n9167) );
  NAND2_X1 U11458 ( .A1(n9168), .A2(n9167), .ZN(n9189) );
  NAND2_X1 U11459 ( .A1(n9190), .A2(n9189), .ZN(n9169) );
  MUX2_X1 U11460 ( .A(n13472), .B(n8614), .S(n9171), .Z(n9174) );
  NAND2_X1 U11461 ( .A1(n9172), .A2(n13472), .ZN(n9173) );
  AND2_X1 U11462 ( .A1(n9174), .A2(n9173), .ZN(n9194) );
  INV_X1 U11463 ( .A(n9175), .ZN(n9182) );
  INV_X1 U11464 ( .A(n9176), .ZN(n9181) );
  INV_X1 U11465 ( .A(n9177), .ZN(n9180) );
  INV_X1 U11466 ( .A(n9178), .ZN(n9179) );
  AOI22_X1 U11467 ( .A1(n9182), .A2(n9181), .B1(n9180), .B2(n9179), .ZN(n9193)
         );
  INV_X1 U11468 ( .A(n9183), .ZN(n9186) );
  INV_X1 U11469 ( .A(n9184), .ZN(n9185) );
  NAND3_X1 U11470 ( .A1(n9187), .A2(n9186), .A3(n9185), .ZN(n9192) );
  INV_X1 U11471 ( .A(n9188), .ZN(n9191) );
  NAND2_X1 U11472 ( .A1(n9171), .A2(n9196), .ZN(n9197) );
  NAND3_X1 U11473 ( .A1(n9197), .A2(n8614), .A3(n13472), .ZN(n9200) );
  INV_X1 U11474 ( .A(n13472), .ZN(n13571) );
  NAND3_X1 U11475 ( .A1(n9171), .A2(n13571), .A3(n9198), .ZN(n9199) );
  OAI21_X1 U11476 ( .B1(n11035), .B2(n10304), .A(n8471), .ZN(n9205) );
  AOI21_X1 U11477 ( .B1(n10305), .B2(n8482), .A(n9205), .ZN(n9206) );
  XNOR2_X1 U11478 ( .A(n13565), .B(n13638), .ZN(n9226) );
  NAND2_X1 U11479 ( .A1(n13660), .A2(n13635), .ZN(n13602) );
  OR2_X1 U11480 ( .A1(n13660), .A2(n13635), .ZN(n9207) );
  NAND2_X1 U11481 ( .A1(n13602), .A2(n9207), .ZN(n13647) );
  INV_X1 U11482 ( .A(n13598), .ZN(n13629) );
  XNOR2_X1 U11483 ( .A(n13705), .B(n13629), .ZN(n13701) );
  XNOR2_X1 U11484 ( .A(n13888), .B(n13625), .ZN(n13712) );
  XNOR2_X1 U11485 ( .A(n13763), .B(n13618), .ZN(n13767) );
  XNOR2_X1 U11486 ( .A(n13915), .B(n13616), .ZN(n13777) );
  XNOR2_X1 U11487 ( .A(n13925), .B(n13611), .ZN(n13809) );
  OR2_X1 U11488 ( .A1(n13920), .A2(n13475), .ZN(n13586) );
  NAND2_X1 U11489 ( .A1(n13920), .A2(n13475), .ZN(n13585) );
  INV_X1 U11490 ( .A(n13581), .ZN(n13610) );
  XNOR2_X1 U11491 ( .A(n13930), .B(n13610), .ZN(n13834) );
  XNOR2_X1 U11492 ( .A(n13607), .B(n13606), .ZN(n11866) );
  INV_X1 U11493 ( .A(n13476), .ZN(n11854) );
  XNOR2_X1 U11494 ( .A(n11863), .B(n11854), .ZN(n11688) );
  OR2_X1 U11495 ( .A1(n14887), .A2(n13477), .ZN(n11684) );
  NAND2_X1 U11496 ( .A1(n14887), .A2(n13477), .ZN(n11686) );
  NAND2_X1 U11497 ( .A1(n11684), .A2(n11686), .ZN(n11680) );
  INV_X1 U11498 ( .A(n13479), .ZN(n11350) );
  OR2_X1 U11499 ( .A1(n13847), .A2(n11350), .ZN(n11347) );
  NAND2_X1 U11500 ( .A1(n13847), .A2(n11350), .ZN(n9208) );
  NAND2_X1 U11501 ( .A1(n11347), .A2(n9208), .ZN(n11346) );
  NAND2_X1 U11502 ( .A1(n11010), .A2(n13481), .ZN(n10927) );
  OR2_X1 U11503 ( .A1(n11010), .A2(n13481), .ZN(n9209) );
  NAND2_X1 U11504 ( .A1(n10927), .A2(n9209), .ZN(n10924) );
  INV_X1 U11505 ( .A(n13484), .ZN(n10354) );
  XNOR2_X1 U11506 ( .A(n15178), .B(n10354), .ZN(n10347) );
  XNOR2_X1 U11507 ( .A(n10334), .B(n13485), .ZN(n10331) );
  INV_X1 U11508 ( .A(n13488), .ZN(n9944) );
  XNOR2_X1 U11509 ( .A(n9210), .B(n10053), .ZN(n9840) );
  NAND2_X1 U11510 ( .A1(n13491), .A2(n10541), .ZN(n9661) );
  OR2_X1 U11511 ( .A1(n13491), .A2(n10541), .ZN(n9212) );
  NAND2_X1 U11512 ( .A1(n9661), .A2(n9212), .ZN(n10545) );
  NAND4_X1 U11513 ( .A1(n9666), .A2(n9840), .A3(n10545), .A4(n9668), .ZN(n9213) );
  NOR2_X1 U11514 ( .A1(n9843), .A2(n9213), .ZN(n9214) );
  XNOR2_X1 U11515 ( .A(n10319), .B(n13486), .ZN(n10099) );
  XNOR2_X1 U11516 ( .A(n10644), .B(n13487), .ZN(n10025) );
  NAND4_X1 U11517 ( .A1(n10331), .A2(n9214), .A3(n10099), .A4(n10025), .ZN(
        n9215) );
  NOR2_X1 U11518 ( .A1(n10347), .A2(n9215), .ZN(n9216) );
  XNOR2_X1 U11519 ( .A(n10723), .B(n13482), .ZN(n10548) );
  XNOR2_X1 U11520 ( .A(n10552), .B(n13483), .ZN(n10357) );
  NAND4_X1 U11521 ( .A1(n10924), .A2(n9216), .A3(n10548), .A4(n10357), .ZN(
        n9217) );
  NOR2_X1 U11522 ( .A1(n11346), .A2(n9217), .ZN(n9218) );
  XNOR2_X1 U11523 ( .A(n11678), .B(n13478), .ZN(n11358) );
  XNOR2_X1 U11524 ( .A(n11412), .B(n13480), .ZN(n10929) );
  NAND4_X1 U11525 ( .A1(n11680), .A2(n9218), .A3(n11358), .A4(n10929), .ZN(
        n9219) );
  OR4_X1 U11526 ( .A1(n13834), .A2(n11866), .A3(n11688), .A4(n9219), .ZN(n9220) );
  OR4_X1 U11527 ( .A1(n13777), .A2(n13809), .A3(n13793), .A4(n9220), .ZN(n9221) );
  NOR2_X1 U11528 ( .A1(n13767), .A2(n9221), .ZN(n9222) );
  XNOR2_X1 U11529 ( .A(n13753), .B(n13592), .ZN(n13748) );
  OR2_X1 U11530 ( .A1(n13964), .A2(n13621), .ZN(n13594) );
  NAND2_X1 U11531 ( .A1(n13964), .A2(n13621), .ZN(n13595) );
  NAND2_X1 U11532 ( .A1(n13594), .A2(n13595), .ZN(n13737) );
  NAND4_X1 U11533 ( .A1(n13712), .A2(n9222), .A3(n13748), .A4(n13737), .ZN(
        n9223) );
  NOR2_X1 U11534 ( .A1(n13701), .A2(n9223), .ZN(n9224) );
  XNOR2_X1 U11535 ( .A(n13871), .B(n13632), .ZN(n13678) );
  XNOR2_X1 U11536 ( .A(n13955), .B(n13630), .ZN(n13685) );
  NAND4_X1 U11537 ( .A1(n13647), .A2(n9224), .A3(n13678), .A4(n13685), .ZN(
        n9225) );
  NOR2_X1 U11538 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  XNOR2_X1 U11539 ( .A(n13864), .B(n13474), .ZN(n13636) );
  NAND3_X1 U11540 ( .A1(n9228), .A2(n9227), .A3(n13636), .ZN(n9229) );
  XNOR2_X1 U11541 ( .A(n9229), .B(n10304), .ZN(n9230) );
  OAI211_X1 U11542 ( .C1(n9252), .C2(n9231), .A(n9230), .B(n11035), .ZN(n9254)
         );
  MUX2_X1 U11543 ( .A(n8466), .B(n9232), .S(n10962), .Z(n9233) );
  OR2_X1 U11544 ( .A1(n9234), .A2(P2_U3088), .ZN(n11664) );
  NAND2_X1 U11545 ( .A1(n9243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9237) );
  INV_X1 U11546 ( .A(n14002), .ZN(n9246) );
  NOR2_X1 U11547 ( .A1(n6578), .A2(n13982), .ZN(n9238) );
  MUX2_X1 U11548 ( .A(n13982), .B(n9238), .S(P2_IR_REG_24__SCAN_IN), .Z(n9239)
         );
  INV_X1 U11549 ( .A(n9239), .ZN(n9240) );
  NAND2_X1 U11550 ( .A1(n9240), .A2(n9241), .ZN(n11744) );
  NAND2_X1 U11551 ( .A1(n9241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9242) );
  MUX2_X1 U11552 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9242), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9244) );
  NAND2_X1 U11553 ( .A1(n9244), .A2(n9243), .ZN(n11807) );
  NOR2_X1 U11554 ( .A1(n11744), .A2(n11807), .ZN(n9245) );
  NAND2_X1 U11555 ( .A1(n9246), .A2(n9245), .ZN(n9342) );
  AND2_X1 U11556 ( .A1(n9234), .A2(n9342), .ZN(n9634) );
  INV_X1 U11557 ( .A(n13996), .ZN(n9425) );
  INV_X1 U11558 ( .A(n9247), .ZN(n9248) );
  NAND4_X1 U11559 ( .A1(n15176), .A2(n9425), .A3(n9621), .A4(n13464), .ZN(
        n9249) );
  OAI211_X1 U11560 ( .C1(n9232), .C2(n11664), .A(n9249), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9250) );
  NAND3_X1 U11561 ( .A1(n7664), .A2(n9254), .A3(n9253), .ZN(n9256) );
  INV_X1 U11562 ( .A(P2_B_REG_SCAN_IN), .ZN(n13568) );
  NAND2_X1 U11563 ( .A1(n11664), .A2(n13568), .ZN(n9255) );
  AND2_X1 U11564 ( .A1(n9256), .A2(n9255), .ZN(P2_U3328) );
  NOR2_X1 U11565 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9258) );
  NOR2_X1 U11566 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9260) );
  NOR2_X1 U11567 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9259) );
  INV_X1 U11568 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9265) );
  OAI21_X1 U11569 ( .B1(n9361), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9266) );
  XNOR2_X1 U11570 ( .A(n9266), .B(P1_IR_REG_23__SCAN_IN), .ZN(n9372) );
  NOR2_X1 U11571 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9268) );
  NOR2_X1 U11572 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9267) );
  NAND3_X1 U11573 ( .A1(n9269), .A2(n9268), .A3(n9267), .ZN(n9369) );
  INV_X1 U11574 ( .A(n9369), .ZN(n9270) );
  NAND2_X1 U11575 ( .A1(n9274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9271) );
  MUX2_X1 U11576 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9271), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9272) );
  NAND2_X1 U11577 ( .A1(n9272), .A2(n9276), .ZN(n11806) );
  NAND2_X1 U11578 ( .A1(n9364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9273) );
  MUX2_X1 U11579 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9273), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9275) );
  NAND2_X1 U11580 ( .A1(n9275), .A2(n9274), .ZN(n11746) );
  NOR2_X1 U11581 ( .A1(n11806), .A2(n11746), .ZN(n9278) );
  NAND2_X1 U11582 ( .A1(n9276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9277) );
  OR2_X2 U11583 ( .A1(n9380), .A2(n9736), .ZN(n14156) );
  INV_X1 U11584 ( .A(n14156), .ZN(P1_U4016) );
  NOR2_X1 U11585 ( .A1(n9716), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13992) );
  INV_X2 U11586 ( .A(n13992), .ZN(n13999) );
  NAND2_X1 U11587 ( .A1(n9716), .A2(P2_U3088), .ZN(n13994) );
  INV_X1 U11588 ( .A(n9959), .ZN(n9291) );
  OAI222_X1 U11589 ( .A1(n13999), .A2(n9279), .B1(n13994), .B2(n9291), .C1(
        P2_U3088), .C2(n13496), .ZN(P2_U3325) );
  NAND2_X1 U11590 ( .A1(n9716), .A2(P1_U3086), .ZN(n14709) );
  INV_X1 U11591 ( .A(n14709), .ZN(n14690) );
  INV_X1 U11592 ( .A(n14690), .ZN(n14701) );
  AND2_X1 U11593 ( .A1(n8598), .A2(P1_U3086), .ZN(n11661) );
  INV_X2 U11594 ( .A(n11661), .ZN(n14707) );
  INV_X1 U11595 ( .A(n9855), .ZN(n9312) );
  NAND2_X1 U11596 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9280) );
  MUX2_X1 U11597 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9280), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9283) );
  INV_X1 U11598 ( .A(n9281), .ZN(n9282) );
  NAND2_X1 U11599 ( .A1(n9283), .A2(n9282), .ZN(n14162) );
  OAI222_X1 U11600 ( .A1(n14701), .A2(n6848), .B1(n14707), .B2(n9312), .C1(
        n14162), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U11601 ( .A(n10111), .ZN(n9286) );
  NAND2_X1 U11602 ( .A1(n9284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9285) );
  XNOR2_X1 U11603 ( .A(n9285), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14184) );
  INV_X1 U11604 ( .A(n14184), .ZN(n9497) );
  OAI222_X1 U11605 ( .A1(n14701), .A2(n10114), .B1(n14707), .B2(n9286), .C1(
        n9497), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U11606 ( .A1(n13999), .A2(n9287), .B1(n13994), .B2(n9286), .C1(
        P2_U3088), .C2(n6886), .ZN(P2_U3324) );
  NOR2_X1 U11607 ( .A1(n9281), .A2(n9306), .ZN(n9288) );
  MUX2_X1 U11608 ( .A(n9306), .B(n9288), .S(P1_IR_REG_2__SCAN_IN), .Z(n9290)
         );
  INV_X1 U11609 ( .A(n9284), .ZN(n9289) );
  NOR2_X1 U11610 ( .A1(n9290), .A2(n9289), .ZN(n14173) );
  INV_X1 U11611 ( .A(n14173), .ZN(n9292) );
  OAI222_X1 U11612 ( .A1(n9292), .A2(P1_U3086), .B1(n14707), .B2(n9291), .C1(
        n9962), .C2(n14701), .ZN(P1_U3353) );
  NAND2_X1 U11613 ( .A1(n9716), .A2(P3_U3151), .ZN(n12420) );
  NAND2_X1 U11614 ( .A1(n8598), .A2(P3_U3151), .ZN(n13303) );
  OAI222_X1 U11615 ( .A1(P3_U3151), .A2(n11393), .B1(n12420), .B2(n9294), .C1(
        n13303), .C2(n9293), .ZN(P3_U3285) );
  OAI222_X1 U11616 ( .A1(P3_U3151), .A2(n11172), .B1(n12420), .B2(n9296), .C1(
        n13303), .C2(n9295), .ZN(P3_U3286) );
  INV_X1 U11617 ( .A(n10227), .ZN(n9301) );
  INV_X1 U11618 ( .A(n9599), .ZN(n9401) );
  OAI222_X1 U11619 ( .A1(n13999), .A2(n9297), .B1(n13994), .B2(n9301), .C1(
        P2_U3088), .C2(n9401), .ZN(P2_U3323) );
  NAND2_X1 U11620 ( .A1(n9298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9299) );
  XNOR2_X1 U11621 ( .A(n9299), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10228) );
  INV_X1 U11622 ( .A(n10228), .ZN(n9302) );
  OAI222_X1 U11623 ( .A1(n9302), .A2(P1_U3086), .B1(n14707), .B2(n9301), .C1(
        n9300), .C2(n14701), .ZN(P1_U3351) );
  OAI222_X1 U11624 ( .A1(P3_U3151), .A2(n11394), .B1(n12420), .B2(n9304), .C1(
        n13303), .C2(n9303), .ZN(P3_U3284) );
  OR2_X1 U11625 ( .A1(n9305), .A2(n9306), .ZN(n9307) );
  XNOR2_X1 U11626 ( .A(n9307), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10233) );
  INV_X1 U11627 ( .A(n10233), .ZN(n9519) );
  INV_X1 U11628 ( .A(n10232), .ZN(n9310) );
  OAI222_X1 U11629 ( .A1(n9519), .A2(P1_U3086), .B1(n14707), .B2(n9310), .C1(
        n9308), .C2(n14701), .ZN(P1_U3350) );
  INV_X1 U11630 ( .A(n9443), .ZN(n9309) );
  OAI222_X1 U11631 ( .A1(n13999), .A2(n9311), .B1(n13994), .B2(n9310), .C1(
        P2_U3088), .C2(n9309), .ZN(P2_U3322) );
  INV_X1 U11632 ( .A(n13994), .ZN(n11663) );
  INV_X1 U11633 ( .A(n11663), .ZN(n14001) );
  OAI222_X1 U11634 ( .A1(n13999), .A2(n9313), .B1(n14001), .B2(n9312), .C1(
        P2_U3088), .C2(n9453), .ZN(P2_U3326) );
  INV_X1 U11635 ( .A(n12420), .ZN(n13301) );
  INV_X1 U11636 ( .A(n13301), .ZN(n11887) );
  OAI222_X1 U11637 ( .A1(P3_U3151), .A2(n11222), .B1(n11887), .B2(n9315), .C1(
        n13303), .C2(n9314), .ZN(P3_U3290) );
  INV_X1 U11638 ( .A(SI_4_), .ZN(n9317) );
  OAI222_X1 U11639 ( .A1(P3_U3151), .A2(n11258), .B1(n11887), .B2(n9317), .C1(
        n13303), .C2(n9316), .ZN(P3_U3291) );
  INV_X1 U11640 ( .A(SI_7_), .ZN(n9319) );
  OAI222_X1 U11641 ( .A1(P3_U3151), .A2(n11152), .B1(n11887), .B2(n9319), .C1(
        n13303), .C2(n9318), .ZN(P3_U3288) );
  INV_X1 U11642 ( .A(n9320), .ZN(n9321) );
  OAI222_X1 U11643 ( .A1(P3_U3151), .A2(n12739), .B1(n12420), .B2(n9322), .C1(
        n13303), .C2(n9321), .ZN(P3_U3283) );
  INV_X1 U11644 ( .A(n10270), .ZN(n9328) );
  INV_X1 U11645 ( .A(n9544), .ZN(n9323) );
  OAI222_X1 U11646 ( .A1(n13999), .A2(n9324), .B1(n13994), .B2(n9328), .C1(
        P2_U3088), .C2(n9323), .ZN(P2_U3321) );
  AND2_X1 U11647 ( .A1(n9305), .A2(n9325), .ZN(n10297) );
  OR2_X1 U11648 ( .A1(n10297), .A2(n9306), .ZN(n9326) );
  XNOR2_X1 U11649 ( .A(n9326), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14205) );
  INV_X1 U11650 ( .A(n14205), .ZN(n9327) );
  OAI222_X1 U11651 ( .A1(n14701), .A2(n9329), .B1(n14707), .B2(n9328), .C1(
        n9327), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U11652 ( .A(n13303), .ZN(n10606) );
  INV_X1 U11653 ( .A(n9330), .ZN(n9332) );
  OAI222_X1 U11654 ( .A1(n11891), .A2(n9332), .B1(n12420), .B2(n9331), .C1(
        P3_U3151), .C2(n11629), .ZN(P3_U3294) );
  INV_X1 U11655 ( .A(SI_8_), .ZN(n9333) );
  OAI222_X1 U11656 ( .A1(n11891), .A2(n9334), .B1(n11887), .B2(n9333), .C1(
        P3_U3151), .C2(n12720), .ZN(P3_U3287) );
  INV_X1 U11657 ( .A(n12705), .ZN(n11141) );
  INV_X1 U11658 ( .A(n9335), .ZN(n9337) );
  INV_X1 U11659 ( .A(SI_6_), .ZN(n9336) );
  OAI222_X1 U11660 ( .A1(P3_U3151), .A2(n11141), .B1(n11891), .B2(n9337), .C1(
        n9336), .C2(n11887), .ZN(P3_U3289) );
  INV_X1 U11661 ( .A(SI_3_), .ZN(n9339) );
  OAI222_X1 U11662 ( .A1(P3_U3151), .A2(n11135), .B1(n11887), .B2(n9339), .C1(
        n11891), .C2(n9338), .ZN(P3_U3292) );
  INV_X1 U11663 ( .A(SI_2_), .ZN(n9341) );
  OAI222_X1 U11664 ( .A1(P3_U3151), .A2(n11299), .B1(n11887), .B2(n9341), .C1(
        n11891), .C2(n9340), .ZN(P3_U3293) );
  INV_X1 U11665 ( .A(n9342), .ZN(n9343) );
  NAND2_X1 U11666 ( .A1(n9343), .A2(n9234), .ZN(n9395) );
  OR2_X2 U11667 ( .A1(n9395), .A2(P2_U3088), .ZN(n13490) );
  INV_X1 U11668 ( .A(n13490), .ZN(P2_U3947) );
  INV_X1 U11669 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U11670 ( .A1(n10297), .A2(n9344), .ZN(n9350) );
  NAND2_X1 U11671 ( .A1(n9350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9345) );
  XNOR2_X1 U11672 ( .A(n9345), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10477) );
  INV_X1 U11673 ( .A(n10477), .ZN(n9524) );
  INV_X1 U11674 ( .A(n10476), .ZN(n9348) );
  OAI222_X1 U11675 ( .A1(n9524), .A2(P1_U3086), .B1(n14707), .B2(n9348), .C1(
        n9346), .C2(n14709), .ZN(P1_U3348) );
  INV_X1 U11676 ( .A(n15124), .ZN(n9347) );
  OAI222_X1 U11677 ( .A1(n13999), .A2(n9349), .B1(n13994), .B2(n9348), .C1(
        P2_U3088), .C2(n9347), .ZN(P2_U3320) );
  NAND2_X1 U11678 ( .A1(n9570), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9384) );
  XNOR2_X1 U11679 ( .A(n9384), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10740) );
  INV_X1 U11680 ( .A(n10740), .ZN(n9352) );
  INV_X1 U11681 ( .A(n10739), .ZN(n9353) );
  OAI222_X1 U11682 ( .A1(n9352), .A2(P1_U3086), .B1(n14707), .B2(n9353), .C1(
        n9351), .C2(n14709), .ZN(P1_U3347) );
  INV_X1 U11683 ( .A(n9807), .ZN(n9542) );
  OAI222_X1 U11684 ( .A1(n13999), .A2(n9354), .B1(n13994), .B2(n9353), .C1(
        P2_U3088), .C2(n9542), .ZN(P2_U3319) );
  OR2_X1 U11685 ( .A1(n9356), .A2(n9355), .ZN(n9360) );
  NOR2_X1 U11686 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  NAND2_X1 U11687 ( .A1(n9755), .A2(n12072), .ZN(n12069) );
  INV_X1 U11688 ( .A(n9372), .ZN(n9720) );
  INV_X1 U11689 ( .A(n9367), .ZN(n9363) );
  NOR2_X1 U11690 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9366) );
  NAND2_X1 U11691 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NOR2_X1 U11692 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  AOI21_X1 U11693 ( .B1(n9871), .B2(n9720), .A(n12022), .ZN(n9489) );
  INV_X1 U11694 ( .A(n9489), .ZN(n9373) );
  NAND2_X1 U11695 ( .A1(n9372), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12256) );
  INV_X1 U11696 ( .A(n12256), .ZN(n12248) );
  OR2_X1 U11697 ( .A1(n10191), .A2(n12248), .ZN(n9490) );
  NOR2_X1 U11698 ( .A1(n14977), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U11699 ( .A1(P3_U3151), .A2(n12771), .B1(n12420), .B2(n9375), .C1(
        n13303), .C2(n9374), .ZN(P3_U3282) );
  NAND2_X1 U11700 ( .A1(n11806), .A2(P1_B_REG_SCAN_IN), .ZN(n9376) );
  MUX2_X1 U11701 ( .A(P1_B_REG_SCAN_IN), .B(n9376), .S(n11746), .Z(n9377) );
  AND2_X2 U11702 ( .A1(n10191), .A2(n9705), .ZN(n15050) );
  INV_X1 U11703 ( .A(n9378), .ZN(n14705) );
  NAND2_X1 U11704 ( .A1(n14705), .A2(n11806), .ZN(n9704) );
  OAI22_X1 U11705 ( .A1(n15050), .A2(P1_D_REG_1__SCAN_IN), .B1(n9380), .B2(
        n9704), .ZN(n9379) );
  INV_X1 U11706 ( .A(n9379), .ZN(P1_U3446) );
  NAND2_X1 U11707 ( .A1(n14705), .A2(n11746), .ZN(n9693) );
  OAI22_X1 U11708 ( .A1(n15050), .A2(P1_D_REG_0__SCAN_IN), .B1(n9380), .B2(
        n9693), .ZN(n9381) );
  INV_X1 U11709 ( .A(n9381), .ZN(P1_U3445) );
  INV_X1 U11710 ( .A(n10820), .ZN(n9390) );
  INV_X1 U11711 ( .A(n9912), .ZN(n9823) );
  OAI222_X1 U11712 ( .A1(n13999), .A2(n9382), .B1(n13994), .B2(n9390), .C1(
        P2_U3088), .C2(n9823), .ZN(P2_U3318) );
  INV_X1 U11713 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11714 ( .A1(n9384), .A2(n9383), .ZN(n9385) );
  NAND2_X1 U11715 ( .A1(n9385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9387) );
  INV_X1 U11716 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U11717 ( .A1(n9387), .A2(n9386), .ZN(n9463) );
  OR2_X1 U11718 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  INV_X1 U11719 ( .A(n10821), .ZN(n9784) );
  OAI222_X1 U11720 ( .A1(n9784), .A2(P1_U3086), .B1(n14707), .B2(n9390), .C1(
        n9389), .C2(n14709), .ZN(P1_U3346) );
  OAI222_X1 U11721 ( .A1(n12796), .A2(P3_U3151), .B1(n13303), .B2(n9392), .C1(
        n9391), .C2(n11887), .ZN(P3_U3281) );
  NAND2_X1 U11722 ( .A1(n9633), .A2(n9234), .ZN(n9394) );
  NAND2_X1 U11723 ( .A1(n9394), .A2(n9393), .ZN(n9396) );
  NAND2_X1 U11724 ( .A1(n9396), .A2(n9395), .ZN(n9410) );
  OR2_X1 U11725 ( .A1(n9410), .A2(P2_U3088), .ZN(n15127) );
  INV_X1 U11726 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10675) );
  AND2_X1 U11727 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9447) );
  NAND2_X1 U11728 ( .A1(n9397), .A2(n9447), .ZN(n9448) );
  OAI21_X1 U11729 ( .B1(n10675), .B2(n9453), .A(n9448), .ZN(n13498) );
  INV_X1 U11730 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9398) );
  MUX2_X1 U11731 ( .A(n9398), .B(P2_REG2_REG_2__SCAN_IN), .S(n13496), .Z(n9399) );
  NAND2_X1 U11732 ( .A1(n13498), .A2(n9399), .ZN(n13514) );
  NAND2_X1 U11733 ( .A1(n9415), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13513) );
  MUX2_X1 U11734 ( .A(n6885), .B(P2_REG2_REG_3__SCAN_IN), .S(n13505), .Z(
        n13512) );
  AOI21_X1 U11735 ( .B1(n13514), .B2(n13513), .A(n13512), .ZN(n13511) );
  INV_X1 U11736 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9400) );
  MUX2_X1 U11737 ( .A(n9400), .B(P2_REG2_REG_4__SCAN_IN), .S(n9599), .Z(n9594)
         );
  NOR2_X1 U11738 ( .A1(n9401), .A2(n9400), .ZN(n9433) );
  INV_X1 U11739 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10318) );
  MUX2_X1 U11740 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10318), .S(n9443), .Z(n9402) );
  NAND2_X1 U11741 ( .A1(n9443), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9406) );
  INV_X1 U11742 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9403) );
  MUX2_X1 U11743 ( .A(n9403), .B(P2_REG2_REG_6__SCAN_IN), .S(n9544), .Z(n9405)
         );
  INV_X1 U11744 ( .A(n9543), .ZN(n9408) );
  NOR2_X1 U11745 ( .A1(n9247), .A2(P2_U3088), .ZN(n13991) );
  NAND2_X1 U11746 ( .A1(n9410), .A2(n13991), .ZN(n9426) );
  INV_X1 U11747 ( .A(n9426), .ZN(n9404) );
  NAND3_X1 U11748 ( .A1(n9436), .A2(n9406), .A3(n9405), .ZN(n9407) );
  NAND3_X1 U11749 ( .A1(n9408), .A2(n15158), .A3(n9407), .ZN(n9432) );
  AND2_X1 U11750 ( .A1(n9247), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9409) );
  NAND2_X1 U11751 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10143) );
  INV_X1 U11752 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9411) );
  MUX2_X1 U11753 ( .A(n9411), .B(P2_REG1_REG_1__SCAN_IN), .S(n9453), .Z(n9412)
         );
  AND2_X1 U11754 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9452) );
  NAND2_X1 U11755 ( .A1(n9412), .A2(n9452), .ZN(n9454) );
  INV_X1 U11756 ( .A(n9453), .ZN(n9460) );
  NAND2_X1 U11757 ( .A1(n9460), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11758 ( .A1(n9454), .A2(n9413), .ZN(n13494) );
  INV_X1 U11759 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U11760 ( .A(n9414), .B(P2_REG1_REG_2__SCAN_IN), .S(n13496), .Z(
        n13495) );
  NAND2_X1 U11761 ( .A1(n13494), .A2(n13495), .ZN(n13507) );
  NAND2_X1 U11762 ( .A1(n9415), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U11763 ( .A1(n13507), .A2(n13506), .ZN(n9417) );
  MUX2_X1 U11764 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8537), .S(n13505), .Z(n9416) );
  NAND2_X1 U11765 ( .A1(n9417), .A2(n9416), .ZN(n13510) );
  NAND2_X1 U11766 ( .A1(n13505), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U11767 ( .A1(n13510), .A2(n9590), .ZN(n9420) );
  INV_X1 U11768 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9418) );
  MUX2_X1 U11769 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9418), .S(n9599), .Z(n9419)
         );
  NAND2_X1 U11770 ( .A1(n9420), .A2(n9419), .ZN(n9592) );
  NAND2_X1 U11771 ( .A1(n9599), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11772 ( .A1(n9592), .A2(n9421), .ZN(n9440) );
  INV_X1 U11773 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9422) );
  MUX2_X1 U11774 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9422), .S(n9443), .Z(n9439)
         );
  NAND2_X1 U11775 ( .A1(n9440), .A2(n9439), .ZN(n9438) );
  NAND2_X1 U11776 ( .A1(n9443), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U11777 ( .A1(n9438), .A2(n9423), .ZN(n9428) );
  INV_X1 U11778 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9424) );
  MUX2_X1 U11779 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9424), .S(n9544), .Z(n9427)
         );
  INV_X1 U11780 ( .A(n13556), .ZN(n15161) );
  NAND2_X1 U11781 ( .A1(n9428), .A2(n9427), .ZN(n9537) );
  OAI211_X1 U11782 ( .C1(n9428), .C2(n9427), .A(n15161), .B(n9537), .ZN(n9429)
         );
  NAND2_X1 U11783 ( .A1(n10143), .A2(n9429), .ZN(n9430) );
  AOI21_X1 U11784 ( .B1(n15155), .B2(n9544), .A(n9430), .ZN(n9431) );
  OAI211_X1 U11785 ( .C1(n15127), .C2(n7360), .A(n9432), .B(n9431), .ZN(
        P2_U3220) );
  INV_X1 U11786 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9446) );
  INV_X1 U11787 ( .A(n9433), .ZN(n9435) );
  MUX2_X1 U11788 ( .A(n10318), .B(P2_REG2_REG_5__SCAN_IN), .S(n9443), .Z(n9434) );
  NAND2_X1 U11789 ( .A1(n9435), .A2(n9434), .ZN(n9437) );
  OAI211_X1 U11790 ( .C1(n9593), .C2(n9437), .A(n15158), .B(n9436), .ZN(n9445)
         );
  NAND2_X1 U11791 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10074) );
  OAI211_X1 U11792 ( .C1(n9440), .C2(n9439), .A(n15161), .B(n9438), .ZN(n9441)
         );
  NAND2_X1 U11793 ( .A1(n10074), .A2(n9441), .ZN(n9442) );
  AOI21_X1 U11794 ( .B1(n15155), .B2(n9443), .A(n9442), .ZN(n9444) );
  OAI211_X1 U11795 ( .C1(n15127), .C2(n9446), .A(n9445), .B(n9444), .ZN(
        P2_U3219) );
  MUX2_X1 U11796 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10675), .S(n9453), .Z(n9451) );
  INV_X1 U11797 ( .A(n9447), .ZN(n9450) );
  INV_X1 U11798 ( .A(n9448), .ZN(n9449) );
  AOI211_X1 U11799 ( .C1(n9451), .C2(n9450), .A(n9449), .B(n15129), .ZN(n9459)
         );
  INV_X1 U11800 ( .A(n9452), .ZN(n9457) );
  MUX2_X1 U11801 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9411), .S(n9453), .Z(n9456)
         );
  INV_X1 U11802 ( .A(n9454), .ZN(n9455) );
  AOI211_X1 U11803 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n13556), .ZN(n9458)
         );
  NOR2_X1 U11804 ( .A1(n9459), .A2(n9458), .ZN(n9462) );
  AOI22_X1 U11805 ( .A1(n15155), .A2(n9460), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3088), .ZN(n9461) );
  OAI211_X1 U11806 ( .C1(n15127), .C2(n7102), .A(n9462), .B(n9461), .ZN(
        P2_U3215) );
  NAND2_X1 U11807 ( .A1(n9463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9464) );
  XNOR2_X1 U11808 ( .A(n9464), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14220) );
  INV_X1 U11809 ( .A(n14220), .ZN(n9466) );
  INV_X1 U11810 ( .A(n10825), .ZN(n9467) );
  OAI222_X1 U11811 ( .A1(n9466), .A2(P1_U3086), .B1(n14707), .B2(n9467), .C1(
        n9465), .C2(n14709), .ZN(P1_U3345) );
  INV_X1 U11812 ( .A(n9994), .ZN(n10003) );
  OAI222_X1 U11813 ( .A1(n13999), .A2(n9468), .B1(n13994), .B2(n9467), .C1(
        P2_U3088), .C2(n10003), .ZN(P2_U3317) );
  AOI22_X1 U11814 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15161), .B1(n15158), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9472) );
  INV_X1 U11815 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9470) );
  OAI21_X1 U11816 ( .B1(n15129), .B2(P2_REG2_REG_0__SCAN_IN), .A(n15143), .ZN(
        n9469) );
  AOI21_X1 U11817 ( .B1(n15161), .B2(n9470), .A(n9469), .ZN(n9471) );
  MUX2_X1 U11818 ( .A(n9472), .B(n9471), .S(P2_IR_REG_0__SCAN_IN), .Z(n9474)
         );
  INV_X1 U11819 ( .A(n15127), .ZN(n15154) );
  AOI22_X1 U11820 ( .A1(n15154), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9473) );
  NAND2_X1 U11821 ( .A1(n9474), .A2(n9473), .ZN(P2_U3214) );
  INV_X1 U11822 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9475) );
  MUX2_X1 U11823 ( .A(n9475), .B(P1_REG1_REG_5__SCAN_IN), .S(n10233), .Z(n9488) );
  INV_X1 U11824 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U11825 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9476), .S(n14173), .Z(
        n14177) );
  INV_X1 U11826 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15112) );
  MUX2_X1 U11827 ( .A(n15112), .B(P1_REG1_REG_1__SCAN_IN), .S(n14162), .Z(
        n9478) );
  AND2_X1 U11828 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9477) );
  NAND2_X1 U11829 ( .A1(n9478), .A2(n9477), .ZN(n14166) );
  OAI21_X1 U11830 ( .B1(n15112), .B2(n14162), .A(n14166), .ZN(n14176) );
  NAND2_X1 U11831 ( .A1(n14177), .A2(n14176), .ZN(n14187) );
  NAND2_X1 U11832 ( .A1(n14173), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14186) );
  NAND2_X1 U11833 ( .A1(n14187), .A2(n14186), .ZN(n9481) );
  INV_X1 U11834 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9479) );
  MUX2_X1 U11835 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9479), .S(n14184), .Z(n9480) );
  NAND2_X1 U11836 ( .A1(n9481), .A2(n9480), .ZN(n14189) );
  NAND2_X1 U11837 ( .A1(n14184), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U11838 ( .A1(n14189), .A2(n9882), .ZN(n9484) );
  INV_X1 U11839 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9482) );
  MUX2_X1 U11840 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9482), .S(n10228), .Z(n9483) );
  NAND2_X1 U11841 ( .A1(n9484), .A2(n9483), .ZN(n9884) );
  NAND2_X1 U11842 ( .A1(n10228), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U11843 ( .A1(n9884), .A2(n9485), .ZN(n9487) );
  OR2_X1 U11844 ( .A1(n9487), .A2(n9488), .ZN(n9506) );
  INV_X1 U11845 ( .A(n9506), .ZN(n9486) );
  AOI21_X1 U11846 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9504) );
  NAND2_X1 U11847 ( .A1(n9490), .A2(n9489), .ZN(n14980) );
  INV_X1 U11848 ( .A(n9491), .ZN(n12253) );
  INV_X1 U11849 ( .A(n14700), .ZN(n9895) );
  INV_X1 U11850 ( .A(n14977), .ZN(n14996) );
  INV_X1 U11851 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U11852 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9492) );
  OAI21_X1 U11853 ( .B1(n14996), .B2(n9493), .A(n9492), .ZN(n9494) );
  AOI21_X1 U11854 ( .B1(n10233), .B2(n14219), .A(n9494), .ZN(n9503) );
  OR3_X1 U11855 ( .A1(n14980), .A2(n9491), .A3(n14700), .ZN(n14983) );
  INV_X1 U11856 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9495) );
  MUX2_X1 U11857 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9495), .S(n14173), .Z(
        n14175) );
  INV_X1 U11858 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9496) );
  MUX2_X1 U11859 ( .A(n9496), .B(P1_REG2_REG_1__SCAN_IN), .S(n14162), .Z(
        n14159) );
  NAND3_X1 U11860 ( .A1(n14159), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG2_REG_0__SCAN_IN), .ZN(n14158) );
  OAI21_X1 U11861 ( .B1(n9496), .B2(n14162), .A(n14158), .ZN(n14174) );
  NAND2_X1 U11862 ( .A1(n14175), .A2(n14174), .ZN(n14193) );
  NAND2_X1 U11863 ( .A1(n14173), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14192) );
  INV_X1 U11864 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U11865 ( .A(n10202), .B(P1_REG2_REG_3__SCAN_IN), .S(n14184), .Z(
        n14191) );
  AOI21_X1 U11866 ( .B1(n14193), .B2(n14192), .A(n14191), .ZN(n14190) );
  NOR2_X1 U11867 ( .A1(n9497), .A2(n10202), .ZN(n9885) );
  INV_X1 U11868 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10466) );
  MUX2_X1 U11869 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10466), .S(n10228), .Z(
        n9498) );
  OAI21_X1 U11870 ( .B1(n14190), .B2(n9885), .A(n9498), .ZN(n9888) );
  NAND2_X1 U11871 ( .A1(n10228), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9500) );
  INV_X1 U11872 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9518) );
  MUX2_X1 U11873 ( .A(n9518), .B(P1_REG2_REG_5__SCAN_IN), .S(n10233), .Z(n9499) );
  AOI21_X1 U11874 ( .B1(n9888), .B2(n9500), .A(n9499), .ZN(n9522) );
  INV_X1 U11875 ( .A(n9522), .ZN(n14208) );
  NAND3_X1 U11876 ( .A1(n9888), .A2(n9500), .A3(n9499), .ZN(n9501) );
  NAND3_X1 U11877 ( .A1(n14243), .A2(n14208), .A3(n9501), .ZN(n9502) );
  OAI211_X1 U11878 ( .C1(n9504), .C2(n14987), .A(n9503), .B(n9502), .ZN(
        P1_U3248) );
  OR2_X1 U11879 ( .A1(n10233), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9505) );
  AND2_X1 U11880 ( .A1(n9506), .A2(n9505), .ZN(n14203) );
  INV_X1 U11881 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9507) );
  MUX2_X1 U11882 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9507), .S(n14205), .Z(
        n14202) );
  NAND2_X1 U11883 ( .A1(n14203), .A2(n14202), .ZN(n14201) );
  NAND2_X1 U11884 ( .A1(n14205), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U11885 ( .A1(n14201), .A2(n9560), .ZN(n9510) );
  INV_X1 U11886 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9508) );
  MUX2_X1 U11887 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9508), .S(n10477), .Z(n9509) );
  NAND2_X1 U11888 ( .A1(n9510), .A2(n9509), .ZN(n9562) );
  NAND2_X1 U11889 ( .A1(n10477), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11890 ( .A1(n9562), .A2(n9511), .ZN(n9577) );
  INV_X1 U11891 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9512) );
  MUX2_X1 U11892 ( .A(n9512), .B(P1_REG1_REG_8__SCAN_IN), .S(n10740), .Z(n9578) );
  OR2_X1 U11893 ( .A1(n9577), .A2(n9578), .ZN(n9575) );
  OR2_X1 U11894 ( .A1(n10740), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U11895 ( .A1(n9575), .A2(n9515), .ZN(n9513) );
  INV_X1 U11896 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15118) );
  MUX2_X1 U11897 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15118), .S(n10821), .Z(
        n9514) );
  NAND2_X1 U11898 ( .A1(n9513), .A2(n9514), .ZN(n9786) );
  INV_X1 U11899 ( .A(n9514), .ZN(n9516) );
  NAND3_X1 U11900 ( .A1(n9575), .A2(n9516), .A3(n9515), .ZN(n9517) );
  AND2_X1 U11901 ( .A1(n9786), .A2(n9517), .ZN(n9535) );
  NOR2_X1 U11902 ( .A1(n9519), .A2(n9518), .ZN(n14204) );
  INV_X1 U11903 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9520) );
  MUX2_X1 U11904 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9520), .S(n14205), .Z(n9521) );
  OAI21_X1 U11905 ( .B1(n9522), .B2(n14204), .A(n9521), .ZN(n14210) );
  NAND2_X1 U11906 ( .A1(n14205), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9555) );
  INV_X1 U11907 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9523) );
  MUX2_X1 U11908 ( .A(n9523), .B(P1_REG2_REG_7__SCAN_IN), .S(n10477), .Z(n9554) );
  AOI21_X1 U11909 ( .B1(n14210), .B2(n9555), .A(n9554), .ZN(n9585) );
  NOR2_X1 U11910 ( .A1(n9524), .A2(n9523), .ZN(n9580) );
  INV_X1 U11911 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9525) );
  MUX2_X1 U11912 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9525), .S(n10740), .Z(n9526) );
  OAI21_X1 U11913 ( .B1(n9585), .B2(n9580), .A(n9526), .ZN(n9583) );
  NAND2_X1 U11914 ( .A1(n10740), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9528) );
  INV_X1 U11915 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9775) );
  MUX2_X1 U11916 ( .A(n9775), .B(P1_REG2_REG_9__SCAN_IN), .S(n10821), .Z(n9527) );
  AOI21_X1 U11917 ( .B1(n9583), .B2(n9528), .A(n9527), .ZN(n14226) );
  INV_X1 U11918 ( .A(n14226), .ZN(n9530) );
  NAND3_X1 U11919 ( .A1(n9583), .A2(n9528), .A3(n9527), .ZN(n9529) );
  NAND3_X1 U11920 ( .A1(n9530), .A2(n14243), .A3(n9529), .ZN(n9534) );
  INV_X1 U11921 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14732) );
  NAND2_X1 U11922 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9531) );
  OAI21_X1 U11923 ( .B1(n14996), .B2(n14732), .A(n9531), .ZN(n9532) );
  AOI21_X1 U11924 ( .B1(n10821), .B2(n14219), .A(n9532), .ZN(n9533) );
  OAI211_X1 U11925 ( .C1(n9535), .C2(n14987), .A(n9534), .B(n9533), .ZN(
        P1_U3252) );
  NAND2_X1 U11926 ( .A1(n9544), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U11927 ( .A1(n9537), .A2(n9536), .ZN(n15136) );
  INV_X1 U11928 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9538) );
  MUX2_X1 U11929 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9538), .S(n15124), .Z(
        n15135) );
  NAND2_X1 U11930 ( .A1(n15136), .A2(n15135), .ZN(n15134) );
  NAND2_X1 U11931 ( .A1(n15124), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9540) );
  INV_X1 U11932 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10374) );
  MUX2_X1 U11933 ( .A(n10374), .B(P2_REG1_REG_8__SCAN_IN), .S(n9807), .Z(n9539) );
  AOI21_X1 U11934 ( .B1(n15134), .B2(n9540), .A(n9539), .ZN(n9806) );
  NAND3_X1 U11935 ( .A1(n15134), .A2(n9540), .A3(n9539), .ZN(n9541) );
  NAND2_X1 U11936 ( .A1(n15161), .A2(n9541), .ZN(n9553) );
  NAND2_X1 U11937 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10440) );
  OAI21_X1 U11938 ( .B1(n15143), .B2(n9542), .A(n10440), .ZN(n9551) );
  AOI21_X1 U11939 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9544), .A(n9543), .ZN(
        n15131) );
  INV_X1 U11940 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9545) );
  MUX2_X1 U11941 ( .A(n9545), .B(P2_REG2_REG_7__SCAN_IN), .S(n15124), .Z(
        n15130) );
  NAND2_X1 U11942 ( .A1(n15124), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9548) );
  INV_X1 U11943 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9546) );
  MUX2_X1 U11944 ( .A(n9546), .B(P2_REG2_REG_8__SCAN_IN), .S(n9807), .Z(n9547)
         );
  AND3_X1 U11945 ( .A1(n15132), .A2(n9548), .A3(n9547), .ZN(n9549) );
  NOR3_X1 U11946 ( .A1(n9805), .A2(n9549), .A3(n15129), .ZN(n9550) );
  AOI211_X1 U11947 ( .C1(n15154), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9551), .B(
        n9550), .ZN(n9552) );
  OAI21_X1 U11948 ( .B1(n9806), .B2(n9553), .A(n9552), .ZN(P2_U3222) );
  NAND3_X1 U11949 ( .A1(n14210), .A2(n9555), .A3(n9554), .ZN(n9556) );
  NAND2_X1 U11950 ( .A1(n14243), .A2(n9556), .ZN(n9565) );
  INV_X1 U11951 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U11952 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10956) );
  OAI21_X1 U11953 ( .B1(n14996), .B2(n9557), .A(n10956), .ZN(n9558) );
  AOI21_X1 U11954 ( .B1(n10477), .B2(n14219), .A(n9558), .ZN(n9564) );
  MUX2_X1 U11955 ( .A(n9508), .B(P1_REG1_REG_7__SCAN_IN), .S(n10477), .Z(n9559) );
  NAND3_X1 U11956 ( .A1(n14201), .A2(n9560), .A3(n9559), .ZN(n9561) );
  NAND3_X1 U11957 ( .A1(n14245), .A2(n9562), .A3(n9561), .ZN(n9563) );
  OAI211_X1 U11958 ( .C1(n9585), .C2(n9565), .A(n9564), .B(n9563), .ZN(
        P1_U3250) );
  INV_X1 U11959 ( .A(n11321), .ZN(n9573) );
  INV_X1 U11960 ( .A(n10006), .ZN(n10173) );
  OAI222_X1 U11961 ( .A1(n13999), .A2(n9566), .B1(n13994), .B2(n9573), .C1(
        P2_U3088), .C2(n10173), .ZN(P2_U3316) );
  INV_X1 U11962 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U11963 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  NOR2_X1 U11964 ( .A1(n9570), .A2(n9569), .ZN(n9762) );
  OR2_X1 U11965 ( .A1(n9762), .A2(n9306), .ZN(n9571) );
  XNOR2_X1 U11966 ( .A(n9571), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11322) );
  INV_X1 U11967 ( .A(n11322), .ZN(n9574) );
  OAI222_X1 U11968 ( .A1(n9574), .A2(P1_U3086), .B1(n14707), .B2(n9573), .C1(
        n9572), .C2(n14709), .ZN(P1_U3344) );
  INV_X1 U11969 ( .A(n9575), .ZN(n9576) );
  AOI21_X1 U11970 ( .B1(n9578), .B2(n9577), .A(n9576), .ZN(n9588) );
  INV_X1 U11971 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14730) );
  NAND2_X1 U11972 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11063) );
  OAI21_X1 U11973 ( .B1(n14996), .B2(n14730), .A(n11063), .ZN(n9579) );
  AOI21_X1 U11974 ( .B1(n10740), .B2(n14219), .A(n9579), .ZN(n9587) );
  MUX2_X1 U11975 ( .A(n9525), .B(P1_REG2_REG_8__SCAN_IN), .S(n10740), .Z(n9582) );
  INV_X1 U11976 ( .A(n9580), .ZN(n9581) );
  NAND2_X1 U11977 ( .A1(n9582), .A2(n9581), .ZN(n9584) );
  OAI211_X1 U11978 ( .C1(n9585), .C2(n9584), .A(n14243), .B(n9583), .ZN(n9586)
         );
  OAI211_X1 U11979 ( .C1(n9588), .C2(n14987), .A(n9587), .B(n9586), .ZN(
        P1_U3251) );
  INV_X1 U11980 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9602) );
  MUX2_X1 U11981 ( .A(n9418), .B(P2_REG1_REG_4__SCAN_IN), .S(n9599), .Z(n9589)
         );
  NAND3_X1 U11982 ( .A1(n13510), .A2(n9590), .A3(n9589), .ZN(n9591) );
  NAND3_X1 U11983 ( .A1(n15161), .A2(n9592), .A3(n9591), .ZN(n9601) );
  NAND2_X1 U11984 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9933) );
  AOI211_X1 U11985 ( .C1(n9595), .C2(n9594), .A(n9593), .B(n15129), .ZN(n9596)
         );
  INV_X1 U11986 ( .A(n9596), .ZN(n9597) );
  NAND2_X1 U11987 ( .A1(n9933), .A2(n9597), .ZN(n9598) );
  AOI21_X1 U11988 ( .B1(n15155), .B2(n9599), .A(n9598), .ZN(n9600) );
  OAI211_X1 U11989 ( .C1(n15127), .C2(n9602), .A(n9601), .B(n9600), .ZN(
        P2_U3218) );
  INV_X1 U11990 ( .A(n12809), .ZN(n12797) );
  INV_X1 U11991 ( .A(n9603), .ZN(n9605) );
  OAI222_X1 U11992 ( .A1(n12797), .A2(P3_U3151), .B1(n11891), .B2(n9605), .C1(
        n9604), .C2(n11887), .ZN(P3_U3280) );
  XNOR2_X1 U11993 ( .A(n11744), .B(P2_B_REG_SCAN_IN), .ZN(n9606) );
  INV_X1 U11994 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U11995 ( .A1(n15167), .A2(n15174), .ZN(n9608) );
  NAND2_X1 U11996 ( .A1(n14002), .A2(n11807), .ZN(n9607) );
  NAND2_X1 U11997 ( .A1(n9608), .A2(n9607), .ZN(n15175) );
  INV_X1 U11998 ( .A(n15175), .ZN(n10301) );
  INV_X1 U11999 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15172) );
  NAND2_X1 U12000 ( .A1(n15167), .A2(n15172), .ZN(n9610) );
  NAND2_X1 U12001 ( .A1(n14002), .A2(n11744), .ZN(n9609) );
  AND2_X1 U12002 ( .A1(n9610), .A2(n9609), .ZN(n15170) );
  NOR4_X1 U12003 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9614) );
  NOR4_X1 U12004 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n9613) );
  NOR4_X1 U12005 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9612) );
  NOR4_X1 U12006 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9611) );
  NAND4_X1 U12007 ( .A1(n9614), .A2(n9613), .A3(n9612), .A4(n9611), .ZN(n9620)
         );
  NOR2_X1 U12008 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n9618) );
  NOR4_X1 U12009 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9617) );
  NOR4_X1 U12010 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9616) );
  NOR4_X1 U12011 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9615) );
  NAND4_X1 U12012 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n9619)
         );
  OAI21_X1 U12013 ( .B1(n9620), .B2(n9619), .A(n15167), .ZN(n9658) );
  NAND3_X1 U12014 ( .A1(n10301), .A2(n15170), .A3(n9658), .ZN(n9632) );
  INV_X1 U12015 ( .A(n15176), .ZN(n15173) );
  OR2_X1 U12016 ( .A1(n9632), .A2(n15173), .ZN(n9630) );
  INV_X1 U12017 ( .A(n9630), .ZN(n9624) );
  INV_X1 U12018 ( .A(n9633), .ZN(n9622) );
  AND2_X1 U12019 ( .A1(n9622), .A2(n11874), .ZN(n9623) );
  OAI21_X1 U12020 ( .B1(n10023), .B2(n9625), .A(n9648), .ZN(n9627) );
  NOR2_X2 U12021 ( .A1(n9630), .A2(n8471), .ZN(n14885) );
  INV_X1 U12022 ( .A(n13570), .ZN(n13455) );
  INV_X1 U12023 ( .A(n13489), .ZN(n9626) );
  NOR2_X1 U12024 ( .A1(n13455), .A2(n9626), .ZN(n9769) );
  AOI22_X1 U12025 ( .A1(n14883), .A2(n9627), .B1(n14885), .B2(n9769), .ZN(
        n9638) );
  OR2_X1 U12026 ( .A1(n10540), .A2(n10962), .ZN(n10308) );
  INV_X1 U12027 ( .A(n9659), .ZN(n9629) );
  NAND2_X1 U12028 ( .A1(n9632), .A2(n9659), .ZN(n9636) );
  NAND2_X1 U12029 ( .A1(n9633), .A2(n8471), .ZN(n9657) );
  AND2_X1 U12030 ( .A1(n9634), .A2(n9657), .ZN(n9635) );
  NAND2_X1 U12031 ( .A1(n9636), .A2(n9635), .ZN(n9829) );
  OR2_X1 U12032 ( .A1(n9829), .A2(P2_U3088), .ZN(n9679) );
  AOI22_X1 U12033 ( .A1(n9631), .A2(n10541), .B1(n9679), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12034 ( .A1(n9638), .A2(n9637), .ZN(P2_U3204) );
  XNOR2_X1 U12035 ( .A(n10908), .B(P3_B_REG_SCAN_IN), .ZN(n9639) );
  AOI21_X2 U12036 ( .B1(n11032), .B2(n9639), .A(n11301), .ZN(n11883) );
  INV_X1 U12037 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12038 ( .A1(n11883), .A2(n9640), .ZN(n9642) );
  NAND2_X1 U12039 ( .A1(n10908), .A2(n11301), .ZN(n9641) );
  NAND2_X1 U12040 ( .A1(n11882), .A2(P3_D_REG_0__SCAN_IN), .ZN(n9643) );
  OAI21_X1 U12041 ( .B1(n10610), .B2(n11882), .A(n9643), .ZN(P3_U3376) );
  NAND2_X1 U12042 ( .A1(n13464), .A2(n13491), .ZN(n9646) );
  NAND2_X1 U12043 ( .A1(n13570), .A2(n9210), .ZN(n9645) );
  NAND2_X1 U12044 ( .A1(n9646), .A2(n9645), .ZN(n9671) );
  AOI22_X1 U12045 ( .A1(n14885), .A2(n9671), .B1(n9679), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9653) );
  INV_X1 U12046 ( .A(n10305), .ZN(n9647) );
  NAND2_X1 U12047 ( .A1(n13489), .A2(n9680), .ZN(n9683) );
  XNOR2_X1 U12048 ( .A(n9685), .B(n9683), .ZN(n9649) );
  OAI21_X1 U12049 ( .B1(n13338), .B2(n10541), .A(n9648), .ZN(n9650) );
  NAND2_X1 U12050 ( .A1(n9649), .A2(n9650), .ZN(n9687) );
  OAI21_X1 U12051 ( .B1(n9649), .B2(n9650), .A(n9687), .ZN(n9651) );
  NAND2_X1 U12052 ( .A1(n14883), .A2(n9651), .ZN(n9652) );
  OAI211_X1 U12053 ( .C1(n13452), .C2(n10049), .A(n9653), .B(n9652), .ZN(
        P2_U3194) );
  INV_X1 U12054 ( .A(n12830), .ZN(n12814) );
  INV_X1 U12055 ( .A(n9654), .ZN(n9656) );
  OAI222_X1 U12056 ( .A1(n12814), .A2(P3_U3151), .B1(n13303), .B2(n9656), .C1(
        n9655), .C2(n11887), .ZN(P3_U3279) );
  AND2_X1 U12057 ( .A1(n15175), .A2(n9659), .ZN(n9767) );
  INV_X1 U12058 ( .A(n9661), .ZN(n9662) );
  NAND2_X1 U12059 ( .A1(n9666), .A2(n9662), .ZN(n9663) );
  NAND2_X1 U12060 ( .A1(n9795), .A2(n9663), .ZN(n10680) );
  INV_X1 U12061 ( .A(n10680), .ZN(n9674) );
  INV_X1 U12062 ( .A(n9665), .ZN(n13891) );
  OR2_X1 U12063 ( .A1(n8482), .A2(n9628), .ZN(n9670) );
  NAND2_X1 U12064 ( .A1(n8466), .A2(n9668), .ZN(n9669) );
  AOI21_X1 U12065 ( .B1(n9672), .B2(n13822), .A(n9671), .ZN(n10682) );
  OAI211_X1 U12066 ( .C1(n10049), .C2(n9673), .A(n10023), .B(n9797), .ZN(
        n10678) );
  OAI211_X1 U12067 ( .C1(n9674), .C2(n15182), .A(n10682), .B(n10678), .ZN(
        n10051) );
  NAND2_X1 U12068 ( .A1(n15190), .A2(n15179), .ZN(n13912) );
  OAI22_X1 U12069 ( .A1(n13912), .A2(n10049), .B1(n15190), .B2(n9411), .ZN(
        n9675) );
  AOI21_X1 U12070 ( .B1(n15190), .B2(n10051), .A(n9675), .ZN(n9676) );
  INV_X1 U12071 ( .A(n9676), .ZN(P2_U3500) );
  INV_X1 U12072 ( .A(n10053), .ZN(n10568) );
  NAND2_X1 U12073 ( .A1(n13464), .A2(n13489), .ZN(n9678) );
  NAND2_X1 U12074 ( .A1(n13570), .A2(n13488), .ZN(n9677) );
  NAND2_X1 U12075 ( .A1(n9678), .A2(n9677), .ZN(n9801) );
  AOI22_X1 U12076 ( .A1(n14885), .A2(n9801), .B1(n9679), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n9692) );
  AND2_X1 U12077 ( .A1(n9210), .A2(n9680), .ZN(n9682) );
  NOR2_X1 U12078 ( .A1(n9681), .A2(n9682), .ZN(n9825) );
  INV_X1 U12079 ( .A(n9683), .ZN(n9684) );
  OR2_X1 U12080 ( .A1(n9685), .A2(n9684), .ZN(n9686) );
  NAND2_X1 U12081 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  OAI21_X1 U12082 ( .B1(n9689), .B2(n9688), .A(n9827), .ZN(n9690) );
  NAND2_X1 U12083 ( .A1(n14883), .A2(n9690), .ZN(n9691) );
  OAI211_X1 U12084 ( .C1(n13452), .C2(n10568), .A(n9692), .B(n9691), .ZN(
        P2_U3209) );
  NOR2_X1 U12085 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n15441) );
  NOR4_X1 U12086 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9696) );
  NOR4_X1 U12087 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9695) );
  NOR4_X1 U12088 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9694) );
  NAND4_X1 U12089 ( .A1(n15441), .A2(n9696), .A3(n9695), .A4(n9694), .ZN(n9702) );
  NOR4_X1 U12090 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9700) );
  NOR4_X1 U12091 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9699) );
  NOR4_X1 U12092 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9698) );
  NOR4_X1 U12093 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9697) );
  NAND4_X1 U12094 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(n9701)
         );
  NOR2_X1 U12095 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  NOR2_X1 U12096 ( .A1(n9705), .A2(n9703), .ZN(n9721) );
  NOR2_X1 U12097 ( .A1(n10203), .A2(n9721), .ZN(n9706) );
  OAI21_X1 U12098 ( .B1(n9705), .B2(P1_D_REG_1__SCAN_IN), .A(n9704), .ZN(
        n10187) );
  INV_X1 U12099 ( .A(n10187), .ZN(n9723) );
  NAND2_X1 U12100 ( .A1(n9706), .A2(n9723), .ZN(n9742) );
  NAND2_X1 U12101 ( .A1(n9707), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9708) );
  MUX2_X1 U12102 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9708), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9710) );
  NAND2_X1 U12103 ( .A1(n9711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U12104 ( .A1(n15016), .A2(n14433), .ZN(n10189) );
  NAND2_X1 U12105 ( .A1(n9742), .A2(n10189), .ZN(n10126) );
  NAND2_X1 U12106 ( .A1(n10126), .A2(n10191), .ZN(n14913) );
  NAND2_X1 U12107 ( .A1(n10923), .A2(n14320), .ZN(n9719) );
  AND2_X1 U12108 ( .A1(n9719), .A2(n9756), .ZN(n9713) );
  INV_X1 U12109 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14164) );
  INV_X1 U12110 ( .A(SI_0_), .ZN(n9715) );
  OAI21_X1 U12111 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9717) );
  NAND2_X1 U12112 ( .A1(n9718), .A2(n9717), .ZN(n14711) );
  NAND2_X1 U12113 ( .A1(n9871), .A2(n9719), .ZN(n9747) );
  NAND3_X1 U12114 ( .A1(n9747), .A2(n9720), .A3(n9736), .ZN(n10124) );
  NOR2_X1 U12115 ( .A1(n10124), .A2(P1_U3086), .ZN(n12254) );
  INV_X1 U12116 ( .A(n9721), .ZN(n9722) );
  NAND2_X1 U12117 ( .A1(n12254), .A2(n9722), .ZN(n10188) );
  INV_X1 U12118 ( .A(n10203), .ZN(n10289) );
  NAND2_X1 U12119 ( .A1(n9723), .A2(n10289), .ZN(n9724) );
  INV_X1 U12120 ( .A(n14111), .ZN(n14143) );
  NAND2_X1 U12121 ( .A1(n9871), .A2(n14700), .ZN(n14527) );
  NAND2_X1 U12122 ( .A1(n14143), .A2(n14509), .ZN(n14120) );
  INV_X1 U12123 ( .A(n14120), .ZN(n14925) );
  NAND2_X1 U12124 ( .A1(n10243), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9728) );
  INV_X1 U12125 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9735) );
  INV_X2 U12126 ( .A(n10783), .ZN(n12404) );
  INV_X1 U12127 ( .A(n14999), .ZN(n9757) );
  NAND2_X1 U12128 ( .A1(n12404), .A2(n9757), .ZN(n9734) );
  NAND2_X1 U12129 ( .A1(n11974), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12130 ( .A1(n10243), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U12131 ( .A1(n10484), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U12132 ( .A1(n15006), .A2(n10039), .ZN(n9733) );
  OAI211_X1 U12133 ( .C1(n9736), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9867)
         );
  INV_X1 U12134 ( .A(n9867), .ZN(n9741) );
  NAND2_X2 U12135 ( .A1(n12404), .A2(n14640), .ZN(n12360) );
  INV_X1 U12136 ( .A(n12360), .ZN(n9737) );
  NAND2_X1 U12137 ( .A1(n15006), .A2(n9737), .ZN(n9740) );
  AOI22_X1 U12138 ( .A1(n9757), .A2(n10039), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9738), .ZN(n9739) );
  NAND2_X1 U12139 ( .A1(n9740), .A2(n9739), .ZN(n9868) );
  XNOR2_X1 U12140 ( .A(n9741), .B(n9868), .ZN(n9894) );
  INV_X1 U12141 ( .A(n9742), .ZN(n9746) );
  INV_X1 U12142 ( .A(n10191), .ZN(n9744) );
  NAND2_X1 U12143 ( .A1(n15072), .A2(n12069), .ZN(n9743) );
  NOR2_X1 U12144 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  AOI22_X1 U12145 ( .A1(n14925), .A2(n15002), .B1(n9894), .B2(n14930), .ZN(
        n9750) );
  INV_X1 U12146 ( .A(n14913), .ZN(n9748) );
  NAND2_X1 U12147 ( .A1(n9748), .A2(n9747), .ZN(n10044) );
  NAND2_X1 U12148 ( .A1(n10044), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9749) );
  OAI211_X1 U12149 ( .C1(n14927), .C2(n14999), .A(n9750), .B(n9749), .ZN(
        P1_U3232) );
  NAND2_X1 U12150 ( .A1(n10189), .A2(n10187), .ZN(n9751) );
  OR2_X1 U12151 ( .A1(n10188), .A2(n9751), .ZN(n10290) );
  NOR2_X1 U12152 ( .A1(n10290), .A2(n10203), .ZN(n9971) );
  AND2_X1 U12153 ( .A1(n12105), .A2(n9752), .ZN(n9753) );
  NOR2_X1 U12154 ( .A1(n10786), .A2(n9753), .ZN(n10193) );
  NAND2_X1 U12155 ( .A1(n10193), .A2(n14320), .ZN(n10242) );
  INV_X1 U12156 ( .A(n12068), .ZN(n9754) );
  NAND2_X1 U12157 ( .A1(n9754), .A2(n14433), .ZN(n15064) );
  NAND2_X1 U12158 ( .A1(n9755), .A2(n12077), .ZN(n12076) );
  NAND2_X1 U12159 ( .A1(n12072), .A2(n14433), .ZN(n12074) );
  INV_X1 U12160 ( .A(n12106), .ZN(n12003) );
  OAI21_X1 U12161 ( .B1(n15108), .B2(n15079), .A(n12003), .ZN(n9759) );
  NAND2_X1 U12162 ( .A1(n14509), .A2(n15002), .ZN(n10524) );
  NAND3_X1 U12163 ( .A1(n9757), .A2(n12075), .A3(n9756), .ZN(n9758) );
  NAND3_X1 U12164 ( .A1(n9759), .A2(n10524), .A3(n9758), .ZN(n10366) );
  NAND2_X1 U12165 ( .A1(n10366), .A2(n15123), .ZN(n9760) );
  OAI21_X1 U12166 ( .B1(n15123), .B2(n9735), .A(n9760), .ZN(P1_U3528) );
  INV_X1 U12167 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U12168 ( .A1(n9762), .A2(n9761), .ZN(n10218) );
  NAND2_X1 U12169 ( .A1(n10218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9898) );
  XNOR2_X1 U12170 ( .A(n9898), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11467) );
  INV_X1 U12171 ( .A(n11467), .ZN(n9986) );
  INV_X1 U12172 ( .A(n11466), .ZN(n9765) );
  OAI222_X1 U12173 ( .A1(P1_U3086), .A2(n9986), .B1(n14707), .B2(n9765), .C1(
        n9763), .C2(n14709), .ZN(P1_U3343) );
  OAI222_X1 U12174 ( .A1(P2_U3088), .A2(n11270), .B1(n13994), .B2(n9765), .C1(
        n9764), .C2(n13999), .ZN(P2_U3315) );
  INV_X1 U12175 ( .A(n10300), .ZN(n9766) );
  NOR2_X1 U12176 ( .A1(n9766), .A2(n15170), .ZN(n9768) );
  INV_X2 U12177 ( .A(n15185), .ZN(n15187) );
  INV_X1 U12178 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9774) );
  AOI21_X1 U12179 ( .B1(n13795), .B2(n9664), .A(n10545), .ZN(n9770) );
  NOR2_X1 U12180 ( .A1(n9770), .A2(n9769), .ZN(n10538) );
  INV_X1 U12181 ( .A(n10540), .ZN(n9771) );
  NAND2_X1 U12182 ( .A1(n9771), .A2(n10541), .ZN(n9772) );
  OAI211_X1 U12183 ( .C1(n10545), .C2(n13891), .A(n10538), .B(n9772), .ZN(
        n13939) );
  NAND2_X1 U12184 ( .A1(n15187), .A2(n13939), .ZN(n9773) );
  OAI21_X1 U12185 ( .B1(n15187), .B2(n9774), .A(n9773), .ZN(P2_U3430) );
  NOR2_X1 U12186 ( .A1(n9784), .A2(n9775), .ZN(n14221) );
  INV_X1 U12187 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9776) );
  MUX2_X1 U12188 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9776), .S(n14220), .Z(
        n9777) );
  OAI21_X1 U12189 ( .B1(n14226), .B2(n14221), .A(n9777), .ZN(n14224) );
  NAND2_X1 U12190 ( .A1(n14220), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9780) );
  INV_X1 U12191 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9778) );
  MUX2_X1 U12192 ( .A(n9778), .B(P1_REG2_REG_11__SCAN_IN), .S(n11322), .Z(
        n9779) );
  AOI21_X1 U12193 ( .B1(n14224), .B2(n9780), .A(n9779), .ZN(n9974) );
  NAND3_X1 U12194 ( .A1(n14224), .A2(n9780), .A3(n9779), .ZN(n9781) );
  NAND2_X1 U12195 ( .A1(n9781), .A2(n14243), .ZN(n9793) );
  INV_X1 U12196 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14736) );
  NAND2_X1 U12197 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14932)
         );
  OAI21_X1 U12198 ( .B1(n14996), .B2(n14736), .A(n14932), .ZN(n9782) );
  AOI21_X1 U12199 ( .B1(n11322), .B2(n14219), .A(n9782), .ZN(n9792) );
  INV_X1 U12200 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9783) );
  MUX2_X1 U12201 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9783), .S(n11322), .Z(
        n9789) );
  NAND2_X1 U12202 ( .A1(n9784), .A2(n15118), .ZN(n9785) );
  NAND2_X1 U12203 ( .A1(n9786), .A2(n9785), .ZN(n14215) );
  INV_X1 U12204 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15121) );
  MUX2_X1 U12205 ( .A(n15121), .B(P1_REG1_REG_10__SCAN_IN), .S(n14220), .Z(
        n14214) );
  OR2_X1 U12206 ( .A1(n14215), .A2(n14214), .ZN(n14216) );
  NAND2_X1 U12207 ( .A1(n14220), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9787) );
  AND2_X1 U12208 ( .A1(n14216), .A2(n9787), .ZN(n9788) );
  NAND2_X1 U12209 ( .A1(n9788), .A2(n9789), .ZN(n9982) );
  OAI21_X1 U12210 ( .B1(n9789), .B2(n9788), .A(n9982), .ZN(n9790) );
  NAND2_X1 U12211 ( .A1(n9790), .A2(n14245), .ZN(n9791) );
  OAI211_X1 U12212 ( .C1(n9974), .C2(n9793), .A(n9792), .B(n9791), .ZN(
        P1_U3254) );
  OR2_X1 U12213 ( .A1(n13489), .A2(n9644), .ZN(n9794) );
  INV_X1 U12214 ( .A(n9840), .ZN(n9796) );
  NAND2_X1 U12215 ( .A1(n9797), .A2(n10053), .ZN(n9798) );
  NAND2_X1 U12216 ( .A1(n10023), .A2(n9798), .ZN(n9799) );
  NOR2_X1 U12217 ( .A1(n9847), .A2(n9799), .ZN(n10571) );
  OR2_X1 U12218 ( .A1(n13489), .A2(n10049), .ZN(n9800) );
  XNOR2_X1 U12219 ( .A(n9841), .B(n9840), .ZN(n9802) );
  AOI21_X1 U12220 ( .B1(n9802), .B2(n13822), .A(n9801), .ZN(n10575) );
  INV_X1 U12221 ( .A(n10575), .ZN(n9803) );
  AOI211_X1 U12222 ( .C1(n13905), .C2(n10572), .A(n10571), .B(n9803), .ZN(
        n10055) );
  AOI22_X1 U12223 ( .A1(n13899), .A2(n10053), .B1(n15188), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n9804) );
  OAI21_X1 U12224 ( .B1(n10055), .B2(n15188), .A(n9804), .ZN(P2_U3501) );
  INV_X1 U12225 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9811) );
  NOR3_X1 U12226 ( .A1(n9813), .A2(n9811), .A3(n15129), .ZN(n9809) );
  AOI21_X1 U12227 ( .B1(n9807), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9806), .ZN(
        n9818) );
  INV_X1 U12228 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10564) );
  NOR3_X1 U12229 ( .A1(n9818), .A2(n10564), .A3(n13556), .ZN(n9808) );
  NOR3_X1 U12230 ( .A1(n9809), .A2(n15155), .A3(n9808), .ZN(n9824) );
  AND2_X1 U12231 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9816) );
  INV_X1 U12232 ( .A(n9813), .ZN(n9810) );
  NAND3_X1 U12233 ( .A1(n9810), .A2(n9823), .A3(n9811), .ZN(n9814) );
  MUX2_X1 U12234 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9811), .S(n9912), .Z(n9812)
         );
  AOI21_X1 U12235 ( .B1(n9814), .B2(n9907), .A(n15129), .ZN(n9815) );
  AOI211_X1 U12236 ( .C1(n15154), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n9816), .B(
        n9815), .ZN(n9822) );
  NOR3_X1 U12237 ( .A1(n9818), .A2(n9912), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9820) );
  MUX2_X1 U12238 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10564), .S(n9912), .Z(n9817) );
  NAND2_X1 U12239 ( .A1(n9818), .A2(n9817), .ZN(n9911) );
  INV_X1 U12240 ( .A(n9911), .ZN(n9819) );
  OAI21_X1 U12241 ( .B1(n9820), .B2(n9819), .A(n15161), .ZN(n9821) );
  OAI211_X1 U12242 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9821), .ZN(
        P2_U3223) );
  INV_X1 U12243 ( .A(n9825), .ZN(n9826) );
  NAND2_X1 U12244 ( .A1(n9827), .A2(n9826), .ZN(n9925) );
  AND2_X1 U12245 ( .A1(n13488), .A2(n13687), .ZN(n9921) );
  XNOR2_X1 U12246 ( .A(n9920), .B(n9921), .ZN(n9924) );
  XNOR2_X1 U12247 ( .A(n9925), .B(n9924), .ZN(n9833) );
  NAND2_X1 U12248 ( .A1(n9829), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14891) );
  AOI22_X1 U12249 ( .A1(n13464), .A2(n9210), .B1(n13570), .B2(n13487), .ZN(
        n9844) );
  NAND2_X1 U12250 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U12251 ( .A1(n9631), .A2(n10684), .ZN(n9830) );
  OAI211_X1 U12252 ( .C1(n13447), .C2(n9844), .A(n13503), .B(n9830), .ZN(n9831) );
  AOI21_X1 U12253 ( .B1(n13449), .B2(n8535), .A(n9831), .ZN(n9832) );
  OAI21_X1 U12254 ( .B1(n9833), .B2(n13470), .A(n9832), .ZN(P2_U3190) );
  INV_X1 U12255 ( .A(n9834), .ZN(n9836) );
  OAI222_X1 U12256 ( .A1(n7368), .A2(P3_U3151), .B1(n11891), .B2(n9836), .C1(
        n9835), .C2(n11887), .ZN(P3_U3278) );
  OR2_X1 U12257 ( .A1(n9210), .A2(n10053), .ZN(n9837) );
  NAND2_X1 U12258 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  NAND2_X1 U12259 ( .A1(n9839), .A2(n9843), .ZN(n9938) );
  OAI21_X1 U12260 ( .B1(n9839), .B2(n9843), .A(n9938), .ZN(n10688) );
  INV_X1 U12261 ( .A(n10688), .ZN(n9848) );
  OR2_X1 U12262 ( .A1(n9210), .A2(n10568), .ZN(n9842) );
  INV_X1 U12263 ( .A(n9843), .ZN(n9942) );
  XNOR2_X1 U12264 ( .A(n9943), .B(n9942), .ZN(n9846) );
  INV_X1 U12265 ( .A(n9844), .ZN(n9845) );
  AOI21_X1 U12266 ( .B1(n9846), .B2(n13822), .A(n9845), .ZN(n10690) );
  OAI211_X1 U12267 ( .C1(n10057), .C2(n9847), .A(n10023), .B(n9940), .ZN(
        n10686) );
  OAI211_X1 U12268 ( .C1(n9848), .C2(n15182), .A(n10690), .B(n10686), .ZN(
        n10059) );
  OAI22_X1 U12269 ( .A1(n13912), .A2(n10057), .B1(n15190), .B2(n8537), .ZN(
        n9849) );
  AOI21_X1 U12270 ( .B1(n10059), .B2(n15190), .A(n9849), .ZN(n9850) );
  INV_X1 U12271 ( .A(n9850), .ZN(P2_U3502) );
  INV_X1 U12272 ( .A(n12404), .ZN(n12350) );
  NAND2_X1 U12273 ( .A1(n9855), .A2(n8598), .ZN(n9852) );
  NAND2_X1 U12274 ( .A1(n9716), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12275 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NAND2_X1 U12276 ( .A1(n9853), .A2(n9895), .ZN(n9858) );
  NAND2_X1 U12277 ( .A1(n9716), .A2(n6848), .ZN(n9854) );
  OAI211_X1 U12278 ( .C1(n9855), .C2(n9716), .A(n12253), .B(n9854), .ZN(n9857)
         );
  INV_X1 U12279 ( .A(n14162), .ZN(n14161) );
  NAND3_X1 U12280 ( .A1(n9491), .A2(n14161), .A3(n14700), .ZN(n9856) );
  NAND2_X1 U12281 ( .A1(n15002), .A2(n10039), .ZN(n9859) );
  OAI21_X1 U12282 ( .B1(n12350), .B2(n15053), .A(n9859), .ZN(n9860) );
  XNOR2_X1 U12283 ( .A(n9860), .B(n10786), .ZN(n9862) );
  INV_X2 U12284 ( .A(n12360), .ZN(n10120) );
  NOR2_X1 U12285 ( .A1(n12361), .A2(n15053), .ZN(n9861) );
  AOI21_X1 U12286 ( .B1(n10120), .B2(n15002), .A(n9861), .ZN(n9863) );
  NAND2_X1 U12287 ( .A1(n9862), .A2(n9863), .ZN(n10036) );
  INV_X1 U12288 ( .A(n9862), .ZN(n9865) );
  NAND2_X1 U12289 ( .A1(n9865), .A2(n9864), .ZN(n9866) );
  MUX2_X1 U12290 ( .A(n10786), .B(n9868), .S(n9867), .Z(n9869) );
  AOI21_X1 U12291 ( .B1(n9870), .B2(n9869), .A(n10038), .ZN(n9880) );
  NOR2_X1 U12292 ( .A1(n14927), .A2(n15053), .ZN(n9878) );
  INV_X1 U12293 ( .A(n15007), .ZN(n14525) );
  NOR2_X2 U12294 ( .A1(n14111), .A2(n14525), .ZN(n14923) );
  INV_X1 U12295 ( .A(n14923), .ZN(n9876) );
  INV_X1 U12296 ( .A(n15006), .ZN(n9875) );
  NAND2_X1 U12297 ( .A1(n10243), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U12298 ( .A1(n10201), .A2(n14527), .ZN(n15011) );
  INV_X1 U12299 ( .A(n15011), .ZN(n9874) );
  OAI22_X1 U12300 ( .A1(n9876), .A2(n9875), .B1(n9874), .B2(n14111), .ZN(n9877) );
  AOI211_X1 U12301 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10044), .A(n9878), .B(
        n9877), .ZN(n9879) );
  OAI21_X1 U12302 ( .B1(n9880), .B2(n14133), .A(n9879), .ZN(P1_U3222) );
  MUX2_X1 U12303 ( .A(n9482), .B(P1_REG1_REG_4__SCAN_IN), .S(n10228), .Z(n9881) );
  NAND3_X1 U12304 ( .A1(n14189), .A2(n9882), .A3(n9881), .ZN(n9883) );
  AND3_X1 U12305 ( .A1(n14245), .A2(n9884), .A3(n9883), .ZN(n9893) );
  INV_X1 U12306 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9891) );
  INV_X1 U12307 ( .A(n9885), .ZN(n9887) );
  MUX2_X1 U12308 ( .A(n10466), .B(P1_REG2_REG_4__SCAN_IN), .S(n10228), .Z(
        n9886) );
  NAND2_X1 U12309 ( .A1(n9887), .A2(n9886), .ZN(n9889) );
  OAI211_X1 U12310 ( .C1(n14190), .C2(n9889), .A(n14243), .B(n9888), .ZN(n9890) );
  NAND2_X1 U12311 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10637) );
  OAI211_X1 U12312 ( .C1(n9891), .C2(n14996), .A(n9890), .B(n10637), .ZN(n9892) );
  AOI211_X1 U12313 ( .C1(n14219), .C2(n10228), .A(n9893), .B(n9892), .ZN(n9897) );
  NAND2_X1 U12314 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14157) );
  MUX2_X1 U12315 ( .A(n9894), .B(n14157), .S(n12253), .Z(n9896) );
  OAI21_X1 U12316 ( .B1(n9491), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9895), .ZN(
        n14971) );
  NAND2_X1 U12317 ( .A1(n14971), .A2(n14164), .ZN(n14974) );
  OAI211_X1 U12318 ( .C1(n9896), .C2(n14700), .A(P1_U4016), .B(n14974), .ZN(
        n14181) );
  NAND2_X1 U12319 ( .A1(n9897), .A2(n14181), .ZN(P1_U3247) );
  INV_X1 U12320 ( .A(n11472), .ZN(n9903) );
  OAI222_X1 U12321 ( .A1(n13999), .A2(n6931), .B1(n14001), .B2(n9903), .C1(
        n15142), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12322 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12323 ( .A1(n9898), .A2(n10216), .ZN(n9899) );
  NAND2_X1 U12324 ( .A1(n9899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9900) );
  INV_X1 U12325 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U12326 ( .A1(n9900), .A2(n10215), .ZN(n10061) );
  OR2_X1 U12327 ( .A1(n9900), .A2(n10215), .ZN(n9901) );
  INV_X1 U12328 ( .A(n11473), .ZN(n10156) );
  OAI222_X1 U12329 ( .A1(P1_U3086), .A2(n10156), .B1(n14707), .B2(n9903), .C1(
        n9902), .C2(n14709), .ZN(P1_U3342) );
  INV_X1 U12330 ( .A(n12876), .ZN(n9906) );
  INV_X1 U12331 ( .A(SI_18_), .ZN(n9905) );
  OAI222_X1 U12332 ( .A1(P3_U3151), .A2(n9906), .B1(n12420), .B2(n9905), .C1(
        n13303), .C2(n9904), .ZN(P3_U3277) );
  OAI21_X1 U12333 ( .B1(n9912), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9907), .ZN(
        n9910) );
  INV_X1 U12334 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9908) );
  MUX2_X1 U12335 ( .A(n9908), .B(P2_REG2_REG_10__SCAN_IN), .S(n9994), .Z(n9909) );
  AOI211_X1 U12336 ( .C1(n9910), .C2(n9909), .A(n15129), .B(n9993), .ZN(n9919)
         );
  OAI21_X1 U12337 ( .B1(n9912), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9911), .ZN(
        n9914) );
  INV_X1 U12338 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10002) );
  MUX2_X1 U12339 ( .A(n10002), .B(P2_REG1_REG_10__SCAN_IN), .S(n9994), .Z(
        n9913) );
  NOR2_X1 U12340 ( .A1(n9914), .A2(n9913), .ZN(n10010) );
  AOI211_X1 U12341 ( .C1(n9914), .C2(n9913), .A(n13556), .B(n10010), .ZN(n9918) );
  INV_X1 U12342 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U12343 ( .A1(n15155), .A2(n9994), .ZN(n9915) );
  NAND2_X1 U12344 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10997)
         );
  OAI211_X1 U12345 ( .C1(n15127), .C2(n9916), .A(n9915), .B(n10997), .ZN(n9917) );
  OR3_X1 U12346 ( .A1(n9919), .A2(n9918), .A3(n9917), .ZN(P2_U3224) );
  INV_X1 U12347 ( .A(n9920), .ZN(n9923) );
  INV_X1 U12348 ( .A(n9921), .ZN(n9922) );
  OAI22_X1 U12349 ( .A1(n9925), .A2(n9924), .B1(n9923), .B2(n9922), .ZN(n9929)
         );
  XNOR2_X1 U12350 ( .A(n10644), .B(n13338), .ZN(n9927) );
  NAND2_X1 U12351 ( .A1(n13487), .A2(n13343), .ZN(n9926) );
  NAND2_X1 U12352 ( .A1(n9927), .A2(n9926), .ZN(n10066) );
  OAI21_X1 U12353 ( .B1(n9927), .B2(n9926), .A(n10066), .ZN(n9928) );
  AOI21_X1 U12354 ( .B1(n9929), .B2(n9928), .A(n10068), .ZN(n9936) );
  INV_X1 U12355 ( .A(n10644), .ZN(n10017) );
  NAND2_X1 U12356 ( .A1(n13464), .A2(n13488), .ZN(n9931) );
  NAND2_X1 U12357 ( .A1(n13570), .A2(n13486), .ZN(n9930) );
  NAND2_X1 U12358 ( .A1(n9931), .A2(n9930), .ZN(n9948) );
  NAND2_X1 U12359 ( .A1(n14885), .A2(n9948), .ZN(n9932) );
  OAI211_X1 U12360 ( .C1(n13452), .C2(n10017), .A(n9933), .B(n9932), .ZN(n9934) );
  AOI21_X1 U12361 ( .B1(n10643), .B2(n13449), .A(n9934), .ZN(n9935) );
  OAI21_X1 U12362 ( .B1(n9936), .B2(n13470), .A(n9935), .ZN(P2_U3202) );
  OR2_X1 U12363 ( .A1(n10684), .A2(n13488), .ZN(n9937) );
  NAND2_X1 U12364 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  INV_X1 U12365 ( .A(n10025), .ZN(n9947) );
  NAND2_X1 U12366 ( .A1(n9939), .A2(n9947), .ZN(n10022) );
  OAI21_X1 U12367 ( .B1(n9939), .B2(n9947), .A(n10022), .ZN(n10650) );
  AOI21_X1 U12368 ( .B1(n9940), .B2(n10644), .A(n13687), .ZN(n9941) );
  AND2_X1 U12369 ( .A1(n9941), .A2(n10024), .ZN(n10642) );
  NAND2_X1 U12370 ( .A1(n10684), .A2(n9944), .ZN(n9945) );
  XNOR2_X1 U12371 ( .A(n10026), .B(n9947), .ZN(n9950) );
  INV_X1 U12372 ( .A(n9948), .ZN(n9949) );
  OAI21_X1 U12373 ( .B1(n9950), .B2(n13795), .A(n9949), .ZN(n10647) );
  AOI211_X1 U12374 ( .C1(n13905), .C2(n10650), .A(n10642), .B(n10647), .ZN(
        n10020) );
  OAI22_X1 U12375 ( .A1(n13912), .A2(n10017), .B1(n15190), .B2(n9418), .ZN(
        n9951) );
  INV_X1 U12376 ( .A(n9951), .ZN(n9952) );
  OAI21_X1 U12377 ( .B1(n10020), .B2(n15188), .A(n9952), .ZN(P2_U3503) );
  INV_X1 U12378 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15337) );
  NAND2_X1 U12379 ( .A1(n12635), .A2(n12692), .ZN(n9953) );
  OAI21_X1 U12380 ( .B1(n12692), .B2(n15337), .A(n9953), .ZN(P3_U3501) );
  INV_X1 U12381 ( .A(n15053), .ZN(n9954) );
  NAND2_X1 U12382 ( .A1(n9955), .A2(n9954), .ZN(n12107) );
  NAND2_X1 U12383 ( .A1(n15002), .A2(n15053), .ZN(n12104) );
  NAND2_X1 U12384 ( .A1(n12107), .A2(n12104), .ZN(n15003) );
  NAND2_X1 U12385 ( .A1(n15003), .A2(n14998), .ZN(n9957) );
  NAND2_X1 U12386 ( .A1(n9955), .A2(n15053), .ZN(n9956) );
  NAND2_X2 U12387 ( .A1(n9958), .A2(n9716), .ZN(n12054) );
  XNOR2_X1 U12388 ( .A(n10195), .B(n12002), .ZN(n10519) );
  NOR2_X1 U12389 ( .A1(n15006), .A2(n14999), .ZN(n12108) );
  NAND2_X1 U12390 ( .A1(n12108), .A2(n12104), .ZN(n12109) );
  NAND2_X1 U12391 ( .A1(n12109), .A2(n12107), .ZN(n10198) );
  XNOR2_X1 U12392 ( .A(n12002), .B(n10198), .ZN(n10522) );
  INV_X1 U12393 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12394 ( .A1(n11974), .A2(n10133), .ZN(n9966) );
  NAND2_X1 U12395 ( .A1(n12059), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12396 ( .A1(n10484), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U12397 ( .A1(n10243), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9963) );
  OR2_X1 U12398 ( .A1(n10225), .A2(n14527), .ZN(n9968) );
  NAND2_X1 U12399 ( .A1(n15002), .A2(n15007), .ZN(n9967) );
  NAND2_X1 U12400 ( .A1(n9968), .A2(n9967), .ZN(n10514) );
  INV_X1 U12401 ( .A(n10514), .ZN(n9969) );
  AND2_X1 U12402 ( .A1(n14999), .A2(n15053), .ZN(n15001) );
  OAI211_X1 U12403 ( .C1(n15001), .C2(n10515), .A(n15016), .B(n10206), .ZN(
        n10513) );
  OAI211_X1 U12404 ( .C1(n10522), .C2(n14936), .A(n9969), .B(n10513), .ZN(
        n9970) );
  AOI21_X1 U12405 ( .B1(n15108), .B2(n10519), .A(n9970), .ZN(n10504) );
  NAND2_X1 U12406 ( .A1(n15123), .A2(n15062), .ZN(n14630) );
  AOI22_X1 U12407 ( .A1(n11847), .A2(n10045), .B1(n15120), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n9972) );
  OAI21_X1 U12408 ( .B1(n10504), .B2(n15120), .A(n9972), .ZN(P1_U3530) );
  INV_X1 U12409 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U12410 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9973), .S(n11467), .Z(
        n9976) );
  AOI21_X1 U12411 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n11322), .A(n9974), .ZN(
        n9975) );
  NAND2_X1 U12412 ( .A1(n9975), .A2(n9976), .ZN(n10079) );
  OAI21_X1 U12413 ( .B1(n9976), .B2(n9975), .A(n10079), .ZN(n9989) );
  OR2_X1 U12414 ( .A1(n11322), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U12415 ( .A1(n9982), .A2(n9980), .ZN(n9978) );
  INV_X1 U12416 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9977) );
  MUX2_X1 U12417 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9977), .S(n11467), .Z(
        n9979) );
  NAND2_X1 U12418 ( .A1(n9978), .A2(n9979), .ZN(n10084) );
  INV_X1 U12419 ( .A(n9979), .ZN(n9981) );
  NAND3_X1 U12420 ( .A1(n9982), .A2(n9981), .A3(n9980), .ZN(n9983) );
  AOI21_X1 U12421 ( .B1(n10084), .B2(n9983), .A(n14987), .ZN(n9988) );
  INV_X1 U12422 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n14039) );
  NOR2_X1 U12423 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14039), .ZN(n9984) );
  AOI21_X1 U12424 ( .B1(n14977), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9984), .ZN(
        n9985) );
  OAI21_X1 U12425 ( .B1(n9986), .B2(n14992), .A(n9985), .ZN(n9987) );
  AOI211_X1 U12426 ( .C1(n9989), .C2(n14243), .A(n9988), .B(n9987), .ZN(n9990)
         );
  INV_X1 U12427 ( .A(n9990), .ZN(P1_U3255) );
  OAI222_X1 U12428 ( .A1(n11891), .A2(n9992), .B1(n11887), .B2(n9991), .C1(
        P3_U3151), .C2(n6688), .ZN(P3_U3276) );
  INV_X1 U12429 ( .A(n9997), .ZN(n10000) );
  INV_X1 U12430 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9995) );
  MUX2_X1 U12431 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9995), .S(n10006), .Z(
        n9996) );
  INV_X1 U12432 ( .A(n9996), .ZN(n9999) );
  INV_X1 U12433 ( .A(n10176), .ZN(n9998) );
  AOI21_X1 U12434 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10013) );
  NAND2_X1 U12435 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11402)
         );
  OAI21_X1 U12436 ( .B1(n15143), .B2(n10173), .A(n11402), .ZN(n10001) );
  AOI21_X1 U12437 ( .B1(n15154), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10001), 
        .ZN(n10012) );
  INV_X1 U12438 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10168) );
  MUX2_X1 U12439 ( .A(n10168), .B(P2_REG1_REG_11__SCAN_IN), .S(n10006), .Z(
        n10005) );
  NOR2_X1 U12440 ( .A1(n10003), .A2(n10002), .ZN(n10008) );
  INV_X1 U12441 ( .A(n10008), .ZN(n10004) );
  NAND2_X1 U12442 ( .A1(n10005), .A2(n10004), .ZN(n10009) );
  MUX2_X1 U12443 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10168), .S(n10006), .Z(
        n10007) );
  OAI21_X1 U12444 ( .B1(n10010), .B2(n10008), .A(n10007), .ZN(n10167) );
  OAI211_X1 U12445 ( .C1(n10010), .C2(n10009), .A(n10167), .B(n15161), .ZN(
        n10011) );
  OAI211_X1 U12446 ( .C1(n10013), .C2(n15129), .A(n10012), .B(n10011), .ZN(
        P2_U3225) );
  INV_X1 U12447 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15395) );
  INV_X1 U12448 ( .A(n13020), .ZN(n12625) );
  NAND2_X1 U12449 ( .A1(n12625), .A2(n12692), .ZN(n10014) );
  OAI21_X1 U12450 ( .B1(n12692), .B2(n15395), .A(n10014), .ZN(P3_U3512) );
  INV_X1 U12451 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15442) );
  NAND2_X1 U12452 ( .A1(n13100), .A2(n12692), .ZN(n10015) );
  OAI21_X1 U12453 ( .B1(n12692), .B2(n15442), .A(n10015), .ZN(P3_U3506) );
  NAND2_X1 U12454 ( .A1(n15187), .A2(n15179), .ZN(n13974) );
  INV_X1 U12455 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10016) );
  OAI22_X1 U12456 ( .A1(n13974), .A2(n10017), .B1(n15187), .B2(n10016), .ZN(
        n10018) );
  INV_X1 U12457 ( .A(n10018), .ZN(n10019) );
  OAI21_X1 U12458 ( .B1(n10020), .B2(n15185), .A(n10019), .ZN(P2_U3442) );
  INV_X1 U12459 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10035) );
  OR2_X1 U12460 ( .A1(n10644), .A2(n13487), .ZN(n10021) );
  NAND2_X1 U12461 ( .A1(n10022), .A2(n10021), .ZN(n10093) );
  XNOR2_X1 U12462 ( .A(n10093), .B(n10099), .ZN(n10326) );
  AOI211_X1 U12463 ( .C1(n10319), .C2(n10024), .A(n13343), .B(n10096), .ZN(
        n10323) );
  AOI21_X1 U12464 ( .B1(n15179), .B2(n10319), .A(n10323), .ZN(n10033) );
  NAND2_X1 U12465 ( .A1(n10026), .A2(n10025), .ZN(n10029) );
  INV_X1 U12466 ( .A(n13487), .ZN(n10027) );
  NAND2_X1 U12467 ( .A1(n10644), .A2(n10027), .ZN(n10028) );
  XNOR2_X1 U12468 ( .A(n10100), .B(n10099), .ZN(n10032) );
  NAND2_X1 U12469 ( .A1(n13464), .A2(n13487), .ZN(n10031) );
  NAND2_X1 U12470 ( .A1(n13570), .A2(n13485), .ZN(n10030) );
  NAND2_X1 U12471 ( .A1(n10031), .A2(n10030), .ZN(n10073) );
  AOI21_X1 U12472 ( .B1(n10032), .B2(n13822), .A(n10073), .ZN(n10317) );
  OAI211_X1 U12473 ( .C1(n15182), .C2(n10326), .A(n10033), .B(n10317), .ZN(
        n13938) );
  NAND2_X1 U12474 ( .A1(n13938), .A2(n15187), .ZN(n10034) );
  OAI21_X1 U12475 ( .B1(n15187), .B2(n10035), .A(n10034), .ZN(P2_U3445) );
  INV_X1 U12476 ( .A(n10036), .ZN(n10037) );
  NAND2_X1 U12477 ( .A1(n12404), .A2(n10045), .ZN(n10040) );
  OAI21_X1 U12478 ( .B1(n10201), .B2(n12361), .A(n10040), .ZN(n10041) );
  XNOR2_X1 U12479 ( .A(n10041), .B(n12292), .ZN(n10115) );
  OAI22_X1 U12480 ( .A1(n12360), .A2(n10201), .B1(n10515), .B2(n12361), .ZN(
        n10116) );
  XNOR2_X1 U12481 ( .A(n10115), .B(n10116), .ZN(n10042) );
  AOI21_X1 U12482 ( .B1(n10043), .B2(n10042), .A(n6591), .ZN(n10048) );
  AOI22_X1 U12483 ( .A1(n10044), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14143), 
        .B2(n10514), .ZN(n10047) );
  NAND2_X1 U12484 ( .A1(n14131), .A2(n10045), .ZN(n10046) );
  OAI211_X1 U12485 ( .C1(n10048), .C2(n14133), .A(n10047), .B(n10046), .ZN(
        P1_U3237) );
  OAI22_X1 U12486 ( .A1(n13974), .A2(n10049), .B1(n15187), .B2(n8476), .ZN(
        n10050) );
  AOI21_X1 U12487 ( .B1(n15187), .B2(n10051), .A(n10050), .ZN(n10052) );
  INV_X1 U12488 ( .A(n10052), .ZN(P2_U3433) );
  INV_X1 U12489 ( .A(n13974), .ZN(n13965) );
  AOI22_X1 U12490 ( .A1(n13965), .A2(n10053), .B1(n15185), .B2(
        P2_REG0_REG_2__SCAN_IN), .ZN(n10054) );
  OAI21_X1 U12491 ( .B1(n10055), .B2(n15185), .A(n10054), .ZN(P2_U3436) );
  INV_X1 U12492 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10056) );
  OAI22_X1 U12493 ( .A1(n13974), .A2(n10057), .B1(n15187), .B2(n10056), .ZN(
        n10058) );
  AOI21_X1 U12494 ( .B1(n10059), .B2(n15187), .A(n10058), .ZN(n10060) );
  INV_X1 U12495 ( .A(n10060), .ZN(P2_U3439) );
  NAND2_X1 U12496 ( .A1(n10061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10062) );
  XNOR2_X1 U12497 ( .A(n10062), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11764) );
  INV_X1 U12498 ( .A(n11764), .ZN(n10972) );
  INV_X1 U12499 ( .A(n11763), .ZN(n10064) );
  OAI222_X1 U12500 ( .A1(P1_U3086), .A2(n10972), .B1(n14707), .B2(n10064), 
        .C1(n10063), .C2(n14709), .ZN(P1_U3341) );
  INV_X1 U12501 ( .A(n13524), .ZN(n11273) );
  OAI222_X1 U12502 ( .A1(n13999), .A2(n10065), .B1(n14001), .B2(n10064), .C1(
        n11273), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U12503 ( .A(n10066), .ZN(n10067) );
  XNOR2_X1 U12504 ( .A(n10319), .B(n13338), .ZN(n10070) );
  NAND2_X1 U12505 ( .A1(n13486), .A2(n13343), .ZN(n10069) );
  NAND2_X1 U12506 ( .A1(n10070), .A2(n10069), .ZN(n10138) );
  OAI21_X1 U12507 ( .B1(n10070), .B2(n10069), .A(n10138), .ZN(n10071) );
  AOI21_X1 U12508 ( .B1(n10072), .B2(n10071), .A(n10140), .ZN(n10078) );
  NAND2_X1 U12509 ( .A1(n14885), .A2(n10073), .ZN(n10075) );
  OAI211_X1 U12510 ( .C1(n14891), .C2(n10320), .A(n10075), .B(n10074), .ZN(
        n10076) );
  AOI21_X1 U12511 ( .B1(n10319), .B2(n9631), .A(n10076), .ZN(n10077) );
  OAI21_X1 U12512 ( .B1(n10078), .B2(n13470), .A(n10077), .ZN(P2_U3199) );
  OAI21_X1 U12513 ( .B1(n11467), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10079), 
        .ZN(n10081) );
  INV_X1 U12514 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10155) );
  MUX2_X1 U12515 ( .A(n10155), .B(P1_REG2_REG_13__SCAN_IN), .S(n11473), .Z(
        n10080) );
  NOR2_X1 U12516 ( .A1(n10081), .A2(n10080), .ZN(n10162) );
  AOI211_X1 U12517 ( .C1(n10081), .C2(n10080), .A(n14983), .B(n10162), .ZN(
        n10082) );
  INV_X1 U12518 ( .A(n10082), .ZN(n10091) );
  NAND2_X1 U12519 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14099)
         );
  OR2_X1 U12520 ( .A1(n11467), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10083) );
  INV_X1 U12521 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10085) );
  MUX2_X1 U12522 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10085), .S(n11473), .Z(
        n10086) );
  NAND2_X1 U12523 ( .A1(n10087), .A2(n10086), .ZN(n10150) );
  OAI211_X1 U12524 ( .C1(n10087), .C2(n10086), .A(n14245), .B(n10150), .ZN(
        n10088) );
  NAND2_X1 U12525 ( .A1(n14099), .A2(n10088), .ZN(n10089) );
  AOI21_X1 U12526 ( .B1(n14977), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10089), 
        .ZN(n10090) );
  OAI211_X1 U12527 ( .C1(n14992), .C2(n10156), .A(n10091), .B(n10090), .ZN(
        P1_U3256) );
  NAND2_X1 U12528 ( .A1(n10319), .A2(n13486), .ZN(n10092) );
  NAND2_X1 U12529 ( .A1(n10093), .A2(n10092), .ZN(n10095) );
  OR2_X1 U12530 ( .A1(n10319), .A2(n13486), .ZN(n10094) );
  NAND2_X1 U12531 ( .A1(n10095), .A2(n10094), .ZN(n10328) );
  XNOR2_X1 U12532 ( .A(n10328), .B(n10331), .ZN(n10316) );
  INV_X1 U12533 ( .A(n10096), .ZN(n10098) );
  INV_X1 U12534 ( .A(n10334), .ZN(n10311) );
  INV_X1 U12535 ( .A(n10338), .ZN(n10097) );
  AOI211_X1 U12536 ( .C1(n10334), .C2(n10098), .A(n13687), .B(n10097), .ZN(
        n10313) );
  AOI21_X1 U12537 ( .B1(n15179), .B2(n10334), .A(n10313), .ZN(n10106) );
  INV_X1 U12538 ( .A(n13486), .ZN(n10101) );
  NAND2_X1 U12539 ( .A1(n10319), .A2(n10101), .ZN(n10102) );
  XNOR2_X1 U12540 ( .A(n10332), .B(n10331), .ZN(n10105) );
  NAND2_X1 U12541 ( .A1(n13464), .A2(n13486), .ZN(n10104) );
  NAND2_X1 U12542 ( .A1(n13570), .A2(n13484), .ZN(n10103) );
  NAND2_X1 U12543 ( .A1(n10104), .A2(n10103), .ZN(n10142) );
  AOI21_X1 U12544 ( .B1(n10105), .B2(n13822), .A(n10142), .ZN(n10307) );
  OAI211_X1 U12545 ( .C1(n15182), .C2(n10316), .A(n10106), .B(n10307), .ZN(
        n10108) );
  NAND2_X1 U12546 ( .A1(n10108), .A2(n15190), .ZN(n10107) );
  OAI21_X1 U12547 ( .B1(n15190), .B2(n9424), .A(n10107), .ZN(P2_U3505) );
  INV_X1 U12548 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U12549 ( .A1(n10108), .A2(n15187), .ZN(n10109) );
  OAI21_X1 U12550 ( .B1(n15187), .B2(n10110), .A(n10109), .ZN(P2_U3448) );
  NAND2_X1 U12551 ( .A1(n10111), .A2(n12041), .ZN(n10113) );
  NAND2_X1 U12552 ( .A1(n12022), .A2(n14184), .ZN(n10112) );
  OAI211_X1 U12553 ( .C1(n12054), .C2(n10114), .A(n10113), .B(n10112), .ZN(
        n15061) );
  INV_X1 U12554 ( .A(n15061), .ZN(n10224) );
  INV_X1 U12555 ( .A(n10115), .ZN(n10118) );
  INV_X1 U12556 ( .A(n10116), .ZN(n10117) );
  OAI22_X1 U12557 ( .A1(n10225), .A2(n12361), .B1(n10224), .B2(n12350), .ZN(
        n10119) );
  XNOR2_X1 U12558 ( .A(n10119), .B(n12292), .ZN(n10628) );
  INV_X1 U12559 ( .A(n10225), .ZN(n14154) );
  AND2_X1 U12560 ( .A1(n10039), .A2(n15061), .ZN(n10121) );
  AOI21_X1 U12561 ( .B1(n10120), .B2(n14154), .A(n10121), .ZN(n10630) );
  XNOR2_X1 U12562 ( .A(n10628), .B(n10630), .ZN(n10122) );
  OAI211_X1 U12563 ( .C1(n10123), .C2(n10122), .A(n10631), .B(n14930), .ZN(
        n10137) );
  INV_X1 U12564 ( .A(n10124), .ZN(n10125) );
  NAND2_X1 U12565 ( .A1(n10126), .A2(n10125), .ZN(n10127) );
  NAND2_X1 U12566 ( .A1(n10127), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14935) );
  AND2_X1 U12567 ( .A1(n14113), .A2(n10133), .ZN(n10135) );
  NAND2_X1 U12568 ( .A1(n12059), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10132) );
  AND2_X1 U12569 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10236) );
  NOR2_X1 U12570 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10128) );
  NOR2_X1 U12571 ( .A1(n10236), .A2(n10128), .ZN(n10639) );
  NAND2_X1 U12572 ( .A1(n11974), .A2(n10639), .ZN(n10131) );
  NAND2_X1 U12573 ( .A1(n12061), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U12574 ( .A1(n10484), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10129) );
  OAI22_X1 U12575 ( .A1(n14120), .A2(n12122), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10133), .ZN(n10134) );
  AOI211_X1 U12576 ( .C1(n14923), .C2(n14155), .A(n10135), .B(n10134), .ZN(
        n10136) );
  OAI211_X1 U12577 ( .C1(n10224), .C2(n14927), .A(n10137), .B(n10136), .ZN(
        P1_U3218) );
  INV_X1 U12578 ( .A(n10138), .ZN(n10139) );
  NAND2_X1 U12579 ( .A1(n13485), .A2(n13343), .ZN(n10260) );
  XNOR2_X1 U12580 ( .A(n10261), .B(n10260), .ZN(n10263) );
  XNOR2_X1 U12581 ( .A(n6584), .B(n10263), .ZN(n10147) );
  INV_X1 U12582 ( .A(n10141), .ZN(n10310) );
  NAND2_X1 U12583 ( .A1(n14885), .A2(n10142), .ZN(n10144) );
  OAI211_X1 U12584 ( .C1(n14891), .C2(n10310), .A(n10144), .B(n10143), .ZN(
        n10145) );
  AOI21_X1 U12585 ( .B1(n10334), .B2(n9631), .A(n10145), .ZN(n10146) );
  OAI21_X1 U12586 ( .B1(n10147), .B2(n13470), .A(n10146), .ZN(P2_U3211) );
  INV_X1 U12587 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10148) );
  MUX2_X1 U12588 ( .A(n10148), .B(P1_REG1_REG_14__SCAN_IN), .S(n11764), .Z(
        n10153) );
  NAND2_X1 U12589 ( .A1(n11473), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U12590 ( .A1(n10150), .A2(n10149), .ZN(n10152) );
  INV_X1 U12591 ( .A(n10979), .ZN(n10151) );
  AOI21_X1 U12592 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10166) );
  INV_X1 U12593 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10154) );
  MUX2_X1 U12594 ( .A(n10154), .B(P1_REG2_REG_14__SCAN_IN), .S(n11764), .Z(
        n10158) );
  NOR2_X1 U12595 ( .A1(n10156), .A2(n10155), .ZN(n10160) );
  INV_X1 U12596 ( .A(n10160), .ZN(n10157) );
  NAND2_X1 U12597 ( .A1(n10158), .A2(n10157), .ZN(n10161) );
  MUX2_X1 U12598 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10154), .S(n11764), .Z(
        n10159) );
  OAI21_X1 U12599 ( .B1(n10162), .B2(n10160), .A(n10159), .ZN(n10971) );
  OAI211_X1 U12600 ( .C1(n10162), .C2(n10161), .A(n10971), .B(n14243), .ZN(
        n10165) );
  INV_X1 U12601 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14713) );
  NAND2_X1 U12602 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14902)
         );
  OAI21_X1 U12603 ( .B1(n14996), .B2(n14713), .A(n14902), .ZN(n10163) );
  AOI21_X1 U12604 ( .B1(n11764), .B2(n14219), .A(n10163), .ZN(n10164) );
  OAI211_X1 U12605 ( .C1(n10166), .C2(n14987), .A(n10165), .B(n10164), .ZN(
        P1_U3257) );
  OAI21_X1 U12606 ( .B1(n10168), .B2(n10173), .A(n10167), .ZN(n10171) );
  INV_X1 U12607 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10169) );
  MUX2_X1 U12608 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10169), .S(n11270), .Z(
        n10170) );
  NOR2_X1 U12609 ( .A1(n10171), .A2(n10170), .ZN(n11269) );
  AOI21_X1 U12610 ( .B1(n10171), .B2(n10170), .A(n11269), .ZN(n10183) );
  INV_X1 U12611 ( .A(n11270), .ZN(n10181) );
  INV_X1 U12612 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U12613 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n10172)
         );
  OAI21_X1 U12614 ( .B1(n15127), .B2(n14954), .A(n10172), .ZN(n10180) );
  NAND2_X1 U12615 ( .A1(n10173), .A2(n9995), .ZN(n10174) );
  INV_X1 U12616 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13843) );
  MUX2_X1 U12617 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n13843), .S(n11270), .Z(
        n10175) );
  INV_X1 U12618 ( .A(n11259), .ZN(n10178) );
  NAND3_X1 U12619 ( .A1(n10176), .A2(n10175), .A3(n10174), .ZN(n10177) );
  AOI21_X1 U12620 ( .B1(n10178), .B2(n10177), .A(n15129), .ZN(n10179) );
  AOI211_X1 U12621 ( .C1(n15155), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10182) );
  OAI21_X1 U12622 ( .B1(n10183), .B2(n13556), .A(n10182), .ZN(P2_U3226) );
  INV_X1 U12623 ( .A(n10184), .ZN(n10186) );
  OAI222_X1 U12624 ( .A1(n11891), .A2(n10186), .B1(n12420), .B2(n10185), .C1(
        P3_U3151), .C2(n10417), .ZN(P3_U3275) );
  NOR2_X1 U12625 ( .A1(n10188), .A2(n10187), .ZN(n10205) );
  NAND2_X1 U12626 ( .A1(n10205), .A2(n10203), .ZN(n10192) );
  INV_X1 U12627 ( .A(n10189), .ZN(n10190) );
  INV_X1 U12628 ( .A(n10193), .ZN(n10194) );
  NAND2_X1 U12629 ( .A1(n10195), .A2(n12002), .ZN(n10197) );
  NAND2_X1 U12630 ( .A1(n10201), .A2(n10515), .ZN(n10196) );
  NAND2_X1 U12631 ( .A1(n10225), .A2(n15061), .ZN(n12118) );
  NAND2_X1 U12632 ( .A1(n10224), .A2(n14154), .ZN(n12119) );
  XNOR2_X1 U12633 ( .A(n10223), .B(n12116), .ZN(n15065) );
  NAND2_X1 U12634 ( .A1(n10198), .A2(n12113), .ZN(n10199) );
  NAND2_X1 U12635 ( .A1(n10199), .A2(n12115), .ZN(n10248) );
  INV_X1 U12636 ( .A(n12116), .ZN(n12001) );
  XNOR2_X1 U12637 ( .A(n10248), .B(n12001), .ZN(n10200) );
  OAI222_X1 U12638 ( .A1(n14527), .A2(n12122), .B1(n14525), .B2(n10201), .C1(
        n10200), .C2(n14936), .ZN(n15059) );
  NAND2_X1 U12639 ( .A1(n12075), .A2(n12077), .ZN(n12091) );
  INV_X1 U12640 ( .A(n14544), .ZN(n15013) );
  AOI22_X1 U12641 ( .A1(n15022), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15013), 
        .B2(n10133), .ZN(n10210) );
  AND2_X1 U12642 ( .A1(n10203), .A2(n14320), .ZN(n10204) );
  NAND2_X1 U12643 ( .A1(n10206), .A2(n15061), .ZN(n10207) );
  NAND2_X1 U12644 ( .A1(n10207), .A2(n15016), .ZN(n10208) );
  NOR2_X1 U12645 ( .A1(n10463), .A2(n10208), .ZN(n15060) );
  NAND2_X1 U12646 ( .A1(n15018), .A2(n15060), .ZN(n10209) );
  OAI211_X1 U12647 ( .C1(n15012), .C2(n10224), .A(n10210), .B(n10209), .ZN(
        n10211) );
  AOI21_X1 U12648 ( .B1(n14541), .B2(n15059), .A(n10211), .ZN(n10212) );
  OAI21_X1 U12649 ( .B1(n14520), .B2(n15065), .A(n10212), .ZN(P1_U3290) );
  INV_X1 U12650 ( .A(n15156), .ZN(n11275) );
  INV_X1 U12651 ( .A(n11787), .ZN(n10221) );
  OAI222_X1 U12652 ( .A1(P2_U3088), .A2(n11275), .B1(n14001), .B2(n10221), 
        .C1(n10213), .C2(n13999), .ZN(P2_U3312) );
  INV_X1 U12653 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10214) );
  NAND3_X1 U12654 ( .A1(n10216), .A2(n10215), .A3(n10214), .ZN(n10217) );
  OAI21_X1 U12655 ( .B1(n10218), .B2(n10217), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10219) );
  XNOR2_X1 U12656 ( .A(n10219), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11788) );
  INV_X1 U12657 ( .A(n11788), .ZN(n14991) );
  OAI222_X1 U12658 ( .A1(P1_U3086), .A2(n14991), .B1(n14707), .B2(n10221), 
        .C1(n10220), .C2(n14709), .ZN(P1_U3340) );
  INV_X1 U12659 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15323) );
  NAND2_X1 U12660 ( .A1(n12527), .A2(n12692), .ZN(n10222) );
  OAI21_X1 U12661 ( .B1(n12692), .B2(n15323), .A(n10222), .ZN(P3_U3515) );
  NAND2_X1 U12662 ( .A1(n10225), .A2(n10224), .ZN(n10226) );
  NAND2_X1 U12663 ( .A1(n10227), .A2(n6429), .ZN(n10230) );
  AOI22_X1 U12664 ( .A1(n12023), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12022), 
        .B2(n10228), .ZN(n10229) );
  AND2_X2 U12665 ( .A1(n10230), .A2(n10229), .ZN(n15073) );
  INV_X1 U12666 ( .A(n15073), .ZN(n12123) );
  OR2_X1 U12667 ( .A1(n14153), .A2(n12123), .ZN(n10459) );
  INV_X1 U12668 ( .A(n10459), .ZN(n10231) );
  NAND2_X1 U12669 ( .A1(n12123), .A2(n14153), .ZN(n10458) );
  NAND2_X1 U12670 ( .A1(n10232), .A2(n6429), .ZN(n10235) );
  AOI22_X1 U12671 ( .A1(n12023), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12022), 
        .B2(n10233), .ZN(n10234) );
  NAND2_X1 U12672 ( .A1(n10236), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10282) );
  OAI21_X1 U12673 ( .B1(n10236), .B2(P1_REG3_REG_5__SCAN_IN), .A(n10282), .ZN(
        n14068) );
  INV_X1 U12674 ( .A(n14068), .ZN(n10237) );
  NAND2_X1 U12675 ( .A1(n11974), .A2(n10237), .ZN(n10241) );
  NAND2_X1 U12676 ( .A1(n12059), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U12677 ( .A1(n12060), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10239) );
  NAND2_X1 U12678 ( .A1(n10243), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10238) );
  OAI21_X1 U12679 ( .B1(n6581), .B2(n10251), .A(n10269), .ZN(n10452) );
  INV_X1 U12680 ( .A(n10452), .ZN(n10259) );
  NAND2_X1 U12681 ( .A1(n12105), .A2(n14433), .ZN(n12070) );
  NOR2_X1 U12682 ( .A1(n15022), .A2(n12070), .ZN(n15019) );
  INV_X1 U12683 ( .A(n15019), .ZN(n11542) );
  XNOR2_X1 U12684 ( .A(n10282), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U12685 ( .A1(n11974), .A2(n10798), .ZN(n10247) );
  NAND2_X1 U12686 ( .A1(n12059), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U12687 ( .A1(n12061), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U12688 ( .A1(n10484), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10244) );
  NAND4_X1 U12689 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n14151) );
  INV_X1 U12690 ( .A(n14151), .ZN(n10473) );
  OAI22_X1 U12691 ( .A1(n10473), .A2(n14527), .B1(n12122), .B2(n14525), .ZN(
        n14066) );
  NOR2_X1 U12692 ( .A1(n14153), .A2(n15073), .ZN(n10249) );
  NAND2_X1 U12693 ( .A1(n14153), .A2(n15073), .ZN(n10250) );
  NAND2_X1 U12694 ( .A1(n10252), .A2(n10251), .ZN(n10253) );
  AOI21_X1 U12695 ( .B1(n10278), .B2(n10253), .A(n14936), .ZN(n10254) );
  AOI211_X1 U12696 ( .C1(n15068), .C2(n10452), .A(n14066), .B(n10254), .ZN(
        n10449) );
  MUX2_X1 U12697 ( .A(n9518), .B(n10449), .S(n14541), .Z(n10258) );
  INV_X1 U12698 ( .A(n10273), .ZN(n10255) );
  AOI211_X1 U12699 ( .C1(n14067), .C2(n10462), .A(n14640), .B(n10255), .ZN(
        n10451) );
  OAI22_X1 U12700 ( .A1(n15012), .A2(n6833), .B1(n14544), .B2(n14068), .ZN(
        n10256) );
  AOI21_X1 U12701 ( .B1(n10451), .B2(n15018), .A(n10256), .ZN(n10257) );
  OAI211_X1 U12702 ( .C1(n10259), .C2(n11542), .A(n10258), .B(n10257), .ZN(
        P1_U3288) );
  INV_X1 U12703 ( .A(n10260), .ZN(n10262) );
  XNOR2_X1 U12704 ( .A(n15178), .B(n13338), .ZN(n10432) );
  NAND2_X1 U12705 ( .A1(n13484), .A2(n13343), .ZN(n10431) );
  XNOR2_X1 U12706 ( .A(n10432), .B(n10431), .ZN(n10433) );
  XNOR2_X1 U12707 ( .A(n10434), .B(n10433), .ZN(n10267) );
  AOI22_X1 U12708 ( .A1(n13570), .A2(n13483), .B1(n13464), .B2(n13485), .ZN(
        n10335) );
  NAND2_X1 U12709 ( .A1(n13449), .A2(n10339), .ZN(n10264) );
  NAND2_X1 U12710 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15125) );
  OAI211_X1 U12711 ( .C1(n13447), .C2(n10335), .A(n10264), .B(n15125), .ZN(
        n10265) );
  AOI21_X1 U12712 ( .B1(n15178), .B2(n9631), .A(n10265), .ZN(n10266) );
  OAI21_X1 U12713 ( .B1(n10267), .B2(n13470), .A(n10266), .ZN(P2_U3185) );
  OR2_X1 U12714 ( .A1(n14067), .A2(n14152), .ZN(n10268) );
  AOI22_X1 U12715 ( .A1(n12023), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12022), 
        .B2(n14205), .ZN(n10271) );
  XNOR2_X1 U12716 ( .A(n12132), .B(n14151), .ZN(n12005) );
  OAI21_X1 U12717 ( .B1(n10272), .B2(n10279), .A(n10492), .ZN(n10511) );
  NAND2_X1 U12718 ( .A1(n10273), .A2(n12132), .ZN(n10274) );
  NAND2_X1 U12719 ( .A1(n10274), .A2(n15016), .ZN(n10275) );
  NOR2_X1 U12720 ( .A1(n10495), .A2(n10275), .ZN(n10505) );
  INV_X1 U12721 ( .A(n14152), .ZN(n10276) );
  NAND2_X1 U12722 ( .A1(n14067), .A2(n10276), .ZN(n10277) );
  NAND2_X1 U12723 ( .A1(n10278), .A2(n10277), .ZN(n10472) );
  XNOR2_X1 U12724 ( .A(n10472), .B(n10279), .ZN(n10288) );
  INV_X1 U12725 ( .A(n10282), .ZN(n10280) );
  AOI21_X1 U12726 ( .B1(n10280), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12727 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n10281) );
  NOR2_X1 U12728 ( .A1(n10282), .A2(n10281), .ZN(n10482) );
  OR2_X1 U12729 ( .A1(n10283), .A2(n10482), .ZN(n10957) );
  INV_X1 U12730 ( .A(n10957), .ZN(n10496) );
  NAND2_X1 U12731 ( .A1(n11974), .A2(n10496), .ZN(n10287) );
  NAND2_X1 U12732 ( .A1(n12059), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U12733 ( .A1(n10484), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U12734 ( .A1(n12061), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10284) );
  NAND4_X1 U12735 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n14150) );
  AOI22_X1 U12736 ( .A1(n14509), .A2(n14150), .B1(n15007), .B2(n14152), .ZN(
        n10796) );
  OAI21_X1 U12737 ( .B1(n10288), .B2(n14936), .A(n10796), .ZN(n10508) );
  AOI211_X1 U12738 ( .C1(n15108), .C2(n10511), .A(n10505), .B(n10508), .ZN(
        n10295) );
  NAND2_X1 U12739 ( .A1(n14655), .A2(n15062), .ZN(n14683) );
  INV_X1 U12740 ( .A(n12132), .ZN(n10801) );
  INV_X1 U12741 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10291) );
  OAI22_X1 U12742 ( .A1(n14683), .A2(n10801), .B1(n14655), .B2(n10291), .ZN(
        n10292) );
  INV_X1 U12743 ( .A(n10292), .ZN(n10293) );
  OAI21_X1 U12744 ( .B1(n10295), .B2(n15109), .A(n10293), .ZN(P1_U3477) );
  AOI22_X1 U12745 ( .A1(n11847), .A2(n12132), .B1(n15120), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n10294) );
  OAI21_X1 U12746 ( .B1(n10295), .B2(n15120), .A(n10294), .ZN(P1_U3534) );
  INV_X1 U12747 ( .A(n12020), .ZN(n10299) );
  OAI222_X1 U12748 ( .A1(P2_U3088), .A2(n11511), .B1(n14001), .B2(n10299), 
        .C1(n10296), .C2(n13999), .ZN(P2_U3311) );
  NAND2_X1 U12749 ( .A1(n10297), .A2(n6570), .ZN(n10529) );
  NAND2_X1 U12750 ( .A1(n10529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10298) );
  XNOR2_X1 U12751 ( .A(n10298), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12021) );
  INV_X1 U12752 ( .A(n12021), .ZN(n11373) );
  OAI222_X1 U12753 ( .A1(P1_U3086), .A2(n11373), .B1(n14707), .B2(n10299), 
        .C1(n15443), .C2(n14709), .ZN(P1_U3339) );
  INV_X1 U12754 ( .A(n15170), .ZN(n10302) );
  NAND3_X1 U12755 ( .A1(n10302), .A2(n10301), .A3(n10300), .ZN(n10303) );
  NAND2_X1 U12756 ( .A1(n10305), .A2(n10304), .ZN(n10535) );
  NAND2_X1 U12757 ( .A1(n9664), .A2(n10535), .ZN(n10306) );
  MUX2_X1 U12758 ( .A(n9403), .B(n10307), .S(n13844), .Z(n10315) );
  INV_X1 U12759 ( .A(n10308), .ZN(n10309) );
  OAI22_X1 U12760 ( .A1(n13816), .A2(n10311), .B1(n13841), .B2(n10310), .ZN(
        n10312) );
  AOI21_X1 U12761 ( .B1(n10313), .B2(n13850), .A(n10312), .ZN(n10314) );
  OAI211_X1 U12762 ( .C1(n13835), .C2(n10316), .A(n10315), .B(n10314), .ZN(
        P2_U3259) );
  MUX2_X1 U12763 ( .A(n10318), .B(n10317), .S(n13844), .Z(n10325) );
  INV_X1 U12764 ( .A(n10319), .ZN(n10321) );
  OAI22_X1 U12765 ( .A1(n13816), .A2(n10321), .B1(n13841), .B2(n10320), .ZN(
        n10322) );
  AOI21_X1 U12766 ( .B1(n10323), .B2(n13850), .A(n10322), .ZN(n10324) );
  OAI211_X1 U12767 ( .C1(n13835), .C2(n10326), .A(n10325), .B(n10324), .ZN(
        P2_U3260) );
  INV_X1 U12768 ( .A(n10331), .ZN(n10327) );
  NAND2_X1 U12769 ( .A1(n10328), .A2(n10327), .ZN(n10330) );
  OR2_X1 U12770 ( .A1(n10334), .A2(n13485), .ZN(n10329) );
  NAND2_X1 U12771 ( .A1(n10330), .A2(n10329), .ZN(n10348) );
  XOR2_X1 U12772 ( .A(n10347), .B(n10348), .Z(n15183) );
  XOR2_X1 U12773 ( .A(n10347), .B(n10353), .Z(n10337) );
  INV_X1 U12774 ( .A(n10335), .ZN(n10336) );
  AOI21_X1 U12775 ( .B1(n10337), .B2(n13822), .A(n10336), .ZN(n15181) );
  MUX2_X1 U12776 ( .A(n9545), .B(n15181), .S(n13844), .Z(n10344) );
  AOI211_X1 U12777 ( .C1(n15178), .C2(n10338), .A(n13343), .B(n7126), .ZN(
        n15177) );
  INV_X1 U12778 ( .A(n15178), .ZN(n10341) );
  INV_X1 U12779 ( .A(n10339), .ZN(n10340) );
  OAI22_X1 U12780 ( .A1(n13816), .A2(n10341), .B1(n13841), .B2(n10340), .ZN(
        n10342) );
  AOI21_X1 U12781 ( .B1(n15177), .B2(n13850), .A(n10342), .ZN(n10343) );
  OAI211_X1 U12782 ( .C1(n13835), .C2(n15183), .A(n10344), .B(n10343), .ZN(
        P2_U3258) );
  INV_X1 U12783 ( .A(n10345), .ZN(n10346) );
  INV_X1 U12784 ( .A(SI_21_), .ZN(n15391) );
  OAI222_X1 U12785 ( .A1(n10416), .A2(P3_U3151), .B1(n11891), .B2(n10346), 
        .C1(n15391), .C2(n11887), .ZN(P3_U3274) );
  OR2_X1 U12786 ( .A1(n15178), .A2(n13484), .ZN(n10349) );
  INV_X1 U12787 ( .A(n10357), .ZN(n10351) );
  OAI21_X1 U12788 ( .B1(n6580), .B2(n10351), .A(n10547), .ZN(n10372) );
  AND2_X1 U12789 ( .A1(n15178), .A2(n10354), .ZN(n10352) );
  OR2_X1 U12790 ( .A1(n15178), .A2(n10354), .ZN(n10355) );
  XOR2_X1 U12791 ( .A(n10357), .B(n10550), .Z(n10359) );
  AOI22_X1 U12792 ( .A1(n13464), .A2(n13484), .B1(n13570), .B2(n13482), .ZN(
        n10442) );
  INV_X1 U12793 ( .A(n10442), .ZN(n10358) );
  AOI21_X1 U12794 ( .B1(n10359), .B2(n13822), .A(n10358), .ZN(n10371) );
  MUX2_X1 U12795 ( .A(n9546), .B(n10371), .S(n13844), .Z(n10365) );
  INV_X1 U12796 ( .A(n10559), .ZN(n10360) );
  AOI211_X1 U12797 ( .C1(n10552), .C2(n10361), .A(n13687), .B(n10360), .ZN(
        n10369) );
  INV_X1 U12798 ( .A(n10439), .ZN(n10362) );
  OAI22_X1 U12799 ( .A1(n7125), .A2(n13816), .B1(n13841), .B2(n10362), .ZN(
        n10363) );
  AOI21_X1 U12800 ( .B1(n10369), .B2(n13850), .A(n10363), .ZN(n10364) );
  OAI211_X1 U12801 ( .C1(n13835), .C2(n10372), .A(n10365), .B(n10364), .ZN(
        P2_U3257) );
  INV_X1 U12802 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U12803 ( .A1(n10366), .A2(n15111), .ZN(n10367) );
  OAI21_X1 U12804 ( .B1(n15111), .B2(n10368), .A(n10367), .ZN(P1_U3459) );
  AOI21_X1 U12805 ( .B1(n15179), .B2(n10552), .A(n10369), .ZN(n10370) );
  OAI211_X1 U12806 ( .C1(n10372), .C2(n15182), .A(n10371), .B(n10370), .ZN(
        n10408) );
  NAND2_X1 U12807 ( .A1(n10408), .A2(n15190), .ZN(n10373) );
  OAI21_X1 U12808 ( .B1(n15190), .B2(n10374), .A(n10373), .ZN(P2_U3507) );
  INV_X1 U12809 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10375) );
  NAND2_X1 U12810 ( .A1(n11883), .A2(n10375), .ZN(n10377) );
  NAND2_X1 U12811 ( .A1(n11032), .A2(n11301), .ZN(n10376) );
  NOR2_X1 U12812 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n10381) );
  NOR4_X1 U12813 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n10380) );
  NOR4_X1 U12814 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n10379) );
  NOR4_X1 U12815 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U12816 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10387) );
  NOR4_X1 U12817 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n10385) );
  NOR4_X1 U12818 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n10384) );
  NOR4_X1 U12819 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10383) );
  NOR4_X1 U12820 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n10382) );
  NAND4_X1 U12821 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10386) );
  OAI21_X1 U12822 ( .B1(n10387), .B2(n10386), .A(n11883), .ZN(n10611) );
  NAND3_X1 U12823 ( .A1(n10620), .A2(n10610), .A3(n10611), .ZN(n10589) );
  NAND2_X1 U12824 ( .A1(n10615), .A2(n12878), .ZN(n10597) );
  OR2_X1 U12825 ( .A1(n10597), .A2(n10414), .ZN(n10587) );
  INV_X1 U12826 ( .A(n10587), .ZN(n10388) );
  NAND2_X1 U12827 ( .A1(n10589), .A2(n10388), .ZN(n10395) );
  NAND2_X1 U12828 ( .A1(n13296), .A2(n10611), .ZN(n10389) );
  NAND2_X1 U12829 ( .A1(n10416), .A2(n10417), .ZN(n10390) );
  XNOR2_X1 U12830 ( .A(n10615), .B(n10390), .ZN(n10392) );
  NAND2_X1 U12831 ( .A1(n10416), .A2(n6688), .ZN(n10391) );
  NAND2_X1 U12832 ( .A1(n10392), .A2(n10391), .ZN(n10766) );
  NAND2_X1 U12833 ( .A1(n10591), .A2(n10766), .ZN(n10393) );
  NAND4_X1 U12834 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10652), .ZN(
        n10396) );
  NAND2_X1 U12835 ( .A1(n10396), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10398) );
  NAND2_X1 U12836 ( .A1(n11070), .A2(n10764), .ZN(n10401) );
  NAND2_X1 U12837 ( .A1(n10589), .A2(n10592), .ZN(n10397) );
  NAND2_X1 U12838 ( .A1(n10398), .A2(n10397), .ZN(n10714) );
  NOR2_X1 U12839 ( .A1(n10714), .A2(n11882), .ZN(n10586) );
  NAND2_X1 U12840 ( .A1(n10766), .A2(n15281), .ZN(n10598) );
  OAI22_X1 U12841 ( .A1(n10589), .A2(n10587), .B1(n10591), .B2(n10598), .ZN(
        n10399) );
  INV_X1 U12842 ( .A(n15232), .ZN(n15242) );
  NAND2_X1 U12843 ( .A1(n10591), .A2(n15242), .ZN(n10400) );
  INV_X1 U12844 ( .A(n10401), .ZN(n10403) );
  NAND2_X1 U12845 ( .A1(n11076), .A2(n11118), .ZN(n10402) );
  NAND2_X1 U12846 ( .A1(n10403), .A2(n15215), .ZN(n10404) );
  OAI22_X1 U12847 ( .A1(n10626), .A2(n12652), .B1(n12666), .B2(n7715), .ZN(
        n10405) );
  AOI21_X1 U12848 ( .B1(n12644), .B2(n10600), .A(n10405), .ZN(n10406) );
  OAI21_X1 U12849 ( .B1(n10586), .B2(n10407), .A(n10406), .ZN(P3_U3172) );
  INV_X1 U12850 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U12851 ( .A1(n10408), .A2(n15187), .ZN(n10409) );
  OAI21_X1 U12852 ( .B1(n15187), .B2(n10410), .A(n10409), .ZN(P2_U3454) );
  INV_X1 U12853 ( .A(n13213), .ZN(n10412) );
  OAI22_X1 U12854 ( .A1(n10712), .A2(n12666), .B1(n12659), .B2(n10412), .ZN(
        n10413) );
  AOI21_X1 U12855 ( .B1(n12672), .B2(n7714), .A(n10413), .ZN(n10430) );
  NAND2_X1 U12856 ( .A1(n10416), .A2(n12878), .ZN(n10418) );
  NAND2_X1 U12857 ( .A1(n10418), .A2(n10417), .ZN(n10419) );
  XNOR2_X1 U12858 ( .A(n10859), .B(n7714), .ZN(n10421) );
  NAND2_X1 U12859 ( .A1(n10421), .A2(n7715), .ZN(n10577) );
  INV_X2 U12860 ( .A(n10859), .ZN(n12503) );
  NAND3_X1 U12861 ( .A1(n12503), .A2(n12693), .A3(n7714), .ZN(n10422) );
  NAND2_X1 U12862 ( .A1(n12503), .A2(n13212), .ZN(n10423) );
  NAND2_X1 U12863 ( .A1(n10424), .A2(n10423), .ZN(n10425) );
  NAND3_X1 U12864 ( .A1(n10769), .A2(n10859), .A3(n13219), .ZN(n10426) );
  OAI211_X1 U12865 ( .C1(n10427), .C2(n13212), .A(n10578), .B(n10426), .ZN(
        n10428) );
  NAND2_X1 U12866 ( .A1(n10428), .A2(n12644), .ZN(n10429) );
  OAI211_X1 U12867 ( .C1(n10586), .C2(n11624), .A(n10430), .B(n10429), .ZN(
        P3_U3162) );
  XNOR2_X1 U12868 ( .A(n10552), .B(n13338), .ZN(n10436) );
  NAND2_X1 U12869 ( .A1(n13483), .A2(n13343), .ZN(n10435) );
  NOR2_X1 U12870 ( .A1(n10436), .A2(n10435), .ZN(n10720) );
  NAND2_X1 U12871 ( .A1(n10436), .A2(n10435), .ZN(n10721) );
  INV_X1 U12872 ( .A(n10721), .ZN(n10437) );
  NOR2_X1 U12873 ( .A1(n10720), .A2(n10437), .ZN(n10438) );
  XNOR2_X1 U12874 ( .A(n10722), .B(n10438), .ZN(n10445) );
  NAND2_X1 U12875 ( .A1(n13449), .A2(n10439), .ZN(n10441) );
  OAI211_X1 U12876 ( .C1(n13447), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10443) );
  AOI21_X1 U12877 ( .B1(n10552), .B2(n9631), .A(n10443), .ZN(n10444) );
  OAI21_X1 U12878 ( .B1(n10445), .B2(n13470), .A(n10444), .ZN(P2_U3193) );
  INV_X1 U12879 ( .A(n10446), .ZN(n10448) );
  OAI22_X1 U12880 ( .A1(n10615), .A2(P3_U3151), .B1(SI_22_), .B2(n11887), .ZN(
        n10447) );
  AOI21_X1 U12881 ( .B1(n10448), .B2(n10606), .A(n10447), .ZN(P3_U3273) );
  INV_X1 U12882 ( .A(n15064), .ZN(n15098) );
  INV_X1 U12883 ( .A(n10449), .ZN(n10450) );
  AOI211_X1 U12884 ( .C1(n15098), .C2(n10452), .A(n10451), .B(n10450), .ZN(
        n10457) );
  INV_X1 U12885 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10453) );
  OAI22_X1 U12886 ( .A1(n14683), .A2(n6833), .B1(n14655), .B2(n10453), .ZN(
        n10454) );
  INV_X1 U12887 ( .A(n10454), .ZN(n10455) );
  OAI21_X1 U12888 ( .B1(n10457), .B2(n15109), .A(n10455), .ZN(P1_U3474) );
  AOI22_X1 U12889 ( .A1(n11847), .A2(n14067), .B1(n15120), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n10456) );
  OAI21_X1 U12890 ( .B1(n10457), .B2(n15120), .A(n10456), .ZN(P1_U3533) );
  NAND2_X1 U12891 ( .A1(n10459), .A2(n10458), .ZN(n12007) );
  XNOR2_X1 U12892 ( .A(n10460), .B(n12007), .ZN(n15075) );
  NOR2_X1 U12893 ( .A1(n15022), .A2(n14936), .ZN(n14518) );
  XNOR2_X1 U12894 ( .A(n10461), .B(n12007), .ZN(n15078) );
  OAI211_X1 U12895 ( .C1(n10463), .C2(n15073), .A(n15016), .B(n10462), .ZN(
        n15071) );
  AOI22_X1 U12896 ( .A1(n14546), .A2(n12123), .B1(n10639), .B2(n15013), .ZN(
        n10468) );
  NAND2_X1 U12897 ( .A1(n14154), .A2(n15007), .ZN(n10465) );
  NAND2_X1 U12898 ( .A1(n14509), .A2(n14152), .ZN(n10464) );
  AND2_X1 U12899 ( .A1(n10465), .A2(n10464), .ZN(n15070) );
  MUX2_X1 U12900 ( .A(n15070), .B(n10466), .S(n15022), .Z(n10467) );
  OAI211_X1 U12901 ( .C1(n15071), .C2(n14537), .A(n10468), .B(n10467), .ZN(
        n10469) );
  AOI21_X1 U12902 ( .B1(n14518), .B2(n15078), .A(n10469), .ZN(n10470) );
  OAI21_X1 U12903 ( .B1(n14520), .B2(n15075), .A(n10470), .ZN(P1_U3289) );
  OR2_X1 U12904 ( .A1(n12132), .A2(n10473), .ZN(n10471) );
  NAND2_X1 U12905 ( .A1(n10472), .A2(n10471), .ZN(n10475) );
  NAND2_X1 U12906 ( .A1(n12132), .A2(n10473), .ZN(n10474) );
  NAND2_X1 U12907 ( .A1(n10475), .A2(n10474), .ZN(n10756) );
  NAND2_X1 U12908 ( .A1(n10476), .A2(n6429), .ZN(n10479) );
  AOI22_X1 U12909 ( .A1(n12023), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12022), 
        .B2(n10477), .ZN(n10478) );
  NAND2_X1 U12910 ( .A1(n10479), .A2(n10478), .ZN(n12135) );
  INV_X1 U12911 ( .A(n14150), .ZN(n10758) );
  XNOR2_X1 U12912 ( .A(n12135), .B(n10758), .ZN(n12009) );
  INV_X1 U12913 ( .A(n12009), .ZN(n10480) );
  XNOR2_X1 U12914 ( .A(n10756), .B(n10480), .ZN(n10481) );
  AND2_X1 U12915 ( .A1(n10481), .A2(n15079), .ZN(n15085) );
  NAND2_X1 U12916 ( .A1(n10482), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10749) );
  OR2_X1 U12917 ( .A1(n10482), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10483) );
  AND2_X1 U12918 ( .A1(n10749), .A2(n10483), .ZN(n11067) );
  NAND2_X1 U12919 ( .A1(n11974), .A2(n11067), .ZN(n10488) );
  NAND2_X1 U12920 ( .A1(n12059), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10487) );
  NAND2_X1 U12921 ( .A1(n10484), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U12922 ( .A1(n12061), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U12923 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n14149) );
  INV_X1 U12924 ( .A(n14149), .ZN(n10874) );
  NAND2_X1 U12925 ( .A1(n14151), .A2(n15007), .ZN(n10489) );
  OAI21_X1 U12926 ( .B1(n10874), .B2(n14527), .A(n10489), .ZN(n15081) );
  NOR2_X1 U12927 ( .A1(n15085), .A2(n15081), .ZN(n10490) );
  MUX2_X1 U12928 ( .A(n9523), .B(n10490), .S(n14541), .Z(n10500) );
  OR2_X1 U12929 ( .A1(n12132), .A2(n14151), .ZN(n10491) );
  NAND2_X1 U12930 ( .A1(n10492), .A2(n10491), .ZN(n10493) );
  NAND2_X1 U12931 ( .A1(n10493), .A2(n12009), .ZN(n10738) );
  OAI21_X1 U12932 ( .B1(n10493), .B2(n12009), .A(n10738), .ZN(n15087) );
  INV_X1 U12933 ( .A(n12135), .ZN(n10494) );
  OAI211_X1 U12934 ( .C1(n10495), .C2(n10494), .A(n15016), .B(n10744), .ZN(
        n15084) );
  AOI22_X1 U12935 ( .A1(n14546), .A2(n12135), .B1(n10496), .B2(n15013), .ZN(
        n10497) );
  OAI21_X1 U12936 ( .B1(n14537), .B2(n15084), .A(n10497), .ZN(n10498) );
  AOI21_X1 U12937 ( .B1(n15087), .B2(n14548), .A(n10498), .ZN(n10499) );
  NAND2_X1 U12938 ( .A1(n10500), .A2(n10499), .ZN(P1_U3286) );
  INV_X1 U12939 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10501) );
  OAI22_X1 U12940 ( .A1(n14683), .A2(n10515), .B1(n15111), .B2(n10501), .ZN(
        n10502) );
  INV_X1 U12941 ( .A(n10502), .ZN(n10503) );
  OAI21_X1 U12942 ( .B1(n10504), .B2(n15109), .A(n10503), .ZN(P1_U3465) );
  INV_X1 U12943 ( .A(n10505), .ZN(n10507) );
  AOI22_X1 U12944 ( .A1(n14546), .A2(n12132), .B1(n10798), .B2(n15013), .ZN(
        n10506) );
  OAI21_X1 U12945 ( .B1(n14537), .B2(n10507), .A(n10506), .ZN(n10510) );
  MUX2_X1 U12946 ( .A(n10508), .B(P1_REG2_REG_6__SCAN_IN), .S(n15022), .Z(
        n10509) );
  AOI211_X1 U12947 ( .C1(n14548), .C2(n10511), .A(n10510), .B(n10509), .ZN(
        n10512) );
  INV_X1 U12948 ( .A(n10512), .ZN(P1_U3287) );
  INV_X1 U12949 ( .A(n14518), .ZN(n14441) );
  INV_X1 U12950 ( .A(n10513), .ZN(n10518) );
  MUX2_X1 U12951 ( .A(n10514), .B(P1_REG2_REG_2__SCAN_IN), .S(n15022), .Z(
        n10517) );
  INV_X1 U12952 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14171) );
  OAI22_X1 U12953 ( .A1(n15012), .A2(n10515), .B1(n14171), .B2(n14544), .ZN(
        n10516) );
  AOI211_X1 U12954 ( .C1(n10518), .C2(n15018), .A(n10517), .B(n10516), .ZN(
        n10521) );
  NAND2_X1 U12955 ( .A1(n14548), .A2(n10519), .ZN(n10520) );
  OAI211_X1 U12956 ( .C1(n10522), .C2(n14441), .A(n10521), .B(n10520), .ZN(
        P1_U3291) );
  INV_X1 U12957 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10523) );
  OAI22_X1 U12958 ( .A1(n15022), .A2(n10524), .B1(n10523), .B2(n14544), .ZN(
        n10526) );
  AND2_X1 U12959 ( .A1(n15018), .A2(n15016), .ZN(n14354) );
  INV_X1 U12960 ( .A(n14354), .ZN(n14516) );
  AOI21_X1 U12961 ( .B1(n14516), .B2(n15012), .A(n14999), .ZN(n10525) );
  AOI211_X1 U12962 ( .C1(n15022), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10526), .B(
        n10525), .ZN(n10528) );
  OAI21_X1 U12963 ( .B1(n14518), .B2(n14548), .A(n12003), .ZN(n10527) );
  NAND2_X1 U12964 ( .A1(n10528), .A2(n10527), .ZN(P1_U3293) );
  OAI21_X1 U12965 ( .B1(n10529), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10530) );
  MUX2_X1 U12966 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10530), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10531) );
  INV_X1 U12967 ( .A(n9371), .ZN(n10812) );
  INV_X1 U12968 ( .A(n11992), .ZN(n11835) );
  INV_X1 U12969 ( .A(n11991), .ZN(n10533) );
  OAI222_X1 U12970 ( .A1(P1_U3086), .A2(n11835), .B1(n14707), .B2(n10533), 
        .C1(n10532), .C2(n14709), .ZN(P1_U3338) );
  OAI222_X1 U12971 ( .A1(n13999), .A2(n10534), .B1(n14001), .B2(n10533), .C1(
        n13537), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U12972 ( .A(n10535), .ZN(n10536) );
  NAND2_X1 U12973 ( .A1(n13844), .A2(n10536), .ZN(n13725) );
  INV_X1 U12974 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10537) );
  OAI22_X1 U12975 ( .A1(n6430), .A2(n10538), .B1(n10537), .B2(n13841), .ZN(
        n10539) );
  AOI21_X1 U12976 ( .B1(n6430), .B2(P2_REG2_REG_0__SCAN_IN), .A(n10539), .ZN(
        n10544) );
  OAI21_X1 U12977 ( .B1(n13766), .B2(n10540), .A(n13816), .ZN(n10542) );
  NAND2_X1 U12978 ( .A1(n10542), .A2(n10541), .ZN(n10543) );
  OAI211_X1 U12979 ( .C1(n13725), .C2(n10545), .A(n10544), .B(n10543), .ZN(
        P2_U3265) );
  NAND2_X1 U12980 ( .A1(n10552), .A2(n13483), .ZN(n10546) );
  OAI21_X1 U12981 ( .B1(n10549), .B2(n10554), .A(n10702), .ZN(n10669) );
  INV_X1 U12982 ( .A(n13483), .ZN(n10551) );
  NAND2_X1 U12983 ( .A1(n10552), .A2(n10551), .ZN(n10553) );
  AOI21_X1 U12984 ( .B1(n10555), .B2(n10554), .A(n13795), .ZN(n10558) );
  NAND2_X1 U12985 ( .A1(n13464), .A2(n13483), .ZN(n10557) );
  NAND2_X1 U12986 ( .A1(n13570), .A2(n13481), .ZN(n10556) );
  NAND2_X1 U12987 ( .A1(n10557), .A2(n10556), .ZN(n10727) );
  AOI21_X1 U12988 ( .B1(n10558), .B2(n10692), .A(n10727), .ZN(n10672) );
  NAND2_X1 U12989 ( .A1(n10723), .A2(n10559), .ZN(n10560) );
  NAND2_X1 U12990 ( .A1(n10560), .A2(n10023), .ZN(n10561) );
  NOR2_X1 U12991 ( .A1(n6434), .A2(n10561), .ZN(n10666) );
  AOI21_X1 U12992 ( .B1(n15179), .B2(n10723), .A(n10666), .ZN(n10562) );
  OAI211_X1 U12993 ( .C1(n10669), .C2(n15182), .A(n10672), .B(n10562), .ZN(
        n10565) );
  NAND2_X1 U12994 ( .A1(n10565), .A2(n15190), .ZN(n10563) );
  OAI21_X1 U12995 ( .B1(n15190), .B2(n10564), .A(n10563), .ZN(P2_U3508) );
  INV_X1 U12996 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U12997 ( .A1(n10565), .A2(n15187), .ZN(n10566) );
  OAI21_X1 U12998 ( .B1(n15187), .B2(n10567), .A(n10566), .ZN(P2_U3457) );
  INV_X1 U12999 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13492) );
  OAI22_X1 U13000 ( .A1(n13844), .A2(n9398), .B1(n13492), .B2(n13841), .ZN(
        n10570) );
  NOR2_X1 U13001 ( .A1(n13816), .A2(n10568), .ZN(n10569) );
  AOI211_X1 U13002 ( .C1(n10571), .C2(n13850), .A(n10570), .B(n10569), .ZN(
        n10574) );
  NAND2_X1 U13003 ( .A1(n13848), .A2(n10572), .ZN(n10573) );
  OAI211_X1 U13004 ( .C1(n6430), .C2(n10575), .A(n10574), .B(n10573), .ZN(
        P2_U3263) );
  INV_X1 U13005 ( .A(n10576), .ZN(n10894) );
  XNOR2_X1 U13006 ( .A(n10894), .B(n10859), .ZN(n10706) );
  XNOR2_X1 U13007 ( .A(n10706), .B(n13214), .ZN(n10580) );
  NAND2_X1 U13008 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  OAI21_X1 U13009 ( .B1(n10580), .B2(n10579), .A(n10711), .ZN(n10581) );
  NAND2_X1 U13010 ( .A1(n10581), .A2(n12644), .ZN(n10584) );
  INV_X1 U13011 ( .A(n12691), .ZN(n10868) );
  OAI22_X1 U13012 ( .A1(n7715), .A2(n12659), .B1(n12666), .B2(n10868), .ZN(
        n10582) );
  AOI21_X1 U13013 ( .B1(n10894), .B2(n12672), .A(n10582), .ZN(n10583) );
  OAI211_X1 U13014 ( .C1(n10586), .C2(n10585), .A(n10584), .B(n10583), .ZN(
        P3_U3177) );
  INV_X1 U13015 ( .A(n10766), .ZN(n10588) );
  OAI22_X1 U13016 ( .A1(n10589), .A2(n10588), .B1(n10591), .B2(n10587), .ZN(
        n10590) );
  NAND2_X1 U13017 ( .A1(n10590), .A2(n11070), .ZN(n10595) );
  INV_X1 U13018 ( .A(n10591), .ZN(n10593) );
  NAND2_X1 U13019 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  NAND2_X1 U13020 ( .A1(n10598), .A2(n14854), .ZN(n10599) );
  NAND2_X1 U13021 ( .A1(n10600), .A2(n10599), .ZN(n10602) );
  NAND2_X1 U13022 ( .A1(n12693), .A2(n15215), .ZN(n10601) );
  NAND2_X1 U13023 ( .A1(n10602), .A2(n10601), .ZN(n10661) );
  INV_X1 U13024 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10603) );
  NOR2_X1 U13025 ( .A1(n15293), .A2(n10603), .ZN(n10604) );
  AOI21_X1 U13026 ( .B1(n15293), .B2(n10661), .A(n10604), .ZN(n10605) );
  OAI21_X1 U13027 ( .B1(n10626), .B2(n13294), .A(n10605), .ZN(P3_U3390) );
  NAND2_X1 U13028 ( .A1(n10607), .A2(n10606), .ZN(n10608) );
  OAI211_X1 U13029 ( .C1(n10609), .C2(n11887), .A(n10608), .B(n11071), .ZN(
        P3_U3272) );
  XNOR2_X1 U13030 ( .A(n13296), .B(n10610), .ZN(n10613) );
  AND2_X1 U13031 ( .A1(n10611), .A2(n11070), .ZN(n10612) );
  AND2_X1 U13032 ( .A1(n10617), .A2(n6688), .ZN(n10614) );
  NAND2_X1 U13033 ( .A1(n10615), .A2(n10614), .ZN(n10767) );
  NAND2_X1 U13034 ( .A1(n10616), .A2(n10767), .ZN(n10654) );
  AND2_X1 U13035 ( .A1(n10652), .A2(n10654), .ZN(n10622) );
  OAI22_X1 U13036 ( .A1(n15281), .A2(n10617), .B1(n12878), .B2(n10777), .ZN(
        n10619) );
  AOI21_X1 U13037 ( .B1(n10619), .B2(n10618), .A(n11074), .ZN(n10621) );
  MUX2_X1 U13038 ( .A(n10622), .B(n10621), .S(n10620), .Z(n10623) );
  NOR2_X1 U13039 ( .A1(n15308), .A2(n11084), .ZN(n10624) );
  AOI21_X1 U13040 ( .B1(n15308), .B2(n10661), .A(n10624), .ZN(n10625) );
  OAI21_X1 U13041 ( .B1(n10626), .B2(n13210), .A(n10625), .ZN(P3_U3459) );
  OAI22_X1 U13042 ( .A1(n15073), .A2(n12350), .B1(n12122), .B2(n12361), .ZN(
        n10627) );
  XOR2_X1 U13043 ( .A(n12292), .B(n10627), .Z(n10635) );
  INV_X1 U13044 ( .A(n10628), .ZN(n10629) );
  OAI22_X1 U13045 ( .A1(n12122), .A2(n12360), .B1(n15073), .B2(n12361), .ZN(
        n10632) );
  OAI21_X1 U13046 ( .B1(n10635), .B2(n10634), .A(n10782), .ZN(n10636) );
  NAND2_X1 U13047 ( .A1(n10636), .A2(n14930), .ZN(n10641) );
  OAI21_X1 U13048 ( .B1(n14111), .B2(n15070), .A(n10637), .ZN(n10638) );
  AOI21_X1 U13049 ( .B1(n14113), .B2(n10639), .A(n10638), .ZN(n10640) );
  OAI211_X1 U13050 ( .C1(n15073), .C2(n14927), .A(n10641), .B(n10640), .ZN(
        P1_U3230) );
  INV_X1 U13051 ( .A(n10642), .ZN(n10646) );
  INV_X1 U13052 ( .A(n13841), .ZN(n13828) );
  AOI22_X1 U13053 ( .A1(n13846), .A2(n10644), .B1(n13828), .B2(n10643), .ZN(
        n10645) );
  OAI21_X1 U13054 ( .B1(n13766), .B2(n10646), .A(n10645), .ZN(n10649) );
  MUX2_X1 U13055 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10647), .S(n13844), .Z(
        n10648) );
  AOI211_X1 U13056 ( .C1(n13848), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10651) );
  INV_X1 U13057 ( .A(n10651), .ZN(P2_U3261) );
  INV_X1 U13058 ( .A(n10652), .ZN(n10653) );
  NOR2_X1 U13059 ( .A1(n13296), .A2(n10653), .ZN(n10655) );
  MUX2_X1 U13060 ( .A(n13296), .B(n10655), .S(n10654), .Z(n10656) );
  NAND2_X1 U13061 ( .A1(n10657), .A2(n10656), .ZN(n10659) );
  OR2_X1 U13062 ( .A1(n10659), .A2(n15232), .ZN(n10917) );
  NAND2_X1 U13063 ( .A1(n13107), .A2(n10660), .ZN(n10663) );
  AOI22_X1 U13064 ( .A1(n15248), .A2(n10661), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15244), .ZN(n10662) );
  OAI211_X1 U13065 ( .C1(n11085), .C2(n15248), .A(n10663), .B(n10662), .ZN(
        P3_U3233) );
  INV_X1 U13066 ( .A(n10731), .ZN(n10664) );
  OAI22_X1 U13067 ( .A1(n13844), .A2(n9811), .B1(n10664), .B2(n13841), .ZN(
        n10665) );
  AOI21_X1 U13068 ( .B1(n10723), .B2(n13846), .A(n10665), .ZN(n10668) );
  NAND2_X1 U13069 ( .A1(n10666), .A2(n13850), .ZN(n10667) );
  OAI211_X1 U13070 ( .C1(n10669), .C2(n13835), .A(n10668), .B(n10667), .ZN(
        n10670) );
  INV_X1 U13071 ( .A(n10670), .ZN(n10671) );
  OAI21_X1 U13072 ( .B1(n6430), .B2(n10672), .A(n10671), .ZN(P2_U3256) );
  NAND2_X1 U13073 ( .A1(n12680), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10673) );
  OAI21_X1 U13074 ( .B1(n12919), .B2(n12680), .A(n10673), .ZN(P3_U3519) );
  INV_X1 U13075 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10674) );
  OAI22_X1 U13076 ( .A1(n13844), .A2(n10675), .B1(n10674), .B2(n13841), .ZN(
        n10676) );
  AOI21_X1 U13077 ( .B1(n13846), .B2(n9644), .A(n10676), .ZN(n10677) );
  OAI21_X1 U13078 ( .B1(n13766), .B2(n10678), .A(n10677), .ZN(n10679) );
  AOI21_X1 U13079 ( .B1(n13848), .B2(n10680), .A(n10679), .ZN(n10681) );
  OAI21_X1 U13080 ( .B1(n6430), .B2(n10682), .A(n10681), .ZN(P2_U3264) );
  OAI22_X1 U13081 ( .A1(n13844), .A2(n6885), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n13841), .ZN(n10683) );
  AOI21_X1 U13082 ( .B1(n13846), .B2(n10684), .A(n10683), .ZN(n10685) );
  OAI21_X1 U13083 ( .B1(n13766), .B2(n10686), .A(n10685), .ZN(n10687) );
  AOI21_X1 U13084 ( .B1(n13848), .B2(n10688), .A(n10687), .ZN(n10689) );
  OAI21_X1 U13085 ( .B1(n6430), .B2(n10690), .A(n10689), .ZN(P2_U3262) );
  INV_X1 U13086 ( .A(n13482), .ZN(n10694) );
  OR2_X1 U13087 ( .A1(n10723), .A2(n10694), .ZN(n10691) );
  NAND2_X1 U13088 ( .A1(n10692), .A2(n10691), .ZN(n10693) );
  NAND2_X1 U13089 ( .A1(n10693), .A2(n10924), .ZN(n10932) );
  OAI211_X1 U13090 ( .C1(n10924), .C2(n10693), .A(n10932), .B(n13822), .ZN(
        n10696) );
  INV_X1 U13091 ( .A(n13480), .ZN(n11343) );
  OAI22_X1 U13092 ( .A1(n11343), .A2(n13455), .B1(n13640), .B2(n10694), .ZN(
        n10996) );
  INV_X1 U13093 ( .A(n10996), .ZN(n10695) );
  NAND2_X1 U13094 ( .A1(n10696), .A2(n10695), .ZN(n10802) );
  INV_X1 U13095 ( .A(n10802), .ZN(n10705) );
  INV_X1 U13096 ( .A(n6434), .ZN(n10699) );
  INV_X1 U13097 ( .A(n11010), .ZN(n10807) );
  INV_X1 U13098 ( .A(n10938), .ZN(n10698) );
  AOI211_X1 U13099 ( .C1(n11010), .C2(n10699), .A(n9680), .B(n10698), .ZN(
        n10803) );
  NOR2_X1 U13100 ( .A1(n10807), .A2(n13816), .ZN(n10701) );
  OAI22_X1 U13101 ( .A1(n13844), .A2(n9908), .B1(n10999), .B2(n13841), .ZN(
        n10700) );
  AOI211_X1 U13102 ( .C1(n10803), .C2(n13850), .A(n10701), .B(n10700), .ZN(
        n10704) );
  XNOR2_X1 U13103 ( .A(n10926), .B(n10924), .ZN(n10804) );
  NAND2_X1 U13104 ( .A1(n10804), .A2(n13848), .ZN(n10703) );
  OAI211_X1 U13105 ( .C1(n10705), .C2(n6430), .A(n10704), .B(n10703), .ZN(
        P2_U3255) );
  NAND2_X1 U13106 ( .A1(n10706), .A2(n10712), .ZN(n10708) );
  INV_X1 U13107 ( .A(n10707), .ZN(n10911) );
  XNOR2_X1 U13108 ( .A(n10859), .B(n10911), .ZN(n10855) );
  XNOR2_X1 U13109 ( .A(n10855), .B(n12691), .ZN(n10709) );
  AOI21_X1 U13110 ( .B1(n10711), .B2(n10708), .A(n10709), .ZN(n10719) );
  AND2_X1 U13111 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  NAND2_X1 U13112 ( .A1(n10858), .A2(n12644), .ZN(n10718) );
  INV_X1 U13113 ( .A(n12690), .ZN(n11019) );
  OAI22_X1 U13114 ( .A1(n10712), .A2(n12659), .B1(n12666), .B2(n11019), .ZN(
        n10716) );
  MUX2_X1 U13115 ( .A(n12656), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n10715) );
  AOI211_X1 U13116 ( .C1(n12672), .C2(n10911), .A(n10716), .B(n10715), .ZN(
        n10717) );
  OAI21_X1 U13117 ( .B1(n10719), .B2(n10718), .A(n10717), .ZN(P3_U3158) );
  INV_X1 U13118 ( .A(n10723), .ZN(n10734) );
  XNOR2_X1 U13119 ( .A(n10723), .B(n9828), .ZN(n11004) );
  NAND2_X1 U13120 ( .A1(n13482), .A2(n13343), .ZN(n11002) );
  XNOR2_X1 U13121 ( .A(n11004), .B(n11002), .ZN(n10724) );
  OAI21_X1 U13122 ( .B1(n10725), .B2(n10724), .A(n11003), .ZN(n10726) );
  NAND2_X1 U13123 ( .A1(n10726), .A2(n14883), .ZN(n10733) );
  NAND2_X1 U13124 ( .A1(n14885), .A2(n10727), .ZN(n10728) );
  OAI21_X1 U13125 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10729), .A(n10728), .ZN(
        n10730) );
  AOI21_X1 U13126 ( .B1(n10731), .B2(n13449), .A(n10730), .ZN(n10732) );
  OAI211_X1 U13127 ( .C1(n10734), .C2(n13452), .A(n10733), .B(n10732), .ZN(
        P2_U3203) );
  NAND2_X1 U13128 ( .A1(n12680), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10735) );
  OAI21_X1 U13129 ( .B1(n12454), .B2(n12680), .A(n10735), .ZN(P3_U3521) );
  NAND2_X1 U13130 ( .A1(n12680), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10736) );
  OAI21_X1 U13131 ( .B1(n12907), .B2(n12680), .A(n10736), .ZN(P3_U3520) );
  OR2_X1 U13132 ( .A1(n12135), .A2(n14150), .ZN(n10737) );
  NAND2_X1 U13133 ( .A1(n10738), .A2(n10737), .ZN(n10743) );
  NAND2_X1 U13134 ( .A1(n10739), .A2(n6429), .ZN(n10742) );
  AOI22_X1 U13135 ( .A1(n12023), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12022), 
        .B2(n10740), .ZN(n10741) );
  NAND2_X1 U13136 ( .A1(n10742), .A2(n10741), .ZN(n12139) );
  XNOR2_X1 U13137 ( .A(n12139), .B(n10874), .ZN(n12010) );
  OAI21_X1 U13138 ( .B1(n10743), .B2(n12010), .A(n10838), .ZN(n15093) );
  INV_X1 U13139 ( .A(n10744), .ZN(n10746) );
  INV_X1 U13140 ( .A(n12139), .ZN(n10745) );
  OAI211_X1 U13141 ( .C1(n10746), .C2(n10745), .A(n15016), .B(n10881), .ZN(
        n15090) );
  AOI22_X1 U13142 ( .A1(n14546), .A2(n12139), .B1(n15013), .B2(n11067), .ZN(
        n10747) );
  OAI21_X1 U13143 ( .B1(n15090), .B2(n14537), .A(n10747), .ZN(n10760) );
  INV_X1 U13144 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13145 ( .A1(n10749), .A2(n10748), .ZN(n10750) );
  AND2_X1 U13146 ( .A1(n10828), .A2(n10750), .ZN(n11757) );
  NAND2_X1 U13147 ( .A1(n11974), .A2(n11757), .ZN(n10754) );
  NAND2_X1 U13148 ( .A1(n12059), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13149 ( .A1(n12060), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U13150 ( .A1(n12061), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10751) );
  NAND4_X1 U13151 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n14909) );
  AND2_X1 U13152 ( .A1(n12135), .A2(n10758), .ZN(n10755) );
  OAI22_X1 U13153 ( .A1(n10756), .A2(n10755), .B1(n10758), .B2(n12135), .ZN(
        n10817) );
  INV_X1 U13154 ( .A(n12010), .ZN(n10816) );
  XNOR2_X1 U13155 ( .A(n10817), .B(n10816), .ZN(n10757) );
  OAI222_X1 U13156 ( .A1(n14527), .A2(n11751), .B1(n14525), .B2(n10758), .C1(
        n10757), .C2(n14936), .ZN(n15091) );
  MUX2_X1 U13157 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n15091), .S(n14541), .Z(
        n10759) );
  AOI211_X1 U13158 ( .C1(n14548), .C2(n15093), .A(n10760), .B(n10759), .ZN(
        n10761) );
  INV_X1 U13159 ( .A(n10761), .ZN(P1_U3285) );
  INV_X1 U13160 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11130) );
  XNOR2_X1 U13161 ( .A(n10763), .B(n10762), .ZN(n15237) );
  AND2_X1 U13162 ( .A1(n15281), .A2(n10764), .ZN(n10765) );
  NAND2_X1 U13163 ( .A1(n10766), .A2(n10765), .ZN(n10768) );
  NAND2_X1 U13164 ( .A1(n15237), .A2(n15201), .ZN(n10776) );
  AOI22_X1 U13165 ( .A1(n15212), .A2(n12693), .B1(n12691), .B2(n15215), .ZN(
        n10775) );
  NAND2_X1 U13166 ( .A1(n13212), .A2(n10769), .ZN(n13211) );
  OR2_X1 U13167 ( .A1(n12693), .A2(n7714), .ZN(n10770) );
  NAND2_X1 U13168 ( .A1(n13211), .A2(n10770), .ZN(n10772) );
  OAI21_X1 U13169 ( .B1(n10772), .B2(n10771), .A(n10897), .ZN(n10773) );
  NAND2_X1 U13170 ( .A1(n10773), .A2(n15218), .ZN(n10774) );
  NAND3_X1 U13171 ( .A1(n10776), .A2(n10775), .A3(n10774), .ZN(n15235) );
  INV_X1 U13172 ( .A(n15237), .ZN(n10778) );
  NAND2_X1 U13173 ( .A1(n10777), .A2(n15232), .ZN(n13143) );
  NAND2_X1 U13174 ( .A1(n10894), .A2(n15287), .ZN(n15233) );
  OAI21_X1 U13175 ( .B1(n10778), .B2(n13143), .A(n15233), .ZN(n10779) );
  NOR2_X1 U13176 ( .A1(n15235), .A2(n10779), .ZN(n15252) );
  MUX2_X1 U13177 ( .A(n11130), .B(n15252), .S(n15308), .Z(n10780) );
  INV_X1 U13178 ( .A(n10780), .ZN(P3_U3461) );
  NAND2_X1 U13179 ( .A1(n14067), .A2(n12404), .ZN(n10785) );
  INV_X2 U13180 ( .A(n12361), .ZN(n12400) );
  NAND2_X1 U13181 ( .A1(n14152), .A2(n12400), .ZN(n10784) );
  NAND2_X1 U13182 ( .A1(n10785), .A2(n10784), .ZN(n10787) );
  XNOR2_X1 U13183 ( .A(n10787), .B(n10786), .ZN(n10789) );
  AOI22_X1 U13184 ( .A1(n14067), .A2(n12400), .B1(n10120), .B2(n14152), .ZN(
        n10788) );
  AND2_X1 U13185 ( .A1(n10789), .A2(n10788), .ZN(n14061) );
  OR2_X1 U13186 ( .A1(n10789), .A2(n10788), .ZN(n14060) );
  NAND2_X1 U13187 ( .A1(n12132), .A2(n12404), .ZN(n10791) );
  NAND2_X1 U13188 ( .A1(n14151), .A2(n12400), .ZN(n10790) );
  NAND2_X1 U13189 ( .A1(n10791), .A2(n10790), .ZN(n10792) );
  XNOR2_X1 U13190 ( .A(n10792), .B(n12292), .ZN(n10945) );
  AOI22_X1 U13191 ( .A1(n12132), .A2(n12400), .B1(n9737), .B2(n14151), .ZN(
        n10946) );
  XNOR2_X1 U13192 ( .A(n10945), .B(n10946), .ZN(n10793) );
  NAND2_X1 U13193 ( .A1(n10794), .A2(n10793), .ZN(n10949) );
  OAI211_X1 U13194 ( .C1(n10794), .C2(n10793), .A(n10949), .B(n14930), .ZN(
        n10800) );
  INV_X1 U13195 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10795) );
  NOR2_X1 U13196 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10795), .ZN(n14200) );
  NOR2_X1 U13197 ( .A1(n14111), .A2(n10796), .ZN(n10797) );
  AOI211_X1 U13198 ( .C1(n14113), .C2(n10798), .A(n14200), .B(n10797), .ZN(
        n10799) );
  OAI211_X1 U13199 ( .C1(n10801), .C2(n14927), .A(n10800), .B(n10799), .ZN(
        P1_U3239) );
  AOI211_X1 U13200 ( .C1(n13905), .C2(n10804), .A(n10803), .B(n10802), .ZN(
        n10810) );
  AOI22_X1 U13201 ( .A1(n11010), .A2(n13899), .B1(n15188), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n10805) );
  OAI21_X1 U13202 ( .B1(n10810), .B2(n15188), .A(n10805), .ZN(P2_U3509) );
  INV_X1 U13203 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10806) );
  OAI22_X1 U13204 ( .A1(n10807), .A2(n13974), .B1(n15187), .B2(n10806), .ZN(
        n10808) );
  INV_X1 U13205 ( .A(n10808), .ZN(n10809) );
  OAI21_X1 U13206 ( .B1(n10810), .B2(n15185), .A(n10809), .ZN(P2_U3460) );
  INV_X1 U13207 ( .A(n13550), .ZN(n13538) );
  INV_X1 U13208 ( .A(n11981), .ZN(n10815) );
  OAI222_X1 U13209 ( .A1(P2_U3088), .A2(n13538), .B1(n14001), .B2(n10815), 
        .C1(n10811), .C2(n13999), .ZN(P2_U3309) );
  NAND2_X1 U13210 ( .A1(n10812), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10813) );
  XNOR2_X1 U13211 ( .A(n10813), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14236) );
  INV_X1 U13212 ( .A(n14236), .ZN(n14230) );
  OAI222_X1 U13213 ( .A1(P1_U3086), .A2(n14230), .B1(n14707), .B2(n10815), 
        .C1(n10814), .C2(n14709), .ZN(P1_U3337) );
  OR2_X1 U13214 ( .A1(n12139), .A2(n10874), .ZN(n10818) );
  NAND2_X1 U13215 ( .A1(n10820), .A2(n6429), .ZN(n10823) );
  AOI22_X1 U13216 ( .A1(n12023), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10821), 
        .B2(n12022), .ZN(n10822) );
  XNOR2_X1 U13217 ( .A(n12148), .B(n11751), .ZN(n12011) );
  NAND2_X1 U13218 ( .A1(n12148), .A2(n11751), .ZN(n10824) );
  NAND2_X1 U13219 ( .A1(n10825), .A2(n6429), .ZN(n10827) );
  AOI22_X1 U13220 ( .A1(n14220), .A2(n12022), .B1(n12023), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10826) );
  AND2_X1 U13221 ( .A1(n10828), .A2(n15349), .ZN(n10829) );
  OR2_X1 U13222 ( .A1(n10829), .A2(n10843), .ZN(n14917) );
  INV_X1 U13223 ( .A(n14917), .ZN(n10830) );
  NAND2_X1 U13224 ( .A1(n11974), .A2(n10830), .ZN(n10834) );
  NAND2_X1 U13225 ( .A1(n12059), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13226 ( .A1(n12060), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U13227 ( .A1(n12061), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10831) );
  NAND4_X1 U13228 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(
        n14922) );
  XNOR2_X1 U13229 ( .A(n14905), .B(n14922), .ZN(n12012) );
  AOI21_X1 U13230 ( .B1(n10835), .B2(n10839), .A(n14936), .ZN(n10836) );
  AOI22_X1 U13231 ( .A1(n10836), .A2(n11336), .B1(n15007), .B2(n14909), .ZN(
        n15105) );
  OR2_X1 U13232 ( .A1(n12139), .A2(n14149), .ZN(n10837) );
  NAND2_X1 U13233 ( .A1(n10840), .A2(n10839), .ZN(n11320) );
  OAI21_X1 U13234 ( .B1(n10840), .B2(n10839), .A(n11320), .ZN(n15107) );
  INV_X1 U13235 ( .A(n10880), .ZN(n10841) );
  AOI21_X1 U13236 ( .B1(n10841), .B2(n14905), .A(n14640), .ZN(n10850) );
  INV_X1 U13237 ( .A(n14905), .ZN(n10842) );
  NOR2_X1 U13238 ( .A1(n10843), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10844) );
  OR2_X1 U13239 ( .A1(n11329), .A2(n10844), .ZN(n14934) );
  INV_X1 U13240 ( .A(n14934), .ZN(n10845) );
  NAND2_X1 U13241 ( .A1(n11974), .A2(n10845), .ZN(n10849) );
  NAND2_X1 U13242 ( .A1(n12059), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U13243 ( .A1(n10484), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13244 ( .A1(n12061), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10846) );
  NAND4_X1 U13245 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n14910) );
  AOI22_X1 U13246 ( .A1(n10850), .A2(n11327), .B1(n14509), .B2(n14910), .ZN(
        n15104) );
  OAI22_X1 U13247 ( .A1(n14541), .A2(n9776), .B1(n14917), .B2(n14544), .ZN(
        n10851) );
  AOI21_X1 U13248 ( .B1(n14546), .B2(n14905), .A(n10851), .ZN(n10852) );
  OAI21_X1 U13249 ( .B1(n15104), .B2(n14537), .A(n10852), .ZN(n10853) );
  AOI21_X1 U13250 ( .B1(n15107), .B2(n14548), .A(n10853), .ZN(n10854) );
  OAI21_X1 U13251 ( .B1(n15105), .B2(n15022), .A(n10854), .ZN(P1_U3283) );
  INV_X1 U13252 ( .A(n10855), .ZN(n10856) );
  NAND2_X1 U13253 ( .A1(n10856), .A2(n12691), .ZN(n10857) );
  INV_X1 U13254 ( .A(n10918), .ZN(n11015) );
  XNOR2_X1 U13255 ( .A(n10859), .B(n11015), .ZN(n10860) );
  NAND2_X1 U13256 ( .A1(n10860), .A2(n11019), .ZN(n10987) );
  INV_X1 U13257 ( .A(n10860), .ZN(n10861) );
  NAND2_X1 U13258 ( .A1(n10861), .A2(n12690), .ZN(n10862) );
  NAND2_X1 U13259 ( .A1(n10987), .A2(n10862), .ZN(n10864) );
  INV_X1 U13260 ( .A(n10988), .ZN(n10863) );
  AOI21_X1 U13261 ( .B1(n10865), .B2(n10864), .A(n10863), .ZN(n10871) );
  INV_X1 U13262 ( .A(n10866), .ZN(n10919) );
  INV_X1 U13263 ( .A(n12666), .ZN(n12655) );
  AOI22_X1 U13264 ( .A1(n11015), .A2(n12672), .B1(n12655), .B2(n15213), .ZN(
        n10867) );
  NAND2_X1 U13265 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11242) );
  OAI211_X1 U13266 ( .C1(n10868), .C2(n12659), .A(n10867), .B(n11242), .ZN(
        n10869) );
  AOI21_X1 U13267 ( .B1(n10919), .B2(n12656), .A(n10869), .ZN(n10870) );
  OAI21_X1 U13268 ( .B1(n10871), .B2(n12674), .A(n10870), .ZN(P3_U3170) );
  OAI21_X1 U13269 ( .B1(n10873), .B2(n12011), .A(n10872), .ZN(n15099) );
  INV_X1 U13270 ( .A(n15099), .ZN(n10887) );
  INV_X1 U13271 ( .A(n14922), .ZN(n12276) );
  OAI22_X1 U13272 ( .A1(n12276), .A2(n14527), .B1(n10874), .B2(n14525), .ZN(
        n10879) );
  NAND2_X1 U13273 ( .A1(n10875), .A2(n12011), .ZN(n10876) );
  AOI21_X1 U13274 ( .B1(n10877), .B2(n10876), .A(n14936), .ZN(n10878) );
  AOI211_X1 U13275 ( .C1(n15068), .C2(n15099), .A(n10879), .B(n10878), .ZN(
        n15101) );
  MUX2_X1 U13276 ( .A(n9775), .B(n15101), .S(n14541), .Z(n10886) );
  AOI211_X1 U13277 ( .C1(n12148), .C2(n10881), .A(n14640), .B(n10880), .ZN(
        n15096) );
  INV_X1 U13278 ( .A(n12148), .ZN(n10883) );
  INV_X1 U13279 ( .A(n11757), .ZN(n10882) );
  OAI22_X1 U13280 ( .A1(n10883), .A2(n15012), .B1(n14544), .B2(n10882), .ZN(
        n10884) );
  AOI21_X1 U13281 ( .B1(n15096), .B2(n15018), .A(n10884), .ZN(n10885) );
  OAI211_X1 U13282 ( .C1(n10887), .C2(n11542), .A(n10886), .B(n10885), .ZN(
        P1_U3284) );
  INV_X1 U13283 ( .A(n11961), .ZN(n10889) );
  OAI222_X1 U13284 ( .A1(P1_U3086), .A2(n14320), .B1(n14707), .B2(n10889), 
        .C1(n10888), .C2(n14701), .ZN(P1_U3336) );
  OAI222_X1 U13285 ( .A1(n13999), .A2(n10890), .B1(n14001), .B2(n10889), .C1(
        n9628), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U13286 ( .A(n10892), .B(n10891), .ZN(n15256) );
  INV_X2 U13287 ( .A(n15250), .ZN(n15248) );
  NAND2_X1 U13288 ( .A1(n10893), .A2(n15232), .ZN(n15202) );
  INV_X1 U13289 ( .A(n15202), .ZN(n15238) );
  NAND2_X1 U13290 ( .A1(n10911), .A2(n15287), .ZN(n15253) );
  OAI22_X1 U13291 ( .A1(n10917), .A2(n15253), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15234), .ZN(n10903) );
  OR2_X1 U13292 ( .A1(n13214), .A2(n10894), .ZN(n10896) );
  AOI21_X1 U13293 ( .B1(n10897), .B2(n10896), .A(n10895), .ZN(n10901) );
  NAND2_X1 U13294 ( .A1(n10913), .A2(n15218), .ZN(n10900) );
  NAND2_X1 U13295 ( .A1(n15256), .A2(n15201), .ZN(n10899) );
  AOI22_X1 U13296 ( .A1(n15212), .A2(n13214), .B1(n12690), .B2(n15215), .ZN(
        n10898) );
  OAI211_X1 U13297 ( .C1(n10901), .C2(n10900), .A(n10899), .B(n10898), .ZN(
        n15254) );
  MUX2_X1 U13298 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15254), .S(n15248), .Z(
        n10902) );
  AOI211_X1 U13299 ( .C1(n15256), .C2(n15246), .A(n10903), .B(n10902), .ZN(
        n10904) );
  INV_X1 U13300 ( .A(n10904), .ZN(P3_U3230) );
  INV_X1 U13301 ( .A(n10905), .ZN(n10907) );
  INV_X1 U13302 ( .A(SI_24_), .ZN(n10906) );
  OAI222_X1 U13303 ( .A1(P3_U3151), .A2(n10908), .B1(n11891), .B2(n10907), 
        .C1(n10906), .C2(n11887), .ZN(P3_U3271) );
  XNOR2_X1 U13304 ( .A(n10910), .B(n10909), .ZN(n15261) );
  INV_X1 U13305 ( .A(n15261), .ZN(n10922) );
  NAND2_X1 U13306 ( .A1(n12691), .A2(n10911), .ZN(n10912) );
  XNOR2_X1 U13307 ( .A(n11014), .B(n11013), .ZN(n10915) );
  AOI22_X1 U13308 ( .A1(n15215), .A2(n15213), .B1(n12691), .B2(n15212), .ZN(
        n10914) );
  OAI21_X1 U13309 ( .B1(n10915), .B2(n14854), .A(n10914), .ZN(n10916) );
  AOI21_X1 U13310 ( .B1(n15261), .B2(n15201), .A(n10916), .ZN(n15258) );
  MUX2_X1 U13311 ( .A(n15315), .B(n15258), .S(n15248), .Z(n10921) );
  NOR2_X1 U13312 ( .A1(n10918), .A2(n15281), .ZN(n15260) );
  AOI22_X1 U13313 ( .A1(n15228), .A2(n15260), .B1(n15244), .B2(n10919), .ZN(
        n10920) );
  OAI211_X1 U13314 ( .C1(n10922), .C2(n12945), .A(n10921), .B(n10920), .ZN(
        P3_U3229) );
  INV_X1 U13315 ( .A(n11970), .ZN(n10961) );
  OAI222_X1 U13316 ( .A1(n10923), .A2(P1_U3086), .B1(n14707), .B2(n10961), 
        .C1(n6945), .C2(n14701), .ZN(P1_U3335) );
  INV_X1 U13317 ( .A(n10924), .ZN(n10925) );
  XNOR2_X1 U13318 ( .A(n11354), .B(n10929), .ZN(n10965) );
  INV_X1 U13319 ( .A(n10965), .ZN(n10944) );
  INV_X1 U13320 ( .A(n13481), .ZN(n10930) );
  OR2_X1 U13321 ( .A1(n11010), .A2(n10930), .ZN(n10931) );
  NAND2_X1 U13322 ( .A1(n10932), .A2(n10931), .ZN(n10935) );
  INV_X1 U13323 ( .A(n11345), .ZN(n10934) );
  AOI21_X1 U13324 ( .B1(n7646), .B2(n10935), .A(n10934), .ZN(n10936) );
  AOI22_X1 U13325 ( .A1(n13570), .A2(n13479), .B1(n13464), .B2(n13481), .ZN(
        n11404) );
  OAI21_X1 U13326 ( .B1(n10936), .B2(n13795), .A(n11404), .ZN(n10963) );
  INV_X1 U13327 ( .A(n11412), .ZN(n10941) );
  INV_X1 U13328 ( .A(n11415), .ZN(n10937) );
  AOI211_X1 U13329 ( .C1(n11412), .C2(n10938), .A(n13343), .B(n10937), .ZN(
        n10964) );
  NAND2_X1 U13330 ( .A1(n10964), .A2(n13850), .ZN(n10940) );
  AOI22_X1 U13331 ( .A1(n6430), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11401), 
        .B2(n13828), .ZN(n10939) );
  OAI211_X1 U13332 ( .C1(n10941), .C2(n13816), .A(n10940), .B(n10939), .ZN(
        n10942) );
  AOI21_X1 U13333 ( .B1(n10963), .B2(n13844), .A(n10942), .ZN(n10943) );
  OAI21_X1 U13334 ( .B1(n10944), .B2(n13835), .A(n10943), .ZN(P2_U3254) );
  NAND2_X1 U13335 ( .A1(n12135), .A2(n15062), .ZN(n15082) );
  NAND2_X1 U13336 ( .A1(n10945), .A2(n10947), .ZN(n10948) );
  NAND2_X1 U13337 ( .A1(n12135), .A2(n12404), .ZN(n10951) );
  NAND2_X1 U13338 ( .A1(n14150), .A2(n12400), .ZN(n10950) );
  NAND2_X1 U13339 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  XNOR2_X1 U13340 ( .A(n10952), .B(n12292), .ZN(n11057) );
  AOI22_X1 U13341 ( .A1(n12135), .A2(n12400), .B1(n9737), .B2(n14150), .ZN(
        n11060) );
  XNOR2_X1 U13342 ( .A(n11057), .B(n11060), .ZN(n10953) );
  OAI211_X1 U13343 ( .C1(n10954), .C2(n10953), .A(n11058), .B(n14930), .ZN(
        n10960) );
  NAND2_X1 U13344 ( .A1(n14143), .A2(n15081), .ZN(n10955) );
  OAI211_X1 U13345 ( .C1(n14935), .C2(n10957), .A(n10956), .B(n10955), .ZN(
        n10958) );
  INV_X1 U13346 ( .A(n10958), .ZN(n10959) );
  OAI211_X1 U13347 ( .C1(n14913), .C2(n15082), .A(n10960), .B(n10959), .ZN(
        P1_U3213) );
  OAI222_X1 U13348 ( .A1(n13999), .A2(n15429), .B1(P2_U3088), .B2(n10962), 
        .C1(n13994), .C2(n10961), .ZN(P2_U3307) );
  AOI211_X1 U13349 ( .C1(n13905), .C2(n10965), .A(n10964), .B(n10963), .ZN(
        n10970) );
  AOI22_X1 U13350 ( .A1(n11412), .A2(n13899), .B1(n15188), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n10966) );
  OAI21_X1 U13351 ( .B1(n10970), .B2(n15188), .A(n10966), .ZN(P2_U3510) );
  INV_X1 U13352 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10967) );
  NOR2_X1 U13353 ( .A1(n15187), .A2(n10967), .ZN(n10968) );
  AOI21_X1 U13354 ( .B1(n11412), .B2(n13965), .A(n10968), .ZN(n10969) );
  OAI21_X1 U13355 ( .B1(n10970), .B2(n15185), .A(n10969), .ZN(P2_U3463) );
  OAI21_X1 U13356 ( .B1(n10972), .B2(n10154), .A(n10971), .ZN(n10973) );
  NOR2_X1 U13357 ( .A1(n11788), .A2(n10973), .ZN(n10974) );
  XNOR2_X1 U13358 ( .A(n10973), .B(n11788), .ZN(n14982) );
  NOR2_X1 U13359 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14982), .ZN(n14981) );
  NOR2_X1 U13360 ( .A1(n10974), .A2(n14981), .ZN(n10977) );
  NOR2_X1 U13361 ( .A1(n12021), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10975) );
  AOI21_X1 U13362 ( .B1(n12021), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10975), 
        .ZN(n10976) );
  NAND2_X1 U13363 ( .A1(n10976), .A2(n10977), .ZN(n11368) );
  OAI211_X1 U13364 ( .C1(n10977), .C2(n10976), .A(n14243), .B(n11368), .ZN(
        n10986) );
  NAND2_X1 U13365 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14054)
         );
  OR2_X1 U13366 ( .A1(n11764), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13367 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  XNOR2_X1 U13368 ( .A(n10980), .B(n14991), .ZN(n14986) );
  NOR2_X1 U13369 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14986), .ZN(n14985) );
  AOI21_X1 U13370 ( .B1(n14991), .B2(n10980), .A(n14985), .ZN(n10982) );
  XNOR2_X1 U13371 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11373), .ZN(n10981) );
  NAND2_X1 U13372 ( .A1(n10981), .A2(n10982), .ZN(n11372) );
  OAI211_X1 U13373 ( .C1(n10982), .C2(n10981), .A(n14245), .B(n11372), .ZN(
        n10983) );
  NAND2_X1 U13374 ( .A1(n14054), .A2(n10983), .ZN(n10984) );
  AOI21_X1 U13375 ( .B1(n14977), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10984), 
        .ZN(n10985) );
  OAI211_X1 U13376 ( .C1(n14992), .C2(n11373), .A(n10986), .B(n10985), .ZN(
        P1_U3259) );
  INV_X1 U13377 ( .A(n12656), .ZN(n12670) );
  XNOR2_X1 U13378 ( .A(n12543), .B(n11040), .ZN(n11223) );
  XNOR2_X1 U13379 ( .A(n11223), .B(n15213), .ZN(n10990) );
  NAND2_X1 U13380 ( .A1(n10989), .A2(n10990), .ZN(n11445) );
  OAI21_X1 U13381 ( .B1(n10990), .B2(n10989), .A(n11445), .ZN(n10991) );
  NAND2_X1 U13382 ( .A1(n10991), .A2(n12644), .ZN(n10995) );
  OAI22_X1 U13383 ( .A1(n12652), .A2(n11024), .B1(n12659), .B2(n11019), .ZN(
        n10993) );
  INV_X1 U13384 ( .A(n12689), .ZN(n11521) );
  OR2_X1 U13385 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7763), .ZN(n11215) );
  OAI21_X1 U13386 ( .B1(n12666), .B2(n11521), .A(n11215), .ZN(n10992) );
  NOR2_X1 U13387 ( .A1(n10993), .A2(n10992), .ZN(n10994) );
  OAI211_X1 U13388 ( .C1(n11025), .C2(n12670), .A(n10995), .B(n10994), .ZN(
        P3_U3167) );
  NAND2_X1 U13389 ( .A1(n14885), .A2(n10996), .ZN(n10998) );
  OAI211_X1 U13390 ( .C1(n14891), .C2(n10999), .A(n10998), .B(n10997), .ZN(
        n11009) );
  XNOR2_X1 U13391 ( .A(n11010), .B(n9828), .ZN(n11001) );
  AND2_X1 U13392 ( .A1(n13481), .A2(n13687), .ZN(n11000) );
  NAND2_X1 U13393 ( .A1(n11001), .A2(n11000), .ZN(n11405) );
  OAI21_X1 U13394 ( .B1(n11001), .B2(n11000), .A(n11405), .ZN(n11007) );
  INV_X1 U13395 ( .A(n11002), .ZN(n11005) );
  AOI211_X1 U13396 ( .C1(n11007), .C2(n11006), .A(n13470), .B(n11407), .ZN(
        n11008) );
  AOI211_X1 U13397 ( .C1(n11010), .C2(n9631), .A(n11009), .B(n11008), .ZN(
        n11011) );
  INV_X1 U13398 ( .A(n11011), .ZN(P2_U3189) );
  XNOR2_X1 U13399 ( .A(n11012), .B(n11039), .ZN(n11023) );
  NAND2_X1 U13400 ( .A1(n12690), .A2(n11015), .ZN(n11016) );
  NAND2_X1 U13401 ( .A1(n11017), .A2(n11016), .ZN(n11044) );
  OR2_X1 U13402 ( .A1(n11044), .A2(n11018), .ZN(n15217) );
  OAI21_X1 U13403 ( .B1(n6670), .B2(n11039), .A(n15217), .ZN(n11021) );
  OAI22_X1 U13404 ( .A1(n11521), .A2(n14859), .B1(n11019), .B2(n14857), .ZN(
        n11020) );
  AOI21_X1 U13405 ( .B1(n11021), .B2(n15218), .A(n11020), .ZN(n11022) );
  OAI21_X1 U13406 ( .B1(n15223), .B2(n11023), .A(n11022), .ZN(n15263) );
  INV_X1 U13407 ( .A(n15263), .ZN(n11030) );
  INV_X1 U13408 ( .A(n11023), .ZN(n15265) );
  NOR2_X1 U13409 ( .A1(n11024), .A2(n15281), .ZN(n15264) );
  INV_X1 U13410 ( .A(n11025), .ZN(n11026) );
  AOI22_X1 U13411 ( .A1(n15228), .A2(n15264), .B1(n15244), .B2(n11026), .ZN(
        n11027) );
  OAI21_X1 U13412 ( .B1(n11102), .B2(n15248), .A(n11027), .ZN(n11028) );
  AOI21_X1 U13413 ( .B1(n15265), .B2(n15246), .A(n11028), .ZN(n11029) );
  OAI21_X1 U13414 ( .B1(n11030), .B2(n15250), .A(n11029), .ZN(P3_U3228) );
  INV_X1 U13415 ( .A(n11031), .ZN(n11034) );
  OAI222_X1 U13416 ( .A1(n11891), .A2(n11034), .B1(n12420), .B2(n11033), .C1(
        P3_U3151), .C2(n11032), .ZN(P3_U3270) );
  INV_X1 U13417 ( .A(n12028), .ZN(n11381) );
  OAI222_X1 U13418 ( .A1(n13999), .A2(n11036), .B1(n14001), .B2(n11381), .C1(
        n11035), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U13419 ( .A(n11037), .B(n11047), .ZN(n15277) );
  INV_X1 U13420 ( .A(n15225), .ZN(n11038) );
  NAND2_X1 U13421 ( .A1(n12689), .A2(n11038), .ZN(n11307) );
  NAND2_X1 U13422 ( .A1(n11039), .A2(n11307), .ZN(n11043) );
  OR2_X1 U13423 ( .A1(n15213), .A2(n11040), .ZN(n15216) );
  NAND2_X1 U13424 ( .A1(n11041), .A2(n15216), .ZN(n11305) );
  AOI21_X1 U13425 ( .B1(n11305), .B2(n11307), .A(n11441), .ZN(n11042) );
  INV_X1 U13426 ( .A(n11522), .ZN(n11045) );
  NAND2_X1 U13427 ( .A1(n15214), .A2(n11045), .ZN(n11046) );
  INV_X1 U13428 ( .A(n11047), .ZN(n11048) );
  XNOR2_X1 U13429 ( .A(n11599), .B(n11048), .ZN(n11050) );
  AOI22_X1 U13430 ( .A1(n15212), .A2(n15214), .B1(n15196), .B2(n15215), .ZN(
        n11049) );
  OAI21_X1 U13431 ( .B1(n11050), .B2(n14854), .A(n11049), .ZN(n11051) );
  AOI21_X1 U13432 ( .B1(n15277), .B2(n15201), .A(n11051), .ZN(n15279) );
  INV_X1 U13433 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11155) );
  AND2_X1 U13434 ( .A1(n11596), .A2(n15287), .ZN(n15276) );
  AOI22_X1 U13435 ( .A1(n15228), .A2(n15276), .B1(n15244), .B2(n11052), .ZN(
        n11053) );
  OAI21_X1 U13436 ( .B1(n11155), .B2(n15248), .A(n11053), .ZN(n11054) );
  AOI21_X1 U13437 ( .B1(n15277), .B2(n15246), .A(n11054), .ZN(n11055) );
  OAI21_X1 U13438 ( .B1(n15279), .B2(n15250), .A(n11055), .ZN(P3_U3225) );
  AOI22_X1 U13439 ( .A1(n12139), .A2(n12404), .B1(n12400), .B2(n14149), .ZN(
        n11056) );
  XNOR2_X1 U13440 ( .A(n11056), .B(n12292), .ZN(n11750) );
  AOI22_X1 U13441 ( .A1(n12139), .A2(n12400), .B1(n10120), .B2(n14149), .ZN(
        n11749) );
  XNOR2_X1 U13442 ( .A(n11750), .B(n11749), .ZN(n11062) );
  INV_X1 U13443 ( .A(n11057), .ZN(n11059) );
  AOI21_X1 U13444 ( .B1(n11062), .B2(n11061), .A(n6582), .ZN(n11069) );
  NAND2_X1 U13445 ( .A1(n14923), .A2(n14150), .ZN(n11064) );
  OAI211_X1 U13446 ( .C1(n14120), .C2(n11751), .A(n11064), .B(n11063), .ZN(
        n11066) );
  NAND2_X1 U13447 ( .A1(n12139), .A2(n15062), .ZN(n15089) );
  NOR2_X1 U13448 ( .A1(n15089), .A2(n14913), .ZN(n11065) );
  AOI211_X1 U13449 ( .C1(n14113), .C2(n11067), .A(n11066), .B(n11065), .ZN(
        n11068) );
  OAI21_X1 U13450 ( .B1(n11069), .B2(n14133), .A(n11068), .ZN(P1_U3221) );
  INV_X1 U13451 ( .A(n11070), .ZN(n11072) );
  NAND2_X1 U13452 ( .A1(n11072), .A2(n11071), .ZN(n11129) );
  NAND2_X1 U13453 ( .A1(n11074), .A2(n11073), .ZN(n11075) );
  NAND2_X1 U13454 ( .A1(n11076), .A2(n11075), .ZN(n11128) );
  INV_X1 U13455 ( .A(n11128), .ZN(n11077) );
  NAND2_X1 U13456 ( .A1(n11129), .A2(n11077), .ZN(n11144) );
  MUX2_X1 U13457 ( .A(n11144), .B(n12680), .S(n12452), .Z(n12881) );
  INV_X1 U13458 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U13459 ( .A1(n11081), .A2(n11080), .ZN(n11295) );
  INV_X1 U13460 ( .A(n11081), .ZN(n11082) );
  NAND2_X1 U13461 ( .A1(n11082), .A2(n11629), .ZN(n11083) );
  NAND2_X1 U13462 ( .A1(n11295), .A2(n11083), .ZN(n11621) );
  OR2_X1 U13463 ( .A1(n11621), .A2(n11620), .ZN(n11618) );
  INV_X1 U13464 ( .A(n11299), .ZN(n11086) );
  NAND2_X1 U13465 ( .A1(n11087), .A2(n11086), .ZN(n11578) );
  INV_X1 U13466 ( .A(n11087), .ZN(n11088) );
  NAND2_X1 U13467 ( .A1(n11088), .A2(n11299), .ZN(n11089) );
  NAND2_X1 U13468 ( .A1(n11578), .A2(n11089), .ZN(n11294) );
  INV_X1 U13469 ( .A(n11578), .ZN(n11095) );
  NAND2_X1 U13470 ( .A1(n11092), .A2(n7384), .ZN(n11253) );
  INV_X1 U13471 ( .A(n11092), .ZN(n11093) );
  NAND2_X1 U13472 ( .A1(n11093), .A2(n11135), .ZN(n11094) );
  NAND2_X1 U13473 ( .A1(n11253), .A2(n11094), .ZN(n11577) );
  INV_X1 U13474 ( .A(n11258), .ZN(n11096) );
  NAND2_X1 U13475 ( .A1(n11097), .A2(n11096), .ZN(n11100) );
  INV_X1 U13476 ( .A(n11097), .ZN(n11098) );
  NAND2_X1 U13477 ( .A1(n11098), .A2(n11258), .ZN(n11099) );
  NAND2_X1 U13478 ( .A1(n11100), .A2(n11099), .ZN(n11252) );
  INV_X1 U13479 ( .A(n11100), .ZN(n11209) );
  NAND2_X1 U13480 ( .A1(n11103), .A2(n11138), .ZN(n12695) );
  INV_X1 U13481 ( .A(n11103), .ZN(n11104) );
  NAND2_X1 U13482 ( .A1(n11104), .A2(n11222), .ZN(n11105) );
  AND2_X1 U13483 ( .A1(n12695), .A2(n11105), .ZN(n11208) );
  NAND2_X1 U13484 ( .A1(n11106), .A2(n12705), .ZN(n11109) );
  INV_X1 U13485 ( .A(n11106), .ZN(n11107) );
  NAND2_X1 U13486 ( .A1(n11107), .A2(n11141), .ZN(n11108) );
  NAND2_X1 U13487 ( .A1(n11109), .A2(n11108), .ZN(n12694) );
  AOI21_X1 U13488 ( .B1(n12696), .B2(n12695), .A(n12694), .ZN(n12698) );
  INV_X1 U13489 ( .A(n11109), .ZN(n11115) );
  NAND2_X1 U13490 ( .A1(n11112), .A2(n11142), .ZN(n12716) );
  INV_X1 U13491 ( .A(n11112), .ZN(n11113) );
  NAND2_X1 U13492 ( .A1(n11113), .A2(n11152), .ZN(n11114) );
  INV_X1 U13493 ( .A(n12717), .ZN(n11117) );
  NOR3_X1 U13494 ( .A1(n12698), .A2(n11115), .A3(n7663), .ZN(n11116) );
  OAI21_X1 U13495 ( .B1(n11117), .B2(n11116), .A(n12890), .ZN(n11151) );
  XNOR2_X1 U13496 ( .A(n11299), .B(n11119), .ZN(n11289) );
  NOR2_X1 U13497 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11085), .ZN(n11654) );
  NAND2_X1 U13498 ( .A1(n11120), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11121) );
  OAI21_X1 U13499 ( .B1(n11629), .B2(n11654), .A(n11121), .ZN(n11617) );
  OR2_X1 U13500 ( .A1(n11617), .A2(n11079), .ZN(n11615) );
  NAND2_X1 U13501 ( .A1(n11615), .A2(n11121), .ZN(n11288) );
  NAND2_X1 U13502 ( .A1(n11289), .A2(n11288), .ZN(n11287) );
  NAND2_X1 U13503 ( .A1(n11299), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U13504 ( .A1(n11287), .A2(n11122), .ZN(n11123) );
  NAND2_X1 U13505 ( .A1(n11123), .A2(n11135), .ZN(n11245) );
  XNOR2_X1 U13506 ( .A(n11258), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11246) );
  AOI21_X1 U13507 ( .B1(n11124), .B2(n11138), .A(n11125), .ZN(n11212) );
  NAND2_X1 U13508 ( .A1(n11212), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n12708) );
  INV_X1 U13509 ( .A(n11125), .ZN(n12706) );
  XNOR2_X1 U13510 ( .A(n12705), .B(n15230), .ZN(n12707) );
  AOI21_X1 U13511 ( .B1(n12708), .B2(n12706), .A(n12707), .ZN(n12710) );
  AOI21_X1 U13512 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n11141), .A(n12710), .ZN(
        n11126) );
  OAI21_X1 U13513 ( .B1(n11127), .B2(P3_REG2_REG_7__SCAN_IN), .A(n12723), .ZN(
        n11149) );
  INV_X1 U13514 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11147) );
  XNOR2_X1 U13515 ( .A(n11299), .B(n11130), .ZN(n11286) );
  NOR2_X1 U13516 ( .A1(n11084), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11131) );
  INV_X1 U13517 ( .A(n11131), .ZN(n11658) );
  NAND2_X1 U13518 ( .A1(n11629), .A2(n11658), .ZN(n11133) );
  NAND2_X1 U13519 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11131), .ZN(n11132) );
  NAND2_X1 U13520 ( .A1(n11133), .A2(n11132), .ZN(n11614) );
  NAND2_X1 U13521 ( .A1(n11614), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11613) );
  NAND2_X1 U13522 ( .A1(n11613), .A2(n7665), .ZN(n11285) );
  NAND2_X1 U13523 ( .A1(n11286), .A2(n11285), .ZN(n11284) );
  NAND2_X1 U13524 ( .A1(n11299), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U13525 ( .A1(n11284), .A2(n11134), .ZN(n11136) );
  NAND2_X1 U13526 ( .A1(n11136), .A2(n11135), .ZN(n11238) );
  OR2_X1 U13527 ( .A1(n11136), .A2(n11135), .ZN(n11137) );
  AOI21_X1 U13528 ( .B1(n11139), .B2(n11138), .A(n11140), .ZN(n11213) );
  NAND2_X1 U13529 ( .A1(n11213), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n12701) );
  INV_X1 U13530 ( .A(n11140), .ZN(n12699) );
  XNOR2_X1 U13531 ( .A(n12705), .B(n15300), .ZN(n12700) );
  OAI21_X1 U13532 ( .B1(n6463), .B2(P3_REG1_REG_7__SCAN_IN), .A(n12730), .ZN(
        n11145) );
  NAND2_X1 U13533 ( .A1(n11145), .A2(n12864), .ZN(n11146) );
  NAND2_X1 U13534 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11523) );
  OAI211_X1 U13535 ( .C1(n12849), .C2(n11147), .A(n11146), .B(n11523), .ZN(
        n11148) );
  AOI21_X1 U13536 ( .B1(n12835), .B2(n11149), .A(n11148), .ZN(n11150) );
  OAI211_X1 U13537 ( .C1(n12881), .C2(n11152), .A(n11151), .B(n11150), .ZN(
        P3_U3189) );
  INV_X1 U13538 ( .A(n12727), .ZN(n11153) );
  XNOR2_X1 U13539 ( .A(n12720), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n12724) );
  NOR2_X1 U13540 ( .A1(n11162), .A2(n11154), .ZN(n11181) );
  AOI21_X1 U13541 ( .B1(n11162), .B2(n11154), .A(n11181), .ZN(n11179) );
  NAND2_X1 U13542 ( .A1(n11157), .A2(n11156), .ZN(n11160) );
  INV_X1 U13543 ( .A(n11157), .ZN(n11158) );
  NAND2_X1 U13544 ( .A1(n11158), .A2(n12720), .ZN(n11159) );
  NAND2_X1 U13545 ( .A1(n11160), .A2(n11159), .ZN(n12715) );
  INV_X1 U13546 ( .A(n11160), .ZN(n11166) );
  NAND2_X1 U13547 ( .A1(n11163), .A2(n7232), .ZN(n11191) );
  INV_X1 U13548 ( .A(n11163), .ZN(n11164) );
  NAND2_X1 U13549 ( .A1(n11164), .A2(n11172), .ZN(n11165) );
  INV_X1 U13550 ( .A(n11192), .ZN(n11168) );
  NOR3_X1 U13551 ( .A1(n12719), .A2(n11166), .A3(n7662), .ZN(n11167) );
  OAI21_X1 U13552 ( .B1(n11168), .B2(n11167), .A(n12890), .ZN(n11178) );
  INV_X1 U13553 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11170) );
  NOR2_X1 U13554 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7838), .ZN(n11458) );
  INV_X1 U13555 ( .A(n11458), .ZN(n11169) );
  OAI21_X1 U13556 ( .B1(n12849), .B2(n11170), .A(n11169), .ZN(n11176) );
  INV_X1 U13557 ( .A(n12732), .ZN(n11171) );
  AOI21_X1 U13558 ( .B1(n11161), .B2(n11173), .A(n11197), .ZN(n11174) );
  NOR2_X1 U13559 ( .A1(n11174), .A2(n12892), .ZN(n11175) );
  AOI211_X1 U13560 ( .C1(n12859), .C2(n7232), .A(n11176), .B(n11175), .ZN(
        n11177) );
  OAI211_X1 U13561 ( .C1(n11179), .C2(n12888), .A(n11178), .B(n11177), .ZN(
        P3_U3191) );
  NOR2_X1 U13562 ( .A1(n7232), .A2(n11180), .ZN(n11182) );
  NAND2_X1 U13563 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11393), .ZN(n11183) );
  OAI21_X1 U13564 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11393), .A(n11183), 
        .ZN(n11184) );
  AOI21_X1 U13565 ( .B1(n11185), .B2(n11184), .A(n11392), .ZN(n11207) );
  INV_X1 U13566 ( .A(n11393), .ZN(n11204) );
  NAND2_X1 U13567 ( .A1(n11187), .A2(n11204), .ZN(n11382) );
  INV_X1 U13568 ( .A(n11187), .ZN(n11188) );
  NAND2_X1 U13569 ( .A1(n11188), .A2(n11393), .ZN(n11189) );
  NAND2_X1 U13570 ( .A1(n11382), .A2(n11189), .ZN(n11190) );
  AND3_X1 U13571 ( .A1(n11192), .A2(n11191), .A3(n11190), .ZN(n11193) );
  OAI21_X1 U13572 ( .B1(n11384), .B2(n11193), .A(n12890), .ZN(n11206) );
  INV_X1 U13573 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11195) );
  INV_X1 U13574 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11194) );
  OR2_X1 U13575 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11194), .ZN(n11569) );
  OAI21_X1 U13576 ( .B1(n12849), .B2(n11195), .A(n11569), .ZN(n11203) );
  NAND2_X1 U13577 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11393), .ZN(n11198) );
  OAI21_X1 U13578 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11393), .A(n11198), 
        .ZN(n11199) );
  AOI21_X1 U13579 ( .B1(n11200), .B2(n11199), .A(n11387), .ZN(n11201) );
  NOR2_X1 U13580 ( .A1(n11201), .A2(n12892), .ZN(n11202) );
  AOI211_X1 U13581 ( .C1(n12859), .C2(n11204), .A(n11203), .B(n11202), .ZN(
        n11205) );
  OAI211_X1 U13582 ( .C1(n11207), .C2(n12888), .A(n11206), .B(n11205), .ZN(
        P3_U3192) );
  INV_X1 U13583 ( .A(n12696), .ZN(n11211) );
  NOR3_X1 U13584 ( .A1(n11255), .A2(n11209), .A3(n11208), .ZN(n11210) );
  OAI21_X1 U13585 ( .B1(n11211), .B2(n11210), .A(n12890), .ZN(n11221) );
  OAI21_X1 U13586 ( .B1(n11212), .B2(P3_REG2_REG_5__SCAN_IN), .A(n12708), .ZN(
        n11219) );
  INV_X1 U13587 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11217) );
  OAI21_X1 U13588 ( .B1(n11213), .B2(P3_REG1_REG_5__SCAN_IN), .A(n12701), .ZN(
        n11214) );
  NAND2_X1 U13589 ( .A1(n12864), .A2(n11214), .ZN(n11216) );
  OAI211_X1 U13590 ( .C1(n12849), .C2(n11217), .A(n11216), .B(n11215), .ZN(
        n11218) );
  AOI21_X1 U13591 ( .B1(n12835), .B2(n11219), .A(n11218), .ZN(n11220) );
  OAI211_X1 U13592 ( .C1(n12881), .C2(n11222), .A(n11221), .B(n11220), .ZN(
        P3_U3187) );
  INV_X1 U13593 ( .A(n15213), .ZN(n11226) );
  NAND2_X1 U13594 ( .A1(n11223), .A2(n11226), .ZN(n11442) );
  AND2_X1 U13595 ( .A1(n11445), .A2(n11442), .ZN(n11225) );
  XNOR2_X1 U13596 ( .A(n12543), .B(n15225), .ZN(n11446) );
  XOR2_X1 U13597 ( .A(n11446), .B(n12689), .Z(n11224) );
  NAND2_X1 U13598 ( .A1(n11225), .A2(n11224), .ZN(n11518) );
  OAI211_X1 U13599 ( .C1(n11225), .C2(n11224), .A(n11518), .B(n12644), .ZN(
        n11236) );
  OAI22_X1 U13600 ( .A1(n15225), .A2(n12652), .B1(n12659), .B2(n11226), .ZN(
        n11234) );
  AND4_X1 U13601 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(
        n11734) );
  INV_X1 U13602 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11231) );
  NOR2_X1 U13603 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11231), .ZN(n12704) );
  INV_X1 U13604 ( .A(n12704), .ZN(n11232) );
  OAI21_X1 U13605 ( .B1(n12666), .B2(n11734), .A(n11232), .ZN(n11233) );
  NOR2_X1 U13606 ( .A1(n11234), .A2(n11233), .ZN(n11235) );
  OAI211_X1 U13607 ( .C1(n15226), .C2(n12670), .A(n11236), .B(n11235), .ZN(
        P3_U3179) );
  INV_X1 U13608 ( .A(n11237), .ZN(n11241) );
  NAND3_X1 U13609 ( .A1(n11584), .A2(n11239), .A3(n11238), .ZN(n11240) );
  NAND2_X1 U13610 ( .A1(n11241), .A2(n11240), .ZN(n11251) );
  NAND2_X1 U13611 ( .A1(n15191), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U13612 ( .A1(n11243), .A2(n11242), .ZN(n11250) );
  INV_X1 U13613 ( .A(n11244), .ZN(n11248) );
  NAND3_X1 U13614 ( .A1(n11587), .A2(n11246), .A3(n11245), .ZN(n11247) );
  AOI21_X1 U13615 ( .B1(n11248), .B2(n11247), .A(n12888), .ZN(n11249) );
  AOI211_X1 U13616 ( .C1(n12864), .C2(n11251), .A(n11250), .B(n11249), .ZN(
        n11257) );
  AND3_X1 U13617 ( .A1(n11581), .A2(n11253), .A3(n11252), .ZN(n11254) );
  OAI21_X1 U13618 ( .B1(n11255), .B2(n11254), .A(n12890), .ZN(n11256) );
  OAI211_X1 U13619 ( .C1(n12881), .C2(n11258), .A(n11257), .B(n11256), .ZN(
        P3_U3186) );
  INV_X1 U13620 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11260) );
  AOI21_X1 U13621 ( .B1(n11270), .B2(n13843), .A(n11259), .ZN(n15147) );
  MUX2_X1 U13622 ( .A(n11260), .B(P2_REG2_REG_13__SCAN_IN), .S(n15142), .Z(
        n15146) );
  NAND2_X1 U13623 ( .A1(n15147), .A2(n15146), .ZN(n15145) );
  OAI21_X1 U13624 ( .B1(n11260), .B2(n15142), .A(n15145), .ZN(n11261) );
  NAND2_X1 U13625 ( .A1(n13524), .A2(n11261), .ZN(n11262) );
  NAND2_X1 U13626 ( .A1(n15156), .A2(n11263), .ZN(n11264) );
  NAND2_X1 U13627 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15159), .ZN(n15157) );
  OR2_X1 U13628 ( .A1(n11511), .A2(n11858), .ZN(n11266) );
  NAND2_X1 U13629 ( .A1(n11511), .A2(n11858), .ZN(n11265) );
  AND2_X1 U13630 ( .A1(n11266), .A2(n11265), .ZN(n11267) );
  OAI211_X1 U13631 ( .C1(n11268), .C2(n11267), .A(n15158), .B(n11506), .ZN(
        n11283) );
  NAND2_X1 U13632 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13409)
         );
  INV_X1 U13633 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11272) );
  XNOR2_X1 U13634 ( .A(n11273), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n13521) );
  INV_X1 U13635 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11271) );
  AOI21_X1 U13636 ( .B1(n10169), .B2(n11270), .A(n11269), .ZN(n15150) );
  MUX2_X1 U13637 ( .A(n11271), .B(P2_REG1_REG_13__SCAN_IN), .S(n15142), .Z(
        n15149) );
  NAND2_X1 U13638 ( .A1(n15150), .A2(n15149), .ZN(n15148) );
  OAI21_X1 U13639 ( .B1(n11271), .B2(n15142), .A(n15148), .ZN(n13522) );
  NAND2_X1 U13640 ( .A1(n13521), .A2(n13522), .ZN(n13520) );
  OAI21_X1 U13641 ( .B1(n11273), .B2(n11272), .A(n13520), .ZN(n11274) );
  NAND2_X1 U13642 ( .A1(n15156), .A2(n11274), .ZN(n11276) );
  XNOR2_X1 U13643 ( .A(n11275), .B(n11274), .ZN(n15162) );
  NAND2_X1 U13644 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15162), .ZN(n15160) );
  NAND2_X1 U13645 ( .A1(n11276), .A2(n15160), .ZN(n11279) );
  INV_X1 U13646 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11877) );
  XNOR2_X1 U13647 ( .A(n11277), .B(n11877), .ZN(n11278) );
  NAND2_X1 U13648 ( .A1(n11278), .A2(n11279), .ZN(n11510) );
  OAI211_X1 U13649 ( .C1(n11279), .C2(n11278), .A(n11510), .B(n15161), .ZN(
        n11280) );
  NAND2_X1 U13650 ( .A1(n13409), .A2(n11280), .ZN(n11281) );
  AOI21_X1 U13651 ( .B1(n15154), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11281), 
        .ZN(n11282) );
  OAI211_X1 U13652 ( .C1(n15143), .C2(n11511), .A(n11283), .B(n11282), .ZN(
        P2_U3230) );
  OAI21_X1 U13653 ( .B1(n11286), .B2(n11285), .A(n11284), .ZN(n11293) );
  OAI21_X1 U13654 ( .B1(n11289), .B2(n11288), .A(n11287), .ZN(n11290) );
  AND2_X1 U13655 ( .A1(n12835), .A2(n11290), .ZN(n11292) );
  OAI22_X1 U13656 ( .A1(n12849), .A2(n15313), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10585), .ZN(n11291) );
  AOI211_X1 U13657 ( .C1(n12864), .C2(n11293), .A(n11292), .B(n11291), .ZN(
        n11298) );
  AND3_X1 U13658 ( .A1(n11618), .A2(n11295), .A3(n11294), .ZN(n11296) );
  OAI21_X1 U13659 ( .B1(n11296), .B2(n11576), .A(n12890), .ZN(n11297) );
  OAI211_X1 U13660 ( .C1(n12881), .C2(n11299), .A(n11298), .B(n11297), .ZN(
        P3_U3184) );
  INV_X1 U13661 ( .A(n11300), .ZN(n11303) );
  OAI222_X1 U13662 ( .A1(n11891), .A2(n11303), .B1(n11887), .B2(n11302), .C1(
        P3_U3151), .C2(n11301), .ZN(P3_U3269) );
  XNOR2_X1 U13663 ( .A(n11304), .B(n11441), .ZN(n15272) );
  NAND2_X1 U13664 ( .A1(n15272), .A2(n15201), .ZN(n11314) );
  INV_X1 U13665 ( .A(n11305), .ZN(n11306) );
  NAND2_X1 U13666 ( .A1(n15217), .A2(n11306), .ZN(n15219) );
  NAND2_X1 U13667 ( .A1(n15219), .A2(n11307), .ZN(n11308) );
  XNOR2_X1 U13668 ( .A(n11308), .B(n11441), .ZN(n11312) );
  NAND2_X1 U13669 ( .A1(n12689), .A2(n15212), .ZN(n11310) );
  NAND2_X1 U13670 ( .A1(n12688), .A2(n15215), .ZN(n11309) );
  NAND2_X1 U13671 ( .A1(n11310), .A2(n11309), .ZN(n11311) );
  AOI21_X1 U13672 ( .B1(n11312), .B2(n15218), .A(n11311), .ZN(n11313) );
  AND2_X1 U13673 ( .A1(n11314), .A2(n11313), .ZN(n15274) );
  NOR2_X1 U13674 ( .A1(n11522), .A2(n15281), .ZN(n15271) );
  INV_X1 U13675 ( .A(n11529), .ZN(n11315) );
  AOI22_X1 U13676 ( .A1(n15228), .A2(n15271), .B1(n15244), .B2(n11315), .ZN(
        n11316) );
  OAI21_X1 U13677 ( .B1(n11111), .B2(n15248), .A(n11316), .ZN(n11317) );
  AOI21_X1 U13678 ( .B1(n15272), .B2(n15246), .A(n11317), .ZN(n11318) );
  OAI21_X1 U13679 ( .B1(n15274), .B2(n15250), .A(n11318), .ZN(P3_U3226) );
  OR2_X1 U13680 ( .A1(n14905), .A2(n14922), .ZN(n11319) );
  NAND2_X1 U13681 ( .A1(n11320), .A2(n11319), .ZN(n11326) );
  NAND2_X1 U13682 ( .A1(n11321), .A2(n6429), .ZN(n11324) );
  AOI22_X1 U13683 ( .A1(n12023), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11322), 
        .B2(n12022), .ZN(n11323) );
  XNOR2_X1 U13684 ( .A(n14547), .B(n14910), .ZN(n12013) );
  INV_X1 U13685 ( .A(n12013), .ZN(n11325) );
  NAND2_X1 U13686 ( .A1(n11326), .A2(n11325), .ZN(n11484) );
  OAI21_X1 U13687 ( .B1(n11326), .B2(n11325), .A(n11484), .ZN(n14549) );
  AOI21_X1 U13688 ( .B1(n11327), .B2(n14547), .A(n14640), .ZN(n11328) );
  AND2_X1 U13689 ( .A1(n11328), .A2(n11537), .ZN(n14550) );
  NAND2_X1 U13690 ( .A1(n11329), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11477) );
  OR2_X1 U13691 ( .A1(n11329), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11330) );
  AND2_X1 U13692 ( .A1(n11477), .A2(n11330), .ZN(n14042) );
  NAND2_X1 U13693 ( .A1(n11974), .A2(n14042), .ZN(n11334) );
  NAND2_X1 U13694 ( .A1(n12059), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11333) );
  INV_X2 U13695 ( .A(n11900), .ZN(n12060) );
  NAND2_X1 U13696 ( .A1(n12060), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U13697 ( .A1(n12061), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U13698 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n14924) );
  INV_X1 U13699 ( .A(n14924), .ZN(n11470) );
  OR2_X1 U13700 ( .A1(n14905), .A2(n12276), .ZN(n11335) );
  XNOR2_X1 U13701 ( .A(n11463), .B(n12013), .ZN(n11337) );
  OAI222_X1 U13702 ( .A1(n14527), .A2(n11470), .B1(n14525), .B2(n12276), .C1(
        n11337), .C2(n14936), .ZN(n14542) );
  AOI211_X1 U13703 ( .C1(n15108), .C2(n14549), .A(n14550), .B(n14542), .ZN(
        n11342) );
  INV_X1 U13704 ( .A(n14547), .ZN(n14928) );
  INV_X1 U13705 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11338) );
  OAI22_X1 U13706 ( .A1(n14928), .A2(n14683), .B1(n14655), .B2(n11338), .ZN(
        n11339) );
  INV_X1 U13707 ( .A(n11339), .ZN(n11340) );
  OAI21_X1 U13708 ( .B1(n11342), .B2(n15109), .A(n11340), .ZN(P1_U3492) );
  AOI22_X1 U13709 ( .A1(n14547), .A2(n11847), .B1(n15120), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11341) );
  OAI21_X1 U13710 ( .B1(n11342), .B2(n15120), .A(n11341), .ZN(P1_U3539) );
  NAND2_X1 U13711 ( .A1(n11412), .A2(n11343), .ZN(n11344) );
  INV_X1 U13712 ( .A(n11358), .ZN(n11348) );
  NAND3_X1 U13713 ( .A1(n11418), .A2(n11348), .A3(n11347), .ZN(n11349) );
  NAND3_X1 U13714 ( .A1(n11668), .A2(n13822), .A3(n11349), .ZN(n11352) );
  INV_X1 U13715 ( .A(n13477), .ZN(n11698) );
  OAI22_X1 U13716 ( .A1(n11698), .A2(n13455), .B1(n11350), .B2(n13640), .ZN(
        n11556) );
  INV_X1 U13717 ( .A(n11556), .ZN(n11351) );
  NAND2_X1 U13718 ( .A1(n11352), .A2(n11351), .ZN(n11544) );
  INV_X1 U13719 ( .A(n11544), .ZN(n11366) );
  OR2_X1 U13720 ( .A1(n11412), .A2(n13480), .ZN(n11353) );
  NAND2_X1 U13721 ( .A1(n11412), .A2(n13480), .ZN(n11355) );
  AND2_X1 U13722 ( .A1(n13847), .A2(n13479), .ZN(n11356) );
  OR2_X1 U13723 ( .A1(n13847), .A2(n13479), .ZN(n11357) );
  XOR2_X1 U13724 ( .A(n11358), .B(n11677), .Z(n11546) );
  NAND2_X1 U13725 ( .A1(n11546), .A2(n13848), .ZN(n11365) );
  INV_X1 U13726 ( .A(n11672), .ZN(n11361) );
  AOI211_X1 U13727 ( .C1(n11678), .C2(n11416), .A(n9680), .B(n11361), .ZN(
        n11545) );
  NOR2_X1 U13728 ( .A1(n11359), .A2(n13816), .ZN(n11363) );
  OAI22_X1 U13729 ( .A1(n13844), .A2(n11260), .B1(n11558), .B2(n13841), .ZN(
        n11362) );
  AOI211_X1 U13730 ( .C1(n11545), .C2(n13850), .A(n11363), .B(n11362), .ZN(
        n11364) );
  OAI211_X1 U13731 ( .C1(n11366), .C2(n6430), .A(n11365), .B(n11364), .ZN(
        P2_U3252) );
  INV_X1 U13732 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11834) );
  NOR2_X1 U13733 ( .A1(n11835), .A2(n11834), .ZN(n11367) );
  AOI21_X1 U13734 ( .B1(n11834), .B2(n11835), .A(n11367), .ZN(n11371) );
  INV_X1 U13735 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11369) );
  OAI21_X1 U13736 ( .B1(n11373), .B2(n11369), .A(n11368), .ZN(n11370) );
  NAND2_X1 U13737 ( .A1(n11371), .A2(n11370), .ZN(n11833) );
  OAI211_X1 U13738 ( .C1(n11371), .C2(n11370), .A(n14243), .B(n11833), .ZN(
        n11380) );
  NAND2_X1 U13739 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14075)
         );
  XNOR2_X1 U13740 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n11835), .ZN(n11376) );
  INV_X1 U13741 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11374) );
  OAI21_X1 U13742 ( .B1(n11374), .B2(n11373), .A(n11372), .ZN(n11375) );
  NAND2_X1 U13743 ( .A1(n11376), .A2(n11375), .ZN(n11836) );
  OAI211_X1 U13744 ( .C1(n11376), .C2(n11375), .A(n11836), .B(n14245), .ZN(
        n11377) );
  NAND2_X1 U13745 ( .A1(n14075), .A2(n11377), .ZN(n11378) );
  AOI21_X1 U13746 ( .B1(n14977), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11378), 
        .ZN(n11379) );
  OAI211_X1 U13747 ( .C1(n14992), .C2(n11835), .A(n11380), .B(n11379), .ZN(
        P1_U3260) );
  INV_X1 U13748 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12029) );
  OAI222_X1 U13749 ( .A1(P1_U3086), .A2(n12075), .B1(n14707), .B2(n11381), 
        .C1(n12029), .C2(n14701), .ZN(P1_U3334) );
  INV_X1 U13750 ( .A(n11382), .ZN(n11383) );
  NOR2_X1 U13751 ( .A1(n11384), .A2(n11383), .ZN(n11386) );
  XNOR2_X1 U13752 ( .A(n11709), .B(n11394), .ZN(n11385) );
  AOI21_X1 U13753 ( .B1(n11386), .B2(n11385), .A(n11710), .ZN(n11400) );
  AOI21_X1 U13754 ( .B1(n7879), .B2(n11388), .A(n11705), .ZN(n11391) );
  AND2_X1 U13755 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12637) );
  AOI21_X1 U13756 ( .B1(n15191), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12637), 
        .ZN(n11390) );
  INV_X1 U13757 ( .A(n11394), .ZN(n11717) );
  NAND2_X1 U13758 ( .A1(n12859), .A2(n11717), .ZN(n11389) );
  OAI211_X1 U13759 ( .C1(n11391), .C2(n12892), .A(n11390), .B(n11389), .ZN(
        n11398) );
  AOI21_X1 U13760 ( .B1(n7880), .B2(n11395), .A(n11718), .ZN(n11396) );
  NOR2_X1 U13761 ( .A1(n11396), .A2(n12888), .ZN(n11397) );
  NOR2_X1 U13762 ( .A1(n11398), .A2(n11397), .ZN(n11399) );
  OAI21_X1 U13763 ( .B1(n11400), .B2(n12868), .A(n11399), .ZN(P3_U3193) );
  NAND2_X1 U13764 ( .A1(n13449), .A2(n11401), .ZN(n11403) );
  OAI211_X1 U13765 ( .C1(n13447), .C2(n11404), .A(n11403), .B(n11402), .ZN(
        n11411) );
  NAND2_X1 U13766 ( .A1(n13480), .A2(n13343), .ZN(n11427) );
  XNOR2_X1 U13767 ( .A(n11412), .B(n9828), .ZN(n11429) );
  XOR2_X1 U13768 ( .A(n11427), .B(n11429), .Z(n11409) );
  INV_X1 U13769 ( .A(n11405), .ZN(n11406) );
  AOI211_X1 U13770 ( .C1(n11409), .C2(n11408), .A(n13470), .B(n11428), .ZN(
        n11410) );
  AOI211_X1 U13771 ( .C1(n11412), .C2(n9631), .A(n11411), .B(n11410), .ZN(
        n11413) );
  INV_X1 U13772 ( .A(n11413), .ZN(P2_U3208) );
  XNOR2_X1 U13773 ( .A(n11414), .B(n11420), .ZN(n13849) );
  AOI21_X1 U13774 ( .B1(n13847), .B2(n11415), .A(n9680), .ZN(n11417) );
  AND2_X1 U13775 ( .A1(n11417), .A2(n11416), .ZN(n13851) );
  OAI211_X1 U13776 ( .C1(n11420), .C2(n11419), .A(n11418), .B(n13822), .ZN(
        n11421) );
  AOI22_X1 U13777 ( .A1(n13478), .A2(n13570), .B1(n13464), .B2(n13480), .ZN(
        n11436) );
  NAND2_X1 U13778 ( .A1(n11421), .A2(n11436), .ZN(n13839) );
  AOI211_X1 U13779 ( .C1(n13849), .C2(n13905), .A(n13851), .B(n13839), .ZN(
        n11426) );
  AOI22_X1 U13780 ( .A1(n13847), .A2(n13899), .B1(n15188), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11422) );
  OAI21_X1 U13781 ( .B1(n11426), .B2(n15188), .A(n11422), .ZN(P2_U3511) );
  INV_X1 U13782 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11423) );
  NOR2_X1 U13783 ( .A1(n15187), .A2(n11423), .ZN(n11424) );
  AOI21_X1 U13784 ( .B1(n13847), .B2(n13965), .A(n11424), .ZN(n11425) );
  OAI21_X1 U13785 ( .B1(n11426), .B2(n15185), .A(n11425), .ZN(P2_U3466) );
  INV_X1 U13786 ( .A(n11427), .ZN(n11430) );
  XNOR2_X1 U13787 ( .A(n13847), .B(n9828), .ZN(n11432) );
  AND2_X1 U13788 ( .A1(n13479), .A2(n13687), .ZN(n11431) );
  NOR2_X1 U13789 ( .A1(n11432), .A2(n11431), .ZN(n11553) );
  INV_X1 U13790 ( .A(n11553), .ZN(n11433) );
  NAND2_X1 U13791 ( .A1(n11432), .A2(n11431), .ZN(n11552) );
  NAND2_X1 U13792 ( .A1(n11433), .A2(n11552), .ZN(n11434) );
  XNOR2_X1 U13793 ( .A(n11554), .B(n11434), .ZN(n11440) );
  OAI22_X1 U13794 ( .A1(n13447), .A2(n11436), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11435), .ZN(n11437) );
  AOI21_X1 U13795 ( .B1(n13840), .B2(n13449), .A(n11437), .ZN(n11439) );
  NAND2_X1 U13796 ( .A1(n13847), .A2(n9631), .ZN(n11438) );
  OAI211_X1 U13797 ( .C1(n11440), .C2(n13470), .A(n11439), .B(n11438), .ZN(
        P2_U3196) );
  XNOR2_X1 U13798 ( .A(n12543), .B(n15282), .ZN(n11562) );
  XNOR2_X1 U13799 ( .A(n11562), .B(n15196), .ZN(n11456) );
  INV_X2 U13800 ( .A(n12503), .ZN(n12543) );
  XNOR2_X1 U13801 ( .A(n11441), .B(n12543), .ZN(n11729) );
  OAI211_X1 U13802 ( .C1(n11446), .C2(n12689), .A(n11729), .B(n11442), .ZN(
        n11443) );
  XNOR2_X1 U13803 ( .A(n10859), .B(n11735), .ZN(n11447) );
  XNOR2_X1 U13804 ( .A(n11447), .B(n12688), .ZN(n11731) );
  NOR2_X1 U13805 ( .A1(n11443), .A2(n11731), .ZN(n11444) );
  NAND2_X1 U13806 ( .A1(n11445), .A2(n11444), .ZN(n11451) );
  NAND2_X1 U13807 ( .A1(n11446), .A2(n12689), .ZN(n11517) );
  OAI21_X1 U13808 ( .B1(n11731), .B2(n11517), .A(n11729), .ZN(n11449) );
  INV_X1 U13809 ( .A(n11729), .ZN(n11519) );
  OAI21_X1 U13810 ( .B1(n11731), .B2(n11734), .A(n11519), .ZN(n11448) );
  AOI22_X1 U13811 ( .A1(n11449), .A2(n11448), .B1(n11447), .B2(n12688), .ZN(
        n11450) );
  NAND2_X1 U13812 ( .A1(n11451), .A2(n11450), .ZN(n11455) );
  INV_X1 U13813 ( .A(n11566), .ZN(n11454) );
  AOI21_X1 U13814 ( .B1(n11456), .B2(n11455), .A(n11454), .ZN(n11462) );
  INV_X1 U13815 ( .A(n12688), .ZN(n11524) );
  OAI22_X1 U13816 ( .A1(n15282), .A2(n12652), .B1(n12659), .B2(n11524), .ZN(
        n11457) );
  AOI211_X1 U13817 ( .C1(n12655), .C2(n12635), .A(n11458), .B(n11457), .ZN(
        n11461) );
  INV_X1 U13818 ( .A(n11606), .ZN(n11459) );
  NAND2_X1 U13819 ( .A1(n12656), .A2(n11459), .ZN(n11460) );
  OAI211_X1 U13820 ( .C1(n11462), .C2(n12674), .A(n11461), .B(n11460), .ZN(
        P3_U3171) );
  NAND2_X1 U13821 ( .A1(n11463), .A2(n12013), .ZN(n11465) );
  INV_X1 U13822 ( .A(n14910), .ZN(n12281) );
  OR2_X1 U13823 ( .A1(n14547), .A2(n12281), .ZN(n11464) );
  NAND2_X1 U13824 ( .A1(n11466), .A2(n6429), .ZN(n11469) );
  AOI22_X1 U13825 ( .A1(n11467), .A2(n12022), .B1(n12023), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11468) );
  XNOR2_X1 U13826 ( .A(n12291), .B(n14924), .ZN(n12015) );
  OR2_X1 U13827 ( .A1(n12291), .A2(n11470), .ZN(n11471) );
  NAND2_X1 U13828 ( .A1(n11472), .A2(n6429), .ZN(n11475) );
  AOI22_X1 U13829 ( .A1(n11473), .A2(n12022), .B1(n12023), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11474) );
  INV_X1 U13830 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U13831 ( .A1(n11477), .A2(n11476), .ZN(n11478) );
  AND2_X1 U13832 ( .A1(n11488), .A2(n11478), .ZN(n14102) );
  NAND2_X1 U13833 ( .A1(n11974), .A2(n14102), .ZN(n11482) );
  NAND2_X1 U13834 ( .A1(n12059), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U13835 ( .A1(n12061), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U13836 ( .A1(n12060), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U13837 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n14897) );
  INV_X1 U13838 ( .A(n14897), .ZN(n12299) );
  XNOR2_X1 U13839 ( .A(n12301), .B(n12299), .ZN(n12018) );
  XNOR2_X1 U13840 ( .A(n11760), .B(n12018), .ZN(n11634) );
  INV_X1 U13841 ( .A(n11634), .ZN(n11505) );
  OR2_X1 U13842 ( .A1(n14547), .A2(n14910), .ZN(n11483) );
  INV_X1 U13843 ( .A(n12015), .ZN(n11531) );
  OAI21_X1 U13844 ( .B1(n11485), .B2(n12018), .A(n11768), .ZN(n11630) );
  AOI21_X1 U13845 ( .B1(n12301), .B2(n11536), .A(n14640), .ZN(n11486) );
  NAND2_X1 U13846 ( .A1(n11486), .A2(n11770), .ZN(n11631) );
  INV_X1 U13847 ( .A(n14102), .ZN(n11497) );
  INV_X1 U13848 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U13849 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  NAND2_X1 U13850 ( .A1(n11773), .A2(n11489), .ZN(n14904) );
  INV_X1 U13851 ( .A(n14904), .ZN(n11490) );
  NAND2_X1 U13852 ( .A1(n11974), .A2(n11490), .ZN(n11494) );
  NAND2_X1 U13853 ( .A1(n12059), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U13854 ( .A1(n10484), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U13855 ( .A1(n12061), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11491) );
  OR2_X1 U13856 ( .A1(n12306), .A2(n14527), .ZN(n11496) );
  NAND2_X1 U13857 ( .A1(n14924), .A2(n15007), .ZN(n11495) );
  AND2_X1 U13858 ( .A1(n11496), .A2(n11495), .ZN(n14100) );
  OAI21_X1 U13859 ( .B1(n14544), .B2(n11497), .A(n14100), .ZN(n11498) );
  INV_X1 U13860 ( .A(n11498), .ZN(n11500) );
  NAND2_X1 U13861 ( .A1(n15022), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11499) );
  OAI21_X1 U13862 ( .B1(n15022), .B2(n11500), .A(n11499), .ZN(n11501) );
  AOI21_X1 U13863 ( .B1(n12301), .B2(n14546), .A(n11501), .ZN(n11502) );
  OAI21_X1 U13864 ( .B1(n11631), .B2(n14537), .A(n11502), .ZN(n11503) );
  AOI21_X1 U13865 ( .B1(n11630), .B2(n14548), .A(n11503), .ZN(n11504) );
  OAI21_X1 U13866 ( .B1(n14441), .B2(n11505), .A(n11504), .ZN(P1_U3280) );
  AOI22_X1 U13867 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n13530), .B1(n13537), 
        .B2(n13831), .ZN(n11508) );
  OAI21_X1 U13868 ( .B1(n11508), .B2(n11507), .A(n13532), .ZN(n11516) );
  NAND2_X1 U13869 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13420)
         );
  OAI21_X1 U13870 ( .B1(n15143), .B2(n13537), .A(n13420), .ZN(n11509) );
  AOI21_X1 U13871 ( .B1(n15154), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n11509), 
        .ZN(n11515) );
  XNOR2_X1 U13872 ( .A(n13537), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11513) );
  OAI21_X1 U13873 ( .B1(n11511), .B2(n11877), .A(n11510), .ZN(n11512) );
  NAND2_X1 U13874 ( .A1(n11513), .A2(n11512), .ZN(n13535) );
  OAI211_X1 U13875 ( .C1(n11513), .C2(n11512), .A(n15161), .B(n13535), .ZN(
        n11514) );
  OAI211_X1 U13876 ( .C1(n11516), .C2(n15129), .A(n11515), .B(n11514), .ZN(
        P2_U3231) );
  NAND2_X1 U13877 ( .A1(n11518), .A2(n11517), .ZN(n11730) );
  XNOR2_X1 U13878 ( .A(n11730), .B(n11519), .ZN(n11520) );
  NAND2_X1 U13879 ( .A1(n11520), .A2(n12644), .ZN(n11528) );
  OAI22_X1 U13880 ( .A1(n12652), .A2(n11522), .B1(n12659), .B2(n11521), .ZN(
        n11526) );
  OAI21_X1 U13881 ( .B1(n12666), .B2(n11524), .A(n11523), .ZN(n11525) );
  NOR2_X1 U13882 ( .A1(n11526), .A2(n11525), .ZN(n11527) );
  OAI211_X1 U13883 ( .C1(n11529), .C2(n12670), .A(n11528), .B(n11527), .ZN(
        P3_U3153) );
  OAI21_X1 U13884 ( .B1(n11532), .B2(n11531), .A(n11530), .ZN(n11642) );
  INV_X1 U13885 ( .A(n11642), .ZN(n11543) );
  XNOR2_X1 U13886 ( .A(n11533), .B(n12015), .ZN(n11535) );
  NAND2_X1 U13887 ( .A1(n11642), .A2(n15068), .ZN(n11534) );
  AOI22_X1 U13888 ( .A1(n14509), .A2(n14897), .B1(n15007), .B2(n14910), .ZN(
        n14040) );
  OAI211_X1 U13889 ( .C1(n14936), .C2(n11535), .A(n11534), .B(n14040), .ZN(
        n11640) );
  NAND2_X1 U13890 ( .A1(n11640), .A2(n14541), .ZN(n11541) );
  AOI211_X1 U13891 ( .C1(n12291), .C2(n11537), .A(n14640), .B(n7283), .ZN(
        n11641) );
  AOI22_X1 U13892 ( .A1(n15022), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14042), 
        .B2(n15013), .ZN(n11538) );
  OAI21_X1 U13893 ( .B1(n6840), .B2(n15012), .A(n11538), .ZN(n11539) );
  AOI21_X1 U13894 ( .B1(n11641), .B2(n15018), .A(n11539), .ZN(n11540) );
  OAI211_X1 U13895 ( .C1(n11543), .C2(n11542), .A(n11541), .B(n11540), .ZN(
        P1_U3281) );
  AOI211_X1 U13896 ( .C1(n11546), .C2(n13905), .A(n11545), .B(n11544), .ZN(
        n11551) );
  AOI22_X1 U13897 ( .A1(n11678), .A2(n13899), .B1(n15188), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11547) );
  OAI21_X1 U13898 ( .B1(n11551), .B2(n15188), .A(n11547), .ZN(P2_U3512) );
  INV_X1 U13899 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11548) );
  NOR2_X1 U13900 ( .A1(n15187), .A2(n11548), .ZN(n11549) );
  AOI21_X1 U13901 ( .B1(n11678), .B2(n13965), .A(n11549), .ZN(n11550) );
  OAI21_X1 U13902 ( .B1(n11551), .B2(n15185), .A(n11550), .ZN(P2_U3469) );
  XNOR2_X1 U13903 ( .A(n11678), .B(n9828), .ZN(n11816) );
  NAND2_X1 U13904 ( .A1(n13478), .A2(n13343), .ZN(n11815) );
  XNOR2_X1 U13905 ( .A(n11816), .B(n11815), .ZN(n11818) );
  XNOR2_X1 U13906 ( .A(n11819), .B(n11818), .ZN(n11561) );
  NOR2_X1 U13907 ( .A1(n11555), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15140) );
  AOI21_X1 U13908 ( .B1(n14885), .B2(n11556), .A(n15140), .ZN(n11557) );
  OAI21_X1 U13909 ( .B1(n11558), .B2(n14891), .A(n11557), .ZN(n11559) );
  AOI21_X1 U13910 ( .B1(n11678), .B2(n9631), .A(n11559), .ZN(n11560) );
  OAI21_X1 U13911 ( .B1(n11561), .B2(n13470), .A(n11560), .ZN(P2_U3206) );
  INV_X1 U13912 ( .A(n11562), .ZN(n11563) );
  INV_X1 U13913 ( .A(n15196), .ZN(n11738) );
  NAND2_X1 U13914 ( .A1(n11563), .A2(n11738), .ZN(n11564) );
  AND2_X1 U13915 ( .A1(n11566), .A2(n11564), .ZN(n11568) );
  INV_X1 U13916 ( .A(n15205), .ZN(n15288) );
  XNOR2_X1 U13917 ( .A(n12543), .B(n15288), .ZN(n12465) );
  XNOR2_X1 U13918 ( .A(n12465), .B(n12635), .ZN(n11567) );
  AND2_X1 U13919 ( .A1(n11567), .A2(n11564), .ZN(n11565) );
  OAI211_X1 U13920 ( .C1(n11568), .C2(n11567), .A(n12644), .B(n12468), .ZN(
        n11573) );
  OAI22_X1 U13921 ( .A1(n15205), .A2(n12652), .B1(n12659), .B2(n11738), .ZN(
        n11571) );
  INV_X1 U13922 ( .A(n15197), .ZN(n12633) );
  OAI21_X1 U13923 ( .B1(n12666), .B2(n12633), .A(n11569), .ZN(n11570) );
  NOR2_X1 U13924 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  OAI211_X1 U13925 ( .C1(n15210), .C2(n12670), .A(n11573), .B(n11572), .ZN(
        P3_U3157) );
  INV_X1 U13926 ( .A(n11574), .ZN(n11575) );
  OAI222_X1 U13927 ( .A1(n13999), .A2(n15351), .B1(n14001), .B2(n11575), .C1(
        n8482), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13928 ( .A(n11576), .ZN(n11579) );
  NAND3_X1 U13929 ( .A1(n11579), .A2(n11578), .A3(n11577), .ZN(n11580) );
  AOI21_X1 U13930 ( .B1(n11581), .B2(n11580), .A(n12868), .ZN(n11593) );
  NAND2_X1 U13931 ( .A1(n11582), .A2(n11090), .ZN(n11583) );
  AND2_X1 U13932 ( .A1(n11584), .A2(n11583), .ZN(n11591) );
  NAND2_X1 U13933 ( .A1(n11585), .A2(n11091), .ZN(n11586) );
  NAND2_X1 U13934 ( .A1(n11587), .A2(n11586), .ZN(n11588) );
  NAND2_X1 U13935 ( .A1(n12835), .A2(n11588), .ZN(n11590) );
  AOI22_X1 U13936 ( .A1(n15191), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11589) );
  OAI211_X1 U13937 ( .C1(n11591), .C2(n12892), .A(n11590), .B(n11589), .ZN(
        n11592) );
  AOI211_X1 U13938 ( .C1(n12859), .C2(n7384), .A(n11593), .B(n11592), .ZN(
        n11594) );
  INV_X1 U13939 ( .A(n11594), .ZN(P3_U3185) );
  INV_X1 U13940 ( .A(n11600), .ZN(n11602) );
  XNOR2_X1 U13941 ( .A(n11595), .B(n11602), .ZN(n15280) );
  AOI22_X1 U13942 ( .A1(n15212), .A2(n12688), .B1(n12635), .B2(n15215), .ZN(
        n11605) );
  AND2_X1 U13943 ( .A1(n12688), .A2(n11596), .ZN(n11598) );
  OR2_X1 U13944 ( .A1(n12688), .A2(n11596), .ZN(n11597) );
  INV_X1 U13945 ( .A(n11601), .ZN(n11603) );
  OAI211_X1 U13946 ( .C1(n11603), .C2(n11602), .A(n15218), .B(n12423), .ZN(
        n11604) );
  OAI211_X1 U13947 ( .C1(n15280), .C2(n15223), .A(n11605), .B(n11604), .ZN(
        n15283) );
  NAND2_X1 U13948 ( .A1(n15283), .A2(n15248), .ZN(n11609) );
  OAI22_X1 U13949 ( .A1(n15248), .A2(n11162), .B1(n11606), .B2(n15234), .ZN(
        n11607) );
  AOI21_X1 U13950 ( .B1(n13107), .B2(n12421), .A(n11607), .ZN(n11608) );
  OAI211_X1 U13951 ( .C1(n15280), .C2(n12945), .A(n11609), .B(n11608), .ZN(
        P3_U3224) );
  INV_X1 U13952 ( .A(n11610), .ZN(n11612) );
  INV_X1 U13953 ( .A(SI_27_), .ZN(n11611) );
  OAI21_X1 U13954 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n11614), .A(n11613), .ZN(
        n11627) );
  INV_X1 U13955 ( .A(n11615), .ZN(n11616) );
  AOI21_X1 U13956 ( .B1(n11079), .B2(n11617), .A(n11616), .ZN(n11623) );
  INV_X1 U13957 ( .A(n11618), .ZN(n11619) );
  AOI21_X1 U13958 ( .B1(n11621), .B2(n11620), .A(n11619), .ZN(n11622) );
  OAI22_X1 U13959 ( .A1(n12888), .A2(n11623), .B1(n11622), .B2(n12868), .ZN(
        n11626) );
  OAI22_X1 U13960 ( .A1(n12849), .A2(n14715), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11624), .ZN(n11625) );
  AOI211_X1 U13961 ( .C1(n12864), .C2(n11627), .A(n11626), .B(n11625), .ZN(
        n11628) );
  OAI21_X1 U13962 ( .B1(n11629), .B2(n12881), .A(n11628), .ZN(P3_U3183) );
  INV_X1 U13963 ( .A(n11630), .ZN(n11632) );
  OAI211_X1 U13964 ( .C1(n11632), .C2(n15074), .A(n14100), .B(n11631), .ZN(
        n11633) );
  AOI21_X1 U13965 ( .B1(n11634), .B2(n15079), .A(n11633), .ZN(n11639) );
  INV_X1 U13966 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11635) );
  OAI22_X1 U13967 ( .A1(n7282), .A2(n14683), .B1(n14655), .B2(n11635), .ZN(
        n11636) );
  INV_X1 U13968 ( .A(n11636), .ZN(n11637) );
  OAI21_X1 U13969 ( .B1(n11639), .B2(n15109), .A(n11637), .ZN(P1_U3498) );
  AOI22_X1 U13970 ( .A1(n12301), .A2(n11847), .B1(n15120), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11638) );
  OAI21_X1 U13971 ( .B1(n11639), .B2(n15120), .A(n11638), .ZN(P1_U3541) );
  AOI211_X1 U13972 ( .C1(n15098), .C2(n11642), .A(n11641), .B(n11640), .ZN(
        n11647) );
  AOI22_X1 U13973 ( .A1(n12291), .A2(n11847), .B1(n15120), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11643) );
  OAI21_X1 U13974 ( .B1(n11647), .B2(n15120), .A(n11643), .ZN(P1_U3540) );
  INV_X1 U13975 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11644) );
  OAI22_X1 U13976 ( .A1(n6840), .A2(n14683), .B1(n14655), .B2(n11644), .ZN(
        n11645) );
  INV_X1 U13977 ( .A(n11645), .ZN(n11646) );
  OAI21_X1 U13978 ( .B1(n11647), .B2(n15109), .A(n11646), .ZN(P1_U3495) );
  INV_X1 U13979 ( .A(n11649), .ZN(n11648) );
  AND2_X1 U13980 ( .A1(n12890), .A2(n11648), .ZN(n11653) );
  NAND3_X1 U13981 ( .A1(n12892), .A2(n12888), .A3(n12868), .ZN(n11650) );
  NAND2_X1 U13982 ( .A1(n11650), .A2(n11649), .ZN(n11651) );
  NAND2_X1 U13983 ( .A1(n11651), .A2(n12881), .ZN(n11652) );
  MUX2_X1 U13984 ( .A(n11653), .B(n11652), .S(P3_IR_REG_0__SCAN_IN), .Z(n11660) );
  NAND2_X1 U13985 ( .A1(n12835), .A2(n11654), .ZN(n11657) );
  NOR2_X1 U13986 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10407), .ZN(n11655) );
  AOI21_X1 U13987 ( .B1(n15191), .B2(P3_ADDR_REG_0__SCAN_IN), .A(n11655), .ZN(
        n11656) );
  OAI211_X1 U13988 ( .C1(n11658), .C2(n12892), .A(n11657), .B(n11656), .ZN(
        n11659) );
  OR2_X1 U13989 ( .A1(n11660), .A2(n11659), .ZN(P3_U3182) );
  INV_X1 U13990 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U13991 ( .A1(n11941), .A2(n11661), .ZN(n11662) );
  OAI211_X1 U13992 ( .C1(n11942), .C2(n14709), .A(n11662), .B(n12256), .ZN(
        P1_U3332) );
  NAND2_X1 U13993 ( .A1(n11941), .A2(n11663), .ZN(n11665) );
  OAI211_X1 U13994 ( .C1(n11666), .C2(n13999), .A(n11665), .B(n11664), .ZN(
        P2_U3304) );
  INV_X1 U13995 ( .A(n13478), .ZN(n11669) );
  OR2_X1 U13996 ( .A1(n11678), .A2(n11669), .ZN(n11667) );
  XOR2_X1 U13997 ( .A(n11695), .B(n11680), .Z(n11670) );
  OAI22_X1 U13998 ( .A1(n11854), .A2(n13455), .B1(n11669), .B2(n13640), .ZN(
        n14886) );
  AOI21_X1 U13999 ( .B1(n11670), .B2(n13822), .A(n14886), .ZN(n13936) );
  INV_X1 U14000 ( .A(n11689), .ZN(n11671) );
  AOI211_X1 U14001 ( .C1(n14887), .C2(n11672), .A(n13687), .B(n11671), .ZN(
        n13934) );
  INV_X1 U14002 ( .A(n14887), .ZN(n11675) );
  INV_X1 U14003 ( .A(n14890), .ZN(n11673) );
  AOI22_X1 U14004 ( .A1(n6430), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11673), 
        .B2(n13828), .ZN(n11674) );
  OAI21_X1 U14005 ( .B1(n11675), .B2(n13816), .A(n11674), .ZN(n11682) );
  NOR2_X1 U14006 ( .A1(n11678), .A2(n13478), .ZN(n11676) );
  NAND2_X1 U14007 ( .A1(n11678), .A2(n13478), .ZN(n11679) );
  XOR2_X1 U14008 ( .A(n11680), .B(n11685), .Z(n13937) );
  NOR2_X1 U14009 ( .A1(n13937), .A2(n13835), .ZN(n11681) );
  AOI211_X1 U14010 ( .C1(n13934), .C2(n13850), .A(n11682), .B(n11681), .ZN(
        n11683) );
  OAI21_X1 U14011 ( .B1(n6430), .B2(n13936), .A(n11683), .ZN(P2_U3251) );
  NAND2_X1 U14012 ( .A1(n11685), .A2(n11684), .ZN(n11687) );
  NAND2_X1 U14013 ( .A1(n11687), .A2(n11686), .ZN(n11862) );
  XNOR2_X1 U14014 ( .A(n11862), .B(n11861), .ZN(n11811) );
  INV_X1 U14015 ( .A(n11811), .ZN(n11703) );
  AOI211_X1 U14016 ( .C1(n11863), .C2(n11689), .A(n9680), .B(n6577), .ZN(
        n11810) );
  INV_X1 U14017 ( .A(n11863), .ZN(n11690) );
  NOR2_X1 U14018 ( .A1(n11690), .A2(n13816), .ZN(n11693) );
  INV_X1 U14019 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11691) );
  OAI22_X1 U14020 ( .A1(n13844), .A2(n11691), .B1(n11829), .B2(n13841), .ZN(
        n11692) );
  AOI211_X1 U14021 ( .C1(n11810), .C2(n13850), .A(n11693), .B(n11692), .ZN(
        n11702) );
  NAND2_X1 U14022 ( .A1(n14887), .A2(n11698), .ZN(n11694) );
  NAND2_X1 U14023 ( .A1(n11695), .A2(n11694), .ZN(n11697) );
  OR2_X1 U14024 ( .A1(n14887), .A2(n11698), .ZN(n11696) );
  XNOR2_X1 U14025 ( .A(n11853), .B(n11861), .ZN(n11700) );
  OAI22_X1 U14026 ( .A1(n13606), .A2(n13455), .B1(n11698), .B2(n13640), .ZN(
        n11827) );
  INV_X1 U14027 ( .A(n11827), .ZN(n11699) );
  OAI21_X1 U14028 ( .B1(n11700), .B2(n13795), .A(n11699), .ZN(n11809) );
  NAND2_X1 U14029 ( .A1(n11809), .A2(n13844), .ZN(n11701) );
  OAI211_X1 U14030 ( .C1(n11703), .C2(n13835), .A(n11702), .B(n11701), .ZN(
        P2_U3250) );
  NOR2_X1 U14031 ( .A1(n11717), .A2(n11704), .ZN(n11706) );
  NAND2_X1 U14032 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12739), .ZN(n12753) );
  OAI21_X1 U14033 ( .B1(n12739), .B2(P3_REG1_REG_12__SCAN_IN), .A(n12753), 
        .ZN(n11707) );
  AOI21_X1 U14034 ( .B1(n11708), .B2(n11707), .A(n12751), .ZN(n11728) );
  INV_X1 U14035 ( .A(n11709), .ZN(n11711) );
  XNOR2_X1 U14036 ( .A(n12740), .B(n11725), .ZN(n11712) );
  OAI211_X1 U14037 ( .C1(n11713), .C2(n11712), .A(n12743), .B(n12890), .ZN(
        n11727) );
  INV_X1 U14038 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n11715) );
  OR2_X1 U14039 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11714), .ZN(n12562) );
  OAI21_X1 U14040 ( .B1(n12849), .B2(n11715), .A(n12562), .ZN(n11724) );
  NOR2_X1 U14041 ( .A1(n11717), .A2(n11716), .ZN(n11719) );
  NAND2_X1 U14042 ( .A1(n12739), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U14043 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12739), .A(n12748), 
        .ZN(n11720) );
  AOI21_X1 U14044 ( .B1(n11721), .B2(n11720), .A(n12746), .ZN(n11722) );
  NOR2_X1 U14045 ( .A1(n11722), .A2(n12888), .ZN(n11723) );
  AOI211_X1 U14046 ( .C1(n12859), .C2(n11725), .A(n11724), .B(n11723), .ZN(
        n11726) );
  OAI211_X1 U14047 ( .C1(n11728), .C2(n12892), .A(n11727), .B(n11726), .ZN(
        P3_U3194) );
  MUX2_X1 U14048 ( .A(n15214), .B(n11730), .S(n11729), .Z(n11732) );
  XNOR2_X1 U14049 ( .A(n11732), .B(n11731), .ZN(n11733) );
  NAND2_X1 U14050 ( .A1(n11733), .A2(n12644), .ZN(n11742) );
  OAI22_X1 U14051 ( .A1(n11735), .A2(n12652), .B1(n12659), .B2(n11734), .ZN(
        n11740) );
  NOR2_X1 U14052 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11736), .ZN(n12722) );
  INV_X1 U14053 ( .A(n12722), .ZN(n11737) );
  OAI21_X1 U14054 ( .B1(n12666), .B2(n11738), .A(n11737), .ZN(n11739) );
  NOR2_X1 U14055 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  OAI211_X1 U14056 ( .C1(n11743), .C2(n12670), .A(n11742), .B(n11741), .ZN(
        P3_U3161) );
  INV_X1 U14057 ( .A(n11931), .ZN(n11747) );
  OAI222_X1 U14058 ( .A1(n13999), .A2(n11745), .B1(n14001), .B2(n11747), .C1(
        n11744), .C2(P2_U3088), .ZN(P2_U3303) );
  OAI222_X1 U14059 ( .A1(n14701), .A2(n11748), .B1(n14707), .B2(n11747), .C1(
        n11746), .C2(P1_U3086), .ZN(P1_U3331) );
  NOR2_X1 U14060 ( .A1(n12360), .A2(n11751), .ZN(n11752) );
  AOI21_X1 U14061 ( .B1(n12148), .B2(n12400), .A(n11752), .ZN(n12270) );
  AOI22_X1 U14062 ( .A1(n12148), .A2(n12404), .B1(n12400), .B2(n14909), .ZN(
        n11753) );
  XNOR2_X1 U14063 ( .A(n11753), .B(n12292), .ZN(n12271) );
  XOR2_X1 U14064 ( .A(n12272), .B(n12271), .Z(n11759) );
  AOI22_X1 U14065 ( .A1(n14923), .A2(n14149), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11754) );
  OAI21_X1 U14066 ( .B1(n12276), .B2(n14120), .A(n11754), .ZN(n11756) );
  NAND2_X1 U14067 ( .A1(n12148), .A2(n15062), .ZN(n15095) );
  NOR2_X1 U14068 ( .A1(n15095), .A2(n14913), .ZN(n11755) );
  AOI211_X1 U14069 ( .C1(n14113), .C2(n11757), .A(n11756), .B(n11755), .ZN(
        n11758) );
  OAI21_X1 U14070 ( .B1(n11759), .B2(n14133), .A(n11758), .ZN(P1_U3231) );
  OR2_X1 U14071 ( .A1(n12301), .A2(n12299), .ZN(n11761) );
  NAND2_X1 U14072 ( .A1(n11762), .A2(n11761), .ZN(n11785) );
  NAND2_X1 U14073 ( .A1(n11763), .A2(n6429), .ZN(n11766) );
  AOI22_X1 U14074 ( .A1(n11764), .A2(n12022), .B1(n12023), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11765) );
  NAND2_X1 U14075 ( .A1(n12308), .A2(n12306), .ZN(n12165) );
  XNOR2_X1 U14076 ( .A(n11785), .B(n12172), .ZN(n14937) );
  OR2_X1 U14077 ( .A1(n12301), .A2(n14897), .ZN(n11767) );
  AOI21_X1 U14078 ( .B1(n12172), .B2(n11769), .A(n6568), .ZN(n14943) );
  AOI21_X1 U14079 ( .B1(n12308), .B2(n11770), .A(n14640), .ZN(n11771) );
  NAND2_X1 U14080 ( .A1(n11771), .A2(n11799), .ZN(n14939) );
  INV_X1 U14081 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11772) );
  AND2_X1 U14082 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  OR2_X1 U14083 ( .A1(n11774), .A2(n11791), .ZN(n14139) );
  NAND2_X1 U14084 ( .A1(n10484), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U14085 ( .A1(n12061), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11775) );
  AND2_X1 U14086 ( .A1(n11776), .A2(n11775), .ZN(n11778) );
  NAND2_X1 U14087 ( .A1(n12059), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11777) );
  OAI211_X1 U14088 ( .C1(n14139), .C2(n11779), .A(n11778), .B(n11777), .ZN(
        n14898) );
  AOI22_X1 U14089 ( .A1(n14509), .A2(n14898), .B1(n15007), .B2(n14897), .ZN(
        n14938) );
  OAI22_X1 U14090 ( .A1(n15022), .A2(n14938), .B1(n14904), .B2(n14544), .ZN(
        n11781) );
  INV_X1 U14091 ( .A(n12308), .ZN(n14940) );
  NOR2_X1 U14092 ( .A1(n14940), .A2(n15012), .ZN(n11780) );
  AOI211_X1 U14093 ( .C1(n15022), .C2(P1_REG2_REG_14__SCAN_IN), .A(n11781), 
        .B(n11780), .ZN(n11782) );
  OAI21_X1 U14094 ( .B1(n14537), .B2(n14939), .A(n11782), .ZN(n11783) );
  AOI21_X1 U14095 ( .B1(n14943), .B2(n14548), .A(n11783), .ZN(n11784) );
  OAI21_X1 U14096 ( .B1(n14937), .B2(n14441), .A(n11784), .ZN(P1_U3279) );
  NAND2_X1 U14097 ( .A1(n11785), .A2(n12172), .ZN(n11786) );
  NAND2_X1 U14098 ( .A1(n11786), .A2(n12174), .ZN(n14288) );
  NAND2_X1 U14099 ( .A1(n11787), .A2(n6429), .ZN(n11790) );
  AOI22_X1 U14100 ( .A1(n11788), .A2(n12022), .B1(n12023), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n11789) );
  INV_X1 U14101 ( .A(n14898), .ZN(n14524) );
  OR2_X1 U14102 ( .A1(n14264), .A2(n14524), .ZN(n14289) );
  NAND2_X1 U14103 ( .A1(n14264), .A2(n14524), .ZN(n12173) );
  NAND2_X1 U14104 ( .A1(n14289), .A2(n12173), .ZN(n12019) );
  XNOR2_X1 U14105 ( .A(n14288), .B(n14287), .ZN(n11798) );
  NAND2_X1 U14106 ( .A1(n11791), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11996) );
  OR2_X1 U14107 ( .A1(n11791), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U14108 ( .A1(n11996), .A2(n11792), .ZN(n14533) );
  AOI22_X1 U14109 ( .A1(n12060), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n12061), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11794) );
  NAND2_X1 U14110 ( .A1(n12059), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11793) );
  OAI211_X1 U14111 ( .C1(n14533), .C2(n11779), .A(n11794), .B(n11793), .ZN(
        n14507) );
  NAND2_X1 U14112 ( .A1(n14507), .A2(n14509), .ZN(n11796) );
  INV_X1 U14113 ( .A(n12306), .ZN(n14148) );
  NAND2_X1 U14114 ( .A1(n14148), .A2(n15007), .ZN(n11795) );
  NAND2_X1 U14115 ( .A1(n11796), .A2(n11795), .ZN(n14142) );
  INV_X1 U14116 ( .A(n14142), .ZN(n11797) );
  OAI21_X1 U14117 ( .B1(n11798), .B2(n14936), .A(n11797), .ZN(n11844) );
  INV_X1 U14118 ( .A(n11844), .ZN(n11805) );
  AOI211_X1 U14119 ( .C1(n14264), .C2(n11799), .A(n14640), .B(n6437), .ZN(
        n11845) );
  NOR2_X1 U14120 ( .A1(n7280), .A2(n15012), .ZN(n11802) );
  INV_X1 U14121 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11800) );
  OAI22_X1 U14122 ( .A1(n14541), .A2(n11800), .B1(n14139), .B2(n14544), .ZN(
        n11801) );
  AOI211_X1 U14123 ( .C1(n11845), .C2(n15018), .A(n11802), .B(n11801), .ZN(
        n11804) );
  XNOR2_X1 U14124 ( .A(n14263), .B(n14287), .ZN(n11846) );
  NAND2_X1 U14125 ( .A1(n11846), .A2(n14548), .ZN(n11803) );
  OAI211_X1 U14126 ( .C1(n11805), .C2(n15022), .A(n11804), .B(n11803), .ZN(
        P1_U3278) );
  INV_X1 U14127 ( .A(n12052), .ZN(n11808) );
  OAI222_X1 U14128 ( .A1(n14701), .A2(n12053), .B1(n14707), .B2(n11808), .C1(
        n11806), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U14129 ( .A1(n13999), .A2(n15327), .B1(n14001), .B2(n11808), .C1(
        n11807), .C2(P2_U3088), .ZN(P2_U3302) );
  AOI211_X1 U14130 ( .C1(n13905), .C2(n11811), .A(n11810), .B(n11809), .ZN(
        n11814) );
  AOI22_X1 U14131 ( .A1(n11863), .A2(n13899), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n15188), .ZN(n11812) );
  OAI21_X1 U14132 ( .B1(n11814), .B2(n15188), .A(n11812), .ZN(P2_U3514) );
  AOI22_X1 U14133 ( .A1(n11863), .A2(n13965), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n15185), .ZN(n11813) );
  OAI21_X1 U14134 ( .B1(n11814), .B2(n15185), .A(n11813), .ZN(P2_U3475) );
  INV_X1 U14135 ( .A(n11815), .ZN(n11817) );
  NAND2_X1 U14136 ( .A1(n13477), .A2(n13343), .ZN(n11820) );
  INV_X1 U14137 ( .A(n11820), .ZN(n11823) );
  XNOR2_X1 U14138 ( .A(n14887), .B(n13338), .ZN(n11821) );
  INV_X1 U14139 ( .A(n11821), .ZN(n11822) );
  AOI21_X1 U14140 ( .B1(n11823), .B2(n11822), .A(n13306), .ZN(n14882) );
  INV_X1 U14141 ( .A(n13306), .ZN(n11824) );
  NAND2_X1 U14142 ( .A1(n14880), .A2(n11824), .ZN(n11826) );
  XNOR2_X1 U14143 ( .A(n11863), .B(n13338), .ZN(n13308) );
  NAND2_X1 U14144 ( .A1(n13476), .A2(n13343), .ZN(n13307) );
  XNOR2_X1 U14145 ( .A(n13308), .B(n13307), .ZN(n11825) );
  XNOR2_X1 U14146 ( .A(n11826), .B(n11825), .ZN(n11832) );
  AOI22_X1 U14147 ( .A1(n14885), .A2(n11827), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11828) );
  OAI21_X1 U14148 ( .B1(n11829), .B2(n14891), .A(n11828), .ZN(n11830) );
  AOI21_X1 U14149 ( .B1(n11863), .B2(n9631), .A(n11830), .ZN(n11831) );
  OAI21_X1 U14150 ( .B1(n11832), .B2(n13470), .A(n11831), .ZN(P2_U3213) );
  OAI21_X1 U14151 ( .B1(n11835), .B2(n11834), .A(n11833), .ZN(n14237) );
  XNOR2_X1 U14152 ( .A(n14237), .B(n14230), .ZN(n14235) );
  XNOR2_X1 U14153 ( .A(n14235), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n11843) );
  NAND2_X1 U14154 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14118)
         );
  INV_X1 U14155 ( .A(n11836), .ZN(n11837) );
  AOI21_X1 U14156 ( .B1(n11992), .B2(P1_REG1_REG_17__SCAN_IN), .A(n11837), 
        .ZN(n14231) );
  XNOR2_X1 U14157 ( .A(n14231), .B(n14236), .ZN(n11838) );
  NAND2_X1 U14158 ( .A1(n11838), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14232) );
  OAI211_X1 U14159 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11838), .A(n14245), 
        .B(n14232), .ZN(n11839) );
  NAND2_X1 U14160 ( .A1(n14118), .A2(n11839), .ZN(n11841) );
  NOR2_X1 U14161 ( .A1(n14992), .A2(n14230), .ZN(n11840) );
  AOI211_X1 U14162 ( .C1(n14977), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n11841), 
        .B(n11840), .ZN(n11842) );
  OAI21_X1 U14163 ( .B1(n11843), .B2(n14983), .A(n11842), .ZN(P1_U3261) );
  AOI211_X1 U14164 ( .C1(n11846), .C2(n15108), .A(n11845), .B(n11844), .ZN(
        n11852) );
  AOI22_X1 U14165 ( .A1(n14264), .A2(n11847), .B1(n15120), .B2(
        P1_REG1_REG_15__SCAN_IN), .ZN(n11848) );
  OAI21_X1 U14166 ( .B1(n11852), .B2(n15120), .A(n11848), .ZN(P1_U3543) );
  INV_X1 U14167 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11849) );
  OAI22_X1 U14168 ( .A1(n7280), .A2(n14683), .B1(n14655), .B2(n11849), .ZN(
        n11850) );
  INV_X1 U14169 ( .A(n11850), .ZN(n11851) );
  OAI21_X1 U14170 ( .B1(n11852), .B2(n15109), .A(n11851), .ZN(P1_U3504) );
  XNOR2_X1 U14171 ( .A(n13605), .B(n11866), .ZN(n11855) );
  NAND2_X1 U14172 ( .A1(n11855), .A2(n13822), .ZN(n11856) );
  AOI22_X1 U14173 ( .A1(n13581), .A2(n13570), .B1(n13464), .B2(n13476), .ZN(
        n13410) );
  NAND2_X1 U14174 ( .A1(n11856), .A2(n13410), .ZN(n11876) );
  INV_X1 U14175 ( .A(n11876), .ZN(n11870) );
  INV_X1 U14176 ( .A(n13412), .ZN(n11857) );
  OAI22_X1 U14177 ( .A1(n13844), .A2(n11858), .B1(n11857), .B2(n13841), .ZN(
        n11860) );
  INV_X1 U14178 ( .A(n13607), .ZN(n13415) );
  OAI211_X1 U14179 ( .C1(n13415), .C2(n6577), .A(n10023), .B(n13824), .ZN(
        n11872) );
  NOR2_X1 U14180 ( .A1(n11872), .A2(n13766), .ZN(n11859) );
  AOI211_X1 U14181 ( .C1(n13846), .C2(n13607), .A(n11860), .B(n11859), .ZN(
        n11869) );
  OR2_X1 U14182 ( .A1(n11863), .A2(n13476), .ZN(n11864) );
  INV_X1 U14183 ( .A(n11866), .ZN(n13604) );
  NAND2_X1 U14184 ( .A1(n11867), .A2(n13604), .ZN(n11871) );
  NAND3_X1 U14185 ( .A1(n13580), .A2(n11871), .A3(n13848), .ZN(n11868) );
  OAI211_X1 U14186 ( .C1(n11870), .C2(n6430), .A(n11869), .B(n11868), .ZN(
        P2_U3249) );
  NAND3_X1 U14187 ( .A1(n13580), .A2(n13905), .A3(n11871), .ZN(n11873) );
  OAI211_X1 U14188 ( .C1(n13415), .C2(n11874), .A(n11873), .B(n11872), .ZN(
        n11875) );
  NOR2_X1 U14189 ( .A1(n11876), .A2(n11875), .ZN(n11879) );
  MUX2_X1 U14190 ( .A(n11877), .B(n11879), .S(n15190), .Z(n11878) );
  INV_X1 U14191 ( .A(n11878), .ZN(P2_U3515) );
  INV_X1 U14192 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n11880) );
  MUX2_X1 U14193 ( .A(n11880), .B(n11879), .S(n15187), .Z(n11881) );
  INV_X1 U14194 ( .A(n11881), .ZN(P2_U3478) );
  AND2_X1 U14195 ( .A1(n15425), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U14196 ( .A1(n15425), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14197 ( .A1(n15425), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14198 ( .A1(n15425), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U14199 ( .A1(n15425), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14200 ( .A1(n15425), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14201 ( .A1(n15425), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U14202 ( .A1(n15425), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14203 ( .A1(n15425), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14204 ( .A1(n15425), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14205 ( .A1(n15425), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14206 ( .A1(n15425), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14207 ( .A1(n15425), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14208 ( .A1(n15425), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14209 ( .A1(n15425), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14210 ( .A1(n15425), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14211 ( .A1(n15425), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14212 ( .A1(n15425), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14213 ( .A1(n15425), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14214 ( .A1(n15425), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14215 ( .A1(n15425), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14216 ( .A1(n15425), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14217 ( .A1(n15425), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14218 ( .A1(n15425), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14219 ( .A1(n15425), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14220 ( .A1(n15425), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14221 ( .A1(n15425), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14222 ( .A1(n15425), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14223 ( .A1(n15425), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U14224 ( .A(SI_30_), .ZN(n11886) );
  INV_X1 U14225 ( .A(n11884), .ZN(n11885) );
  OAI222_X1 U14226 ( .A1(n7685), .A2(P3_U3151), .B1(n11887), .B2(n11886), .C1(
        n13303), .C2(n11885), .ZN(P3_U3265) );
  INV_X1 U14227 ( .A(n11888), .ZN(n11890) );
  OAI222_X1 U14228 ( .A1(n11891), .A2(n11890), .B1(n12420), .B2(n11889), .C1(
        P3_U3151), .C2(n8404), .ZN(P3_U3267) );
  NAND2_X1 U14229 ( .A1(n11892), .A2(n6429), .ZN(n11894) );
  NAND2_X1 U14230 ( .A1(n12023), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U14231 ( .A1(n12059), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11897) );
  NAND2_X1 U14232 ( .A1(n10484), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U14233 ( .A1(n12061), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11895) );
  AND3_X1 U14234 ( .A1(n11897), .A2(n11896), .A3(n11895), .ZN(n12099) );
  XNOR2_X1 U14235 ( .A(n14251), .B(n12099), .ZN(n12241) );
  INV_X1 U14236 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U14237 ( .A1(n12059), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U14238 ( .A1(n10243), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11898) );
  OAI211_X1 U14239 ( .C1(n11900), .C2(n14258), .A(n11899), .B(n11898), .ZN(
        n14316) );
  OR2_X1 U14240 ( .A1(n12054), .A2(n15339), .ZN(n11901) );
  NAND2_X1 U14241 ( .A1(n13987), .A2(n6429), .ZN(n11904) );
  NAND2_X1 U14242 ( .A1(n12023), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11903) );
  NAND2_X1 U14243 ( .A1(n12059), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11913) );
  INV_X1 U14244 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11995) );
  INV_X1 U14245 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n15413) );
  AND2_X1 U14246 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n11905) );
  NAND2_X1 U14247 ( .A1(n12034), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11953) );
  INV_X1 U14248 ( .A(n11953), .ZN(n11906) );
  NAND2_X1 U14249 ( .A1(n11906), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11935) );
  INV_X1 U14250 ( .A(n11935), .ZN(n11945) );
  NAND2_X1 U14251 ( .A1(n11945), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12058) );
  INV_X1 U14252 ( .A(n12058), .ZN(n11934) );
  NAND2_X1 U14253 ( .A1(n11934), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11923) );
  INV_X1 U14254 ( .A(n11923), .ZN(n12057) );
  NAND2_X1 U14255 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n12057), .ZN(n12045) );
  INV_X1 U14256 ( .A(n12045), .ZN(n11907) );
  NAND2_X1 U14257 ( .A1(n11907), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12047) );
  INV_X1 U14258 ( .A(n12047), .ZN(n11908) );
  NAND2_X1 U14259 ( .A1(n11908), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14318) );
  INV_X1 U14260 ( .A(n14318), .ZN(n11909) );
  NAND2_X1 U14261 ( .A1(n11974), .A2(n11909), .ZN(n11912) );
  NAND2_X1 U14262 ( .A1(n12061), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U14263 ( .A1(n12060), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11910) );
  XNOR2_X1 U14264 ( .A(n14321), .B(n12409), .ZN(n14312) );
  NAND2_X1 U14265 ( .A1(n13990), .A2(n6429), .ZN(n11915) );
  OR2_X1 U14266 ( .A1(n12054), .A2(n14698), .ZN(n11914) );
  NAND2_X1 U14267 ( .A1(n12059), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11920) );
  INV_X1 U14268 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n15354) );
  NAND2_X1 U14269 ( .A1(n12047), .A2(n15354), .ZN(n11916) );
  NAND2_X1 U14270 ( .A1(n11974), .A2(n14330), .ZN(n11919) );
  NAND2_X1 U14271 ( .A1(n12061), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U14272 ( .A1(n12060), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11917) );
  NAND4_X1 U14273 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n14315) );
  XNOR2_X1 U14274 ( .A(n14335), .B(n14315), .ZN(n14337) );
  NAND2_X1 U14275 ( .A1(n13998), .A2(n6429), .ZN(n11922) );
  OR2_X1 U14276 ( .A1(n12054), .A2(n14708), .ZN(n11921) );
  INV_X1 U14277 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U14278 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  AND2_X1 U14279 ( .A1(n11925), .A2(n12045), .ZN(n14365) );
  NAND2_X1 U14280 ( .A1(n11974), .A2(n14365), .ZN(n11929) );
  NAND2_X1 U14281 ( .A1(n12059), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14282 ( .A1(n12060), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U14283 ( .A1(n12061), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11926) );
  NAND4_X1 U14284 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n14281) );
  INV_X1 U14285 ( .A(n14281), .ZN(n14349) );
  NAND2_X1 U14286 ( .A1(n14583), .A2(n14349), .ZN(n14346) );
  OR2_X1 U14287 ( .A1(n14583), .A2(n14349), .ZN(n11930) );
  NAND2_X1 U14288 ( .A1(n14346), .A2(n11930), .ZN(n14361) );
  NAND2_X1 U14289 ( .A1(n11931), .A2(n6429), .ZN(n11933) );
  NAND2_X1 U14290 ( .A1(n12023), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11932) );
  INV_X1 U14291 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n11936) );
  AOI21_X1 U14292 ( .B1(n11936), .B2(n11935), .A(n11934), .ZN(n14406) );
  NAND2_X1 U14293 ( .A1(n11974), .A2(n14406), .ZN(n11940) );
  NAND2_X1 U14294 ( .A1(n12059), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U14295 ( .A1(n12060), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U14296 ( .A1(n12061), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11937) );
  NAND4_X1 U14297 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n14278) );
  INV_X1 U14298 ( .A(n14278), .ZN(n14305) );
  XNOR2_X1 U14299 ( .A(n14593), .B(n14305), .ZN(n14394) );
  NAND2_X1 U14300 ( .A1(n11941), .A2(n6429), .ZN(n11944) );
  OR2_X1 U14301 ( .A1(n12054), .A2(n11942), .ZN(n11943) );
  INV_X1 U14302 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14013) );
  AOI21_X1 U14303 ( .B1(n14013), .B2(n11953), .A(n11945), .ZN(n14420) );
  NAND2_X1 U14304 ( .A1(n11974), .A2(n14420), .ZN(n11949) );
  NAND2_X1 U14305 ( .A1(n12059), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14306 ( .A1(n12060), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11947) );
  NAND2_X1 U14307 ( .A1(n12061), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U14308 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n14398) );
  XNOR2_X1 U14309 ( .A(n11952), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14710) );
  OR2_X1 U14310 ( .A1(n12034), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11954) );
  AND2_X1 U14311 ( .A1(n11954), .A2(n11953), .ZN(n14436) );
  NAND2_X1 U14312 ( .A1(n14436), .A2(n11974), .ZN(n11960) );
  INV_X1 U14313 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U14314 ( .A1(n12060), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U14315 ( .A1(n12061), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11955) );
  OAI211_X1 U14316 ( .C1(n11957), .C2(n12037), .A(n11956), .B(n11955), .ZN(
        n11958) );
  INV_X1 U14317 ( .A(n11958), .ZN(n11959) );
  NAND2_X1 U14318 ( .A1(n11960), .A2(n11959), .ZN(n14275) );
  INV_X1 U14319 ( .A(n14275), .ZN(n14301) );
  XNOR2_X1 U14320 ( .A(n14606), .B(n14301), .ZN(n14427) );
  NAND2_X1 U14321 ( .A1(n11961), .A2(n6429), .ZN(n11963) );
  AOI22_X1 U14322 ( .A1(n12023), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14433), 
        .B2(n12022), .ZN(n11962) );
  INV_X1 U14323 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11964) );
  XNOR2_X1 U14324 ( .A(n11984), .B(n11964), .ZN(n14478) );
  NAND2_X1 U14325 ( .A1(n14478), .A2(n11974), .ZN(n11969) );
  INV_X1 U14326 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U14327 ( .A1(n10484), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U14328 ( .A1(n12061), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11965) );
  OAI211_X1 U14329 ( .C1(n14628), .C2(n12037), .A(n11966), .B(n11965), .ZN(
        n11967) );
  INV_X1 U14330 ( .A(n11967), .ZN(n11968) );
  XNOR2_X1 U14331 ( .A(n14475), .B(n14297), .ZN(n14296) );
  NAND2_X1 U14332 ( .A1(n11970), .A2(n6429), .ZN(n11972) );
  OR2_X1 U14333 ( .A1(n12054), .A2(n6945), .ZN(n11971) );
  AOI21_X1 U14334 ( .B1(n11984), .B2(P1_REG3_REG_19__SCAN_IN), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n11973) );
  NOR2_X1 U14335 ( .A1(n12032), .A2(n11973), .ZN(n14457) );
  NAND2_X1 U14336 ( .A1(n14457), .A2(n11974), .ZN(n11979) );
  INV_X1 U14337 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14623) );
  NAND2_X1 U14338 ( .A1(n12060), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U14339 ( .A1(n12061), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11975) );
  OAI211_X1 U14340 ( .C1(n14623), .C2(n12037), .A(n11976), .B(n11975), .ZN(
        n11977) );
  INV_X1 U14341 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U14342 ( .A1(n14464), .A2(n14471), .ZN(n11980) );
  NAND2_X1 U14343 ( .A1(n14298), .A2(n11980), .ZN(n14271) );
  NAND2_X1 U14344 ( .A1(n11981), .A2(n6429), .ZN(n11983) );
  AOI22_X1 U14345 ( .A1(n12023), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12022), 
        .B2(n14236), .ZN(n11982) );
  AND2_X1 U14346 ( .A1(n11998), .A2(n15413), .ZN(n11985) );
  OR2_X1 U14347 ( .A1(n11985), .A2(n11984), .ZN(n14495) );
  INV_X1 U14348 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11988) );
  NAND2_X1 U14349 ( .A1(n12061), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11987) );
  NAND2_X1 U14350 ( .A1(n10484), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11986) );
  OAI211_X1 U14351 ( .C1(n11988), .C2(n12037), .A(n11987), .B(n11986), .ZN(
        n11989) );
  INV_X1 U14352 ( .A(n11989), .ZN(n11990) );
  OAI21_X1 U14353 ( .B1(n14495), .B2(n11779), .A(n11990), .ZN(n14510) );
  INV_X1 U14354 ( .A(n14510), .ZN(n14472) );
  XNOR2_X1 U14355 ( .A(n14633), .B(n14472), .ZN(n14484) );
  NAND2_X1 U14356 ( .A1(n11991), .A2(n6429), .ZN(n11994) );
  AOI22_X1 U14357 ( .A1(n12023), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12022), 
        .B2(n11992), .ZN(n11993) );
  NAND2_X1 U14358 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  NAND2_X1 U14359 ( .A1(n11998), .A2(n11997), .ZN(n14511) );
  AOI22_X1 U14360 ( .A1(n12060), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n12061), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n12000) );
  NAND2_X1 U14361 ( .A1(n12059), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11999) );
  OAI211_X1 U14362 ( .C1(n14511), .C2(n11779), .A(n12000), .B(n11999), .ZN(
        n14488) );
  XNOR2_X1 U14363 ( .A(n14637), .B(n14488), .ZN(n14501) );
  INV_X1 U14364 ( .A(n12172), .ZN(n12017) );
  NOR4_X1 U14365 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n15003), .ZN(
        n12006) );
  NAND4_X1 U14366 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(
        n12008) );
  NOR4_X1 U14367 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12014) );
  NAND4_X1 U14368 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12016) );
  NOR4_X1 U14369 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12026) );
  NAND2_X1 U14370 ( .A1(n12020), .A2(n6429), .ZN(n12025) );
  AOI22_X1 U14371 ( .A1(n12023), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12022), 
        .B2(n12021), .ZN(n12024) );
  XNOR2_X1 U14372 ( .A(n14535), .B(n14507), .ZN(n14521) );
  NAND3_X1 U14373 ( .A1(n14501), .A2(n12026), .A3(n14521), .ZN(n12027) );
  NOR4_X1 U14374 ( .A1(n14296), .A2(n14271), .A3(n14484), .A4(n12027), .ZN(
        n12040) );
  NAND2_X1 U14375 ( .A1(n12028), .A2(n6429), .ZN(n12031) );
  OR2_X1 U14376 ( .A1(n12054), .A2(n12029), .ZN(n12030) );
  NOR2_X1 U14377 ( .A1(n12032), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12033) );
  OR2_X1 U14378 ( .A1(n12034), .A2(n12033), .ZN(n14444) );
  INV_X1 U14379 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U14380 ( .A1(n12060), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U14381 ( .A1(n12061), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12035) );
  OAI211_X1 U14382 ( .C1(n14616), .C2(n12037), .A(n12036), .B(n12035), .ZN(
        n12038) );
  INV_X1 U14383 ( .A(n12038), .ZN(n12039) );
  OAI21_X1 U14384 ( .B1(n14444), .B2(n11779), .A(n12039), .ZN(n14299) );
  XNOR2_X1 U14385 ( .A(n14443), .B(n14299), .ZN(n14448) );
  NAND2_X1 U14386 ( .A1(n13995), .A2(n6429), .ZN(n12043) );
  OR2_X1 U14387 ( .A1(n12054), .A2(n14702), .ZN(n12042) );
  NAND2_X1 U14388 ( .A1(n12059), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12051) );
  INV_X1 U14389 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U14390 ( .A1(n12045), .A2(n12044), .ZN(n12046) );
  NAND2_X1 U14391 ( .A1(n11974), .A2(n14355), .ZN(n12050) );
  NAND2_X1 U14392 ( .A1(n12061), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U14393 ( .A1(n10484), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12048) );
  NAND4_X1 U14394 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n14284) );
  XNOR2_X1 U14395 ( .A(n14576), .B(n14284), .ZN(n14344) );
  NAND2_X1 U14396 ( .A1(n12052), .A2(n6429), .ZN(n12056) );
  OR2_X1 U14397 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  INV_X1 U14398 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14047) );
  AOI21_X1 U14399 ( .B1(n14047), .B2(n12058), .A(n12057), .ZN(n14385) );
  NAND2_X1 U14400 ( .A1(n11974), .A2(n14385), .ZN(n12065) );
  NAND2_X1 U14401 ( .A1(n12059), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U14402 ( .A1(n12060), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12063) );
  NAND2_X1 U14403 ( .A1(n12061), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12062) );
  NAND4_X1 U14404 ( .A1(n12065), .A2(n12064), .A3(n12063), .A4(n12062), .ZN(
        n14399) );
  XNOR2_X1 U14405 ( .A(n14389), .B(n14399), .ZN(n14379) );
  NAND4_X1 U14406 ( .A1(n14337), .A2(n12066), .A3(n14344), .A4(n14379), .ZN(
        n12067) );
  NAND2_X1 U14407 ( .A1(n12069), .A2(n12068), .ZN(n12071) );
  NAND2_X1 U14408 ( .A1(n12071), .A2(n12070), .ZN(n12090) );
  NAND2_X1 U14409 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  NAND2_X1 U14410 ( .A1(n14251), .A2(n12229), .ZN(n12089) );
  XOR2_X1 U14411 ( .A(n12090), .B(n12089), .Z(n12080) );
  INV_X1 U14412 ( .A(n12099), .ZN(n14254) );
  NOR2_X1 U14413 ( .A1(n12080), .A2(n14254), .ZN(n12085) );
  NOR2_X1 U14414 ( .A1(n14251), .A2(n12229), .ZN(n12081) );
  NAND2_X1 U14415 ( .A1(n12081), .A2(n14254), .ZN(n12093) );
  INV_X1 U14416 ( .A(n12081), .ZN(n12082) );
  NAND3_X1 U14417 ( .A1(n12082), .A2(n14254), .A3(n12090), .ZN(n12083) );
  OAI211_X1 U14418 ( .C1(n12093), .C2(n12090), .A(n12091), .B(n12083), .ZN(
        n12084) );
  INV_X1 U14419 ( .A(n12243), .ZN(n12103) );
  NAND2_X1 U14420 ( .A1(n12229), .A2(n14254), .ZN(n12087) );
  INV_X1 U14421 ( .A(n14316), .ZN(n12097) );
  AOI21_X1 U14422 ( .B1(n12087), .B2(n12086), .A(n12097), .ZN(n12088) );
  AOI21_X1 U14423 ( .B1(n14261), .B2(n12236), .A(n12088), .ZN(n12246) );
  AND2_X1 U14424 ( .A1(n12246), .A2(n12248), .ZN(n12251) );
  INV_X1 U14425 ( .A(n12089), .ZN(n12096) );
  INV_X1 U14426 ( .A(n12090), .ZN(n12242) );
  INV_X1 U14427 ( .A(n12091), .ZN(n12092) );
  NOR2_X1 U14428 ( .A1(n12242), .A2(n12092), .ZN(n12245) );
  INV_X1 U14429 ( .A(n12245), .ZN(n12095) );
  INV_X1 U14430 ( .A(n12093), .ZN(n12094) );
  AOI211_X1 U14431 ( .C1(n12099), .C2(n12096), .A(n12095), .B(n12094), .ZN(
        n12252) );
  INV_X1 U14432 ( .A(n12252), .ZN(n12101) );
  AOI21_X1 U14433 ( .B1(n12099), .B2(n12098), .A(n12097), .ZN(n12100) );
  MUX2_X1 U14434 ( .A(n12100), .B(n14261), .S(n12229), .Z(n12250) );
  INV_X1 U14435 ( .A(n12250), .ZN(n12249) );
  NOR3_X1 U14436 ( .A1(n12101), .A2(n12249), .A3(n12256), .ZN(n12102) );
  AOI21_X1 U14437 ( .B1(n12103), .B2(n12251), .A(n12102), .ZN(n12267) );
  MUX2_X1 U14438 ( .A(n12409), .B(n14564), .S(n12131), .Z(n12238) );
  INV_X1 U14439 ( .A(n12108), .ZN(n12111) );
  NAND2_X1 U14440 ( .A1(n12109), .A2(n12131), .ZN(n12110) );
  MUX2_X1 U14441 ( .A(n12115), .B(n12114), .S(n12236), .Z(n12117) );
  MUX2_X1 U14442 ( .A(n12119), .B(n12118), .S(n12236), .Z(n12120) );
  MUX2_X1 U14443 ( .A(n15073), .B(n12122), .S(n12236), .Z(n12125) );
  MUX2_X1 U14444 ( .A(n14153), .B(n12123), .S(n12236), .Z(n12124) );
  OAI21_X1 U14445 ( .B1(n12126), .B2(n12125), .A(n12124), .ZN(n12128) );
  NAND2_X1 U14446 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  MUX2_X1 U14447 ( .A(n14152), .B(n14067), .S(n12236), .Z(n12130) );
  MUX2_X1 U14448 ( .A(n14152), .B(n14067), .S(n12131), .Z(n12129) );
  MUX2_X1 U14449 ( .A(n14151), .B(n12132), .S(n12131), .Z(n12134) );
  MUX2_X1 U14450 ( .A(n14151), .B(n12132), .S(n12236), .Z(n12133) );
  MUX2_X1 U14451 ( .A(n14150), .B(n12135), .S(n12228), .Z(n12138) );
  MUX2_X1 U14452 ( .A(n14150), .B(n12135), .S(n12229), .Z(n12136) );
  MUX2_X1 U14453 ( .A(n14149), .B(n12139), .S(n12229), .Z(n12143) );
  NAND2_X1 U14454 ( .A1(n12142), .A2(n12143), .ZN(n12141) );
  MUX2_X1 U14455 ( .A(n14149), .B(n12139), .S(n12236), .Z(n12140) );
  NAND2_X1 U14456 ( .A1(n12141), .A2(n12140), .ZN(n12147) );
  INV_X1 U14457 ( .A(n12143), .ZN(n12144) );
  NAND2_X1 U14458 ( .A1(n12145), .A2(n12144), .ZN(n12146) );
  MUX2_X1 U14459 ( .A(n14909), .B(n12148), .S(n12228), .Z(n12150) );
  MUX2_X1 U14460 ( .A(n14909), .B(n12148), .S(n12229), .Z(n12149) );
  MUX2_X1 U14461 ( .A(n14922), .B(n14905), .S(n12229), .Z(n12153) );
  MUX2_X1 U14462 ( .A(n14922), .B(n14905), .S(n12236), .Z(n12151) );
  INV_X1 U14463 ( .A(n12153), .ZN(n12154) );
  MUX2_X1 U14464 ( .A(n14910), .B(n14547), .S(n12228), .Z(n12158) );
  MUX2_X1 U14465 ( .A(n14910), .B(n14547), .S(n12131), .Z(n12155) );
  NAND2_X1 U14466 ( .A1(n12156), .A2(n12155), .ZN(n12162) );
  INV_X1 U14467 ( .A(n12157), .ZN(n12160) );
  INV_X1 U14468 ( .A(n12158), .ZN(n12159) );
  NAND2_X1 U14469 ( .A1(n12160), .A2(n12159), .ZN(n12161) );
  MUX2_X1 U14470 ( .A(n14924), .B(n12291), .S(n12229), .Z(n12164) );
  MUX2_X1 U14471 ( .A(n14924), .B(n12291), .S(n12228), .Z(n12163) );
  MUX2_X1 U14472 ( .A(n14897), .B(n12301), .S(n12228), .Z(n12170) );
  NAND2_X1 U14473 ( .A1(n12169), .A2(n12170), .ZN(n12168) );
  NAND3_X1 U14474 ( .A1(n12168), .A2(n12172), .A3(n12301), .ZN(n12166) );
  NAND3_X1 U14475 ( .A1(n12166), .A2(n12173), .A3(n12165), .ZN(n12167) );
  INV_X1 U14476 ( .A(n12168), .ZN(n12179) );
  NAND4_X1 U14477 ( .A1(n12173), .A2(n12172), .A3(n12228), .A4(n14897), .ZN(
        n12178) );
  INV_X1 U14478 ( .A(n12170), .ZN(n12171) );
  AOI21_X1 U14479 ( .B1(n12174), .B2(n14524), .A(n12229), .ZN(n12176) );
  OAI21_X1 U14480 ( .B1(n12174), .B2(n14524), .A(n14264), .ZN(n12175) );
  MUX2_X1 U14481 ( .A(n14507), .B(n14535), .S(n12228), .Z(n12183) );
  INV_X1 U14482 ( .A(n14507), .ZN(n14291) );
  MUX2_X1 U14483 ( .A(n14291), .B(n14647), .S(n12229), .Z(n12182) );
  AND2_X1 U14484 ( .A1(n14488), .A2(n12131), .ZN(n12185) );
  OAI21_X1 U14485 ( .B1(n12131), .B2(n14488), .A(n14637), .ZN(n12184) );
  OAI21_X1 U14486 ( .B1(n12185), .B2(n14637), .A(n12184), .ZN(n12186) );
  XNOR2_X1 U14487 ( .A(n14510), .B(n12229), .ZN(n12188) );
  AOI21_X1 U14488 ( .B1(n12189), .B2(n12188), .A(n14296), .ZN(n12191) );
  XNOR2_X1 U14489 ( .A(n14633), .B(n12236), .ZN(n12187) );
  OAI21_X1 U14490 ( .B1(n12189), .B2(n12188), .A(n12187), .ZN(n12190) );
  NAND2_X1 U14491 ( .A1(n12191), .A2(n12190), .ZN(n12195) );
  NAND2_X1 U14492 ( .A1(n14489), .A2(n12236), .ZN(n12193) );
  OR2_X1 U14493 ( .A1(n14489), .A2(n12228), .ZN(n12192) );
  MUX2_X1 U14494 ( .A(n12193), .B(n12192), .S(n14475), .Z(n12194) );
  NAND2_X1 U14495 ( .A1(n12195), .A2(n12194), .ZN(n12198) );
  MUX2_X1 U14496 ( .A(n14471), .B(n14679), .S(n12228), .Z(n12197) );
  INV_X1 U14497 ( .A(n14471), .ZN(n14147) );
  MUX2_X1 U14498 ( .A(n14147), .B(n14464), .S(n12131), .Z(n12196) );
  OAI21_X1 U14499 ( .B1(n12198), .B2(n12197), .A(n12196), .ZN(n12200) );
  NAND2_X1 U14500 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  MUX2_X1 U14501 ( .A(n14299), .B(n14443), .S(n12131), .Z(n12202) );
  MUX2_X1 U14502 ( .A(n14299), .B(n14443), .S(n12228), .Z(n12201) );
  MUX2_X1 U14503 ( .A(n14275), .B(n6457), .S(n12228), .Z(n12204) );
  MUX2_X1 U14504 ( .A(n6457), .B(n14275), .S(n12228), .Z(n12203) );
  MUX2_X1 U14505 ( .A(n14398), .B(n14600), .S(n12229), .Z(n12207) );
  MUX2_X1 U14506 ( .A(n14398), .B(n14600), .S(n12228), .Z(n12205) );
  MUX2_X1 U14507 ( .A(n14278), .B(n14593), .S(n12228), .Z(n12211) );
  MUX2_X1 U14508 ( .A(n14278), .B(n14593), .S(n12229), .Z(n12208) );
  NAND2_X1 U14509 ( .A1(n12209), .A2(n12208), .ZN(n12215) );
  INV_X1 U14510 ( .A(n12210), .ZN(n12213) );
  INV_X1 U14511 ( .A(n12211), .ZN(n12212) );
  NAND2_X1 U14512 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  MUX2_X1 U14513 ( .A(n14399), .B(n14389), .S(n12229), .Z(n12217) );
  MUX2_X1 U14514 ( .A(n14399), .B(n14389), .S(n12228), .Z(n12216) );
  MUX2_X1 U14515 ( .A(n14281), .B(n14583), .S(n12228), .Z(n12221) );
  NAND2_X1 U14516 ( .A1(n12220), .A2(n12221), .ZN(n12219) );
  MUX2_X1 U14517 ( .A(n14281), .B(n14583), .S(n12229), .Z(n12218) );
  NAND2_X1 U14518 ( .A1(n12219), .A2(n12218), .ZN(n12225) );
  INV_X1 U14519 ( .A(n12220), .ZN(n12223) );
  INV_X1 U14520 ( .A(n12221), .ZN(n12222) );
  NAND2_X1 U14521 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  MUX2_X1 U14522 ( .A(n14284), .B(n14576), .S(n12131), .Z(n12227) );
  MUX2_X1 U14523 ( .A(n14284), .B(n14576), .S(n12228), .Z(n12226) );
  MUX2_X1 U14524 ( .A(n14315), .B(n14335), .S(n12228), .Z(n12232) );
  NAND2_X1 U14525 ( .A1(n12233), .A2(n12232), .ZN(n12231) );
  MUX2_X1 U14526 ( .A(n14315), .B(n14335), .S(n12229), .Z(n12230) );
  NAND2_X1 U14527 ( .A1(n12231), .A2(n12230), .ZN(n12235) );
  INV_X1 U14528 ( .A(n12409), .ZN(n14146) );
  MUX2_X1 U14529 ( .A(n14146), .B(n14321), .S(n12236), .Z(n12237) );
  INV_X1 U14530 ( .A(n12241), .ZN(n12244) );
  NAND2_X1 U14531 ( .A1(n12244), .A2(n12242), .ZN(n12259) );
  AOI211_X1 U14532 ( .C1(n12246), .C2(n12250), .A(n12256), .B(n12259), .ZN(
        n12264) );
  INV_X1 U14533 ( .A(n12246), .ZN(n12247) );
  NAND3_X1 U14534 ( .A1(n12249), .A2(n12248), .A3(n12247), .ZN(n12260) );
  NAND3_X1 U14535 ( .A1(n12252), .A2(n12251), .A3(n12250), .ZN(n12258) );
  NAND3_X1 U14536 ( .A1(n12254), .A2(n12253), .A3(n15007), .ZN(n12255) );
  OAI211_X1 U14537 ( .C1(n12072), .C2(n12256), .A(n12255), .B(P1_B_REG_SCAN_IN), .ZN(n12257) );
  OAI211_X1 U14538 ( .C1(n12260), .C2(n12259), .A(n12258), .B(n12257), .ZN(
        n12261) );
  AOI21_X1 U14539 ( .B1(n12266), .B2(n12264), .A(n12263), .ZN(n12265) );
  OAI21_X1 U14540 ( .B1(n12267), .B2(n12266), .A(n12265), .ZN(P1_U3242) );
  INV_X1 U14541 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U14542 ( .A1(n14905), .A2(n12404), .ZN(n12274) );
  NAND2_X1 U14543 ( .A1(n14922), .A2(n12400), .ZN(n12273) );
  NAND2_X1 U14544 ( .A1(n12274), .A2(n12273), .ZN(n12275) );
  XNOR2_X1 U14545 ( .A(n12275), .B(n12292), .ZN(n12283) );
  NOR2_X1 U14546 ( .A1(n12360), .A2(n12276), .ZN(n12277) );
  AOI21_X1 U14547 ( .B1(n14905), .B2(n12400), .A(n12277), .ZN(n12284) );
  XNOR2_X1 U14548 ( .A(n12283), .B(n12284), .ZN(n14907) );
  NAND2_X1 U14549 ( .A1(n14547), .A2(n12404), .ZN(n12279) );
  NAND2_X1 U14550 ( .A1(n14910), .A2(n12400), .ZN(n12278) );
  NAND2_X1 U14551 ( .A1(n12279), .A2(n12278), .ZN(n12280) );
  XNOR2_X1 U14552 ( .A(n12280), .B(n12292), .ZN(n12287) );
  NOR2_X1 U14553 ( .A1(n12360), .A2(n12281), .ZN(n12282) );
  AOI21_X1 U14554 ( .B1(n14547), .B2(n12400), .A(n12282), .ZN(n12288) );
  XNOR2_X1 U14555 ( .A(n12287), .B(n12288), .ZN(n14920) );
  INV_X1 U14556 ( .A(n12283), .ZN(n12285) );
  OR2_X1 U14557 ( .A1(n12285), .A2(n12284), .ZN(n14918) );
  INV_X1 U14558 ( .A(n12287), .ZN(n12289) );
  NAND2_X1 U14559 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  AOI22_X1 U14560 ( .A1(n12291), .A2(n12400), .B1(n10120), .B2(n14924), .ZN(
        n12295) );
  AOI22_X1 U14561 ( .A1(n12291), .A2(n12404), .B1(n12400), .B2(n14924), .ZN(
        n12293) );
  XNOR2_X1 U14562 ( .A(n12293), .B(n12292), .ZN(n12294) );
  XOR2_X1 U14563 ( .A(n12295), .B(n12294), .Z(n14037) );
  INV_X1 U14564 ( .A(n12294), .ZN(n12297) );
  INV_X1 U14565 ( .A(n12295), .ZN(n12296) );
  NOR2_X1 U14566 ( .A1(n12360), .A2(n12299), .ZN(n12300) );
  AOI21_X1 U14567 ( .B1(n12301), .B2(n10039), .A(n12300), .ZN(n12309) );
  AOI22_X1 U14568 ( .A1(n12301), .A2(n12404), .B1(n12400), .B2(n14897), .ZN(
        n12302) );
  XNOR2_X1 U14569 ( .A(n12302), .B(n12292), .ZN(n12310) );
  XOR2_X1 U14570 ( .A(n12309), .B(n12310), .Z(n14097) );
  NAND2_X1 U14571 ( .A1(n12308), .A2(n12404), .ZN(n12304) );
  OR2_X1 U14572 ( .A1(n12306), .A2(n12361), .ZN(n12303) );
  NAND2_X1 U14573 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  XNOR2_X1 U14574 ( .A(n12305), .B(n12292), .ZN(n12314) );
  NOR2_X1 U14575 ( .A1(n12360), .A2(n12306), .ZN(n12307) );
  AOI21_X1 U14576 ( .B1(n12308), .B2(n10039), .A(n12307), .ZN(n12312) );
  XNOR2_X1 U14577 ( .A(n12314), .B(n12312), .ZN(n14895) );
  OR2_X1 U14578 ( .A1(n12310), .A2(n12309), .ZN(n14892) );
  INV_X1 U14579 ( .A(n12312), .ZN(n12313) );
  NAND2_X1 U14580 ( .A1(n14264), .A2(n12404), .ZN(n12317) );
  NAND2_X1 U14581 ( .A1(n14898), .A2(n12400), .ZN(n12316) );
  NAND2_X1 U14582 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  XNOR2_X1 U14583 ( .A(n12318), .B(n12292), .ZN(n12319) );
  AOI22_X1 U14584 ( .A1(n14264), .A2(n12400), .B1(n10120), .B2(n14898), .ZN(
        n14137) );
  INV_X1 U14585 ( .A(n12319), .ZN(n12320) );
  OAI22_X1 U14586 ( .A1(n14647), .A2(n12361), .B1(n14291), .B2(n12360), .ZN(
        n12326) );
  NAND2_X1 U14587 ( .A1(n14535), .A2(n12404), .ZN(n12323) );
  NAND2_X1 U14588 ( .A1(n14507), .A2(n12400), .ZN(n12322) );
  NAND2_X1 U14589 ( .A1(n12323), .A2(n12322), .ZN(n12324) );
  XNOR2_X1 U14590 ( .A(n12324), .B(n12292), .ZN(n12325) );
  XOR2_X1 U14591 ( .A(n12326), .B(n12325), .Z(n14052) );
  INV_X1 U14592 ( .A(n12325), .ZN(n12328) );
  INV_X1 U14593 ( .A(n12326), .ZN(n12327) );
  NAND2_X1 U14594 ( .A1(n12328), .A2(n12327), .ZN(n12329) );
  NAND2_X1 U14595 ( .A1(n14637), .A2(n12404), .ZN(n12331) );
  NAND2_X1 U14596 ( .A1(n14488), .A2(n12400), .ZN(n12330) );
  NAND2_X1 U14597 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  XNOR2_X1 U14598 ( .A(n12332), .B(n12292), .ZN(n12333) );
  AOI22_X1 U14599 ( .A1(n14637), .A2(n12400), .B1(n9737), .B2(n14488), .ZN(
        n12334) );
  XNOR2_X1 U14600 ( .A(n12333), .B(n12334), .ZN(n14074) );
  NAND2_X1 U14601 ( .A1(n14073), .A2(n14074), .ZN(n12337) );
  INV_X1 U14602 ( .A(n12333), .ZN(n12335) );
  NAND2_X1 U14603 ( .A1(n12335), .A2(n12334), .ZN(n12336) );
  NAND2_X1 U14604 ( .A1(n14633), .A2(n12404), .ZN(n12339) );
  NAND2_X1 U14605 ( .A1(n14510), .A2(n12400), .ZN(n12338) );
  NAND2_X1 U14606 ( .A1(n12339), .A2(n12338), .ZN(n12340) );
  XNOR2_X1 U14607 ( .A(n12340), .B(n12292), .ZN(n12341) );
  AOI22_X1 U14608 ( .A1(n14633), .A2(n12400), .B1(n10120), .B2(n14510), .ZN(
        n12342) );
  XNOR2_X1 U14609 ( .A(n12341), .B(n12342), .ZN(n14117) );
  INV_X1 U14610 ( .A(n12341), .ZN(n12343) );
  NAND2_X1 U14611 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  AOI22_X1 U14612 ( .A1(n14475), .A2(n12404), .B1(n10039), .B2(n14489), .ZN(
        n12345) );
  XNOR2_X1 U14613 ( .A(n12345), .B(n12292), .ZN(n12346) );
  AOI22_X1 U14614 ( .A1(n14475), .A2(n12400), .B1(n9737), .B2(n14489), .ZN(
        n12347) );
  XNOR2_X1 U14615 ( .A(n12346), .B(n12347), .ZN(n14018) );
  INV_X1 U14616 ( .A(n12346), .ZN(n12349) );
  INV_X1 U14617 ( .A(n12347), .ZN(n12348) );
  OAI22_X1 U14618 ( .A1(n14679), .A2(n12361), .B1(n14471), .B2(n12360), .ZN(
        n12352) );
  OAI22_X1 U14619 ( .A1(n14679), .A2(n12350), .B1(n14471), .B2(n12361), .ZN(
        n12351) );
  XNOR2_X1 U14620 ( .A(n12351), .B(n12292), .ZN(n12353) );
  XOR2_X1 U14621 ( .A(n12352), .B(n12353), .Z(n14089) );
  NAND2_X1 U14622 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  AOI22_X1 U14623 ( .A1(n14443), .A2(n12404), .B1(n10039), .B2(n14299), .ZN(
        n12355) );
  XNOR2_X1 U14624 ( .A(n12355), .B(n12292), .ZN(n12358) );
  AOI22_X1 U14625 ( .A1(n14443), .A2(n12400), .B1(n10120), .B2(n14299), .ZN(
        n12357) );
  XNOR2_X1 U14626 ( .A(n12358), .B(n12357), .ZN(n14029) );
  INV_X1 U14627 ( .A(n14029), .ZN(n12356) );
  NAND2_X1 U14628 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  NAND2_X1 U14629 ( .A1(n14026), .A2(n12359), .ZN(n14106) );
  OAI22_X1 U14630 ( .A1(n14606), .A2(n12361), .B1(n14301), .B2(n12360), .ZN(
        n12366) );
  NAND2_X1 U14631 ( .A1(n6457), .A2(n12404), .ZN(n12363) );
  NAND2_X1 U14632 ( .A1(n14275), .A2(n12400), .ZN(n12362) );
  NAND2_X1 U14633 ( .A1(n12363), .A2(n12362), .ZN(n12364) );
  XNOR2_X1 U14634 ( .A(n12364), .B(n12292), .ZN(n12365) );
  XOR2_X1 U14635 ( .A(n12366), .B(n12365), .Z(n14107) );
  INV_X1 U14636 ( .A(n12365), .ZN(n12368) );
  INV_X1 U14637 ( .A(n12366), .ZN(n12367) );
  NAND2_X1 U14638 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  NAND2_X1 U14639 ( .A1(n14600), .A2(n12404), .ZN(n12371) );
  NAND2_X1 U14640 ( .A1(n14398), .A2(n12400), .ZN(n12370) );
  NAND2_X1 U14641 ( .A1(n12371), .A2(n12370), .ZN(n12372) );
  XNOR2_X1 U14642 ( .A(n12372), .B(n12292), .ZN(n12373) );
  AOI22_X1 U14643 ( .A1(n14600), .A2(n12400), .B1(n10120), .B2(n14398), .ZN(
        n12374) );
  XNOR2_X1 U14644 ( .A(n12373), .B(n12374), .ZN(n14012) );
  INV_X1 U14645 ( .A(n12373), .ZN(n12375) );
  NAND2_X1 U14646 ( .A1(n14593), .A2(n12404), .ZN(n12377) );
  NAND2_X1 U14647 ( .A1(n14278), .A2(n12400), .ZN(n12376) );
  NAND2_X1 U14648 ( .A1(n12377), .A2(n12376), .ZN(n12378) );
  XNOR2_X1 U14649 ( .A(n12378), .B(n12292), .ZN(n12379) );
  AOI22_X1 U14650 ( .A1(n14593), .A2(n12400), .B1(n10120), .B2(n14278), .ZN(
        n12380) );
  XNOR2_X1 U14651 ( .A(n12379), .B(n12380), .ZN(n14082) );
  INV_X1 U14652 ( .A(n12379), .ZN(n12381) );
  NAND2_X1 U14653 ( .A1(n14389), .A2(n12404), .ZN(n12383) );
  NAND2_X1 U14654 ( .A1(n14399), .A2(n12400), .ZN(n12382) );
  NAND2_X1 U14655 ( .A1(n12383), .A2(n12382), .ZN(n12384) );
  XNOR2_X1 U14656 ( .A(n12384), .B(n12292), .ZN(n12385) );
  AOI22_X1 U14657 ( .A1(n14389), .A2(n12400), .B1(n9737), .B2(n14399), .ZN(
        n12386) );
  XNOR2_X1 U14658 ( .A(n12385), .B(n12386), .ZN(n14046) );
  NAND2_X1 U14659 ( .A1(n14045), .A2(n14046), .ZN(n12389) );
  INV_X1 U14660 ( .A(n12385), .ZN(n12387) );
  NAND2_X1 U14661 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U14662 ( .A1(n14583), .A2(n12404), .ZN(n12391) );
  NAND2_X1 U14663 ( .A1(n14281), .A2(n12400), .ZN(n12390) );
  NAND2_X1 U14664 ( .A1(n12391), .A2(n12390), .ZN(n12392) );
  XNOR2_X1 U14665 ( .A(n12392), .B(n12292), .ZN(n12393) );
  AOI22_X1 U14666 ( .A1(n14583), .A2(n12400), .B1(n9737), .B2(n14281), .ZN(
        n12394) );
  XNOR2_X1 U14667 ( .A(n12393), .B(n12394), .ZN(n14126) );
  INV_X1 U14668 ( .A(n12393), .ZN(n12395) );
  NAND2_X1 U14669 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  NAND2_X1 U14670 ( .A1(n14576), .A2(n12404), .ZN(n12398) );
  NAND2_X1 U14671 ( .A1(n14284), .A2(n12400), .ZN(n12397) );
  NAND2_X1 U14672 ( .A1(n12398), .A2(n12397), .ZN(n12399) );
  XNOR2_X1 U14673 ( .A(n12399), .B(n12292), .ZN(n12401) );
  AOI22_X1 U14674 ( .A1(n14576), .A2(n12400), .B1(n10120), .B2(n14284), .ZN(
        n12402) );
  XNOR2_X1 U14675 ( .A(n12401), .B(n12402), .ZN(n14005) );
  INV_X1 U14676 ( .A(n12401), .ZN(n12403) );
  AOI22_X1 U14677 ( .A1(n14335), .A2(n12400), .B1(n10120), .B2(n14315), .ZN(
        n12407) );
  AOI22_X1 U14678 ( .A1(n14335), .A2(n12404), .B1(n10039), .B2(n14315), .ZN(
        n12405) );
  XNOR2_X1 U14679 ( .A(n12405), .B(n12292), .ZN(n12406) );
  XOR2_X1 U14680 ( .A(n12407), .B(n12406), .Z(n12408) );
  OR2_X1 U14681 ( .A1(n12409), .A2(n14527), .ZN(n12411) );
  NAND2_X1 U14682 ( .A1(n14284), .A2(n15007), .ZN(n12410) );
  AND2_X1 U14683 ( .A1(n12411), .A2(n12410), .ZN(n14569) );
  OAI22_X1 U14684 ( .A1(n14111), .A2(n14569), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15354), .ZN(n12413) );
  NOR2_X1 U14685 ( .A1(n14662), .A2(n14927), .ZN(n12412) );
  AOI211_X1 U14686 ( .C1(n14330), .C2(n14113), .A(n12413), .B(n12412), .ZN(
        n12414) );
  OAI21_X1 U14687 ( .B1(n12415), .B2(n14133), .A(n12414), .ZN(P1_U3220) );
  INV_X1 U14688 ( .A(n12416), .ZN(n12418) );
  OAI222_X1 U14689 ( .A1(n12420), .A2(n12419), .B1(n13303), .B2(n12418), .C1(
        n12417), .C2(P3_U3151), .ZN(P3_U3266) );
  NAND2_X1 U14690 ( .A1(n15196), .A2(n12421), .ZN(n12422) );
  OAI21_X1 U14691 ( .B1(n14853), .B2(n15197), .A(n14861), .ZN(n12425) );
  NAND2_X1 U14692 ( .A1(n14853), .A2(n15197), .ZN(n12424) );
  NAND2_X1 U14693 ( .A1(n12425), .A2(n12424), .ZN(n14836) );
  NAND2_X1 U14694 ( .A1(n14836), .A2(n12426), .ZN(n12428) );
  INV_X1 U14695 ( .A(n14846), .ZN(n12473) );
  NAND2_X1 U14696 ( .A1(n12687), .A2(n12473), .ZN(n12427) );
  AND2_X1 U14697 ( .A1(n12621), .A2(n14838), .ZN(n12430) );
  INV_X1 U14698 ( .A(n14838), .ZN(n12563) );
  NAND2_X1 U14699 ( .A1(n12563), .A2(n13293), .ZN(n12429) );
  OR2_X1 U14700 ( .A1(n13289), .A2(n13119), .ZN(n12431) );
  NAND2_X1 U14701 ( .A1(n13089), .A2(n13100), .ZN(n12432) );
  NAND2_X1 U14702 ( .A1(n12433), .A2(n12432), .ZN(n13071) );
  NAND2_X1 U14703 ( .A1(n13071), .A2(n13072), .ZN(n12435) );
  INV_X1 U14704 ( .A(n13085), .ZN(n12685) );
  NAND2_X1 U14705 ( .A1(n13076), .A2(n12685), .ZN(n12434) );
  NAND2_X1 U14706 ( .A1(n12435), .A2(n12434), .ZN(n13056) );
  INV_X1 U14707 ( .A(n13075), .ZN(n12684) );
  NAND2_X1 U14708 ( .A1(n12584), .A2(n12684), .ZN(n12436) );
  OR2_X1 U14709 ( .A1(n12643), .A2(n12683), .ZN(n12437) );
  NAND2_X1 U14710 ( .A1(n13045), .A2(n12437), .ZN(n13027) );
  INV_X1 U14711 ( .A(n13027), .ZN(n12438) );
  NAND2_X1 U14712 ( .A1(n12438), .A2(n13036), .ZN(n13030) );
  OR2_X1 U14713 ( .A1(n13269), .A2(n13049), .ZN(n12439) );
  NAND2_X1 U14714 ( .A1(n13030), .A2(n12439), .ZN(n13018) );
  NAND2_X1 U14715 ( .A1(n12605), .A2(n12681), .ZN(n12440) );
  OR2_X1 U14716 ( .A1(n13170), .A2(n12625), .ZN(n12442) );
  NAND2_X1 U14717 ( .A1(n13003), .A2(n12442), .ZN(n12987) );
  NAND2_X1 U14718 ( .A1(n12996), .A2(n12443), .ZN(n12444) );
  NAND2_X1 U14719 ( .A1(n12987), .A2(n12444), .ZN(n12446) );
  INV_X1 U14720 ( .A(n12942), .ZN(n13241) );
  NOR2_X1 U14721 ( .A1(n12918), .A2(n12448), .ZN(n12904) );
  NAND2_X1 U14722 ( .A1(n12904), .A2(n12903), .ZN(n12909) );
  INV_X1 U14723 ( .A(n13139), .ZN(n12913) );
  NAND2_X1 U14724 ( .A1(n12909), .A2(n12450), .ZN(n12451) );
  XNOR2_X1 U14725 ( .A(n12451), .B(n8230), .ZN(n12456) );
  NAND2_X1 U14726 ( .A1(n12452), .A2(P3_B_REG_SCAN_IN), .ZN(n12453) );
  NAND2_X1 U14727 ( .A1(n15215), .A2(n12453), .ZN(n12894) );
  OAI22_X1 U14728 ( .A1(n12919), .A2(n14857), .B1(n12454), .B2(n12894), .ZN(
        n12455) );
  NAND2_X1 U14729 ( .A1(n12457), .A2(n15244), .ZN(n12896) );
  OAI21_X1 U14730 ( .B1(n15248), .B2(n12458), .A(n12896), .ZN(n12462) );
  XNOR2_X1 U14731 ( .A(n12460), .B(n12459), .ZN(n13135) );
  NAND2_X1 U14732 ( .A1(n15223), .A2(n15202), .ZN(n14860) );
  NOR2_X1 U14733 ( .A1(n13135), .A2(n13125), .ZN(n12461) );
  AOI211_X1 U14734 ( .C1(n13107), .C2(n13133), .A(n12462), .B(n12461), .ZN(
        n12463) );
  OAI21_X1 U14735 ( .B1(n13138), .B2(n15250), .A(n12463), .ZN(P3_U3204) );
  XNOR2_X1 U14736 ( .A(n12464), .B(n12543), .ZN(n12540) );
  XNOR2_X1 U14737 ( .A(n12540), .B(n12677), .ZN(n12541) );
  INV_X1 U14738 ( .A(n12465), .ZN(n12466) );
  NAND2_X1 U14739 ( .A1(n12466), .A2(n12635), .ZN(n12467) );
  XNOR2_X1 U14740 ( .A(n12543), .B(n12636), .ZN(n12469) );
  NAND2_X1 U14741 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  NAND2_X1 U14742 ( .A1(n12632), .A2(n12633), .ZN(n12631) );
  NAND2_X1 U14743 ( .A1(n12631), .A2(n12472), .ZN(n12560) );
  XNOR2_X1 U14744 ( .A(n10859), .B(n12473), .ZN(n12558) );
  INV_X1 U14745 ( .A(n12687), .ZN(n14858) );
  AND2_X1 U14746 ( .A1(n12558), .A2(n14858), .ZN(n12474) );
  XNOR2_X1 U14747 ( .A(n10859), .B(n12621), .ZN(n12475) );
  NAND2_X1 U14748 ( .A1(n12475), .A2(n12563), .ZN(n12614) );
  INV_X1 U14749 ( .A(n12475), .ZN(n12476) );
  NAND2_X1 U14750 ( .A1(n12476), .A2(n14838), .ZN(n12615) );
  XNOR2_X1 U14751 ( .A(n13289), .B(n12503), .ZN(n12517) );
  INV_X1 U14752 ( .A(n12517), .ZN(n12477) );
  NAND2_X1 U14753 ( .A1(n12477), .A2(n12686), .ZN(n12478) );
  XNOR2_X1 U14754 ( .A(n13089), .B(n12543), .ZN(n12480) );
  XNOR2_X1 U14755 ( .A(n12480), .B(n13100), .ZN(n12663) );
  NAND2_X1 U14756 ( .A1(n12664), .A2(n12663), .ZN(n12483) );
  INV_X1 U14757 ( .A(n12480), .ZN(n12481) );
  NAND2_X1 U14758 ( .A1(n12481), .A2(n13100), .ZN(n12482) );
  XNOR2_X1 U14759 ( .A(n13076), .B(n12503), .ZN(n12576) );
  AND2_X1 U14760 ( .A1(n12576), .A2(n12685), .ZN(n12484) );
  INV_X1 U14761 ( .A(n12576), .ZN(n12485) );
  NAND2_X1 U14762 ( .A1(n12485), .A2(n13085), .ZN(n12486) );
  XNOR2_X1 U14763 ( .A(n12584), .B(n12543), .ZN(n12487) );
  XNOR2_X1 U14764 ( .A(n12487), .B(n13075), .ZN(n12585) );
  INV_X1 U14765 ( .A(n12487), .ZN(n12488) );
  NAND2_X1 U14766 ( .A1(n12488), .A2(n12684), .ZN(n12489) );
  XNOR2_X1 U14767 ( .A(n12643), .B(n12543), .ZN(n12490) );
  XNOR2_X1 U14768 ( .A(n12490), .B(n12683), .ZN(n12646) );
  NAND2_X1 U14769 ( .A1(n12647), .A2(n12646), .ZN(n12645) );
  INV_X1 U14770 ( .A(n12490), .ZN(n12491) );
  NAND2_X1 U14771 ( .A1(n12491), .A2(n12683), .ZN(n12492) );
  NAND2_X1 U14772 ( .A1(n12645), .A2(n12492), .ZN(n12535) );
  XNOR2_X1 U14773 ( .A(n13269), .B(n12543), .ZN(n12493) );
  XNOR2_X1 U14774 ( .A(n12493), .B(n13049), .ZN(n12534) );
  NAND2_X1 U14775 ( .A1(n12535), .A2(n12534), .ZN(n12533) );
  NAND2_X1 U14776 ( .A1(n12493), .A2(n12682), .ZN(n12494) );
  NAND2_X1 U14777 ( .A1(n12533), .A2(n12494), .ZN(n12608) );
  XNOR2_X1 U14778 ( .A(n12605), .B(n10859), .ZN(n12495) );
  XNOR2_X1 U14779 ( .A(n12495), .B(n12681), .ZN(n12607) );
  INV_X1 U14780 ( .A(n12495), .ZN(n12496) );
  NAND2_X1 U14781 ( .A1(n12496), .A2(n12681), .ZN(n12497) );
  XNOR2_X1 U14782 ( .A(n13170), .B(n12543), .ZN(n12498) );
  XNOR2_X1 U14783 ( .A(n12498), .B(n13020), .ZN(n12552) );
  XNOR2_X1 U14784 ( .A(n13257), .B(n12543), .ZN(n12499) );
  INV_X1 U14785 ( .A(n12499), .ZN(n12500) );
  AND2_X1 U14786 ( .A1(n12501), .A2(n12500), .ZN(n12502) );
  XNOR2_X1 U14787 ( .A(n12967), .B(n12543), .ZN(n12597) );
  XNOR2_X1 U14788 ( .A(n12974), .B(n12503), .ZN(n12594) );
  INV_X1 U14789 ( .A(n12594), .ZN(n12504) );
  OAI22_X1 U14790 ( .A1(n12597), .A2(n12978), .B1(n12965), .B2(n12504), .ZN(
        n12508) );
  OAI21_X1 U14791 ( .B1(n12594), .B2(n12988), .A(n12527), .ZN(n12506) );
  NOR2_X1 U14792 ( .A1(n12527), .A2(n12988), .ZN(n12505) );
  AOI22_X1 U14793 ( .A1(n12597), .A2(n12506), .B1(n12505), .B2(n12504), .ZN(
        n12507) );
  XNOR2_X1 U14794 ( .A(n12954), .B(n12543), .ZN(n12509) );
  XNOR2_X1 U14795 ( .A(n12509), .B(n12679), .ZN(n12570) );
  XNOR2_X1 U14796 ( .A(n12942), .B(n12543), .ZN(n12510) );
  XNOR2_X1 U14797 ( .A(n12510), .B(n12948), .ZN(n12654) );
  INV_X1 U14798 ( .A(n12510), .ZN(n12511) );
  XOR2_X1 U14799 ( .A(n12541), .B(n12542), .Z(n12516) );
  AOI22_X1 U14800 ( .A1(n12678), .A2(n12668), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12512) );
  OAI21_X1 U14801 ( .B1(n12919), .B2(n12666), .A(n12512), .ZN(n12514) );
  NOR2_X1 U14802 ( .A1(n13238), .A2(n12652), .ZN(n12513) );
  AOI211_X1 U14803 ( .C1(n12926), .C2(n12656), .A(n12514), .B(n12513), .ZN(
        n12515) );
  OAI21_X1 U14804 ( .B1(n12516), .B2(n12674), .A(n12515), .ZN(P3_U3154) );
  XNOR2_X1 U14805 ( .A(n12517), .B(n12686), .ZN(n12518) );
  XNOR2_X1 U14806 ( .A(n12519), .B(n12518), .ZN(n12526) );
  INV_X1 U14807 ( .A(n13289), .ZN(n13106) );
  INV_X1 U14808 ( .A(n13103), .ZN(n12520) );
  NAND2_X1 U14809 ( .A1(n12656), .A2(n12520), .ZN(n12523) );
  INV_X1 U14810 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12521) );
  NOR2_X1 U14811 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12521), .ZN(n12768) );
  AOI21_X1 U14812 ( .B1(n12668), .B2(n14838), .A(n12768), .ZN(n12522) );
  OAI211_X1 U14813 ( .C1(n13074), .C2(n12666), .A(n12523), .B(n12522), .ZN(
        n12524) );
  AOI21_X1 U14814 ( .B1(n13106), .B2(n12672), .A(n12524), .ZN(n12525) );
  OAI21_X1 U14815 ( .B1(n12526), .B2(n12674), .A(n12525), .ZN(P3_U3155) );
  XNOR2_X1 U14816 ( .A(n12595), .B(n12594), .ZN(n12596) );
  XNOR2_X1 U14817 ( .A(n12596), .B(n12965), .ZN(n12532) );
  NAND2_X1 U14818 ( .A1(n12656), .A2(n12981), .ZN(n12529) );
  AOI22_X1 U14819 ( .A1(n12527), .A2(n12655), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12528) );
  OAI211_X1 U14820 ( .C1(n13004), .C2(n12659), .A(n12529), .B(n12528), .ZN(
        n12530) );
  AOI21_X1 U14821 ( .B1(n12974), .B2(n12672), .A(n12530), .ZN(n12531) );
  OAI21_X1 U14822 ( .B1(n12532), .B2(n12674), .A(n12531), .ZN(P3_U3156) );
  OAI211_X1 U14823 ( .C1(n12535), .C2(n12534), .A(n12533), .B(n12644), .ZN(
        n12539) );
  NAND2_X1 U14824 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12886)
         );
  OAI21_X1 U14825 ( .B1(n12666), .B2(n13028), .A(n12886), .ZN(n12537) );
  NOR2_X1 U14826 ( .A1(n12670), .A2(n13032), .ZN(n12536) );
  AOI211_X1 U14827 ( .C1(n12668), .C2(n12683), .A(n12537), .B(n12536), .ZN(
        n12538) );
  OAI211_X1 U14828 ( .C1(n12652), .C2(n13269), .A(n12539), .B(n12538), .ZN(
        P3_U3159) );
  AOI22_X1 U14829 ( .A1(n12542), .A2(n12541), .B1(n12934), .B2(n12540), .ZN(
        n12545) );
  XNOR2_X1 U14830 ( .A(n12905), .B(n12543), .ZN(n12544) );
  XNOR2_X1 U14831 ( .A(n12545), .B(n12544), .ZN(n12550) );
  AOI22_X1 U14832 ( .A1(n12677), .A2(n12668), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12546) );
  OAI21_X1 U14833 ( .B1(n12907), .B2(n12666), .A(n12546), .ZN(n12548) );
  NOR2_X1 U14834 ( .A1(n12913), .A2(n12652), .ZN(n12547) );
  AOI211_X1 U14835 ( .C1(n12911), .C2(n12656), .A(n12548), .B(n12547), .ZN(
        n12549) );
  OAI21_X1 U14836 ( .B1(n12550), .B2(n12674), .A(n12549), .ZN(P3_U3160) );
  AOI21_X1 U14837 ( .B1(n12552), .B2(n12551), .A(n6511), .ZN(n12557) );
  NAND2_X1 U14838 ( .A1(n12656), .A2(n13007), .ZN(n12554) );
  AOI22_X1 U14839 ( .A1(n12668), .A2(n12681), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12553) );
  OAI211_X1 U14840 ( .C1(n13004), .C2(n12666), .A(n12554), .B(n12553), .ZN(
        n12555) );
  AOI21_X1 U14841 ( .B1(n13170), .B2(n12672), .A(n12555), .ZN(n12556) );
  OAI21_X1 U14842 ( .B1(n12557), .B2(n12674), .A(n12556), .ZN(P3_U3163) );
  XNOR2_X1 U14843 ( .A(n12558), .B(n12687), .ZN(n12559) );
  XNOR2_X1 U14844 ( .A(n12560), .B(n12559), .ZN(n12561) );
  NAND2_X1 U14845 ( .A1(n12561), .A2(n12644), .ZN(n12567) );
  OAI22_X1 U14846 ( .A1(n14846), .A2(n12652), .B1(n12659), .B2(n12633), .ZN(
        n12565) );
  OAI21_X1 U14847 ( .B1(n12666), .B2(n12563), .A(n12562), .ZN(n12564) );
  NOR2_X1 U14848 ( .A1(n12565), .A2(n12564), .ZN(n12566) );
  OAI211_X1 U14849 ( .C1(n12568), .C2(n12670), .A(n12567), .B(n12566), .ZN(
        P3_U3164) );
  XOR2_X1 U14850 ( .A(n12570), .B(n12569), .Z(n12575) );
  NAND2_X1 U14851 ( .A1(n12656), .A2(n12955), .ZN(n12572) );
  AOI22_X1 U14852 ( .A1(n12678), .A2(n12655), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12571) );
  OAI211_X1 U14853 ( .C1(n12978), .C2(n12659), .A(n12572), .B(n12571), .ZN(
        n12573) );
  AOI21_X1 U14854 ( .B1(n12954), .B2(n12672), .A(n12573), .ZN(n12574) );
  OAI21_X1 U14855 ( .B1(n12575), .B2(n12674), .A(n12574), .ZN(P3_U3165) );
  XNOR2_X1 U14856 ( .A(n12576), .B(n13085), .ZN(n12577) );
  XNOR2_X1 U14857 ( .A(n12578), .B(n12577), .ZN(n12583) );
  NAND2_X1 U14858 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12821)
         );
  OAI21_X1 U14859 ( .B1(n12666), .B2(n13075), .A(n12821), .ZN(n12579) );
  AOI21_X1 U14860 ( .B1(n12668), .B2(n13100), .A(n12579), .ZN(n12580) );
  OAI21_X1 U14861 ( .B1(n12670), .B2(n13077), .A(n12580), .ZN(n12581) );
  AOI21_X1 U14862 ( .B1(n12672), .B2(n13076), .A(n12581), .ZN(n12582) );
  OAI21_X1 U14863 ( .B1(n12583), .B2(n12674), .A(n12582), .ZN(P3_U3166) );
  INV_X1 U14864 ( .A(n12584), .ZN(n13277) );
  AOI21_X1 U14865 ( .B1(n12586), .B2(n12585), .A(n12674), .ZN(n12588) );
  NAND2_X1 U14866 ( .A1(n12588), .A2(n12587), .ZN(n12593) );
  INV_X1 U14867 ( .A(n13063), .ZN(n12591) );
  OR2_X1 U14868 ( .A1(n12659), .A2(n13085), .ZN(n12589) );
  NAND2_X1 U14869 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12836)
         );
  OAI211_X1 U14870 ( .C1(n13059), .C2(n12666), .A(n12589), .B(n12836), .ZN(
        n12590) );
  AOI21_X1 U14871 ( .B1(n12656), .B2(n12591), .A(n12590), .ZN(n12592) );
  OAI211_X1 U14872 ( .C1(n13277), .C2(n12652), .A(n12593), .B(n12592), .ZN(
        P3_U3168) );
  OAI22_X1 U14873 ( .A1(n12596), .A2(n12988), .B1(n12595), .B2(n12594), .ZN(
        n12599) );
  XNOR2_X1 U14874 ( .A(n12597), .B(n12978), .ZN(n12598) );
  XNOR2_X1 U14875 ( .A(n12599), .B(n12598), .ZN(n12604) );
  NAND2_X1 U14876 ( .A1(n12656), .A2(n12968), .ZN(n12601) );
  AOI22_X1 U14877 ( .A1(n12655), .A2(n12679), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12600) );
  OAI211_X1 U14878 ( .C1(n12965), .C2(n12659), .A(n12601), .B(n12600), .ZN(
        n12602) );
  AOI21_X1 U14879 ( .B1(n12967), .B2(n12672), .A(n12602), .ZN(n12603) );
  OAI21_X1 U14880 ( .B1(n12604), .B2(n12674), .A(n12603), .ZN(P3_U3169) );
  INV_X1 U14881 ( .A(n12605), .ZN(n13265) );
  OAI211_X1 U14882 ( .C1(n12608), .C2(n12607), .A(n12606), .B(n12644), .ZN(
        n12613) );
  INV_X1 U14883 ( .A(n12609), .ZN(n13021) );
  AOI22_X1 U14884 ( .A1(n12655), .A2(n12625), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12610) );
  OAI21_X1 U14885 ( .B1(n13049), .B2(n12659), .A(n12610), .ZN(n12611) );
  AOI21_X1 U14886 ( .B1(n13021), .B2(n12656), .A(n12611), .ZN(n12612) );
  OAI211_X1 U14887 ( .C1(n13265), .C2(n12652), .A(n12613), .B(n12612), .ZN(
        P3_U3173) );
  NAND2_X1 U14888 ( .A1(n12615), .A2(n12614), .ZN(n12617) );
  XOR2_X1 U14889 ( .A(n12617), .B(n12616), .Z(n12623) );
  AND2_X1 U14890 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12757) );
  NOR2_X1 U14891 ( .A1(n12666), .A2(n13119), .ZN(n12618) );
  AOI211_X1 U14892 ( .C1(n12668), .C2(n12687), .A(n12757), .B(n12618), .ZN(
        n12619) );
  OAI21_X1 U14893 ( .B1(n13120), .B2(n12670), .A(n12619), .ZN(n12620) );
  AOI21_X1 U14894 ( .B1(n12621), .B2(n12672), .A(n12620), .ZN(n12622) );
  OAI21_X1 U14895 ( .B1(n12623), .B2(n12674), .A(n12622), .ZN(P3_U3174) );
  XNOR2_X1 U14896 ( .A(n12624), .B(n12443), .ZN(n12630) );
  NAND2_X1 U14897 ( .A1(n12656), .A2(n12992), .ZN(n12627) );
  AOI22_X1 U14898 ( .A1(n12668), .A2(n12625), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12626) );
  OAI211_X1 U14899 ( .C1(n12965), .C2(n12666), .A(n12627), .B(n12626), .ZN(
        n12628) );
  AOI21_X1 U14900 ( .B1(n12996), .B2(n12672), .A(n12628), .ZN(n12629) );
  OAI21_X1 U14901 ( .B1(n12630), .B2(n12674), .A(n12629), .ZN(P3_U3175) );
  OAI21_X1 U14902 ( .B1(n12633), .B2(n12632), .A(n12631), .ZN(n12634) );
  NAND2_X1 U14903 ( .A1(n12634), .A2(n12644), .ZN(n12642) );
  INV_X1 U14904 ( .A(n12635), .ZN(n14856) );
  OAI22_X1 U14905 ( .A1(n12636), .A2(n12652), .B1(n12659), .B2(n14856), .ZN(
        n12640) );
  INV_X1 U14906 ( .A(n12637), .ZN(n12638) );
  OAI21_X1 U14907 ( .B1(n12666), .B2(n14858), .A(n12638), .ZN(n12639) );
  NOR2_X1 U14908 ( .A1(n12640), .A2(n12639), .ZN(n12641) );
  OAI211_X1 U14909 ( .C1(n14862), .C2(n12670), .A(n12642), .B(n12641), .ZN(
        P3_U3176) );
  INV_X1 U14910 ( .A(n12643), .ZN(n13273) );
  OAI211_X1 U14911 ( .C1(n12647), .C2(n12646), .A(n12645), .B(n12644), .ZN(
        n12651) );
  NAND2_X1 U14912 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12848)
         );
  OAI21_X1 U14913 ( .B1(n12666), .B2(n13049), .A(n12848), .ZN(n12649) );
  NOR2_X1 U14914 ( .A1(n12670), .A2(n13050), .ZN(n12648) );
  AOI211_X1 U14915 ( .C1(n12668), .C2(n12684), .A(n12649), .B(n12648), .ZN(
        n12650) );
  OAI211_X1 U14916 ( .C1(n13273), .C2(n12652), .A(n12651), .B(n12650), .ZN(
        P3_U3178) );
  XOR2_X1 U14917 ( .A(n12654), .B(n12653), .Z(n12662) );
  AOI22_X1 U14918 ( .A1(n12677), .A2(n12655), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12658) );
  NAND2_X1 U14919 ( .A1(n12656), .A2(n12938), .ZN(n12657) );
  OAI211_X1 U14920 ( .C1(n12964), .C2(n12659), .A(n12658), .B(n12657), .ZN(
        n12660) );
  AOI21_X1 U14921 ( .B1(n12942), .B2(n12672), .A(n12660), .ZN(n12661) );
  OAI21_X1 U14922 ( .B1(n12662), .B2(n12674), .A(n12661), .ZN(P3_U3180) );
  XNOR2_X1 U14923 ( .A(n12664), .B(n12663), .ZN(n12675) );
  NAND2_X1 U14924 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12791)
         );
  OAI21_X1 U14925 ( .B1(n12666), .B2(n13085), .A(n12791), .ZN(n12667) );
  AOI21_X1 U14926 ( .B1(n12668), .B2(n12686), .A(n12667), .ZN(n12669) );
  OAI21_X1 U14927 ( .B1(n12670), .B2(n13090), .A(n12669), .ZN(n12671) );
  AOI21_X1 U14928 ( .B1(n12672), .B2(n13089), .A(n12671), .ZN(n12673) );
  OAI21_X1 U14929 ( .B1(n12675), .B2(n12674), .A(n12673), .ZN(P3_U3181) );
  MUX2_X1 U14930 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12676), .S(n12692), .Z(
        P3_U3522) );
  MUX2_X1 U14931 ( .A(n12677), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12680), .Z(
        P3_U3518) );
  MUX2_X1 U14932 ( .A(n12678), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12680), .Z(
        P3_U3517) );
  MUX2_X1 U14933 ( .A(n12679), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12680), .Z(
        P3_U3516) );
  MUX2_X1 U14934 ( .A(n12988), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12680), .Z(
        P3_U3514) );
  MUX2_X1 U14935 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12443), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14936 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12681), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14937 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12682), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14938 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12683), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14939 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12684), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14940 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12685), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14941 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12686), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14942 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14838), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14943 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12687), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14944 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n15197), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14945 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n15196), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14946 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12688), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14947 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n15214), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14948 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12689), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14949 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n15213), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14950 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12690), .S(n12692), .Z(
        P3_U3495) );
  MUX2_X1 U14951 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12691), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14952 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13214), .S(n12692), .Z(
        P3_U3493) );
  MUX2_X1 U14953 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12693), .S(n12692), .Z(
        P3_U3492) );
  MUX2_X1 U14954 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13213), .S(P3_U3897), .Z(
        P3_U3491) );
  AND3_X1 U14955 ( .A1(n12696), .A2(n12695), .A3(n12694), .ZN(n12697) );
  OAI21_X1 U14956 ( .B1(n12698), .B2(n12697), .A(n12890), .ZN(n12714) );
  NAND3_X1 U14957 ( .A1(n12701), .A2(n12700), .A3(n12699), .ZN(n12702) );
  AOI21_X1 U14958 ( .B1(n6590), .B2(n12702), .A(n12892), .ZN(n12703) );
  AOI211_X1 U14959 ( .C1(n15191), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n12704), .B(
        n12703), .ZN(n12713) );
  NAND2_X1 U14960 ( .A1(n12859), .A2(n12705), .ZN(n12712) );
  AND3_X1 U14961 ( .A1(n12708), .A2(n12707), .A3(n12706), .ZN(n12709) );
  OAI21_X1 U14962 ( .B1(n12710), .B2(n12709), .A(n12835), .ZN(n12711) );
  NAND4_X1 U14963 ( .A1(n12714), .A2(n12713), .A3(n12712), .A4(n12711), .ZN(
        P3_U3188) );
  AND3_X1 U14964 ( .A1(n12717), .A2(n12716), .A3(n12715), .ZN(n12718) );
  OAI21_X1 U14965 ( .B1(n12719), .B2(n12718), .A(n12890), .ZN(n12738) );
  NOR2_X1 U14966 ( .A1(n12881), .A2(n12720), .ZN(n12721) );
  AOI211_X1 U14967 ( .C1(n15191), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n12722), .B(
        n12721), .ZN(n12737) );
  INV_X1 U14968 ( .A(n12723), .ZN(n12726) );
  INV_X1 U14969 ( .A(n12724), .ZN(n12725) );
  NOR3_X1 U14970 ( .A1(n12727), .A2(n12726), .A3(n12725), .ZN(n12728) );
  OAI21_X1 U14971 ( .B1(n12729), .B2(n12728), .A(n12835), .ZN(n12736) );
  INV_X1 U14972 ( .A(n12730), .ZN(n12731) );
  NOR3_X1 U14973 ( .A1(n12732), .A2(n12731), .A3(n6594), .ZN(n12733) );
  OAI21_X1 U14974 ( .B1(n12734), .B2(n12733), .A(n12864), .ZN(n12735) );
  NAND4_X1 U14975 ( .A1(n12738), .A2(n12737), .A3(n12736), .A4(n12735), .ZN(
        P3_U3190) );
  NAND2_X1 U14976 ( .A1(n12740), .A2(n12739), .ZN(n12742) );
  XOR2_X1 U14977 ( .A(n12771), .B(n12772), .Z(n12741) );
  INV_X1 U14978 ( .A(n12770), .ZN(n12745) );
  AOI21_X1 U14979 ( .B1(n12743), .B2(n12742), .A(n12741), .ZN(n12744) );
  OAI21_X1 U14980 ( .B1(n12745), .B2(n12744), .A(n12890), .ZN(n12762) );
  AOI21_X1 U14981 ( .B1(n6576), .B2(n15428), .A(n6456), .ZN(n12750) );
  NOR2_X1 U14982 ( .A1(n12888), .A2(n12750), .ZN(n12760) );
  INV_X1 U14983 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14740) );
  NOR2_X1 U14984 ( .A1(n12849), .A2(n14740), .ZN(n12759) );
  NAND2_X1 U14985 ( .A1(n12753), .A2(n12752), .ZN(n12754) );
  AOI21_X1 U14986 ( .B1(n12755), .B2(n13208), .A(n12764), .ZN(n12756) );
  NOR2_X1 U14987 ( .A1(n12892), .A2(n12756), .ZN(n12758) );
  NOR4_X1 U14988 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  OAI211_X1 U14989 ( .C1(n12881), .C2(n12771), .A(n12762), .B(n12761), .ZN(
        P3_U3195) );
  XNOR2_X1 U14990 ( .A(n12796), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12794) );
  XNOR2_X1 U14991 ( .A(n12795), .B(n12794), .ZN(n12778) );
  XNOR2_X1 U14992 ( .A(n12796), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12773) );
  AOI21_X1 U14993 ( .B1(n12773), .B2(n12765), .A(n12784), .ZN(n12766) );
  NOR2_X1 U14994 ( .A1(n12892), .A2(n12766), .ZN(n12767) );
  AOI211_X1 U14995 ( .C1(n15191), .C2(P3_ADDR_REG_14__SCAN_IN), .A(n12768), 
        .B(n12767), .ZN(n12769) );
  OAI21_X1 U14996 ( .B1(n12796), .B2(n12881), .A(n12769), .ZN(n12777) );
  NOR2_X1 U14997 ( .A1(n12775), .A2(n12774), .ZN(n12780) );
  AOI211_X1 U14998 ( .C1(n12775), .C2(n12774), .A(n12868), .B(n12780), .ZN(
        n12776) );
  AOI211_X1 U14999 ( .C1(n12778), .C2(n12835), .A(n12777), .B(n12776), .ZN(
        n12779) );
  INV_X1 U15000 ( .A(n12779), .ZN(P3_U3196) );
  AOI21_X1 U15001 ( .B1(n12796), .B2(n12781), .A(n12780), .ZN(n12810) );
  AOI21_X1 U15002 ( .B1(n12783), .B2(n12782), .A(n12808), .ZN(n12804) );
  NAND2_X1 U15003 ( .A1(n12796), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12786) );
  NAND2_X1 U15004 ( .A1(n12786), .A2(n12785), .ZN(n12788) );
  AOI21_X1 U15005 ( .B1(n12789), .B2(n13199), .A(n12805), .ZN(n12790) );
  NOR2_X1 U15006 ( .A1(n12892), .A2(n12790), .ZN(n12793) );
  INV_X1 U15007 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14743) );
  OAI21_X1 U15008 ( .B1(n12849), .B2(n14743), .A(n12791), .ZN(n12792) );
  AOI211_X1 U15009 ( .C1(n12859), .C2(n12809), .A(n12793), .B(n12792), .ZN(
        n12803) );
  NAND2_X1 U15010 ( .A1(n12798), .A2(n12797), .ZN(n12815) );
  OAI21_X1 U15011 ( .B1(n12798), .B2(n12797), .A(n12815), .ZN(n12800) );
  INV_X1 U15012 ( .A(n12800), .ZN(n12799) );
  NOR2_X1 U15013 ( .A1(n12799), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n12801) );
  NOR2_X1 U15014 ( .A1(n13091), .A2(n12800), .ZN(n12816) );
  OAI21_X1 U15015 ( .B1(n12801), .B2(n12816), .A(n12835), .ZN(n12802) );
  OAI211_X1 U15016 ( .C1(n12804), .C2(n12868), .A(n12803), .B(n12802), .ZN(
        P3_U3197) );
  AOI22_X1 U15017 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12830), .B1(n12814), 
        .B2(n13195), .ZN(n12806) );
  AOI21_X1 U15018 ( .B1(n12807), .B2(n12806), .A(n6690), .ZN(n12826) );
  NAND2_X1 U15019 ( .A1(n12811), .A2(n12830), .ZN(n12837) );
  NAND2_X1 U15020 ( .A1(n6586), .A2(n12837), .ZN(n12812) );
  XNOR2_X1 U15021 ( .A(n12838), .B(n12812), .ZN(n12813) );
  NAND2_X1 U15022 ( .A1(n12813), .A2(n12890), .ZN(n12825) );
  AOI22_X1 U15023 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12830), .B1(n12814), 
        .B2(n13078), .ZN(n12819) );
  INV_X1 U15024 ( .A(n12815), .ZN(n12817) );
  AOI21_X1 U15025 ( .B1(n12819), .B2(n12818), .A(n12831), .ZN(n12820) );
  NOR2_X1 U15026 ( .A1(n12888), .A2(n12820), .ZN(n12823) );
  INV_X1 U15027 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14746) );
  OAI21_X1 U15028 ( .B1(n12849), .B2(n14746), .A(n12821), .ZN(n12822) );
  AOI211_X1 U15029 ( .C1(n12859), .C2(n12830), .A(n12823), .B(n12822), .ZN(
        n12824) );
  OAI211_X1 U15030 ( .C1(n12826), .C2(n12892), .A(n12825), .B(n12824), .ZN(
        P3_U3198) );
  NOR2_X1 U15031 ( .A1(n12830), .A2(n13195), .ZN(n12827) );
  INV_X1 U15032 ( .A(n12863), .ZN(n12828) );
  AOI21_X1 U15033 ( .B1(n13191), .B2(n12829), .A(n12828), .ZN(n12843) );
  INV_X1 U15034 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14805) );
  OR2_X1 U15035 ( .A1(n12830), .A2(n13078), .ZN(n12832) );
  NAND2_X1 U15036 ( .A1(n12833), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U15037 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12833), .A(n12854), 
        .ZN(n12834) );
  XOR2_X1 U15038 ( .A(n12845), .B(n12842), .Z(n12840) );
  NOR2_X1 U15039 ( .A1(n12839), .A2(n12840), .ZN(n12844) );
  AOI211_X1 U15040 ( .C1(n12840), .C2(n12839), .A(n12868), .B(n12844), .ZN(
        n12841) );
  AOI21_X1 U15041 ( .B1(n12845), .B2(n7368), .A(n12844), .ZN(n12877) );
  XNOR2_X1 U15042 ( .A(n12877), .B(n12876), .ZN(n12846) );
  NOR2_X1 U15043 ( .A1(n12846), .A2(n12847), .ZN(n12875) );
  AOI21_X1 U15044 ( .B1(n12847), .B2(n12846), .A(n12875), .ZN(n12869) );
  INV_X1 U15045 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14830) );
  OAI21_X1 U15046 ( .B1(n12849), .B2(n14830), .A(n12848), .ZN(n12858) );
  INV_X1 U15047 ( .A(n12850), .ZN(n12853) );
  OR2_X1 U15048 ( .A1(n12876), .A2(n13051), .ZN(n12882) );
  NAND2_X1 U15049 ( .A1(n12876), .A2(n13051), .ZN(n12851) );
  NAND2_X1 U15050 ( .A1(n12882), .A2(n12851), .ZN(n12852) );
  AOI21_X1 U15051 ( .B1(n12854), .B2(n12853), .A(n12852), .ZN(n12883) );
  INV_X1 U15052 ( .A(n12883), .ZN(n12856) );
  NAND3_X1 U15053 ( .A1(n12854), .A2(n12853), .A3(n12852), .ZN(n12855) );
  AOI21_X1 U15054 ( .B1(n12856), .B2(n12855), .A(n12888), .ZN(n12857) );
  AOI211_X1 U15055 ( .C1(n12859), .C2(n12876), .A(n12858), .B(n12857), .ZN(
        n12867) );
  INV_X1 U15056 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13187) );
  OR2_X1 U15057 ( .A1(n12876), .A2(n13187), .ZN(n12870) );
  NAND2_X1 U15058 ( .A1(n12876), .A2(n13187), .ZN(n12860) );
  NAND2_X1 U15059 ( .A1(n12870), .A2(n12860), .ZN(n12861) );
  AND3_X1 U15060 ( .A1(n12863), .A2(n12862), .A3(n12861), .ZN(n12865) );
  OAI21_X1 U15061 ( .B1(n12872), .B2(n12865), .A(n12864), .ZN(n12866) );
  OAI211_X1 U15062 ( .C1(n12869), .C2(n12868), .A(n12867), .B(n12866), .ZN(
        P3_U3200) );
  INV_X1 U15063 ( .A(n12870), .ZN(n12871) );
  NOR2_X1 U15064 ( .A1(n12872), .A2(n12871), .ZN(n12874) );
  XNOR2_X1 U15065 ( .A(n12878), .B(n13183), .ZN(n12879) );
  INV_X1 U15066 ( .A(n12879), .ZN(n12873) );
  XNOR2_X1 U15067 ( .A(n12874), .B(n12873), .ZN(n12893) );
  XNOR2_X1 U15068 ( .A(n12878), .B(n13033), .ZN(n12884) );
  NOR2_X1 U15069 ( .A1(n12881), .A2(n6688), .ZN(n12889) );
  INV_X1 U15070 ( .A(n12884), .ZN(n12885) );
  NAND2_X1 U15071 ( .A1(n15191), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12887) );
  OAI21_X1 U15072 ( .B1(n12893), .B2(n12892), .A(n12891), .ZN(P3_U3201) );
  INV_X1 U15073 ( .A(n13225), .ZN(n12898) );
  OAI21_X1 U15074 ( .B1(n13126), .B2(n15250), .A(n12896), .ZN(n12899) );
  AOI21_X1 U15075 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15250), .A(n12899), 
        .ZN(n12897) );
  OAI21_X1 U15076 ( .B1(n12898), .B2(n15206), .A(n12897), .ZN(P3_U3202) );
  AOI21_X1 U15077 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15250), .A(n12899), 
        .ZN(n12900) );
  OAI21_X1 U15078 ( .B1(n12901), .B2(n15206), .A(n12900), .ZN(P3_U3203) );
  XOR2_X1 U15079 ( .A(n12903), .B(n12902), .Z(n13142) );
  INV_X1 U15080 ( .A(n12904), .ZN(n12906) );
  AOI21_X1 U15081 ( .B1(n12906), .B2(n12905), .A(n14854), .ZN(n12910) );
  OAI22_X1 U15082 ( .A1(n12907), .A2(n14859), .B1(n12934), .B2(n14857), .ZN(
        n12908) );
  AOI21_X1 U15083 ( .B1(n12910), .B2(n12909), .A(n12908), .ZN(n13141) );
  INV_X1 U15084 ( .A(n13141), .ZN(n12915) );
  AOI22_X1 U15085 ( .A1(n15244), .A2(n12911), .B1(n15250), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12912) );
  OAI21_X1 U15086 ( .B1(n12913), .B2(n15206), .A(n12912), .ZN(n12914) );
  AOI21_X1 U15087 ( .B1(n12915), .B2(n15248), .A(n12914), .ZN(n12916) );
  OAI21_X1 U15088 ( .B1(n13142), .B2(n13125), .A(n12916), .ZN(P3_U3205) );
  AOI21_X1 U15089 ( .B1(n12921), .B2(n12917), .A(n12918), .ZN(n12925) );
  OAI22_X1 U15090 ( .A1(n12919), .A2(n14859), .B1(n12948), .B2(n14857), .ZN(
        n12920) );
  INV_X1 U15091 ( .A(n12920), .ZN(n12924) );
  OAI211_X1 U15092 ( .C1(n12925), .C2(n14854), .A(n12924), .B(n12923), .ZN(
        n13144) );
  INV_X1 U15093 ( .A(n13144), .ZN(n12930) );
  AOI22_X1 U15094 ( .A1(n15250), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15244), 
        .B2(n12926), .ZN(n12927) );
  OAI21_X1 U15095 ( .B1(n13238), .B2(n15206), .A(n12927), .ZN(n12928) );
  AOI21_X1 U15096 ( .B1(n13145), .B2(n15246), .A(n12928), .ZN(n12929) );
  OAI21_X1 U15097 ( .B1(n12930), .B2(n15250), .A(n12929), .ZN(P3_U3206) );
  XNOR2_X1 U15098 ( .A(n12932), .B(n12933), .ZN(n12936) );
  OAI22_X1 U15099 ( .A1(n12934), .A2(n14859), .B1(n12964), .B2(n14857), .ZN(
        n12935) );
  AOI21_X1 U15100 ( .B1(n12936), .B2(n15218), .A(n12935), .ZN(n12937) );
  NAND2_X1 U15101 ( .A1(n13149), .A2(n15248), .ZN(n12944) );
  INV_X1 U15102 ( .A(n12938), .ZN(n12939) );
  OAI22_X1 U15103 ( .A1(n15248), .A2(n12940), .B1(n12939), .B2(n15234), .ZN(
        n12941) );
  AOI21_X1 U15104 ( .B1(n12942), .B2(n13107), .A(n12941), .ZN(n12943) );
  OAI211_X1 U15105 ( .C1(n12945), .C2(n13148), .A(n12944), .B(n12943), .ZN(
        P3_U3207) );
  AOI211_X1 U15106 ( .C1(n12952), .C2(n12947), .A(n14854), .B(n12946), .ZN(
        n12950) );
  OAI22_X1 U15107 ( .A1(n12948), .A2(n14859), .B1(n12978), .B2(n14857), .ZN(
        n12949) );
  OR2_X1 U15108 ( .A1(n12950), .A2(n12949), .ZN(n13153) );
  INV_X1 U15109 ( .A(n13153), .ZN(n12959) );
  OAI21_X1 U15110 ( .B1(n12953), .B2(n12952), .A(n12951), .ZN(n13154) );
  INV_X1 U15111 ( .A(n12954), .ZN(n13245) );
  AOI22_X1 U15112 ( .A1(n15250), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15244), 
        .B2(n12955), .ZN(n12956) );
  OAI21_X1 U15113 ( .B1(n13245), .B2(n15206), .A(n12956), .ZN(n12957) );
  AOI21_X1 U15114 ( .B1(n13154), .B2(n14847), .A(n12957), .ZN(n12958) );
  OAI21_X1 U15115 ( .B1(n12959), .B2(n15250), .A(n12958), .ZN(P3_U3208) );
  OAI21_X1 U15116 ( .B1(n6547), .B2(n12961), .A(n12960), .ZN(n12962) );
  INV_X1 U15117 ( .A(n12962), .ZN(n12963) );
  OAI222_X1 U15118 ( .A1(n14857), .A2(n12965), .B1(n14859), .B2(n12964), .C1(
        n14854), .C2(n12963), .ZN(n13157) );
  INV_X1 U15119 ( .A(n13157), .ZN(n12972) );
  OAI21_X1 U15120 ( .B1(n6542), .B2(n8104), .A(n12966), .ZN(n13158) );
  INV_X1 U15121 ( .A(n12967), .ZN(n13249) );
  AOI22_X1 U15122 ( .A1(n15250), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15244), 
        .B2(n12968), .ZN(n12969) );
  OAI21_X1 U15123 ( .B1(n13249), .B2(n15206), .A(n12969), .ZN(n12970) );
  AOI21_X1 U15124 ( .B1(n13158), .B2(n14847), .A(n12970), .ZN(n12971) );
  OAI21_X1 U15125 ( .B1(n12972), .B2(n15250), .A(n12971), .ZN(P3_U3209) );
  XOR2_X1 U15126 ( .A(n12977), .B(n12973), .Z(n13162) );
  INV_X1 U15127 ( .A(n12974), .ZN(n13253) );
  AOI211_X1 U15128 ( .C1(n12977), .C2(n12976), .A(n14854), .B(n12975), .ZN(
        n12980) );
  OAI22_X1 U15129 ( .A1(n12978), .A2(n14859), .B1(n13004), .B2(n14857), .ZN(
        n12979) );
  OR2_X1 U15130 ( .A1(n12980), .A2(n12979), .ZN(n13161) );
  NAND2_X1 U15131 ( .A1(n13161), .A2(n15248), .ZN(n12983) );
  AOI22_X1 U15132 ( .A1(n15250), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15244), 
        .B2(n12981), .ZN(n12982) );
  OAI211_X1 U15133 ( .C1(n13253), .C2(n15206), .A(n12983), .B(n12982), .ZN(
        n12984) );
  AOI21_X1 U15134 ( .B1(n13162), .B2(n14847), .A(n12984), .ZN(n12985) );
  INV_X1 U15135 ( .A(n12985), .ZN(P3_U3210) );
  INV_X1 U15136 ( .A(n12986), .ZN(n12997) );
  XNOR2_X1 U15137 ( .A(n12987), .B(n12997), .ZN(n12991) );
  NAND2_X1 U15138 ( .A1(n12988), .A2(n15215), .ZN(n12989) );
  OAI21_X1 U15139 ( .B1(n13020), .B2(n14857), .A(n12989), .ZN(n12990) );
  AOI21_X1 U15140 ( .B1(n12991), .B2(n15218), .A(n12990), .ZN(n13167) );
  INV_X1 U15141 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12994) );
  INV_X1 U15142 ( .A(n12992), .ZN(n12993) );
  OAI22_X1 U15143 ( .A1(n15248), .A2(n12994), .B1(n12993), .B2(n15234), .ZN(
        n12995) );
  AOI21_X1 U15144 ( .B1(n12996), .B2(n13107), .A(n12995), .ZN(n13000) );
  XNOR2_X1 U15145 ( .A(n12998), .B(n12997), .ZN(n13165) );
  NAND2_X1 U15146 ( .A1(n13165), .A2(n14847), .ZN(n12999) );
  OAI211_X1 U15147 ( .C1(n13167), .C2(n15250), .A(n13000), .B(n12999), .ZN(
        P3_U3211) );
  NAND2_X1 U15148 ( .A1(n13001), .A2(n13011), .ZN(n13002) );
  NAND2_X1 U15149 ( .A1(n13003), .A2(n13002), .ZN(n13006) );
  OAI22_X1 U15150 ( .A1(n13004), .A2(n14859), .B1(n13028), .B2(n14857), .ZN(
        n13005) );
  AOI21_X1 U15151 ( .B1(n13006), .B2(n15218), .A(n13005), .ZN(n13173) );
  INV_X1 U15152 ( .A(n13007), .ZN(n13008) );
  OAI22_X1 U15153 ( .A1(n15248), .A2(n13009), .B1(n13008), .B2(n15234), .ZN(
        n13010) );
  AOI21_X1 U15154 ( .B1(n13170), .B2(n13107), .A(n13010), .ZN(n13014) );
  XNOR2_X1 U15155 ( .A(n13012), .B(n12441), .ZN(n13171) );
  NAND2_X1 U15156 ( .A1(n13171), .A2(n14847), .ZN(n13013) );
  OAI211_X1 U15157 ( .C1(n13173), .C2(n15250), .A(n13014), .B(n13013), .ZN(
        P3_U3212) );
  XNOR2_X1 U15158 ( .A(n13016), .B(n13015), .ZN(n13177) );
  INV_X1 U15159 ( .A(n13177), .ZN(n13025) );
  XNOR2_X1 U15160 ( .A(n13018), .B(n13017), .ZN(n13019) );
  OAI222_X1 U15161 ( .A1(n14859), .A2(n13020), .B1(n14857), .B2(n13049), .C1(
        n13019), .C2(n14854), .ZN(n13176) );
  AOI22_X1 U15162 ( .A1(n15250), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15244), 
        .B2(n13021), .ZN(n13022) );
  OAI21_X1 U15163 ( .B1(n13265), .B2(n15206), .A(n13022), .ZN(n13023) );
  AOI21_X1 U15164 ( .B1(n13176), .B2(n15248), .A(n13023), .ZN(n13024) );
  OAI21_X1 U15165 ( .B1(n13125), .B2(n13025), .A(n13024), .ZN(P3_U3213) );
  AOI21_X1 U15166 ( .B1(n13027), .B2(n13026), .A(n14854), .ZN(n13031) );
  OAI22_X1 U15167 ( .A1(n13059), .A2(n14857), .B1(n13028), .B2(n14859), .ZN(
        n13029) );
  AOI21_X1 U15168 ( .B1(n13031), .B2(n13030), .A(n13029), .ZN(n13182) );
  INV_X1 U15169 ( .A(n13269), .ZN(n13035) );
  OAI22_X1 U15170 ( .A1(n15248), .A2(n13033), .B1(n13032), .B2(n15234), .ZN(
        n13034) );
  AOI21_X1 U15171 ( .B1(n13035), .B2(n13107), .A(n13034), .ZN(n13039) );
  XNOR2_X1 U15172 ( .A(n13037), .B(n13036), .ZN(n13180) );
  NAND2_X1 U15173 ( .A1(n13180), .A2(n14847), .ZN(n13038) );
  OAI211_X1 U15174 ( .C1(n13182), .C2(n15250), .A(n13039), .B(n13038), .ZN(
        P3_U3214) );
  INV_X1 U15175 ( .A(n13040), .ZN(n13043) );
  AOI21_X1 U15176 ( .B1(n13060), .B2(n13041), .A(n13047), .ZN(n13042) );
  NOR2_X1 U15177 ( .A1(n13043), .A2(n13042), .ZN(n13186) );
  INV_X1 U15178 ( .A(n13186), .ZN(n13055) );
  INV_X1 U15179 ( .A(n13045), .ZN(n13046) );
  AOI21_X1 U15180 ( .B1(n13047), .B2(n13044), .A(n13046), .ZN(n13048) );
  OAI222_X1 U15181 ( .A1(n14859), .A2(n13049), .B1(n14857), .B2(n13075), .C1(
        n14854), .C2(n13048), .ZN(n13185) );
  NOR2_X1 U15182 ( .A1(n13273), .A2(n15206), .ZN(n13053) );
  OAI22_X1 U15183 ( .A1(n15248), .A2(n13051), .B1(n13050), .B2(n15234), .ZN(
        n13052) );
  AOI211_X1 U15184 ( .C1(n13185), .C2(n15248), .A(n13053), .B(n13052), .ZN(
        n13054) );
  OAI21_X1 U15185 ( .B1(n13125), .B2(n13055), .A(n13054), .ZN(P3_U3215) );
  XNOR2_X1 U15186 ( .A(n13056), .B(n13057), .ZN(n13058) );
  OAI222_X1 U15187 ( .A1(n14859), .A2(n13059), .B1(n14857), .B2(n13085), .C1(
        n13058), .C2(n14854), .ZN(n13189) );
  INV_X1 U15188 ( .A(n13189), .ZN(n13068) );
  OAI21_X1 U15189 ( .B1(n13062), .B2(n13061), .A(n13060), .ZN(n13190) );
  NOR2_X1 U15190 ( .A1(n15206), .A2(n13277), .ZN(n13066) );
  INV_X1 U15191 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13064) );
  OAI22_X1 U15192 ( .A1(n15248), .A2(n13064), .B1(n13063), .B2(n15234), .ZN(
        n13065) );
  AOI211_X1 U15193 ( .C1(n13190), .C2(n14847), .A(n13066), .B(n13065), .ZN(
        n13067) );
  OAI21_X1 U15194 ( .B1(n13068), .B2(n15250), .A(n13067), .ZN(P3_U3216) );
  XNOR2_X1 U15195 ( .A(n13070), .B(n13069), .ZN(n13194) );
  INV_X1 U15196 ( .A(n13194), .ZN(n13082) );
  XNOR2_X1 U15197 ( .A(n13071), .B(n13072), .ZN(n13073) );
  OAI222_X1 U15198 ( .A1(n14859), .A2(n13075), .B1(n14857), .B2(n13074), .C1(
        n13073), .C2(n14854), .ZN(n13193) );
  INV_X1 U15199 ( .A(n13076), .ZN(n13281) );
  NOR2_X1 U15200 ( .A1(n15206), .A2(n13281), .ZN(n13080) );
  OAI22_X1 U15201 ( .A1(n15248), .A2(n13078), .B1(n13077), .B2(n15234), .ZN(
        n13079) );
  AOI211_X1 U15202 ( .C1(n13193), .C2(n15248), .A(n13080), .B(n13079), .ZN(
        n13081) );
  OAI21_X1 U15203 ( .B1(n13125), .B2(n13082), .A(n13081), .ZN(P3_U3217) );
  XNOR2_X1 U15204 ( .A(n13083), .B(n7198), .ZN(n13084) );
  OAI222_X1 U15205 ( .A1(n14859), .A2(n13085), .B1(n14857), .B2(n13119), .C1(
        n13084), .C2(n14854), .ZN(n13197) );
  INV_X1 U15206 ( .A(n13197), .ZN(n13095) );
  OAI21_X1 U15207 ( .B1(n13088), .B2(n13087), .A(n13086), .ZN(n13198) );
  INV_X1 U15208 ( .A(n13089), .ZN(n13285) );
  NOR2_X1 U15209 ( .A1(n15206), .A2(n13285), .ZN(n13093) );
  OAI22_X1 U15210 ( .A1(n15248), .A2(n13091), .B1(n13090), .B2(n15234), .ZN(
        n13092) );
  AOI211_X1 U15211 ( .C1(n13198), .C2(n14847), .A(n13093), .B(n13092), .ZN(
        n13094) );
  OAI21_X1 U15212 ( .B1(n13095), .B2(n15250), .A(n13094), .ZN(P3_U3218) );
  NAND2_X1 U15213 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NAND3_X1 U15214 ( .A1(n13096), .A2(n15218), .A3(n13099), .ZN(n13102) );
  AOI22_X1 U15215 ( .A1(n15215), .A2(n13100), .B1(n14838), .B2(n15212), .ZN(
        n13101) );
  OAI22_X1 U15216 ( .A1(n15248), .A2(n13104), .B1(n13103), .B2(n15234), .ZN(
        n13105) );
  AOI21_X1 U15217 ( .B1(n13107), .B2(n13106), .A(n13105), .ZN(n13113) );
  NAND2_X1 U15218 ( .A1(n13109), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U15219 ( .A1(n13111), .A2(n13110), .ZN(n13201) );
  NAND2_X1 U15220 ( .A1(n13201), .A2(n14847), .ZN(n13112) );
  OAI211_X1 U15221 ( .C1(n13202), .C2(n15250), .A(n13113), .B(n13112), .ZN(
        P3_U3219) );
  XNOR2_X1 U15222 ( .A(n13115), .B(n13114), .ZN(n13207) );
  INV_X1 U15223 ( .A(n13207), .ZN(n13124) );
  XNOR2_X1 U15224 ( .A(n13117), .B(n13116), .ZN(n13118) );
  OAI222_X1 U15225 ( .A1(n14857), .A2(n14858), .B1(n14859), .B2(n13119), .C1(
        n13118), .C2(n14854), .ZN(n13206) );
  NOR2_X1 U15226 ( .A1(n15206), .A2(n13293), .ZN(n13122) );
  OAI22_X1 U15227 ( .A1(n15248), .A2(n15428), .B1(n13120), .B2(n15234), .ZN(
        n13121) );
  AOI211_X1 U15228 ( .C1(n13206), .C2(n15248), .A(n13122), .B(n13121), .ZN(
        n13123) );
  OAI21_X1 U15229 ( .B1(n13125), .B2(n13124), .A(n13123), .ZN(P3_U3220) );
  INV_X1 U15230 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13128) );
  INV_X1 U15231 ( .A(n13210), .ZN(n13129) );
  NAND2_X1 U15232 ( .A1(n13225), .A2(n13129), .ZN(n13127) );
  INV_X1 U15233 ( .A(n13126), .ZN(n13226) );
  NAND2_X1 U15234 ( .A1(n13226), .A2(n15308), .ZN(n13130) );
  OAI211_X1 U15235 ( .C1(n15308), .C2(n13128), .A(n13127), .B(n13130), .ZN(
        P3_U3490) );
  INV_X1 U15236 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n13132) );
  NAND2_X1 U15237 ( .A1(n13229), .A2(n13129), .ZN(n13131) );
  OAI211_X1 U15238 ( .C1(n15308), .C2(n13132), .A(n13131), .B(n13130), .ZN(
        P3_U3489) );
  AND2_X1 U15239 ( .A1(n15223), .A2(n13143), .ZN(n13152) );
  NAND2_X1 U15240 ( .A1(n13133), .A2(n15287), .ZN(n13134) );
  OAI21_X1 U15241 ( .B1(n13135), .B2(n13152), .A(n13134), .ZN(n13136) );
  INV_X1 U15242 ( .A(n13136), .ZN(n13137) );
  NAND2_X1 U15243 ( .A1(n13138), .A2(n13137), .ZN(n13233) );
  MUX2_X1 U15244 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n13233), .S(n15308), .Z(
        P3_U3488) );
  NAND2_X1 U15245 ( .A1(n13139), .A2(n15287), .ZN(n13140) );
  OAI211_X1 U15246 ( .C1(n13152), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        n13234) );
  MUX2_X1 U15247 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13234), .S(n15308), .Z(
        P3_U3487) );
  INV_X1 U15248 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13146) );
  AOI21_X1 U15249 ( .B1(n15289), .B2(n13145), .A(n13144), .ZN(n13235) );
  MUX2_X1 U15250 ( .A(n13146), .B(n13235), .S(n15308), .Z(n13147) );
  OAI21_X1 U15251 ( .B1(n13238), .B2(n13210), .A(n13147), .ZN(P3_U3486) );
  INV_X1 U15252 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13150) );
  MUX2_X1 U15253 ( .A(n13150), .B(n13239), .S(n15308), .Z(n13151) );
  OAI21_X1 U15254 ( .B1(n13241), .B2(n13210), .A(n13151), .ZN(P3_U3485) );
  INV_X1 U15255 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13155) );
  AOI21_X1 U15256 ( .B1(n14874), .B2(n13154), .A(n13153), .ZN(n13242) );
  MUX2_X1 U15257 ( .A(n13155), .B(n13242), .S(n15308), .Z(n13156) );
  OAI21_X1 U15258 ( .B1(n13245), .B2(n13210), .A(n13156), .ZN(P3_U3484) );
  INV_X1 U15259 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13159) );
  AOI21_X1 U15260 ( .B1(n14874), .B2(n13158), .A(n13157), .ZN(n13246) );
  MUX2_X1 U15261 ( .A(n13159), .B(n13246), .S(n15308), .Z(n13160) );
  OAI21_X1 U15262 ( .B1(n13249), .B2(n13210), .A(n13160), .ZN(P3_U3483) );
  INV_X1 U15263 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13163) );
  AOI21_X1 U15264 ( .B1(n13162), .B2(n14874), .A(n13161), .ZN(n13250) );
  MUX2_X1 U15265 ( .A(n13163), .B(n13250), .S(n15308), .Z(n13164) );
  OAI21_X1 U15266 ( .B1(n13253), .B2(n13210), .A(n13164), .ZN(P3_U3482) );
  INV_X1 U15267 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U15268 ( .A1(n13165), .A2(n14874), .ZN(n13166) );
  AND2_X1 U15269 ( .A1(n13167), .A2(n13166), .ZN(n13254) );
  MUX2_X1 U15270 ( .A(n13168), .B(n13254), .S(n15308), .Z(n13169) );
  OAI21_X1 U15271 ( .B1(n13257), .B2(n13210), .A(n13169), .ZN(P3_U3481) );
  INV_X1 U15272 ( .A(n13170), .ZN(n13261) );
  NAND2_X1 U15273 ( .A1(n13171), .A2(n14874), .ZN(n13172) );
  AND2_X1 U15274 ( .A1(n13173), .A2(n13172), .ZN(n13258) );
  MUX2_X1 U15275 ( .A(n13174), .B(n13258), .S(n15308), .Z(n13175) );
  OAI21_X1 U15276 ( .B1(n13261), .B2(n13210), .A(n13175), .ZN(P3_U3480) );
  AOI21_X1 U15277 ( .B1(n13177), .B2(n14874), .A(n13176), .ZN(n13262) );
  MUX2_X1 U15278 ( .A(n13178), .B(n13262), .S(n15308), .Z(n13179) );
  OAI21_X1 U15279 ( .B1(n13265), .B2(n13210), .A(n13179), .ZN(P3_U3479) );
  NAND2_X1 U15280 ( .A1(n13180), .A2(n14874), .ZN(n13181) );
  AND2_X1 U15281 ( .A1(n13182), .A2(n13181), .ZN(n13266) );
  MUX2_X1 U15282 ( .A(n13183), .B(n13266), .S(n15308), .Z(n13184) );
  OAI21_X1 U15283 ( .B1(n13210), .B2(n13269), .A(n13184), .ZN(P3_U3478) );
  AOI21_X1 U15284 ( .B1(n13186), .B2(n14874), .A(n13185), .ZN(n13270) );
  MUX2_X1 U15285 ( .A(n13187), .B(n13270), .S(n15308), .Z(n13188) );
  OAI21_X1 U15286 ( .B1(n13273), .B2(n13210), .A(n13188), .ZN(P3_U3477) );
  AOI21_X1 U15287 ( .B1(n14874), .B2(n13190), .A(n13189), .ZN(n13274) );
  MUX2_X1 U15288 ( .A(n13191), .B(n13274), .S(n15308), .Z(n13192) );
  OAI21_X1 U15289 ( .B1(n13277), .B2(n13210), .A(n13192), .ZN(P3_U3476) );
  AOI21_X1 U15290 ( .B1(n13194), .B2(n14874), .A(n13193), .ZN(n13278) );
  MUX2_X1 U15291 ( .A(n13195), .B(n13278), .S(n15308), .Z(n13196) );
  OAI21_X1 U15292 ( .B1(n13281), .B2(n13210), .A(n13196), .ZN(P3_U3475) );
  AOI21_X1 U15293 ( .B1(n14874), .B2(n13198), .A(n13197), .ZN(n13282) );
  MUX2_X1 U15294 ( .A(n13199), .B(n13282), .S(n15308), .Z(n13200) );
  OAI21_X1 U15295 ( .B1(n13285), .B2(n13210), .A(n13200), .ZN(P3_U3474) );
  NAND2_X1 U15296 ( .A1(n13201), .A2(n14874), .ZN(n13203) );
  MUX2_X1 U15297 ( .A(n13287), .B(n13204), .S(n15306), .Z(n13205) );
  OAI21_X1 U15298 ( .B1(n13210), .B2(n13289), .A(n13205), .ZN(P3_U3473) );
  AOI21_X1 U15299 ( .B1(n13207), .B2(n14874), .A(n13206), .ZN(n13290) );
  MUX2_X1 U15300 ( .A(n13208), .B(n13290), .S(n15308), .Z(n13209) );
  OAI21_X1 U15301 ( .B1(n13210), .B2(n13293), .A(n13209), .ZN(P3_U3472) );
  OAI21_X1 U15302 ( .B1(n10769), .B2(n13212), .A(n13211), .ZN(n13218) );
  NAND2_X1 U15303 ( .A1(n13213), .A2(n15212), .ZN(n13216) );
  NAND2_X1 U15304 ( .A1(n13214), .A2(n15215), .ZN(n13215) );
  NAND2_X1 U15305 ( .A1(n13216), .A2(n13215), .ZN(n13217) );
  AOI21_X1 U15306 ( .B1(n13218), .B2(n15218), .A(n13217), .ZN(n13221) );
  XNOR2_X1 U15307 ( .A(n10769), .B(n13219), .ZN(n15245) );
  NAND2_X1 U15308 ( .A1(n15245), .A2(n15201), .ZN(n13220) );
  AND2_X1 U15309 ( .A1(n13221), .A2(n13220), .ZN(n15240) );
  NOR2_X1 U15310 ( .A1(n13222), .A2(n15281), .ZN(n15243) );
  AOI21_X1 U15311 ( .B1(n15245), .B2(n15289), .A(n15243), .ZN(n13223) );
  AND2_X1 U15312 ( .A1(n15240), .A2(n13223), .ZN(n15251) );
  INV_X1 U15313 ( .A(n15251), .ZN(n13224) );
  MUX2_X1 U15314 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n13224), .S(n15308), .Z(
        P3_U3460) );
  INV_X1 U15315 ( .A(n13294), .ZN(n13228) );
  NAND2_X1 U15316 ( .A1(n13225), .A2(n13228), .ZN(n13227) );
  NAND2_X1 U15317 ( .A1(n13226), .A2(n15293), .ZN(n13230) );
  OAI211_X1 U15318 ( .C1(n8183), .C2(n15293), .A(n13227), .B(n13230), .ZN(
        P3_U3458) );
  INV_X1 U15319 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U15320 ( .A1(n13229), .A2(n13228), .ZN(n13231) );
  OAI211_X1 U15321 ( .C1(n13232), .C2(n15293), .A(n13231), .B(n13230), .ZN(
        P3_U3457) );
  MUX2_X1 U15322 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n13233), .S(n15293), .Z(
        P3_U3456) );
  MUX2_X1 U15323 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13234), .S(n15293), .Z(
        P3_U3455) );
  INV_X1 U15324 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13236) );
  MUX2_X1 U15325 ( .A(n13236), .B(n13235), .S(n15293), .Z(n13237) );
  OAI21_X1 U15326 ( .B1(n13238), .B2(n13294), .A(n13237), .ZN(P3_U3454) );
  INV_X1 U15327 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13240) );
  INV_X1 U15328 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13243) );
  MUX2_X1 U15329 ( .A(n13243), .B(n13242), .S(n15293), .Z(n13244) );
  OAI21_X1 U15330 ( .B1(n13245), .B2(n13294), .A(n13244), .ZN(P3_U3452) );
  INV_X1 U15331 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13247) );
  MUX2_X1 U15332 ( .A(n13247), .B(n13246), .S(n15293), .Z(n13248) );
  OAI21_X1 U15333 ( .B1(n13249), .B2(n13294), .A(n13248), .ZN(P3_U3451) );
  MUX2_X1 U15334 ( .A(n13251), .B(n13250), .S(n15293), .Z(n13252) );
  OAI21_X1 U15335 ( .B1(n13253), .B2(n13294), .A(n13252), .ZN(P3_U3450) );
  MUX2_X1 U15336 ( .A(n13255), .B(n13254), .S(n15293), .Z(n13256) );
  OAI21_X1 U15337 ( .B1(n13257), .B2(n13294), .A(n13256), .ZN(P3_U3449) );
  MUX2_X1 U15338 ( .A(n13259), .B(n13258), .S(n15293), .Z(n13260) );
  OAI21_X1 U15339 ( .B1(n13261), .B2(n13294), .A(n13260), .ZN(P3_U3448) );
  MUX2_X1 U15340 ( .A(n13263), .B(n13262), .S(n15293), .Z(n13264) );
  OAI21_X1 U15341 ( .B1(n13265), .B2(n13294), .A(n13264), .ZN(P3_U3447) );
  INV_X1 U15342 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13267) );
  MUX2_X1 U15343 ( .A(n13267), .B(n13266), .S(n15293), .Z(n13268) );
  OAI21_X1 U15344 ( .B1(n13294), .B2(n13269), .A(n13268), .ZN(P3_U3446) );
  MUX2_X1 U15345 ( .A(n13271), .B(n13270), .S(n15293), .Z(n13272) );
  OAI21_X1 U15346 ( .B1(n13273), .B2(n13294), .A(n13272), .ZN(P3_U3444) );
  MUX2_X1 U15347 ( .A(n13275), .B(n13274), .S(n15293), .Z(n13276) );
  OAI21_X1 U15348 ( .B1(n13277), .B2(n13294), .A(n13276), .ZN(P3_U3441) );
  INV_X1 U15349 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13279) );
  MUX2_X1 U15350 ( .A(n13279), .B(n13278), .S(n15293), .Z(n13280) );
  OAI21_X1 U15351 ( .B1(n13281), .B2(n13294), .A(n13280), .ZN(P3_U3438) );
  INV_X1 U15352 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13283) );
  MUX2_X1 U15353 ( .A(n13283), .B(n13282), .S(n15293), .Z(n13284) );
  OAI21_X1 U15354 ( .B1(n13285), .B2(n13294), .A(n13284), .ZN(P3_U3435) );
  INV_X1 U15355 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13286) );
  MUX2_X1 U15356 ( .A(n13287), .B(n13286), .S(n15295), .Z(n13288) );
  OAI21_X1 U15357 ( .B1(n13294), .B2(n13289), .A(n13288), .ZN(P3_U3432) );
  INV_X1 U15358 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13291) );
  MUX2_X1 U15359 ( .A(n13291), .B(n13290), .S(n15293), .Z(n13292) );
  OAI21_X1 U15360 ( .B1(n13294), .B2(n13293), .A(n13292), .ZN(P3_U3429) );
  MUX2_X1 U15361 ( .A(P3_D_REG_1__SCAN_IN), .B(n13296), .S(n13295), .Z(
        P3_U3377) );
  INV_X1 U15362 ( .A(n13297), .ZN(n13304) );
  NOR4_X1 U15363 ( .A1(n13299), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13298), .A4(
        P3_U3151), .ZN(n13300) );
  AOI21_X1 U15364 ( .B1(SI_31_), .B2(n13301), .A(n13300), .ZN(n13302) );
  OAI21_X1 U15365 ( .B1(n13304), .B2(n13303), .A(n13302), .ZN(P3_U3264) );
  MUX2_X1 U15366 ( .A(n13305), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15367 ( .A(n13871), .ZN(n13357) );
  XNOR2_X1 U15368 ( .A(n13763), .B(n9828), .ZN(n13326) );
  NAND2_X1 U15369 ( .A1(n13590), .A2(n13343), .ZN(n13327) );
  AOI21_X1 U15370 ( .B1(n13308), .B2(n13307), .A(n13306), .ZN(n13311) );
  INV_X1 U15371 ( .A(n13307), .ZN(n13310) );
  INV_X1 U15372 ( .A(n13308), .ZN(n13309) );
  AND2_X1 U15373 ( .A1(n13578), .A2(n13687), .ZN(n13313) );
  XNOR2_X1 U15374 ( .A(n13607), .B(n9828), .ZN(n13312) );
  NOR2_X1 U15375 ( .A1(n13312), .A2(n13313), .ZN(n13314) );
  AOI21_X1 U15376 ( .B1(n13313), .B2(n13312), .A(n13314), .ZN(n13407) );
  INV_X1 U15377 ( .A(n13314), .ZN(n13315) );
  NAND2_X1 U15378 ( .A1(n13405), .A2(n13315), .ZN(n13417) );
  AND2_X1 U15379 ( .A1(n13581), .A2(n13687), .ZN(n13317) );
  XNOR2_X1 U15380 ( .A(n13930), .B(n9828), .ZN(n13316) );
  NOR2_X1 U15381 ( .A1(n13316), .A2(n13317), .ZN(n13318) );
  AOI21_X1 U15382 ( .B1(n13317), .B2(n13316), .A(n13318), .ZN(n13418) );
  INV_X1 U15383 ( .A(n13318), .ZN(n13319) );
  NAND2_X1 U15384 ( .A1(n13583), .A2(n13343), .ZN(n13321) );
  XNOR2_X1 U15385 ( .A(n13925), .B(n9828), .ZN(n13320) );
  XOR2_X1 U15386 ( .A(n13321), .B(n13320), .Z(n13453) );
  NAND2_X1 U15387 ( .A1(n13475), .A2(n13343), .ZN(n13322) );
  XNOR2_X1 U15388 ( .A(n13915), .B(n9828), .ZN(n13325) );
  AND2_X1 U15389 ( .A1(n13588), .A2(n13687), .ZN(n13324) );
  NOR2_X1 U15390 ( .A1(n13325), .A2(n13324), .ZN(n13435) );
  NAND2_X1 U15391 ( .A1(n13325), .A2(n13324), .ZN(n13436) );
  XNOR2_X1 U15392 ( .A(n13326), .B(n13327), .ZN(n13388) );
  NAND2_X1 U15393 ( .A1(n13389), .A2(n13388), .ZN(n13387) );
  XNOR2_X1 U15394 ( .A(n13753), .B(n9828), .ZN(n13330) );
  INV_X1 U15395 ( .A(n13592), .ZN(n13620) );
  NOR2_X1 U15396 ( .A1(n13620), .A2(n10023), .ZN(n13445) );
  XNOR2_X1 U15397 ( .A(n13964), .B(n9828), .ZN(n13334) );
  NAND2_X1 U15398 ( .A1(n13621), .A2(n13343), .ZN(n13363) );
  INV_X1 U15399 ( .A(n13363), .ZN(n13331) );
  XNOR2_X1 U15400 ( .A(n13888), .B(n13338), .ZN(n13336) );
  NAND2_X1 U15401 ( .A1(n13625), .A2(n13343), .ZN(n13335) );
  NOR2_X1 U15402 ( .A1(n13336), .A2(n13335), .ZN(n13337) );
  AOI21_X1 U15403 ( .B1(n13336), .B2(n13335), .A(n13337), .ZN(n13427) );
  XNOR2_X1 U15404 ( .A(n13705), .B(n13338), .ZN(n13340) );
  NAND2_X1 U15405 ( .A1(n13598), .A2(n13343), .ZN(n13339) );
  NOR2_X1 U15406 ( .A1(n13340), .A2(n13339), .ZN(n13341) );
  AOI21_X1 U15407 ( .B1(n13340), .B2(n13339), .A(n13341), .ZN(n13399) );
  INV_X1 U15408 ( .A(n13341), .ZN(n13342) );
  NAND2_X1 U15409 ( .A1(n13630), .A2(n13343), .ZN(n13345) );
  XNOR2_X1 U15410 ( .A(n13955), .B(n9828), .ZN(n13344) );
  XOR2_X1 U15411 ( .A(n13345), .B(n13344), .Z(n13463) );
  INV_X1 U15412 ( .A(n13344), .ZN(n13346) );
  NAND2_X1 U15413 ( .A1(n13346), .A2(n13345), .ZN(n13347) );
  XNOR2_X1 U15414 ( .A(n13871), .B(n9828), .ZN(n13349) );
  AND2_X1 U15415 ( .A1(n13632), .A2(n13687), .ZN(n13348) );
  NAND2_X1 U15416 ( .A1(n13349), .A2(n13348), .ZN(n13374) );
  OAI21_X1 U15417 ( .B1(n13349), .B2(n13348), .A(n13374), .ZN(n13350) );
  INV_X1 U15418 ( .A(n13673), .ZN(n13354) );
  AOI22_X1 U15419 ( .A1(n13570), .A2(n13635), .B1(n13464), .B2(n13630), .ZN(
        n13667) );
  INV_X1 U15420 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13352) );
  OAI22_X1 U15421 ( .A1(n13447), .A2(n13667), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13352), .ZN(n13353) );
  AOI21_X1 U15422 ( .B1(n13354), .B2(n13449), .A(n13353), .ZN(n13355) );
  OAI211_X1 U15423 ( .C1(n13357), .C2(n13452), .A(n13356), .B(n13355), .ZN(
        P2_U3186) );
  NAND2_X1 U15424 ( .A1(n13570), .A2(n13625), .ZN(n13359) );
  NAND2_X1 U15425 ( .A1(n13464), .A2(n13592), .ZN(n13358) );
  NAND2_X1 U15426 ( .A1(n13359), .A2(n13358), .ZN(n13741) );
  AOI22_X1 U15427 ( .A1(n14885), .A2(n13741), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13360) );
  OAI21_X1 U15428 ( .B1(n13733), .B2(n14891), .A(n13360), .ZN(n13366) );
  INV_X1 U15429 ( .A(n13361), .ZN(n13362) );
  AOI211_X1 U15430 ( .C1(n13364), .C2(n13363), .A(n13470), .B(n13362), .ZN(
        n13365) );
  AOI211_X1 U15431 ( .C1(n13964), .C2(n9631), .A(n13366), .B(n13365), .ZN(
        n13367) );
  INV_X1 U15432 ( .A(n13367), .ZN(P2_U3188) );
  AOI21_X1 U15433 ( .B1(n13369), .B2(n13368), .A(n6566), .ZN(n13373) );
  AOI22_X1 U15434 ( .A1(n13588), .A2(n13570), .B1(n13464), .B2(n13583), .ZN(
        n13794) );
  NAND2_X1 U15435 ( .A1(n13449), .A2(n13800), .ZN(n13370) );
  NAND2_X1 U15436 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13563)
         );
  OAI211_X1 U15437 ( .C1(n13794), .C2(n13447), .A(n13370), .B(n13563), .ZN(
        n13371) );
  AOI21_X1 U15438 ( .B1(n13920), .B2(n9631), .A(n13371), .ZN(n13372) );
  OAI21_X1 U15439 ( .B1(n13373), .B2(n13470), .A(n13372), .ZN(P2_U3191) );
  NAND2_X1 U15440 ( .A1(n13635), .A2(n13343), .ZN(n13376) );
  XNOR2_X1 U15441 ( .A(n9828), .B(n13376), .ZN(n13377) );
  XNOR2_X1 U15442 ( .A(n13660), .B(n13377), .ZN(n13378) );
  XNOR2_X1 U15443 ( .A(n13379), .B(n13378), .ZN(n13386) );
  INV_X1 U15444 ( .A(n13653), .ZN(n13383) );
  NAND2_X1 U15445 ( .A1(n13570), .A2(n13474), .ZN(n13381) );
  NAND2_X1 U15446 ( .A1(n13464), .A2(n13632), .ZN(n13380) );
  NAND2_X1 U15447 ( .A1(n13381), .A2(n13380), .ZN(n13650) );
  AOI22_X1 U15448 ( .A1(n14885), .A2(n13650), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13382) );
  OAI21_X1 U15449 ( .B1(n13383), .B2(n14891), .A(n13382), .ZN(n13384) );
  AOI21_X1 U15450 ( .B1(n13660), .B2(n9631), .A(n13384), .ZN(n13385) );
  OAI21_X1 U15451 ( .B1(n13386), .B2(n13470), .A(n13385), .ZN(P2_U3192) );
  OAI211_X1 U15452 ( .C1(n13389), .C2(n13388), .A(n13387), .B(n14883), .ZN(
        n13396) );
  NAND2_X1 U15453 ( .A1(n13588), .A2(n13464), .ZN(n13391) );
  NAND2_X1 U15454 ( .A1(n13570), .A2(n13592), .ZN(n13390) );
  NAND2_X1 U15455 ( .A1(n13391), .A2(n13390), .ZN(n13770) );
  INV_X1 U15456 ( .A(n13770), .ZN(n13393) );
  INV_X1 U15457 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13392) );
  OAI22_X1 U15458 ( .A1(n13393), .A2(n13447), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13392), .ZN(n13394) );
  AOI21_X1 U15459 ( .B1(n13762), .B2(n13449), .A(n13394), .ZN(n13395) );
  OAI211_X1 U15460 ( .C1(n13975), .C2(n13452), .A(n13396), .B(n13395), .ZN(
        P2_U3195) );
  OAI211_X1 U15461 ( .C1(n13397), .C2(n13399), .A(n13398), .B(n14883), .ZN(
        n13404) );
  INV_X1 U15462 ( .A(n13400), .ZN(n13706) );
  AOI22_X1 U15463 ( .A1(n13464), .A2(n13625), .B1(n13570), .B2(n13630), .ZN(
        n13698) );
  INV_X1 U15464 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13401) );
  OAI22_X1 U15465 ( .A1(n13447), .A2(n13698), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13401), .ZN(n13402) );
  AOI21_X1 U15466 ( .B1(n13706), .B2(n13449), .A(n13402), .ZN(n13403) );
  OAI211_X1 U15467 ( .C1(n13960), .C2(n13452), .A(n13404), .B(n13403), .ZN(
        P2_U3197) );
  OAI21_X1 U15468 ( .B1(n13407), .B2(n13406), .A(n13405), .ZN(n13408) );
  NAND2_X1 U15469 ( .A1(n13408), .A2(n14883), .ZN(n13414) );
  OAI21_X1 U15470 ( .B1(n13447), .B2(n13410), .A(n13409), .ZN(n13411) );
  AOI21_X1 U15471 ( .B1(n13412), .B2(n13449), .A(n13411), .ZN(n13413) );
  OAI211_X1 U15472 ( .C1(n13415), .C2(n13452), .A(n13414), .B(n13413), .ZN(
        P2_U3198) );
  INV_X1 U15473 ( .A(n13930), .ZN(n13425) );
  OAI21_X1 U15474 ( .B1(n13418), .B2(n13417), .A(n13416), .ZN(n13419) );
  NAND2_X1 U15475 ( .A1(n13419), .A2(n14883), .ZN(n13424) );
  OAI22_X1 U15476 ( .A1(n13611), .A2(n13455), .B1(n13606), .B2(n13640), .ZN(
        n13821) );
  INV_X1 U15477 ( .A(n13821), .ZN(n13421) );
  OAI21_X1 U15478 ( .B1(n13447), .B2(n13421), .A(n13420), .ZN(n13422) );
  AOI21_X1 U15479 ( .B1(n13827), .B2(n13449), .A(n13422), .ZN(n13423) );
  OAI211_X1 U15480 ( .C1(n13425), .C2(n13452), .A(n13424), .B(n13423), .ZN(
        P2_U3200) );
  INV_X1 U15481 ( .A(n13888), .ZN(n13723) );
  OAI211_X1 U15482 ( .C1(n13428), .C2(n13427), .A(n13426), .B(n14883), .ZN(
        n13434) );
  NAND2_X1 U15483 ( .A1(n13464), .A2(n13621), .ZN(n13430) );
  NAND2_X1 U15484 ( .A1(n13570), .A2(n13598), .ZN(n13429) );
  AND2_X1 U15485 ( .A1(n13430), .A2(n13429), .ZN(n13716) );
  OAI22_X1 U15486 ( .A1(n13447), .A2(n13716), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13431), .ZN(n13432) );
  AOI21_X1 U15487 ( .B1(n13721), .B2(n13449), .A(n13432), .ZN(n13433) );
  OAI211_X1 U15488 ( .C1(n13723), .C2(n13452), .A(n13434), .B(n13433), .ZN(
        P2_U3201) );
  NAND2_X1 U15489 ( .A1(n7323), .A2(n13436), .ZN(n13437) );
  XNOR2_X1 U15490 ( .A(n13438), .B(n13437), .ZN(n13443) );
  AOI22_X1 U15491 ( .A1(n13590), .A2(n13570), .B1(n13464), .B2(n13475), .ZN(
        n13779) );
  INV_X1 U15492 ( .A(n13779), .ZN(n13439) );
  AOI22_X1 U15493 ( .A1(n13439), .A2(n14885), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13440) );
  OAI21_X1 U15494 ( .B1(n13784), .B2(n14891), .A(n13440), .ZN(n13441) );
  AOI21_X1 U15495 ( .B1(n13915), .B2(n9631), .A(n13441), .ZN(n13442) );
  OAI21_X1 U15496 ( .B1(n13443), .B2(n13470), .A(n13442), .ZN(P2_U3205) );
  OAI211_X1 U15497 ( .C1(n13446), .C2(n13445), .A(n13444), .B(n14883), .ZN(
        n13451) );
  AOI22_X1 U15498 ( .A1(n13590), .A2(n13464), .B1(n13570), .B2(n13621), .ZN(
        n13746) );
  OAI22_X1 U15499 ( .A1(n13746), .A2(n13447), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15379), .ZN(n13448) );
  AOI21_X1 U15500 ( .B1(n13754), .B2(n13449), .A(n13448), .ZN(n13450) );
  OAI211_X1 U15501 ( .C1(n13970), .C2(n13452), .A(n13451), .B(n13450), .ZN(
        P2_U3207) );
  XNOR2_X1 U15502 ( .A(n13454), .B(n13453), .ZN(n13459) );
  INV_X1 U15503 ( .A(n13475), .ZN(n13614) );
  OAI22_X1 U15504 ( .A1(n13614), .A2(n13455), .B1(n13610), .B2(n13640), .ZN(
        n13806) );
  AOI22_X1 U15505 ( .A1(n13806), .A2(n14885), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13456) );
  OAI21_X1 U15506 ( .B1(n13812), .B2(n14891), .A(n13456), .ZN(n13457) );
  AOI21_X1 U15507 ( .B1(n13925), .B2(n9631), .A(n13457), .ZN(n13458) );
  OAI21_X1 U15508 ( .B1(n13459), .B2(n13470), .A(n13458), .ZN(P2_U3210) );
  INV_X1 U15509 ( .A(n13460), .ZN(n13461) );
  AOI21_X1 U15510 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n13471) );
  NAND2_X1 U15511 ( .A1(n13464), .A2(n13598), .ZN(n13466) );
  NAND2_X1 U15512 ( .A1(n13570), .A2(n13632), .ZN(n13465) );
  NAND2_X1 U15513 ( .A1(n13466), .A2(n13465), .ZN(n13683) );
  AOI22_X1 U15514 ( .A1(n14885), .A2(n13683), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13467) );
  OAI21_X1 U15515 ( .B1(n13690), .B2(n14891), .A(n13467), .ZN(n13468) );
  AOI21_X1 U15516 ( .B1(n13955), .B2(n9631), .A(n13468), .ZN(n13469) );
  OAI21_X1 U15517 ( .B1(n13471), .B2(n13470), .A(n13469), .ZN(P2_U3212) );
  MUX2_X1 U15518 ( .A(n13472), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13490), .Z(
        P2_U3562) );
  MUX2_X1 U15519 ( .A(n13473), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13490), .Z(
        P2_U3561) );
  MUX2_X1 U15520 ( .A(n13474), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13490), .Z(
        P2_U3560) );
  MUX2_X1 U15521 ( .A(n13635), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13490), .Z(
        P2_U3559) );
  MUX2_X1 U15522 ( .A(n13632), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13490), .Z(
        P2_U3558) );
  MUX2_X1 U15523 ( .A(n13630), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13490), .Z(
        P2_U3557) );
  MUX2_X1 U15524 ( .A(n13598), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13490), .Z(
        P2_U3556) );
  MUX2_X1 U15525 ( .A(n13625), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13490), .Z(
        P2_U3555) );
  MUX2_X1 U15526 ( .A(n13621), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13490), .Z(
        P2_U3554) );
  MUX2_X1 U15527 ( .A(n13592), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13490), .Z(
        P2_U3553) );
  MUX2_X1 U15528 ( .A(n13590), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13490), .Z(
        P2_U3552) );
  MUX2_X1 U15529 ( .A(n13588), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13490), .Z(
        P2_U3551) );
  MUX2_X1 U15530 ( .A(n13475), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13490), .Z(
        P2_U3550) );
  MUX2_X1 U15531 ( .A(n13583), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13490), .Z(
        P2_U3549) );
  MUX2_X1 U15532 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13581), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15533 ( .A(n13578), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13490), .Z(
        P2_U3547) );
  MUX2_X1 U15534 ( .A(n13476), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13490), .Z(
        P2_U3546) );
  MUX2_X1 U15535 ( .A(n13477), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13490), .Z(
        P2_U3545) );
  MUX2_X1 U15536 ( .A(n13478), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13490), .Z(
        P2_U3544) );
  MUX2_X1 U15537 ( .A(n13479), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13490), .Z(
        P2_U3543) );
  MUX2_X1 U15538 ( .A(n13480), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13490), .Z(
        P2_U3542) );
  MUX2_X1 U15539 ( .A(n13481), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13490), .Z(
        P2_U3541) );
  MUX2_X1 U15540 ( .A(n13482), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13490), .Z(
        P2_U3540) );
  MUX2_X1 U15541 ( .A(n13483), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13490), .Z(
        P2_U3539) );
  MUX2_X1 U15542 ( .A(n13484), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13490), .Z(
        P2_U3538) );
  MUX2_X1 U15543 ( .A(n13485), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13490), .Z(
        P2_U3537) );
  MUX2_X1 U15544 ( .A(n13486), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13490), .Z(
        P2_U3536) );
  MUX2_X1 U15545 ( .A(n13487), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13490), .Z(
        P2_U3535) );
  MUX2_X1 U15546 ( .A(n13488), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13490), .Z(
        P2_U3534) );
  MUX2_X1 U15547 ( .A(n9210), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13490), .Z(
        P2_U3533) );
  MUX2_X1 U15548 ( .A(n13489), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13490), .Z(
        P2_U3532) );
  MUX2_X1 U15549 ( .A(n13491), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13490), .Z(
        P2_U3531) );
  OAI22_X1 U15550 ( .A1(n15143), .A2(n13496), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13492), .ZN(n13493) );
  AOI21_X1 U15551 ( .B1(n15154), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n13493), .ZN(
        n13502) );
  OAI211_X1 U15552 ( .C1(n13495), .C2(n13494), .A(n15161), .B(n13507), .ZN(
        n13501) );
  MUX2_X1 U15553 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9398), .S(n13496), .Z(
        n13497) );
  INV_X1 U15554 ( .A(n13497), .ZN(n13499) );
  OAI211_X1 U15555 ( .C1(n13499), .C2(n13498), .A(n15158), .B(n13514), .ZN(
        n13500) );
  NAND3_X1 U15556 ( .A1(n13502), .A2(n13501), .A3(n13500), .ZN(P2_U3216) );
  OAI21_X1 U15557 ( .B1(n15143), .B2(n6886), .A(n13503), .ZN(n13504) );
  AOI21_X1 U15558 ( .B1(n15154), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13504), .ZN(
        n13519) );
  MUX2_X1 U15559 ( .A(n8537), .B(P2_REG1_REG_3__SCAN_IN), .S(n13505), .Z(
        n13508) );
  NAND3_X1 U15560 ( .A1(n13508), .A2(n13507), .A3(n13506), .ZN(n13509) );
  NAND3_X1 U15561 ( .A1(n15161), .A2(n13510), .A3(n13509), .ZN(n13518) );
  INV_X1 U15562 ( .A(n13511), .ZN(n13516) );
  NAND3_X1 U15563 ( .A1(n13514), .A2(n13513), .A3(n13512), .ZN(n13515) );
  NAND3_X1 U15564 ( .A1(n15158), .A2(n13516), .A3(n13515), .ZN(n13517) );
  NAND3_X1 U15565 ( .A1(n13519), .A2(n13518), .A3(n13517), .ZN(P2_U3217) );
  NAND2_X1 U15566 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14888)
         );
  OAI211_X1 U15567 ( .C1(n13522), .C2(n13521), .A(n15161), .B(n13520), .ZN(
        n13523) );
  AND2_X1 U15568 ( .A1(n14888), .A2(n13523), .ZN(n13529) );
  AOI22_X1 U15569 ( .A1(n15154), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n15155), 
        .B2(n13524), .ZN(n13528) );
  OAI211_X1 U15570 ( .C1(n13526), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15158), 
        .B(n13525), .ZN(n13527) );
  NAND3_X1 U15571 ( .A1(n13529), .A2(n13528), .A3(n13527), .ZN(P2_U3228) );
  NAND2_X1 U15572 ( .A1(n13530), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13531) );
  AOI21_X1 U15573 ( .B1(n13534), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13547), 
        .ZN(n13545) );
  INV_X1 U15574 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13536) );
  OAI21_X1 U15575 ( .B1(n13537), .B2(n13536), .A(n13535), .ZN(n13551) );
  XNOR2_X1 U15576 ( .A(n13551), .B(n13538), .ZN(n13549) );
  XNOR2_X1 U15577 ( .A(n13549), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n13542) );
  NOR2_X1 U15578 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15444), .ZN(n13539) );
  AOI21_X1 U15579 ( .B1(n15154), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13539), 
        .ZN(n13541) );
  NAND2_X1 U15580 ( .A1(n15155), .A2(n13550), .ZN(n13540) );
  OAI211_X1 U15581 ( .C1(n13542), .C2(n13556), .A(n13541), .B(n13540), .ZN(
        n13543) );
  INV_X1 U15582 ( .A(n13543), .ZN(n13544) );
  OAI21_X1 U15583 ( .B1(n13545), .B2(n15129), .A(n13544), .ZN(P2_U3232) );
  XOR2_X1 U15584 ( .A(n13548), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13560) );
  INV_X1 U15585 ( .A(n13560), .ZN(n13558) );
  NAND2_X1 U15586 ( .A1(n13549), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U15587 ( .A1(n13551), .A2(n13550), .ZN(n13552) );
  NAND2_X1 U15588 ( .A1(n13553), .A2(n13552), .ZN(n13555) );
  INV_X1 U15589 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13554) );
  XNOR2_X1 U15590 ( .A(n13555), .B(n13554), .ZN(n13559) );
  NOR2_X1 U15591 ( .A1(n13559), .A2(n13556), .ZN(n13557) );
  AOI211_X1 U15592 ( .C1(n13558), .C2(n15158), .A(n15155), .B(n13557), .ZN(
        n13562) );
  AOI22_X1 U15593 ( .A1(n13560), .A2(n15158), .B1(n15161), .B2(n13559), .ZN(
        n13561) );
  MUX2_X1 U15594 ( .A(n13562), .B(n13561), .S(n9628), .Z(n13564) );
  OAI211_X1 U15595 ( .C1(n7695), .C2(n15127), .A(n13564), .B(n13563), .ZN(
        P2_U3233) );
  NOR2_X1 U15596 ( .A1(n13731), .A2(n13888), .ZN(n13720) );
  NAND2_X1 U15597 ( .A1(n13720), .A2(n13960), .ZN(n13702) );
  NOR2_X2 U15598 ( .A1(n13702), .A2(n13955), .ZN(n13670) );
  OR2_X1 U15599 ( .A1(n13996), .A2(n13568), .ZN(n13569) );
  NAND2_X1 U15600 ( .A1(n13570), .A2(n13569), .ZN(n13639) );
  OR2_X1 U15601 ( .A1(n13639), .A2(n13571), .ZN(n13858) );
  NOR2_X1 U15602 ( .A1(n6430), .A2(n13858), .ZN(n13576) );
  INV_X1 U15603 ( .A(n9171), .ZN(n13942) );
  NOR2_X1 U15604 ( .A1(n13942), .A2(n13816), .ZN(n13572) );
  AOI211_X1 U15605 ( .C1(n6430), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13576), .B(
        n13572), .ZN(n13573) );
  OAI21_X1 U15606 ( .B1(n13856), .B2(n13766), .A(n13573), .ZN(P2_U3234) );
  OAI211_X1 U15607 ( .C1(n13946), .C2(n13641), .A(n10023), .B(n13574), .ZN(
        n13859) );
  NOR2_X1 U15608 ( .A1(n13946), .A2(n13816), .ZN(n13575) );
  AOI211_X1 U15609 ( .C1(n6430), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13576), .B(
        n13575), .ZN(n13577) );
  OAI21_X1 U15610 ( .B1(n13766), .B2(n13859), .A(n13577), .ZN(P2_U3235) );
  NAND2_X1 U15611 ( .A1(n13607), .A2(n13578), .ZN(n13579) );
  NAND2_X1 U15612 ( .A1(n13930), .A2(n13581), .ZN(n13582) );
  OR2_X1 U15613 ( .A1(n13925), .A2(n13583), .ZN(n13584) );
  NAND2_X1 U15614 ( .A1(n13915), .A2(n13588), .ZN(n13587) );
  OR2_X1 U15615 ( .A1(n13915), .A2(n13588), .ZN(n13589) );
  OR2_X1 U15616 ( .A1(n13763), .A2(n13590), .ZN(n13591) );
  NAND2_X1 U15617 ( .A1(n13753), .A2(n13592), .ZN(n13593) );
  INV_X1 U15618 ( .A(n13712), .ZN(n13714) );
  NAND2_X1 U15619 ( .A1(n13713), .A2(n13714), .ZN(n13597) );
  NAND2_X1 U15620 ( .A1(n13888), .A2(n13625), .ZN(n13596) );
  INV_X1 U15621 ( .A(n13701), .ZN(n13628) );
  OR2_X1 U15622 ( .A1(n13705), .A2(n13598), .ZN(n13599) );
  NAND2_X1 U15623 ( .A1(n13955), .A2(n13630), .ZN(n13600) );
  OR2_X1 U15624 ( .A1(n13955), .A2(n13630), .ZN(n13601) );
  INV_X1 U15625 ( .A(n13647), .ZN(n13654) );
  NAND2_X1 U15626 ( .A1(n13655), .A2(n13654), .ZN(n13657) );
  NAND2_X1 U15627 ( .A1(n13657), .A2(n13602), .ZN(n13603) );
  INV_X1 U15628 ( .A(n13660), .ZN(n13951) );
  OR2_X1 U15629 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  NOR2_X1 U15630 ( .A1(n13930), .A2(n13610), .ZN(n13609) );
  AND2_X1 U15631 ( .A1(n13925), .A2(n13611), .ZN(n13612) );
  OAI22_X1 U15632 ( .A1(n13805), .A2(n13612), .B1(n13611), .B2(n13925), .ZN(
        n13792) );
  NOR2_X1 U15633 ( .A1(n13920), .A2(n13614), .ZN(n13613) );
  NAND2_X1 U15634 ( .A1(n13920), .A2(n13614), .ZN(n13615) );
  INV_X1 U15635 ( .A(n13777), .ZN(n13775) );
  NAND2_X1 U15636 ( .A1(n13915), .A2(n13616), .ZN(n13617) );
  AND2_X1 U15637 ( .A1(n13763), .A2(n13618), .ZN(n13619) );
  INV_X1 U15638 ( .A(n13621), .ZN(n13623) );
  NOR2_X1 U15639 ( .A1(n13964), .A2(n13623), .ZN(n13622) );
  NAND2_X1 U15640 ( .A1(n13964), .A2(n13623), .ZN(n13624) );
  INV_X1 U15641 ( .A(n13625), .ZN(n13626) );
  NAND2_X1 U15642 ( .A1(n13888), .A2(n13626), .ZN(n13627) );
  INV_X1 U15643 ( .A(n13630), .ZN(n13631) );
  INV_X1 U15644 ( .A(n13632), .ZN(n13633) );
  AND2_X1 U15645 ( .A1(n13871), .A2(n13633), .ZN(n13634) );
  NAND2_X1 U15646 ( .A1(n13862), .A2(n13844), .ZN(n13646) );
  AOI211_X1 U15647 ( .C1(n13864), .C2(n13658), .A(n13687), .B(n13641), .ZN(
        n13863) );
  AOI22_X1 U15648 ( .A1(n6430), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13642), 
        .B2(n13828), .ZN(n13643) );
  OAI21_X1 U15649 ( .B1(n7123), .B2(n13816), .A(n13643), .ZN(n13644) );
  AOI21_X1 U15650 ( .B1(n13863), .B2(n13850), .A(n13644), .ZN(n13645) );
  OAI211_X1 U15651 ( .C1(n13865), .C2(n13835), .A(n13646), .B(n13645), .ZN(
        P2_U3236) );
  INV_X1 U15652 ( .A(n13650), .ZN(n13651) );
  INV_X1 U15653 ( .A(n13867), .ZN(n13652) );
  AOI21_X1 U15654 ( .B1(n13653), .B2(n13828), .A(n13652), .ZN(n13665) );
  OR2_X1 U15655 ( .A1(n13655), .A2(n13654), .ZN(n13656) );
  NAND2_X1 U15656 ( .A1(n13657), .A2(n13656), .ZN(n13868) );
  INV_X1 U15657 ( .A(n13868), .ZN(n13663) );
  AOI21_X1 U15658 ( .B1(n13660), .B2(n13671), .A(n13687), .ZN(n13659) );
  NAND2_X1 U15659 ( .A1(n13659), .A2(n13658), .ZN(n13866) );
  AOI22_X1 U15660 ( .A1(n13660), .A2(n13846), .B1(n6430), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13661) );
  OAI21_X1 U15661 ( .B1(n13866), .B2(n13766), .A(n13661), .ZN(n13662) );
  AOI21_X1 U15662 ( .B1(n13663), .B2(n13848), .A(n13662), .ZN(n13664) );
  OAI21_X1 U15663 ( .B1(n13665), .B2(n6430), .A(n13664), .ZN(P2_U3237) );
  XNOR2_X1 U15664 ( .A(n13666), .B(n13678), .ZN(n13669) );
  INV_X1 U15665 ( .A(n13667), .ZN(n13668) );
  AOI21_X1 U15666 ( .B1(n13669), .B2(n13822), .A(n13668), .ZN(n13877) );
  INV_X1 U15667 ( .A(n13670), .ZN(n13688) );
  AOI21_X1 U15668 ( .B1(n13871), .B2(n13688), .A(n13687), .ZN(n13672) );
  NAND2_X1 U15669 ( .A1(n13672), .A2(n13671), .ZN(n13874) );
  INV_X1 U15670 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13674) );
  OAI22_X1 U15671 ( .A1(n13844), .A2(n13674), .B1(n13673), .B2(n13841), .ZN(
        n13675) );
  AOI21_X1 U15672 ( .B1(n13871), .B2(n13846), .A(n13675), .ZN(n13676) );
  OAI21_X1 U15673 ( .B1(n13874), .B2(n13766), .A(n13676), .ZN(n13677) );
  INV_X1 U15674 ( .A(n13677), .ZN(n13681) );
  NAND2_X1 U15675 ( .A1(n13679), .A2(n13678), .ZN(n13872) );
  NAND3_X1 U15676 ( .A1(n13873), .A2(n13848), .A3(n13872), .ZN(n13680) );
  OAI211_X1 U15677 ( .C1(n13877), .C2(n6430), .A(n13681), .B(n13680), .ZN(
        P2_U3238) );
  XNOR2_X1 U15678 ( .A(n13682), .B(n13685), .ZN(n13684) );
  AOI21_X1 U15679 ( .B1(n13684), .B2(n13822), .A(n13683), .ZN(n13879) );
  XNOR2_X1 U15680 ( .A(n13686), .B(n13685), .ZN(n13880) );
  INV_X1 U15681 ( .A(n13880), .ZN(n13695) );
  AOI21_X1 U15682 ( .B1(n13702), .B2(n13955), .A(n13687), .ZN(n13689) );
  NAND2_X1 U15683 ( .A1(n13689), .A2(n13688), .ZN(n13878) );
  INV_X1 U15684 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13691) );
  OAI22_X1 U15685 ( .A1(n13844), .A2(n13691), .B1(n13690), .B2(n13841), .ZN(
        n13692) );
  AOI21_X1 U15686 ( .B1(n13955), .B2(n13846), .A(n13692), .ZN(n13693) );
  OAI21_X1 U15687 ( .B1(n13878), .B2(n13766), .A(n13693), .ZN(n13694) );
  AOI21_X1 U15688 ( .B1(n13695), .B2(n13848), .A(n13694), .ZN(n13696) );
  OAI21_X1 U15689 ( .B1(n6430), .B2(n13879), .A(n13696), .ZN(P2_U3239) );
  XNOR2_X1 U15690 ( .A(n13697), .B(n13701), .ZN(n13699) );
  OAI21_X1 U15691 ( .B1(n13699), .B2(n13795), .A(n13698), .ZN(n13883) );
  INV_X1 U15692 ( .A(n13883), .ZN(n13711) );
  OAI21_X1 U15693 ( .B1(n6485), .B2(n13701), .A(n13700), .ZN(n13885) );
  INV_X1 U15694 ( .A(n13720), .ZN(n13704) );
  INV_X1 U15695 ( .A(n13702), .ZN(n13703) );
  AOI211_X1 U15696 ( .C1(n13705), .C2(n13704), .A(n13687), .B(n13703), .ZN(
        n13884) );
  NAND2_X1 U15697 ( .A1(n13884), .A2(n13850), .ZN(n13708) );
  AOI22_X1 U15698 ( .A1(n6430), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13706), 
        .B2(n13828), .ZN(n13707) );
  OAI211_X1 U15699 ( .C1(n13960), .C2(n13816), .A(n13708), .B(n13707), .ZN(
        n13709) );
  AOI21_X1 U15700 ( .B1(n13848), .B2(n13885), .A(n13709), .ZN(n13710) );
  OAI21_X1 U15701 ( .B1(n6430), .B2(n13711), .A(n13710), .ZN(P2_U3240) );
  INV_X1 U15702 ( .A(n9664), .ZN(n13719) );
  XNOR2_X1 U15703 ( .A(n13713), .B(n13712), .ZN(n13724) );
  XNOR2_X1 U15704 ( .A(n13715), .B(n13714), .ZN(n13717) );
  OAI21_X1 U15705 ( .B1(n13717), .B2(n13795), .A(n13716), .ZN(n13718) );
  AOI21_X1 U15706 ( .B1(n13719), .B2(n13724), .A(n13718), .ZN(n13890) );
  AOI211_X1 U15707 ( .C1(n13888), .C2(n13731), .A(n13343), .B(n13720), .ZN(
        n13887) );
  AOI22_X1 U15708 ( .A1(n6430), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13721), 
        .B2(n13828), .ZN(n13722) );
  OAI21_X1 U15709 ( .B1(n13723), .B2(n13816), .A(n13722), .ZN(n13727) );
  INV_X1 U15710 ( .A(n13724), .ZN(n13892) );
  NOR2_X1 U15711 ( .A1(n13892), .A2(n13725), .ZN(n13726) );
  AOI211_X1 U15712 ( .C1(n13887), .C2(n13850), .A(n13727), .B(n13726), .ZN(
        n13728) );
  OAI21_X1 U15713 ( .B1(n6430), .B2(n13890), .A(n13728), .ZN(P2_U3241) );
  XNOR2_X1 U15714 ( .A(n13729), .B(n13737), .ZN(n13893) );
  AOI21_X1 U15715 ( .B1(n13964), .B2(n13752), .A(n13687), .ZN(n13732) );
  NAND2_X1 U15716 ( .A1(n13732), .A2(n13731), .ZN(n13894) );
  INV_X1 U15717 ( .A(n13733), .ZN(n13734) );
  AOI22_X1 U15718 ( .A1(n6430), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13734), 
        .B2(n13828), .ZN(n13736) );
  NAND2_X1 U15719 ( .A1(n13964), .A2(n13846), .ZN(n13735) );
  OAI211_X1 U15720 ( .C1(n13894), .C2(n13766), .A(n13736), .B(n13735), .ZN(
        n13743) );
  INV_X1 U15721 ( .A(n13737), .ZN(n13738) );
  XNOR2_X1 U15722 ( .A(n13739), .B(n13738), .ZN(n13740) );
  NAND2_X1 U15723 ( .A1(n13740), .A2(n13822), .ZN(n13895) );
  INV_X1 U15724 ( .A(n13741), .ZN(n13896) );
  AOI21_X1 U15725 ( .B1(n13895), .B2(n13896), .A(n6430), .ZN(n13742) );
  AOI211_X1 U15726 ( .C1(n13848), .C2(n13893), .A(n13743), .B(n13742), .ZN(
        n13744) );
  INV_X1 U15727 ( .A(n13744), .ZN(P2_U3242) );
  XNOR2_X1 U15728 ( .A(n13745), .B(n13748), .ZN(n13747) );
  OAI21_X1 U15729 ( .B1(n13747), .B2(n13795), .A(n13746), .ZN(n13902) );
  INV_X1 U15730 ( .A(n13902), .ZN(n13759) );
  NAND2_X1 U15731 ( .A1(n13749), .A2(n13748), .ZN(n13750) );
  AND2_X1 U15732 ( .A1(n13751), .A2(n13750), .ZN(n13903) );
  AOI211_X1 U15733 ( .C1(n13753), .C2(n13761), .A(n13687), .B(n13730), .ZN(
        n13901) );
  NAND2_X1 U15734 ( .A1(n13901), .A2(n13850), .ZN(n13756) );
  AOI22_X1 U15735 ( .A1(n6430), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13754), 
        .B2(n13828), .ZN(n13755) );
  OAI211_X1 U15736 ( .C1(n13970), .C2(n13816), .A(n13756), .B(n13755), .ZN(
        n13757) );
  AOI21_X1 U15737 ( .B1(n13848), .B2(n13903), .A(n13757), .ZN(n13758) );
  OAI21_X1 U15738 ( .B1(n6430), .B2(n13759), .A(n13758), .ZN(P2_U3243) );
  XNOR2_X1 U15739 ( .A(n13760), .B(n13767), .ZN(n13906) );
  OAI211_X1 U15740 ( .C1(n13783), .C2(n13975), .A(n10023), .B(n13761), .ZN(
        n13907) );
  AOI22_X1 U15741 ( .A1(n6430), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13762), 
        .B2(n13828), .ZN(n13765) );
  NAND2_X1 U15742 ( .A1(n13763), .A2(n13846), .ZN(n13764) );
  OAI211_X1 U15743 ( .C1(n13907), .C2(n13766), .A(n13765), .B(n13764), .ZN(
        n13773) );
  INV_X1 U15744 ( .A(n13767), .ZN(n13768) );
  XNOR2_X1 U15745 ( .A(n13769), .B(n13768), .ZN(n13771) );
  AOI21_X1 U15746 ( .B1(n13771), .B2(n13822), .A(n13770), .ZN(n13909) );
  NOR2_X1 U15747 ( .A1(n13909), .A2(n6430), .ZN(n13772) );
  AOI211_X1 U15748 ( .C1(n13906), .C2(n13848), .A(n13773), .B(n13772), .ZN(
        n13774) );
  INV_X1 U15749 ( .A(n13774), .ZN(P2_U3244) );
  XNOR2_X1 U15750 ( .A(n13776), .B(n13775), .ZN(n13917) );
  XNOR2_X1 U15751 ( .A(n13778), .B(n13777), .ZN(n13780) );
  OAI21_X1 U15752 ( .B1(n13780), .B2(n13795), .A(n13779), .ZN(n13913) );
  NAND2_X1 U15753 ( .A1(n13798), .A2(n13915), .ZN(n13781) );
  NAND2_X1 U15754 ( .A1(n13781), .A2(n10023), .ZN(n13782) );
  NOR2_X1 U15755 ( .A1(n13783), .A2(n13782), .ZN(n13914) );
  NAND2_X1 U15756 ( .A1(n13914), .A2(n13850), .ZN(n13788) );
  INV_X1 U15757 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13785) );
  OAI22_X1 U15758 ( .A1(n13844), .A2(n13785), .B1(n13784), .B2(n13841), .ZN(
        n13786) );
  AOI21_X1 U15759 ( .B1(n13915), .B2(n13846), .A(n13786), .ZN(n13787) );
  NAND2_X1 U15760 ( .A1(n13788), .A2(n13787), .ZN(n13789) );
  AOI21_X1 U15761 ( .B1(n13913), .B2(n13844), .A(n13789), .ZN(n13790) );
  OAI21_X1 U15762 ( .B1(n13835), .B2(n13917), .A(n13790), .ZN(P2_U3245) );
  XOR2_X1 U15763 ( .A(n13793), .B(n13791), .Z(n13922) );
  XOR2_X1 U15764 ( .A(n13793), .B(n13792), .Z(n13796) );
  OAI21_X1 U15765 ( .B1(n13796), .B2(n13795), .A(n13794), .ZN(n13918) );
  INV_X1 U15766 ( .A(n13797), .ZN(n13811) );
  AOI21_X1 U15767 ( .B1(n13920), .B2(n13811), .A(n13687), .ZN(n13799) );
  AND2_X1 U15768 ( .A1(n13799), .A2(n13798), .ZN(n13919) );
  NAND2_X1 U15769 ( .A1(n13919), .A2(n13850), .ZN(n13802) );
  AOI22_X1 U15770 ( .A1(n6430), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13800), 
        .B2(n13828), .ZN(n13801) );
  OAI211_X1 U15771 ( .C1(n13566), .C2(n13816), .A(n13802), .B(n13801), .ZN(
        n13803) );
  AOI21_X1 U15772 ( .B1(n13918), .B2(n13844), .A(n13803), .ZN(n13804) );
  OAI21_X1 U15773 ( .B1(n13835), .B2(n13922), .A(n13804), .ZN(P2_U3246) );
  XOR2_X1 U15774 ( .A(n13809), .B(n13805), .Z(n13807) );
  AOI21_X1 U15775 ( .B1(n13807), .B2(n13822), .A(n13806), .ZN(n13926) );
  OAI21_X1 U15776 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n13923) );
  INV_X1 U15777 ( .A(n13925), .ZN(n13817) );
  AOI211_X1 U15778 ( .C1(n13925), .C2(n13825), .A(n13343), .B(n13797), .ZN(
        n13924) );
  NAND2_X1 U15779 ( .A1(n13924), .A2(n13850), .ZN(n13815) );
  INV_X1 U15780 ( .A(n13812), .ZN(n13813) );
  AOI22_X1 U15781 ( .A1(n6430), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13813), 
        .B2(n13828), .ZN(n13814) );
  OAI211_X1 U15782 ( .C1(n13817), .C2(n13816), .A(n13815), .B(n13814), .ZN(
        n13818) );
  AOI21_X1 U15783 ( .B1(n13848), .B2(n13923), .A(n13818), .ZN(n13819) );
  OAI21_X1 U15784 ( .B1(n6430), .B2(n13926), .A(n13819), .ZN(P2_U3247) );
  XNOR2_X1 U15785 ( .A(n13820), .B(n13834), .ZN(n13823) );
  AOI21_X1 U15786 ( .B1(n13823), .B2(n13822), .A(n13821), .ZN(n13932) );
  AOI21_X1 U15787 ( .B1(n13824), .B2(n13930), .A(n13343), .ZN(n13826) );
  AND2_X1 U15788 ( .A1(n13826), .A2(n13825), .ZN(n13929) );
  NAND2_X1 U15789 ( .A1(n13930), .A2(n13846), .ZN(n13830) );
  NAND2_X1 U15790 ( .A1(n13828), .A2(n13827), .ZN(n13829) );
  OAI211_X1 U15791 ( .C1(n13844), .C2(n13831), .A(n13830), .B(n13829), .ZN(
        n13837) );
  OAI21_X1 U15792 ( .B1(n13834), .B2(n13833), .A(n13832), .ZN(n13933) );
  NOR2_X1 U15793 ( .A1(n13933), .A2(n13835), .ZN(n13836) );
  AOI211_X1 U15794 ( .C1(n13929), .C2(n13850), .A(n13837), .B(n13836), .ZN(
        n13838) );
  OAI21_X1 U15795 ( .B1(n6430), .B2(n13932), .A(n13838), .ZN(P2_U3248) );
  NAND2_X1 U15796 ( .A1(n13839), .A2(n13844), .ZN(n13855) );
  INV_X1 U15797 ( .A(n13840), .ZN(n13842) );
  OAI22_X1 U15798 ( .A1(n13844), .A2(n13843), .B1(n13842), .B2(n13841), .ZN(
        n13845) );
  AOI21_X1 U15799 ( .B1(n13847), .B2(n13846), .A(n13845), .ZN(n13854) );
  NAND2_X1 U15800 ( .A1(n13849), .A2(n13848), .ZN(n13853) );
  NAND2_X1 U15801 ( .A1(n13851), .A2(n13850), .ZN(n13852) );
  NAND4_X1 U15802 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        P2_U3253) );
  MUX2_X1 U15803 ( .A(n15445), .B(n13940), .S(n15190), .Z(n13857) );
  OAI21_X1 U15804 ( .B1(n13942), .B2(n13912), .A(n13857), .ZN(P2_U3530) );
  INV_X1 U15805 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13860) );
  AND2_X1 U15806 ( .A1(n13859), .A2(n13858), .ZN(n13943) );
  MUX2_X1 U15807 ( .A(n13860), .B(n13943), .S(n15190), .Z(n13861) );
  OAI21_X1 U15808 ( .B1(n13946), .B2(n13912), .A(n13861), .ZN(P2_U3529) );
  MUX2_X1 U15809 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13948), .S(n15190), .Z(
        n13869) );
  INV_X1 U15810 ( .A(n13869), .ZN(n13870) );
  OAI21_X1 U15811 ( .B1(n13951), .B2(n13912), .A(n13870), .ZN(P2_U3527) );
  NAND2_X1 U15812 ( .A1(n13871), .A2(n15179), .ZN(n13876) );
  NAND3_X1 U15813 ( .A1(n13873), .A2(n13905), .A3(n13872), .ZN(n13875) );
  NAND4_X1 U15814 ( .A1(n13877), .A2(n13876), .A3(n13875), .A4(n13874), .ZN(
        n13952) );
  MUX2_X1 U15815 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13952), .S(n15190), .Z(
        P2_U3526) );
  OAI211_X1 U15816 ( .C1(n13880), .C2(n15182), .A(n13879), .B(n13878), .ZN(
        n13953) );
  MUX2_X1 U15817 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13953), .S(n15190), .Z(
        n13881) );
  AOI21_X1 U15818 ( .B1(n13899), .B2(n13955), .A(n13881), .ZN(n13882) );
  INV_X1 U15819 ( .A(n13882), .ZN(P2_U3525) );
  INV_X1 U15820 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15447) );
  AOI211_X1 U15821 ( .C1(n13905), .C2(n13885), .A(n13884), .B(n13883), .ZN(
        n13957) );
  MUX2_X1 U15822 ( .A(n15447), .B(n13957), .S(n15190), .Z(n13886) );
  OAI21_X1 U15823 ( .B1(n13960), .B2(n13912), .A(n13886), .ZN(P2_U3524) );
  AOI21_X1 U15824 ( .B1(n15179), .B2(n13888), .A(n13887), .ZN(n13889) );
  OAI211_X1 U15825 ( .C1(n13892), .C2(n13891), .A(n13890), .B(n13889), .ZN(
        n13961) );
  MUX2_X1 U15826 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13961), .S(n15190), .Z(
        P2_U3523) );
  NAND2_X1 U15827 ( .A1(n13893), .A2(n13905), .ZN(n13897) );
  NAND4_X1 U15828 ( .A1(n13897), .A2(n13896), .A3(n13895), .A4(n13894), .ZN(
        n13962) );
  MUX2_X1 U15829 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13962), .S(n15190), .Z(
        n13898) );
  AOI21_X1 U15830 ( .B1(n13899), .B2(n13964), .A(n13898), .ZN(n13900) );
  INV_X1 U15831 ( .A(n13900), .ZN(P2_U3522) );
  INV_X1 U15832 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15446) );
  AOI211_X1 U15833 ( .C1(n13903), .C2(n13905), .A(n13902), .B(n13901), .ZN(
        n13967) );
  MUX2_X1 U15834 ( .A(n15446), .B(n13967), .S(n15190), .Z(n13904) );
  OAI21_X1 U15835 ( .B1(n13970), .B2(n13912), .A(n13904), .ZN(P2_U3521) );
  INV_X1 U15836 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13910) );
  NAND2_X1 U15837 ( .A1(n13906), .A2(n13905), .ZN(n13908) );
  AND3_X1 U15838 ( .A1(n13909), .A2(n13908), .A3(n13907), .ZN(n13971) );
  MUX2_X1 U15839 ( .A(n13910), .B(n13971), .S(n15190), .Z(n13911) );
  OAI21_X1 U15840 ( .B1(n13975), .B2(n13912), .A(n13911), .ZN(P2_U3520) );
  AOI211_X1 U15841 ( .C1(n15179), .C2(n13915), .A(n13914), .B(n13913), .ZN(
        n13916) );
  OAI21_X1 U15842 ( .B1(n15182), .B2(n13917), .A(n13916), .ZN(n13976) );
  MUX2_X1 U15843 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13976), .S(n15190), .Z(
        P2_U3519) );
  AOI211_X1 U15844 ( .C1(n15179), .C2(n13920), .A(n13919), .B(n13918), .ZN(
        n13921) );
  OAI21_X1 U15845 ( .B1(n15182), .B2(n13922), .A(n13921), .ZN(n13977) );
  MUX2_X1 U15846 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13977), .S(n15190), .Z(
        P2_U3518) );
  INV_X1 U15847 ( .A(n13923), .ZN(n13928) );
  AOI21_X1 U15848 ( .B1(n15179), .B2(n13925), .A(n13924), .ZN(n13927) );
  OAI211_X1 U15849 ( .C1(n15182), .C2(n13928), .A(n13927), .B(n13926), .ZN(
        n13978) );
  MUX2_X1 U15850 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13978), .S(n15190), .Z(
        P2_U3517) );
  AOI21_X1 U15851 ( .B1(n15179), .B2(n13930), .A(n13929), .ZN(n13931) );
  OAI211_X1 U15852 ( .C1(n13933), .C2(n15182), .A(n13932), .B(n13931), .ZN(
        n13979) );
  MUX2_X1 U15853 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13979), .S(n15190), .Z(
        P2_U3516) );
  AOI21_X1 U15854 ( .B1(n15179), .B2(n14887), .A(n13934), .ZN(n13935) );
  OAI211_X1 U15855 ( .C1(n15182), .C2(n13937), .A(n13936), .B(n13935), .ZN(
        n13980) );
  MUX2_X1 U15856 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13980), .S(n15190), .Z(
        P2_U3513) );
  MUX2_X1 U15857 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n13938), .S(n15190), .Z(
        P2_U3504) );
  MUX2_X1 U15858 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n13939), .S(n15190), .Z(
        P2_U3499) );
  INV_X1 U15859 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13941) );
  INV_X1 U15860 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13944) );
  MUX2_X1 U15861 ( .A(n13944), .B(n13943), .S(n15187), .Z(n13945) );
  OAI21_X1 U15862 ( .B1(n13946), .B2(n13974), .A(n13945), .ZN(P2_U3497) );
  MUX2_X1 U15863 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13948), .S(n15187), .Z(
        n13949) );
  INV_X1 U15864 ( .A(n13949), .ZN(n13950) );
  OAI21_X1 U15865 ( .B1(n13951), .B2(n13974), .A(n13950), .ZN(P2_U3495) );
  MUX2_X1 U15866 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13952), .S(n15187), .Z(
        P2_U3494) );
  MUX2_X1 U15867 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13953), .S(n15187), .Z(
        n13954) );
  AOI21_X1 U15868 ( .B1(n13965), .B2(n13955), .A(n13954), .ZN(n13956) );
  INV_X1 U15869 ( .A(n13956), .ZN(P2_U3493) );
  INV_X1 U15870 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13958) );
  MUX2_X1 U15871 ( .A(n13958), .B(n13957), .S(n15187), .Z(n13959) );
  OAI21_X1 U15872 ( .B1(n13960), .B2(n13974), .A(n13959), .ZN(P2_U3492) );
  MUX2_X1 U15873 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13961), .S(n15187), .Z(
        P2_U3491) );
  MUX2_X1 U15874 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13962), .S(n15187), .Z(
        n13963) );
  AOI21_X1 U15875 ( .B1(n13965), .B2(n13964), .A(n13963), .ZN(n13966) );
  INV_X1 U15876 ( .A(n13966), .ZN(P2_U3490) );
  INV_X1 U15877 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13968) );
  MUX2_X1 U15878 ( .A(n13968), .B(n13967), .S(n15187), .Z(n13969) );
  OAI21_X1 U15879 ( .B1(n13970), .B2(n13974), .A(n13969), .ZN(P2_U3489) );
  MUX2_X1 U15880 ( .A(n13972), .B(n13971), .S(n15187), .Z(n13973) );
  OAI21_X1 U15881 ( .B1(n13975), .B2(n13974), .A(n13973), .ZN(P2_U3488) );
  MUX2_X1 U15882 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13976), .S(n15187), .Z(
        P2_U3487) );
  MUX2_X1 U15883 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13977), .S(n15187), .Z(
        P2_U3486) );
  MUX2_X1 U15884 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13978), .S(n15187), .Z(
        P2_U3484) );
  MUX2_X1 U15885 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13979), .S(n15187), .Z(
        P2_U3481) );
  MUX2_X1 U15886 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13980), .S(n15187), .Z(
        P2_U3472) );
  INV_X1 U15887 ( .A(n11892), .ZN(n14692) );
  NOR4_X1 U15888 ( .A1(n13981), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13982), .A4(
        P2_U3088), .ZN(n13983) );
  AOI21_X1 U15889 ( .B1(n13992), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13983), 
        .ZN(n13984) );
  OAI21_X1 U15890 ( .B1(n14692), .B2(n13994), .A(n13984), .ZN(P2_U3296) );
  OAI222_X1 U15891 ( .A1(n14001), .A2(n14694), .B1(P2_U3088), .B2(n13986), 
        .C1(n13985), .C2(n13999), .ZN(P2_U3297) );
  INV_X1 U15892 ( .A(n13987), .ZN(n14696) );
  OAI222_X1 U15893 ( .A1(n14001), .A2(n14696), .B1(P2_U3088), .B2(n13988), 
        .C1(n13989), .C2(n13999), .ZN(P2_U3298) );
  INV_X1 U15894 ( .A(n13990), .ZN(n14699) );
  AOI21_X1 U15895 ( .B1(n13992), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13991), 
        .ZN(n13993) );
  OAI21_X1 U15896 ( .B1(n14699), .B2(n13994), .A(n13993), .ZN(P2_U3299) );
  INV_X1 U15897 ( .A(n13995), .ZN(n14703) );
  OAI222_X1 U15898 ( .A1(n13999), .A2(n13997), .B1(n14001), .B2(n14703), .C1(
        n13996), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15899 ( .A(n13998), .ZN(n14706) );
  OAI222_X1 U15900 ( .A1(n14002), .A2(P2_U3088), .B1(n14001), .B2(n14706), 
        .C1(n14000), .C2(n13999), .ZN(P2_U3301) );
  INV_X1 U15901 ( .A(n14003), .ZN(n14004) );
  MUX2_X1 U15902 ( .A(n14004), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15903 ( .A(n14315), .ZN(n14350) );
  AOI22_X1 U15904 ( .A1(n14923), .A2(n14281), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14007) );
  NAND2_X1 U15905 ( .A1(n14113), .A2(n14355), .ZN(n14006) );
  OAI211_X1 U15906 ( .C1(n14350), .C2(n14120), .A(n14007), .B(n14006), .ZN(
        n14008) );
  AOI21_X1 U15907 ( .B1(n14576), .B2(n14131), .A(n14008), .ZN(n14009) );
  OAI21_X1 U15908 ( .B1(n14010), .B2(n14133), .A(n14009), .ZN(P1_U3214) );
  XOR2_X1 U15909 ( .A(n14012), .B(n14011), .Z(n14017) );
  AOI22_X1 U15910 ( .A1(n14275), .A2(n15007), .B1(n14509), .B2(n14278), .ZN(
        n14413) );
  OAI22_X1 U15911 ( .A1(n14413), .A2(n14111), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14013), .ZN(n14014) );
  AOI21_X1 U15912 ( .B1(n14420), .B2(n14113), .A(n14014), .ZN(n14016) );
  NAND2_X1 U15913 ( .A1(n14600), .A2(n14131), .ZN(n14015) );
  OAI211_X1 U15914 ( .C1(n14017), .C2(n14133), .A(n14016), .B(n14015), .ZN(
        P1_U3216) );
  INV_X1 U15915 ( .A(n14475), .ZN(n14684) );
  AOI21_X1 U15916 ( .B1(n14019), .B2(n14018), .A(n14133), .ZN(n14021) );
  NAND2_X1 U15917 ( .A1(n14021), .A2(n14020), .ZN(n14025) );
  NAND2_X1 U15918 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14249)
         );
  NAND2_X1 U15919 ( .A1(n14923), .A2(n14510), .ZN(n14022) );
  OAI211_X1 U15920 ( .C1(n14471), .C2(n14120), .A(n14249), .B(n14022), .ZN(
        n14023) );
  AOI21_X1 U15921 ( .B1(n14478), .B2(n14113), .A(n14023), .ZN(n14024) );
  OAI211_X1 U15922 ( .C1(n14684), .C2(n14927), .A(n14025), .B(n14024), .ZN(
        P1_U3219) );
  INV_X1 U15923 ( .A(n14026), .ZN(n14027) );
  AOI21_X1 U15924 ( .B1(n14029), .B2(n14028), .A(n14027), .ZN(n14035) );
  NAND2_X1 U15925 ( .A1(n14275), .A2(n14509), .ZN(n14031) );
  OR2_X1 U15926 ( .A1(n14471), .A2(n14525), .ZN(n14030) );
  NAND2_X1 U15927 ( .A1(n14031), .A2(n14030), .ZN(n14612) );
  AOI22_X1 U15928 ( .A1(n14612), .A2(n14143), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14032) );
  OAI21_X1 U15929 ( .B1(n14444), .B2(n14935), .A(n14032), .ZN(n14033) );
  AOI21_X1 U15930 ( .B1(n14443), .B2(n14131), .A(n14033), .ZN(n14034) );
  OAI21_X1 U15931 ( .B1(n14035), .B2(n14133), .A(n14034), .ZN(P1_U3223) );
  OAI211_X1 U15932 ( .C1(n14038), .C2(n14037), .A(n14036), .B(n14930), .ZN(
        n14044) );
  OAI22_X1 U15933 ( .A1(n14111), .A2(n14040), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14039), .ZN(n14041) );
  AOI21_X1 U15934 ( .B1(n14113), .B2(n14042), .A(n14041), .ZN(n14043) );
  OAI211_X1 U15935 ( .C1(n6840), .C2(n14927), .A(n14044), .B(n14043), .ZN(
        P1_U3224) );
  XOR2_X1 U15936 ( .A(n14046), .B(n14045), .Z(n14051) );
  AOI22_X1 U15937 ( .A1(n14509), .A2(n14281), .B1(n15007), .B2(n14278), .ZN(
        n14381) );
  OAI22_X1 U15938 ( .A1(n14111), .A2(n14381), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14047), .ZN(n14049) );
  NOR2_X1 U15939 ( .A1(n14668), .A2(n14927), .ZN(n14048) );
  AOI211_X1 U15940 ( .C1(n14113), .C2(n14385), .A(n14049), .B(n14048), .ZN(
        n14050) );
  OAI21_X1 U15941 ( .B1(n14051), .B2(n14133), .A(n14050), .ZN(P1_U3225) );
  XOR2_X1 U15942 ( .A(n14053), .B(n14052), .Z(n14059) );
  INV_X1 U15943 ( .A(n14488), .ZN(n14526) );
  OAI21_X1 U15944 ( .B1(n14120), .B2(n14526), .A(n14054), .ZN(n14055) );
  AOI21_X1 U15945 ( .B1(n14923), .B2(n14898), .A(n14055), .ZN(n14056) );
  OAI21_X1 U15946 ( .B1(n14533), .B2(n14935), .A(n14056), .ZN(n14057) );
  AOI21_X1 U15947 ( .B1(n14535), .B2(n14131), .A(n14057), .ZN(n14058) );
  OAI21_X1 U15948 ( .B1(n14059), .B2(n14133), .A(n14058), .ZN(P1_U3226) );
  INV_X1 U15949 ( .A(n14060), .ZN(n14062) );
  NOR2_X1 U15950 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  XNOR2_X1 U15951 ( .A(n14064), .B(n14063), .ZN(n14065) );
  NAND2_X1 U15952 ( .A1(n14065), .A2(n14930), .ZN(n14072) );
  AOI22_X1 U15953 ( .A1(n14143), .A2(n14066), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14071) );
  NAND2_X1 U15954 ( .A1(n14131), .A2(n14067), .ZN(n14070) );
  OR2_X1 U15955 ( .A1(n14935), .A2(n14068), .ZN(n14069) );
  NAND4_X1 U15956 ( .A1(n14072), .A2(n14071), .A3(n14070), .A4(n14069), .ZN(
        P1_U3227) );
  XOR2_X1 U15957 ( .A(n14073), .B(n14074), .Z(n14080) );
  NOR2_X1 U15958 ( .A1(n14935), .A2(n14511), .ZN(n14078) );
  NAND2_X1 U15959 ( .A1(n14923), .A2(n14507), .ZN(n14076) );
  OAI211_X1 U15960 ( .C1(n14120), .C2(n14472), .A(n14076), .B(n14075), .ZN(
        n14077) );
  AOI211_X1 U15961 ( .C1(n14637), .C2(n14131), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI21_X1 U15962 ( .B1(n14080), .B2(n14133), .A(n14079), .ZN(P1_U3228) );
  XOR2_X1 U15963 ( .A(n14082), .B(n14081), .Z(n14087) );
  INV_X1 U15964 ( .A(n14399), .ZN(n14307) );
  AOI22_X1 U15965 ( .A1(n14923), .A2(n14398), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14084) );
  NAND2_X1 U15966 ( .A1(n14113), .A2(n14406), .ZN(n14083) );
  OAI211_X1 U15967 ( .C1(n14307), .C2(n14120), .A(n14084), .B(n14083), .ZN(
        n14085) );
  AOI21_X1 U15968 ( .B1(n14593), .B2(n14131), .A(n14085), .ZN(n14086) );
  OAI21_X1 U15969 ( .B1(n14087), .B2(n14133), .A(n14086), .ZN(P1_U3229) );
  OAI211_X1 U15970 ( .C1(n14090), .C2(n14089), .A(n14088), .B(n14930), .ZN(
        n14096) );
  NAND2_X1 U15971 ( .A1(n14299), .A2(n14509), .ZN(n14092) );
  OR2_X1 U15972 ( .A1(n14297), .A2(n14525), .ZN(n14091) );
  AND2_X1 U15973 ( .A1(n14092), .A2(n14091), .ZN(n14619) );
  INV_X1 U15974 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14093) );
  OAI22_X1 U15975 ( .A1(n14619), .A2(n14111), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14093), .ZN(n14094) );
  AOI21_X1 U15976 ( .B1(n14457), .B2(n14113), .A(n14094), .ZN(n14095) );
  OAI211_X1 U15977 ( .C1(n14679), .C2(n14927), .A(n14096), .B(n14095), .ZN(
        P1_U3233) );
  OAI211_X1 U15978 ( .C1(n14098), .C2(n14097), .A(n14893), .B(n14930), .ZN(
        n14104) );
  OAI21_X1 U15979 ( .B1(n14111), .B2(n14100), .A(n14099), .ZN(n14101) );
  AOI21_X1 U15980 ( .B1(n14113), .B2(n14102), .A(n14101), .ZN(n14103) );
  OAI211_X1 U15981 ( .C1(n7282), .C2(n14927), .A(n14104), .B(n14103), .ZN(
        P1_U3234) );
  OAI21_X1 U15982 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(n14108) );
  NAND2_X1 U15983 ( .A1(n14108), .A2(n14930), .ZN(n14115) );
  INV_X1 U15984 ( .A(n14398), .ZN(n14304) );
  NOR2_X1 U15985 ( .A1(n14304), .A2(n14527), .ZN(n14109) );
  AOI21_X1 U15986 ( .B1(n14299), .B2(n15007), .A(n14109), .ZN(n14604) );
  INV_X1 U15987 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14110) );
  OAI22_X1 U15988 ( .A1(n14604), .A2(n14111), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14110), .ZN(n14112) );
  AOI21_X1 U15989 ( .B1(n14436), .B2(n14113), .A(n14112), .ZN(n14114) );
  OAI211_X1 U15990 ( .C1(n14927), .C2(n14606), .A(n14115), .B(n14114), .ZN(
        P1_U3235) );
  XOR2_X1 U15991 ( .A(n14116), .B(n14117), .Z(n14124) );
  NOR2_X1 U15992 ( .A1(n14935), .A2(n14495), .ZN(n14122) );
  NAND2_X1 U15993 ( .A1(n14923), .A2(n14488), .ZN(n14119) );
  OAI211_X1 U15994 ( .C1(n14120), .C2(n14297), .A(n14119), .B(n14118), .ZN(
        n14121) );
  AOI211_X1 U15995 ( .C1(n14633), .C2(n14131), .A(n14122), .B(n14121), .ZN(
        n14123) );
  OAI21_X1 U15996 ( .B1(n14124), .B2(n14133), .A(n14123), .ZN(P1_U3238) );
  XOR2_X1 U15997 ( .A(n14126), .B(n14125), .Z(n14134) );
  INV_X1 U15998 ( .A(n14365), .ZN(n14129) );
  INV_X1 U15999 ( .A(n14284), .ZN(n14309) );
  NAND2_X1 U16000 ( .A1(n14399), .A2(n15007), .ZN(n14127) );
  OAI21_X1 U16001 ( .B1(n14309), .B2(n14527), .A(n14127), .ZN(n14582) );
  AOI22_X1 U16002 ( .A1(n14143), .A2(n14582), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14128) );
  OAI21_X1 U16003 ( .B1(n14129), .B2(n14935), .A(n14128), .ZN(n14130) );
  AOI21_X1 U16004 ( .B1(n14583), .B2(n14131), .A(n14130), .ZN(n14132) );
  OAI21_X1 U16005 ( .B1(n14134), .B2(n14133), .A(n14132), .ZN(P1_U3240) );
  OAI21_X1 U16006 ( .B1(n14137), .B2(n14136), .A(n14135), .ZN(n14138) );
  NAND2_X1 U16007 ( .A1(n14138), .A2(n14930), .ZN(n14145) );
  NAND2_X1 U16008 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14994)
         );
  INV_X1 U16009 ( .A(n14994), .ZN(n14141) );
  NOR2_X1 U16010 ( .A1(n14935), .A2(n14139), .ZN(n14140) );
  AOI211_X1 U16011 ( .C1(n14143), .C2(n14142), .A(n14141), .B(n14140), .ZN(
        n14144) );
  OAI211_X1 U16012 ( .C1(n7280), .C2(n14927), .A(n14145), .B(n14144), .ZN(
        P1_U3241) );
  MUX2_X1 U16013 ( .A(n14254), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14156), .Z(
        P1_U3591) );
  MUX2_X1 U16014 ( .A(n14316), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14156), .Z(
        P1_U3590) );
  MUX2_X1 U16015 ( .A(n14146), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14156), .Z(
        P1_U3589) );
  MUX2_X1 U16016 ( .A(n14315), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14156), .Z(
        P1_U3588) );
  MUX2_X1 U16017 ( .A(n14284), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14156), .Z(
        P1_U3587) );
  MUX2_X1 U16018 ( .A(n14281), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14156), .Z(
        P1_U3586) );
  MUX2_X1 U16019 ( .A(n14399), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14156), .Z(
        P1_U3585) );
  MUX2_X1 U16020 ( .A(n14278), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14156), .Z(
        P1_U3584) );
  MUX2_X1 U16021 ( .A(n14398), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14156), .Z(
        P1_U3583) );
  MUX2_X1 U16022 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14275), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16023 ( .A(n14299), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14156), .Z(
        P1_U3581) );
  MUX2_X1 U16024 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14147), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16025 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14489), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16026 ( .A(n14510), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14156), .Z(
        P1_U3578) );
  MUX2_X1 U16027 ( .A(n14488), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14156), .Z(
        P1_U3577) );
  MUX2_X1 U16028 ( .A(n14507), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14156), .Z(
        P1_U3576) );
  MUX2_X1 U16029 ( .A(n14898), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14156), .Z(
        P1_U3575) );
  MUX2_X1 U16030 ( .A(n14148), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14156), .Z(
        P1_U3574) );
  MUX2_X1 U16031 ( .A(n14897), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14156), .Z(
        P1_U3573) );
  MUX2_X1 U16032 ( .A(n14924), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14156), .Z(
        P1_U3572) );
  MUX2_X1 U16033 ( .A(n14910), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14156), .Z(
        P1_U3571) );
  MUX2_X1 U16034 ( .A(n14922), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14156), .Z(
        P1_U3570) );
  MUX2_X1 U16035 ( .A(n14909), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14156), .Z(
        P1_U3569) );
  MUX2_X1 U16036 ( .A(n14149), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14156), .Z(
        P1_U3568) );
  MUX2_X1 U16037 ( .A(n14150), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14156), .Z(
        P1_U3567) );
  MUX2_X1 U16038 ( .A(n14151), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14156), .Z(
        P1_U3566) );
  MUX2_X1 U16039 ( .A(n14152), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14156), .Z(
        P1_U3565) );
  MUX2_X1 U16040 ( .A(n14153), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14156), .Z(
        P1_U3564) );
  MUX2_X1 U16041 ( .A(n14154), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14156), .Z(
        P1_U3563) );
  MUX2_X1 U16042 ( .A(n14155), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14156), .Z(
        P1_U3562) );
  MUX2_X1 U16043 ( .A(n15002), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14156), .Z(
        P1_U3561) );
  MUX2_X1 U16044 ( .A(n15006), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14156), .Z(
        P1_U3560) );
  INV_X1 U16045 ( .A(n14157), .ZN(n14160) );
  OAI211_X1 U16046 ( .C1(n14160), .C2(n14159), .A(n14243), .B(n14158), .ZN(
        n14170) );
  AOI22_X1 U16047 ( .A1(n14977), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14169) );
  NAND2_X1 U16048 ( .A1(n14219), .A2(n14161), .ZN(n14168) );
  MUX2_X1 U16049 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n15112), .S(n14162), .Z(
        n14163) );
  OAI21_X1 U16050 ( .B1(n9735), .B2(n14164), .A(n14163), .ZN(n14165) );
  NAND3_X1 U16051 ( .A1(n14245), .A2(n14166), .A3(n14165), .ZN(n14167) );
  NAND4_X1 U16052 ( .A1(n14170), .A2(n14169), .A3(n14168), .A4(n14167), .ZN(
        P1_U3244) );
  OAI22_X1 U16053 ( .A1(n14996), .A2(n7359), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14171), .ZN(n14172) );
  AOI21_X1 U16054 ( .B1(n14173), .B2(n14219), .A(n14172), .ZN(n14180) );
  OAI211_X1 U16055 ( .C1(n14175), .C2(n14174), .A(n14243), .B(n14193), .ZN(
        n14179) );
  OAI211_X1 U16056 ( .C1(n14177), .C2(n14176), .A(n14245), .B(n14187), .ZN(
        n14178) );
  NAND4_X1 U16057 ( .A1(n14181), .A2(n14180), .A3(n14179), .A4(n14178), .ZN(
        P1_U3245) );
  INV_X1 U16058 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14182) );
  OAI22_X1 U16059 ( .A1(n14996), .A2(n14182), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10133), .ZN(n14183) );
  AOI21_X1 U16060 ( .B1(n14184), .B2(n14219), .A(n14183), .ZN(n14198) );
  MUX2_X1 U16061 ( .A(n9479), .B(P1_REG1_REG_3__SCAN_IN), .S(n14184), .Z(
        n14185) );
  NAND3_X1 U16062 ( .A1(n14187), .A2(n14186), .A3(n14185), .ZN(n14188) );
  NAND3_X1 U16063 ( .A1(n14245), .A2(n14189), .A3(n14188), .ZN(n14197) );
  INV_X1 U16064 ( .A(n14190), .ZN(n14195) );
  NAND3_X1 U16065 ( .A1(n14193), .A2(n14192), .A3(n14191), .ZN(n14194) );
  NAND3_X1 U16066 ( .A1(n14243), .A2(n14195), .A3(n14194), .ZN(n14196) );
  NAND3_X1 U16067 ( .A1(n14198), .A2(n14197), .A3(n14196), .ZN(P1_U3246) );
  NOR2_X1 U16068 ( .A1(n14996), .A2(n14725), .ZN(n14199) );
  AOI211_X1 U16069 ( .C1(n14219), .C2(n14205), .A(n14200), .B(n14199), .ZN(
        n14213) );
  OAI211_X1 U16070 ( .C1(n14203), .C2(n14202), .A(n14245), .B(n14201), .ZN(
        n14212) );
  INV_X1 U16071 ( .A(n14204), .ZN(n14207) );
  MUX2_X1 U16072 ( .A(n9520), .B(P1_REG2_REG_6__SCAN_IN), .S(n14205), .Z(
        n14206) );
  NAND3_X1 U16073 ( .A1(n14208), .A2(n14207), .A3(n14206), .ZN(n14209) );
  NAND3_X1 U16074 ( .A1(n14243), .A2(n14210), .A3(n14209), .ZN(n14211) );
  NAND3_X1 U16075 ( .A1(n14213), .A2(n14212), .A3(n14211), .ZN(P1_U3249) );
  NAND2_X1 U16076 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n14915)
         );
  AOI21_X1 U16077 ( .B1(n14215), .B2(n14214), .A(n14987), .ZN(n14217) );
  NAND2_X1 U16078 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  AND2_X1 U16079 ( .A1(n14915), .A2(n14218), .ZN(n14229) );
  AOI22_X1 U16080 ( .A1(n14219), .A2(n14220), .B1(n14977), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n14228) );
  MUX2_X1 U16081 ( .A(n9776), .B(P1_REG2_REG_10__SCAN_IN), .S(n14220), .Z(
        n14223) );
  INV_X1 U16082 ( .A(n14221), .ZN(n14222) );
  NAND2_X1 U16083 ( .A1(n14223), .A2(n14222), .ZN(n14225) );
  OAI211_X1 U16084 ( .C1(n14226), .C2(n14225), .A(n14224), .B(n14243), .ZN(
        n14227) );
  NAND3_X1 U16085 ( .A1(n14229), .A2(n14228), .A3(n14227), .ZN(P1_U3253) );
  OR2_X1 U16086 ( .A1(n14231), .A2(n14230), .ZN(n14233) );
  NAND2_X1 U16087 ( .A1(n14233), .A2(n14232), .ZN(n14234) );
  XNOR2_X1 U16088 ( .A(n14628), .B(n14234), .ZN(n14246) );
  INV_X1 U16089 ( .A(n14246), .ZN(n14242) );
  NAND2_X1 U16090 ( .A1(n14235), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14239) );
  NAND2_X1 U16091 ( .A1(n14237), .A2(n14236), .ZN(n14238) );
  NAND2_X1 U16092 ( .A1(n14239), .A2(n14238), .ZN(n14240) );
  XOR2_X1 U16093 ( .A(n14240), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14244) );
  OAI21_X1 U16094 ( .B1(n14244), .B2(n14983), .A(n14992), .ZN(n14241) );
  AOI21_X1 U16095 ( .B1(n14245), .B2(n14242), .A(n14241), .ZN(n14248) );
  AOI22_X1 U16096 ( .A1(n14246), .A2(n14245), .B1(n14244), .B2(n14243), .ZN(
        n14247) );
  MUX2_X1 U16097 ( .A(n14248), .B(n14247), .S(n14320), .Z(n14250) );
  OAI211_X1 U16098 ( .C1(n7001), .C2(n14996), .A(n14250), .B(n14249), .ZN(
        P1_U3262) );
  NAND2_X1 U16099 ( .A1(n14463), .A2(n14679), .ZN(n14462) );
  NAND2_X1 U16100 ( .A1(n14662), .A2(n14353), .ZN(n14329) );
  NAND2_X1 U16101 ( .A1(n14659), .A2(n14314), .ZN(n14257) );
  XOR2_X1 U16102 ( .A(n14257), .B(n14251), .Z(n14556) );
  NAND2_X1 U16103 ( .A1(n14556), .A2(n14354), .ZN(n14256) );
  INV_X1 U16104 ( .A(P1_B_REG_SCAN_IN), .ZN(n14252) );
  NOR2_X1 U16105 ( .A1(n9491), .A2(n14252), .ZN(n14253) );
  NOR2_X1 U16106 ( .A1(n14527), .A2(n14253), .ZN(n14317) );
  AND2_X1 U16107 ( .A1(n14317), .A2(n14254), .ZN(n14555) );
  INV_X1 U16108 ( .A(n14555), .ZN(n14559) );
  NOR2_X1 U16109 ( .A1(n15022), .A2(n14559), .ZN(n14259) );
  AOI21_X1 U16110 ( .B1(n15022), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14259), 
        .ZN(n14255) );
  OAI211_X1 U16111 ( .C1(n14654), .C2(n15012), .A(n14256), .B(n14255), .ZN(
        P1_U3263) );
  OAI211_X1 U16112 ( .C1(n14659), .C2(n14314), .A(n15016), .B(n14257), .ZN(
        n14560) );
  NOR2_X1 U16113 ( .A1(n14541), .A2(n14258), .ZN(n14260) );
  AOI211_X1 U16114 ( .C1(n14261), .C2(n14546), .A(n14260), .B(n14259), .ZN(
        n14262) );
  OAI21_X1 U16115 ( .B1(n14560), .B2(n14537), .A(n14262), .ZN(P1_U3264) );
  OR2_X1 U16116 ( .A1(n14264), .A2(n14898), .ZN(n14265) );
  INV_X1 U16117 ( .A(n14521), .ZN(n14529) );
  OR2_X1 U16118 ( .A1(n14535), .A2(n14507), .ZN(n14267) );
  NAND2_X1 U16119 ( .A1(n14637), .A2(n14488), .ZN(n14268) );
  OR2_X1 U16120 ( .A1(n14475), .A2(n14489), .ZN(n14269) );
  OR2_X1 U16121 ( .A1(n14679), .A2(n14471), .ZN(n14272) );
  OR2_X1 U16122 ( .A1(n14443), .A2(n14299), .ZN(n14273) );
  NAND2_X1 U16123 ( .A1(n14274), .A2(n14273), .ZN(n14431) );
  INV_X1 U16124 ( .A(n14427), .ZN(n14430) );
  NAND2_X1 U16125 ( .A1(n14431), .A2(n14430), .ZN(n14429) );
  OR2_X1 U16126 ( .A1(n6457), .A2(n14275), .ZN(n14276) );
  NAND2_X1 U16127 ( .A1(n14600), .A2(n14398), .ZN(n14277) );
  OR2_X1 U16128 ( .A1(n14593), .A2(n14278), .ZN(n14279) );
  INV_X1 U16129 ( .A(n14379), .ZN(n14376) );
  NAND2_X1 U16130 ( .A1(n14389), .A2(n14399), .ZN(n14280) );
  NAND2_X1 U16131 ( .A1(n14362), .A2(n14361), .ZN(n14283) );
  NAND2_X1 U16132 ( .A1(n14583), .A2(n14281), .ZN(n14282) );
  OR2_X1 U16133 ( .A1(n14576), .A2(n14284), .ZN(n14285) );
  XNOR2_X1 U16134 ( .A(n14286), .B(n14312), .ZN(n14568) );
  NAND2_X1 U16135 ( .A1(n14288), .A2(n14287), .ZN(n14290) );
  NAND2_X1 U16136 ( .A1(n14535), .A2(n14291), .ZN(n14292) );
  OR2_X1 U16137 ( .A1(n14637), .A2(n14526), .ZN(n14293) );
  NAND2_X1 U16138 ( .A1(n14503), .A2(n14293), .ZN(n14487) );
  INV_X1 U16139 ( .A(n14484), .ZN(n14486) );
  NAND2_X1 U16140 ( .A1(n14487), .A2(n14486), .ZN(n14295) );
  OR2_X1 U16141 ( .A1(n14633), .A2(n14472), .ZN(n14294) );
  INV_X1 U16142 ( .A(n14299), .ZN(n14300) );
  NAND2_X1 U16143 ( .A1(n6457), .A2(n14301), .ZN(n14302) );
  OR2_X1 U16144 ( .A1(n14593), .A2(n14305), .ZN(n14306) );
  INV_X1 U16145 ( .A(n14361), .ZN(n14371) );
  NAND2_X1 U16146 ( .A1(n14372), .A2(n14371), .ZN(n14370) );
  NAND2_X1 U16147 ( .A1(n14370), .A2(n14346), .ZN(n14308) );
  NAND2_X1 U16148 ( .A1(n14308), .A2(n14344), .ZN(n14348) );
  NAND2_X1 U16149 ( .A1(n14576), .A2(n14309), .ZN(n14310) );
  NAND2_X1 U16150 ( .A1(n14348), .A2(n14310), .ZN(n14326) );
  NAND2_X1 U16151 ( .A1(n14662), .A2(n14315), .ZN(n14311) );
  AOI22_X1 U16152 ( .A1(n14326), .A2(n14311), .B1(n14350), .B2(n14335), .ZN(
        n14313) );
  AOI22_X1 U16153 ( .A1(n14317), .A2(n14316), .B1(n15007), .B2(n14315), .ZN(
        n14563) );
  OAI21_X1 U16154 ( .B1(n14318), .B2(n14544), .A(n14563), .ZN(n14319) );
  AOI21_X1 U16155 ( .B1(n14565), .B2(n14320), .A(n14319), .ZN(n14323) );
  AOI22_X1 U16156 ( .A1(n14321), .A2(n14546), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n15022), .ZN(n14322) );
  OAI21_X1 U16157 ( .B1(n14323), .B2(n15022), .A(n14322), .ZN(n14324) );
  AOI21_X1 U16158 ( .B1(n14518), .B2(n14567), .A(n14324), .ZN(n14325) );
  OAI21_X1 U16159 ( .B1(n14568), .B2(n14520), .A(n14325), .ZN(P1_U3356) );
  XNOR2_X1 U16160 ( .A(n14326), .B(n14337), .ZN(n14571) );
  INV_X1 U16161 ( .A(n14353), .ZN(n14327) );
  AOI21_X1 U16162 ( .B1(n14335), .B2(n14327), .A(n14640), .ZN(n14328) );
  NAND2_X1 U16163 ( .A1(n14329), .A2(n14328), .ZN(n14570) );
  NAND2_X1 U16164 ( .A1(n15022), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14333) );
  INV_X1 U16165 ( .A(n14330), .ZN(n14331) );
  OR2_X1 U16166 ( .A1(n14544), .A2(n14331), .ZN(n14332) );
  OAI211_X1 U16167 ( .C1(n15022), .C2(n14569), .A(n14333), .B(n14332), .ZN(
        n14334) );
  AOI21_X1 U16168 ( .B1(n14335), .B2(n14546), .A(n14334), .ZN(n14336) );
  OAI21_X1 U16169 ( .B1(n14570), .B2(n14537), .A(n14336), .ZN(n14342) );
  NAND2_X1 U16170 ( .A1(n14338), .A2(n14337), .ZN(n14340) );
  NAND2_X1 U16171 ( .A1(n14340), .A2(n14339), .ZN(n14574) );
  NOR2_X1 U16172 ( .A1(n14574), .A2(n14520), .ZN(n14341) );
  INV_X1 U16173 ( .A(n14343), .ZN(P1_U3265) );
  OAI21_X1 U16174 ( .B1(n6488), .B2(n7620), .A(n14345), .ZN(n14575) );
  NAND3_X1 U16175 ( .A1(n14370), .A2(n7620), .A3(n14346), .ZN(n14347) );
  AOI21_X1 U16176 ( .B1(n14348), .B2(n14347), .A(n14936), .ZN(n14352) );
  OAI22_X1 U16177 ( .A1(n14350), .A2(n14527), .B1(n14349), .B2(n14525), .ZN(
        n14351) );
  INV_X1 U16178 ( .A(n14576), .ZN(n14358) );
  AOI21_X1 U16179 ( .B1(n14576), .B2(n14363), .A(n14353), .ZN(n14577) );
  NAND2_X1 U16180 ( .A1(n14577), .A2(n14354), .ZN(n14357) );
  AOI22_X1 U16181 ( .A1(n15022), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14355), 
        .B2(n15013), .ZN(n14356) );
  OAI211_X1 U16182 ( .C1(n14358), .C2(n15012), .A(n14357), .B(n14356), .ZN(
        n14359) );
  AOI21_X1 U16183 ( .B1(n14575), .B2(n15019), .A(n14359), .ZN(n14360) );
  OAI21_X1 U16184 ( .B1(n14579), .B2(n15022), .A(n14360), .ZN(P1_U3266) );
  XNOR2_X1 U16185 ( .A(n14362), .B(n14361), .ZN(n14587) );
  INV_X1 U16186 ( .A(n14363), .ZN(n14364) );
  AOI211_X1 U16187 ( .C1(n14583), .C2(n14384), .A(n14640), .B(n14364), .ZN(
        n14581) );
  INV_X1 U16188 ( .A(n14583), .ZN(n14368) );
  AOI22_X1 U16189 ( .A1(n14541), .A2(n14582), .B1(n14365), .B2(n15013), .ZN(
        n14367) );
  NAND2_X1 U16190 ( .A1(n15022), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n14366) );
  OAI211_X1 U16191 ( .C1(n14368), .C2(n15012), .A(n14367), .B(n14366), .ZN(
        n14369) );
  AOI21_X1 U16192 ( .B1(n14581), .B2(n15018), .A(n14369), .ZN(n14374) );
  OAI21_X1 U16193 ( .B1(n14372), .B2(n14371), .A(n14370), .ZN(n14584) );
  NAND2_X1 U16194 ( .A1(n14584), .A2(n14518), .ZN(n14373) );
  OAI211_X1 U16195 ( .C1(n14587), .C2(n14520), .A(n14374), .B(n14373), .ZN(
        P1_U3267) );
  OAI21_X1 U16196 ( .B1(n14377), .B2(n14376), .A(n14375), .ZN(n14590) );
  OAI21_X1 U16197 ( .B1(n14380), .B2(n14379), .A(n14378), .ZN(n14383) );
  INV_X1 U16198 ( .A(n14381), .ZN(n14382) );
  AOI21_X1 U16199 ( .B1(n14383), .B2(n15079), .A(n14382), .ZN(n14589) );
  INV_X1 U16200 ( .A(n14589), .ZN(n14388) );
  OAI211_X1 U16201 ( .C1(n14404), .C2(n14668), .A(n15016), .B(n14384), .ZN(
        n14588) );
  INV_X1 U16202 ( .A(n14385), .ZN(n14386) );
  OAI22_X1 U16203 ( .A1(n14588), .A2(n14433), .B1(n14544), .B2(n14386), .ZN(
        n14387) );
  OAI21_X1 U16204 ( .B1(n14388), .B2(n14387), .A(n14541), .ZN(n14391) );
  AOI22_X1 U16205 ( .A1(n14389), .A2(n14546), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15022), .ZN(n14390) );
  OAI211_X1 U16206 ( .C1(n14590), .C2(n14520), .A(n14391), .B(n14390), .ZN(
        P1_U3268) );
  OAI21_X1 U16207 ( .B1(n14393), .B2(n14394), .A(n14392), .ZN(n14596) );
  NAND2_X1 U16208 ( .A1(n14395), .A2(n14394), .ZN(n14396) );
  NAND3_X1 U16209 ( .A1(n14397), .A2(n15079), .A3(n14396), .ZN(n14401) );
  AOI22_X1 U16210 ( .A1(n14509), .A2(n14399), .B1(n15007), .B2(n14398), .ZN(
        n14400) );
  NAND2_X1 U16211 ( .A1(n14401), .A2(n14400), .ZN(n14402) );
  AOI21_X1 U16212 ( .B1(n14596), .B2(n15068), .A(n14402), .ZN(n14598) );
  NAND2_X1 U16213 ( .A1(n14419), .A2(n14593), .ZN(n14403) );
  NAND2_X1 U16214 ( .A1(n14403), .A2(n15016), .ZN(n14405) );
  OR2_X1 U16215 ( .A1(n14405), .A2(n14404), .ZN(n14594) );
  AOI22_X1 U16216 ( .A1(n15022), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14406), 
        .B2(n15013), .ZN(n14408) );
  NAND2_X1 U16217 ( .A1(n14593), .A2(n14546), .ZN(n14407) );
  OAI211_X1 U16218 ( .C1(n14594), .C2(n14537), .A(n14408), .B(n14407), .ZN(
        n14409) );
  AOI21_X1 U16219 ( .B1(n14596), .B2(n15019), .A(n14409), .ZN(n14410) );
  OAI21_X1 U16220 ( .B1(n14598), .B2(n15022), .A(n14410), .ZN(P1_U3269) );
  OAI21_X1 U16221 ( .B1(n14412), .B2(n14416), .A(n14411), .ZN(n14415) );
  INV_X1 U16222 ( .A(n14413), .ZN(n14414) );
  AOI21_X1 U16223 ( .B1(n14415), .B2(n15079), .A(n14414), .ZN(n14602) );
  OAI21_X1 U16224 ( .B1(n6475), .B2(n7628), .A(n14417), .ZN(n14603) );
  INV_X1 U16225 ( .A(n14603), .ZN(n14425) );
  INV_X1 U16226 ( .A(n14600), .ZN(n14423) );
  NAND2_X1 U16227 ( .A1(n14432), .A2(n14600), .ZN(n14418) );
  AND3_X1 U16228 ( .A1(n14419), .A2(n15016), .A3(n14418), .ZN(n14599) );
  NAND2_X1 U16229 ( .A1(n14599), .A2(n15018), .ZN(n14422) );
  AOI22_X1 U16230 ( .A1(n15022), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14420), 
        .B2(n15013), .ZN(n14421) );
  OAI211_X1 U16231 ( .C1(n14423), .C2(n15012), .A(n14422), .B(n14421), .ZN(
        n14424) );
  AOI21_X1 U16232 ( .B1(n14425), .B2(n14548), .A(n14424), .ZN(n14426) );
  OAI21_X1 U16233 ( .B1(n15022), .B2(n14602), .A(n14426), .ZN(P1_U3270) );
  XNOR2_X1 U16234 ( .A(n14428), .B(n14427), .ZN(n14610) );
  OAI21_X1 U16235 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14608) );
  INV_X1 U16236 ( .A(n14604), .ZN(n14435) );
  OAI211_X1 U16237 ( .C1(n14606), .C2(n7285), .A(n15016), .B(n14432), .ZN(
        n14605) );
  NOR2_X1 U16238 ( .A1(n14605), .A2(n14433), .ZN(n14434) );
  AOI211_X1 U16239 ( .C1(n15013), .C2(n14436), .A(n14435), .B(n14434), .ZN(
        n14438) );
  AOI22_X1 U16240 ( .A1(n6457), .A2(n14546), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15022), .ZN(n14437) );
  OAI21_X1 U16241 ( .B1(n14438), .B2(n15022), .A(n14437), .ZN(n14439) );
  AOI21_X1 U16242 ( .B1(n14548), .B2(n14608), .A(n14439), .ZN(n14440) );
  OAI21_X1 U16243 ( .B1(n14610), .B2(n14441), .A(n14440), .ZN(P1_U3271) );
  XOR2_X1 U16244 ( .A(n14448), .B(n14442), .Z(n14611) );
  AOI211_X1 U16245 ( .C1(n14443), .C2(n14462), .A(n14640), .B(n7285), .ZN(
        n14613) );
  INV_X1 U16246 ( .A(n14443), .ZN(n14675) );
  INV_X1 U16247 ( .A(n14444), .ZN(n14445) );
  AOI22_X1 U16248 ( .A1(n15022), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14445), 
        .B2(n15013), .ZN(n14446) );
  OAI21_X1 U16249 ( .B1(n14675), .B2(n15012), .A(n14446), .ZN(n14447) );
  AOI21_X1 U16250 ( .B1(n14613), .B2(n15018), .A(n14447), .ZN(n14452) );
  XNOR2_X1 U16251 ( .A(n14449), .B(n14448), .ZN(n14450) );
  NOR2_X1 U16252 ( .A1(n14450), .A2(n14936), .ZN(n14614) );
  OAI21_X1 U16253 ( .B1(n14614), .B2(n14612), .A(n14541), .ZN(n14451) );
  OAI211_X1 U16254 ( .C1(n14611), .C2(n14520), .A(n14452), .B(n14451), .ZN(
        P1_U3272) );
  INV_X1 U16255 ( .A(n14619), .ZN(n14456) );
  OAI211_X1 U16256 ( .C1(n14454), .C2(n14461), .A(n14453), .B(n15079), .ZN(
        n14620) );
  INV_X1 U16257 ( .A(n14620), .ZN(n14455) );
  AOI211_X1 U16258 ( .C1(n15013), .C2(n14457), .A(n14456), .B(n14455), .ZN(
        n14468) );
  INV_X1 U16259 ( .A(n14458), .ZN(n14459) );
  AOI21_X1 U16260 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(n14622) );
  OAI211_X1 U16261 ( .C1(n14463), .C2(n14679), .A(n15016), .B(n14462), .ZN(
        n14618) );
  AOI22_X1 U16262 ( .A1(n14464), .A2(n14546), .B1(n15022), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14465) );
  OAI21_X1 U16263 ( .B1(n14618), .B2(n14537), .A(n14465), .ZN(n14466) );
  AOI21_X1 U16264 ( .B1(n14622), .B2(n14548), .A(n14466), .ZN(n14467) );
  OAI21_X1 U16265 ( .B1(n14468), .B2(n15022), .A(n14467), .ZN(P1_U3273) );
  XNOR2_X1 U16266 ( .A(n14469), .B(n14473), .ZN(n14470) );
  OAI222_X1 U16267 ( .A1(n14525), .A2(n14472), .B1(n14527), .B2(n14471), .C1(
        n14470), .C2(n14936), .ZN(n14625) );
  INV_X1 U16268 ( .A(n14625), .ZN(n14483) );
  XNOR2_X1 U16269 ( .A(n14474), .B(n14473), .ZN(n14627) );
  AOI21_X1 U16270 ( .B1(n14475), .B2(n14493), .A(n14640), .ZN(n14477) );
  AND2_X1 U16271 ( .A1(n14477), .A2(n14476), .ZN(n14626) );
  NAND2_X1 U16272 ( .A1(n14626), .A2(n15018), .ZN(n14480) );
  AOI22_X1 U16273 ( .A1(n15022), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14478), 
        .B2(n15013), .ZN(n14479) );
  OAI211_X1 U16274 ( .C1(n14684), .C2(n15012), .A(n14480), .B(n14479), .ZN(
        n14481) );
  AOI21_X1 U16275 ( .B1(n14627), .B2(n14548), .A(n14481), .ZN(n14482) );
  OAI21_X1 U16276 ( .B1(n14483), .B2(n15022), .A(n14482), .ZN(P1_U3274) );
  XNOR2_X1 U16277 ( .A(n14485), .B(n14484), .ZN(n14631) );
  XNOR2_X1 U16278 ( .A(n14487), .B(n14486), .ZN(n14491) );
  AOI22_X1 U16279 ( .A1(n14489), .A2(n14509), .B1(n15007), .B2(n14488), .ZN(
        n14490) );
  OAI21_X1 U16280 ( .B1(n14491), .B2(n14936), .A(n14490), .ZN(n14492) );
  AOI21_X1 U16281 ( .B1(n14631), .B2(n15068), .A(n14492), .ZN(n14635) );
  INV_X1 U16282 ( .A(n14493), .ZN(n14494) );
  AOI211_X1 U16283 ( .C1(n14633), .C2(n6563), .A(n14640), .B(n14494), .ZN(
        n14632) );
  NAND2_X1 U16284 ( .A1(n14632), .A2(n15018), .ZN(n14498) );
  INV_X1 U16285 ( .A(n14495), .ZN(n14496) );
  AOI22_X1 U16286 ( .A1(n15022), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14496), 
        .B2(n15013), .ZN(n14497) );
  OAI211_X1 U16287 ( .C1(n7286), .C2(n15012), .A(n14498), .B(n14497), .ZN(
        n14499) );
  AOI21_X1 U16288 ( .B1(n15019), .B2(n14631), .A(n14499), .ZN(n14500) );
  OAI21_X1 U16289 ( .B1(n15022), .B2(n14635), .A(n14500), .ZN(P1_U3275) );
  XNOR2_X1 U16290 ( .A(n14502), .B(n14501), .ZN(n14645) );
  INV_X1 U16291 ( .A(n14503), .ZN(n14504) );
  AOI21_X1 U16292 ( .B1(n7420), .B2(n14505), .A(n14504), .ZN(n14643) );
  INV_X1 U16293 ( .A(n14531), .ZN(n14506) );
  INV_X1 U16294 ( .A(n14637), .ZN(n14512) );
  OAI21_X1 U16295 ( .B1(n14506), .B2(n14512), .A(n6563), .ZN(n14641) );
  AND2_X1 U16296 ( .A1(n14507), .A2(n15007), .ZN(n14508) );
  AOI21_X1 U16297 ( .B1(n14510), .B2(n14509), .A(n14508), .ZN(n14639) );
  OAI22_X1 U16298 ( .A1(n15022), .A2(n14639), .B1(n14511), .B2(n14544), .ZN(
        n14514) );
  NOR2_X1 U16299 ( .A1(n14512), .A2(n15012), .ZN(n14513) );
  AOI211_X1 U16300 ( .C1(n15022), .C2(P1_REG2_REG_17__SCAN_IN), .A(n14514), 
        .B(n14513), .ZN(n14515) );
  OAI21_X1 U16301 ( .B1(n14516), .B2(n14641), .A(n14515), .ZN(n14517) );
  AOI21_X1 U16302 ( .B1(n14643), .B2(n14518), .A(n14517), .ZN(n14519) );
  OAI21_X1 U16303 ( .B1(n14520), .B2(n14645), .A(n14519), .ZN(P1_U3276) );
  XNOR2_X1 U16304 ( .A(n14522), .B(n14521), .ZN(n14523) );
  OAI222_X1 U16305 ( .A1(n14527), .A2(n14526), .B1(n14525), .B2(n14524), .C1(
        n14523), .C2(n14936), .ZN(n14648) );
  INV_X1 U16306 ( .A(n14648), .ZN(n14540) );
  OAI21_X1 U16307 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n14650) );
  OAI211_X1 U16308 ( .C1(n14647), .C2(n6437), .A(n15016), .B(n14531), .ZN(
        n14646) );
  NAND2_X1 U16309 ( .A1(n15022), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14532) );
  OAI21_X1 U16310 ( .B1(n14544), .B2(n14533), .A(n14532), .ZN(n14534) );
  AOI21_X1 U16311 ( .B1(n14535), .B2(n14546), .A(n14534), .ZN(n14536) );
  OAI21_X1 U16312 ( .B1(n14646), .B2(n14537), .A(n14536), .ZN(n14538) );
  AOI21_X1 U16313 ( .B1(n14650), .B2(n14548), .A(n14538), .ZN(n14539) );
  OAI21_X1 U16314 ( .B1(n14540), .B2(n15022), .A(n14539), .ZN(P1_U3277) );
  NAND2_X1 U16315 ( .A1(n14542), .A2(n14541), .ZN(n14554) );
  NAND2_X1 U16316 ( .A1(n15022), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n14543) );
  OAI21_X1 U16317 ( .B1(n14544), .B2(n14934), .A(n14543), .ZN(n14545) );
  AOI21_X1 U16318 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n14553) );
  NAND2_X1 U16319 ( .A1(n14549), .A2(n14548), .ZN(n14552) );
  NAND2_X1 U16320 ( .A1(n14550), .A2(n15018), .ZN(n14551) );
  NAND4_X1 U16321 ( .A1(n14554), .A2(n14553), .A3(n14552), .A4(n14551), .ZN(
        P1_U3282) );
  INV_X1 U16322 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14557) );
  AOI21_X1 U16323 ( .B1(n14556), .B2(n15016), .A(n14555), .ZN(n14652) );
  MUX2_X1 U16324 ( .A(n14557), .B(n14652), .S(n15123), .Z(n14558) );
  OAI21_X1 U16325 ( .B1(n14654), .B2(n14630), .A(n14558), .ZN(P1_U3559) );
  INV_X1 U16326 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14561) );
  AND2_X1 U16327 ( .A1(n14560), .A2(n14559), .ZN(n14656) );
  MUX2_X1 U16328 ( .A(n14561), .B(n14656), .S(n9971), .Z(n14562) );
  OAI21_X1 U16329 ( .B1(n14659), .B2(n14630), .A(n14562), .ZN(P1_U3558) );
  OAI21_X1 U16330 ( .B1(n14564), .B2(n15072), .A(n14563), .ZN(n14566) );
  MUX2_X1 U16331 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14660), .S(n9971), .Z(
        P1_U3557) );
  AND2_X1 U16332 ( .A1(n14570), .A2(n14569), .ZN(n14573) );
  NAND2_X1 U16333 ( .A1(n14571), .A2(n15079), .ZN(n14572) );
  INV_X1 U16334 ( .A(n14575), .ZN(n14580) );
  AOI22_X1 U16335 ( .A1(n14577), .A2(n15016), .B1(n15062), .B2(n14576), .ZN(
        n14578) );
  OAI211_X1 U16336 ( .C1(n14580), .C2(n15064), .A(n14579), .B(n14578), .ZN(
        n14663) );
  MUX2_X1 U16337 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14663), .S(n15123), .Z(
        P1_U3555) );
  AOI211_X1 U16338 ( .C1(n15062), .C2(n14583), .A(n14582), .B(n14581), .ZN(
        n14586) );
  NAND2_X1 U16339 ( .A1(n14584), .A2(n15079), .ZN(n14585) );
  OAI211_X1 U16340 ( .C1(n14587), .C2(n15074), .A(n14586), .B(n14585), .ZN(
        n14664) );
  MUX2_X1 U16341 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14664), .S(n15123), .Z(
        P1_U3554) );
  OAI211_X1 U16342 ( .C1(n14590), .C2(n15074), .A(n14589), .B(n14588), .ZN(
        n14665) );
  MUX2_X1 U16343 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14665), .S(n15123), .Z(
        n14591) );
  INV_X1 U16344 ( .A(n14591), .ZN(n14592) );
  OAI21_X1 U16345 ( .B1(n14668), .B2(n14630), .A(n14592), .ZN(P1_U3553) );
  OAI21_X1 U16346 ( .B1(n6832), .B2(n15072), .A(n14594), .ZN(n14595) );
  AOI21_X1 U16347 ( .B1(n14596), .B2(n15098), .A(n14595), .ZN(n14597) );
  NAND2_X1 U16348 ( .A1(n14598), .A2(n14597), .ZN(n14669) );
  MUX2_X1 U16349 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14669), .S(n15123), .Z(
        P1_U3552) );
  AOI21_X1 U16350 ( .B1(n15062), .B2(n14600), .A(n14599), .ZN(n14601) );
  OAI211_X1 U16351 ( .C1(n14603), .C2(n15074), .A(n14602), .B(n14601), .ZN(
        n14670) );
  MUX2_X1 U16352 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14670), .S(n9971), .Z(
        P1_U3551) );
  OAI211_X1 U16353 ( .C1(n15072), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14607) );
  AOI21_X1 U16354 ( .B1(n14608), .B2(n15108), .A(n14607), .ZN(n14609) );
  OAI21_X1 U16355 ( .B1(n14936), .B2(n14610), .A(n14609), .ZN(n14671) );
  MUX2_X1 U16356 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14671), .S(n9971), .Z(
        P1_U3550) );
  NOR2_X1 U16357 ( .A1(n14611), .A2(n15074), .ZN(n14615) );
  NOR4_X1 U16358 ( .A1(n14615), .A2(n14614), .A3(n14613), .A4(n14612), .ZN(
        n14672) );
  MUX2_X1 U16359 ( .A(n14616), .B(n14672), .S(n9971), .Z(n14617) );
  OAI21_X1 U16360 ( .B1(n14675), .B2(n14630), .A(n14617), .ZN(P1_U3549) );
  NAND3_X1 U16361 ( .A1(n14620), .A2(n14619), .A3(n14618), .ZN(n14621) );
  AOI21_X1 U16362 ( .B1(n14622), .B2(n15108), .A(n14621), .ZN(n14676) );
  MUX2_X1 U16363 ( .A(n14623), .B(n14676), .S(n9971), .Z(n14624) );
  OAI21_X1 U16364 ( .B1(n14679), .B2(n14630), .A(n14624), .ZN(P1_U3548) );
  AOI211_X1 U16365 ( .C1(n15108), .C2(n14627), .A(n14626), .B(n14625), .ZN(
        n14680) );
  MUX2_X1 U16366 ( .A(n14628), .B(n14680), .S(n15123), .Z(n14629) );
  OAI21_X1 U16367 ( .B1(n14684), .B2(n14630), .A(n14629), .ZN(P1_U3547) );
  INV_X1 U16368 ( .A(n14631), .ZN(n14636) );
  AOI21_X1 U16369 ( .B1(n15062), .B2(n14633), .A(n14632), .ZN(n14634) );
  OAI211_X1 U16370 ( .C1(n15064), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14685) );
  MUX2_X1 U16371 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14685), .S(n9971), .Z(
        P1_U3546) );
  NAND2_X1 U16372 ( .A1(n14637), .A2(n15062), .ZN(n14638) );
  OAI211_X1 U16373 ( .C1(n14641), .C2(n14640), .A(n14639), .B(n14638), .ZN(
        n14642) );
  AOI21_X1 U16374 ( .B1(n14643), .B2(n15079), .A(n14642), .ZN(n14644) );
  OAI21_X1 U16375 ( .B1(n15074), .B2(n14645), .A(n14644), .ZN(n14686) );
  MUX2_X1 U16376 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14686), .S(n15123), .Z(
        P1_U3545) );
  OAI21_X1 U16377 ( .B1(n14647), .B2(n15072), .A(n14646), .ZN(n14649) );
  AOI211_X1 U16378 ( .C1(n15108), .C2(n14650), .A(n14649), .B(n14648), .ZN(
        n14651) );
  INV_X1 U16379 ( .A(n14651), .ZN(n14687) );
  MUX2_X1 U16380 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14687), .S(n15123), .Z(
        P1_U3544) );
  INV_X1 U16381 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15412) );
  MUX2_X1 U16382 ( .A(n15412), .B(n14652), .S(n15111), .Z(n14653) );
  OAI21_X1 U16383 ( .B1(n14654), .B2(n14683), .A(n14653), .ZN(P1_U3527) );
  INV_X1 U16384 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14657) );
  MUX2_X1 U16385 ( .A(n14657), .B(n14656), .S(n14655), .Z(n14658) );
  OAI21_X1 U16386 ( .B1(n14659), .B2(n14683), .A(n14658), .ZN(P1_U3526) );
  MUX2_X1 U16387 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14660), .S(n15111), .Z(
        P1_U3525) );
  MUX2_X1 U16388 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14663), .S(n15111), .Z(
        P1_U3523) );
  MUX2_X1 U16389 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14664), .S(n15111), .Z(
        P1_U3522) );
  MUX2_X1 U16390 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14665), .S(n15111), .Z(
        n14666) );
  INV_X1 U16391 ( .A(n14666), .ZN(n14667) );
  OAI21_X1 U16392 ( .B1(n14668), .B2(n14683), .A(n14667), .ZN(P1_U3521) );
  MUX2_X1 U16393 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14669), .S(n15111), .Z(
        P1_U3520) );
  MUX2_X1 U16394 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14670), .S(n15111), .Z(
        P1_U3519) );
  MUX2_X1 U16395 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14671), .S(n15111), .Z(
        P1_U3518) );
  INV_X1 U16396 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14673) );
  MUX2_X1 U16397 ( .A(n14673), .B(n14672), .S(n15111), .Z(n14674) );
  OAI21_X1 U16398 ( .B1(n14675), .B2(n14683), .A(n14674), .ZN(P1_U3517) );
  INV_X1 U16399 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14677) );
  MUX2_X1 U16400 ( .A(n14677), .B(n14676), .S(n15111), .Z(n14678) );
  OAI21_X1 U16401 ( .B1(n14679), .B2(n14683), .A(n14678), .ZN(P1_U3516) );
  INV_X1 U16402 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14681) );
  MUX2_X1 U16403 ( .A(n14681), .B(n14680), .S(n15111), .Z(n14682) );
  OAI21_X1 U16404 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(P1_U3515) );
  MUX2_X1 U16405 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14685), .S(n15111), .Z(
        P1_U3513) );
  MUX2_X1 U16406 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14686), .S(n15111), .Z(
        P1_U3510) );
  MUX2_X1 U16407 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14687), .S(n15111), .Z(
        P1_U3507) );
  NOR4_X1 U16408 ( .A1(n14688), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9306), .A4(
        P1_U3086), .ZN(n14689) );
  AOI21_X1 U16409 ( .B1(n14690), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14689), 
        .ZN(n14691) );
  OAI21_X1 U16410 ( .B1(n14692), .B2(n14707), .A(n14691), .ZN(P1_U3324) );
  OAI222_X1 U16411 ( .A1(n14701), .A2(n15339), .B1(n14707), .B2(n14694), .C1(
        n14693), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U16412 ( .A1(n14697), .A2(P1_U3086), .B1(n14707), .B2(n14696), 
        .C1(n14695), .C2(n14709), .ZN(P1_U3326) );
  OAI222_X1 U16413 ( .A1(P1_U3086), .A2(n14700), .B1(n14707), .B2(n14699), 
        .C1(n14698), .C2(n14701), .ZN(P1_U3327) );
  OAI222_X1 U16414 ( .A1(n9491), .A2(P1_U3086), .B1(n14707), .B2(n14703), .C1(
        n14702), .C2(n14701), .ZN(P1_U3328) );
  OAI222_X1 U16415 ( .A1(n14709), .A2(n14708), .B1(n14707), .B2(n14706), .C1(
        P1_U3086), .C2(n14705), .ZN(P1_U3329) );
  MUX2_X1 U16416 ( .A(n12072), .B(n14710), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16417 ( .A(n14711), .ZN(n14712) );
  MUX2_X1 U16418 ( .A(n14712), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16419 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14742) );
  XOR2_X1 U16420 ( .A(n14742), .B(n14713), .Z(n14753) );
  INV_X1 U16421 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14738) );
  INV_X1 U16422 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14714) );
  XNOR2_X1 U16423 ( .A(n14714), .B(n14736), .ZN(n14793) );
  XNOR2_X1 U16424 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14758) );
  XNOR2_X1 U16425 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14761) );
  NAND2_X1 U16426 ( .A1(n14761), .A2(n14762), .ZN(n14716) );
  NAND2_X1 U16427 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14717), .ZN(n14718) );
  NAND2_X1 U16428 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14719), .ZN(n14720) );
  NAND2_X1 U16429 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14721), .ZN(n14723) );
  NAND2_X1 U16430 ( .A1(n14726), .A2(n11147), .ZN(n14728) );
  XNOR2_X1 U16431 ( .A(n14726), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14781) );
  NAND2_X1 U16432 ( .A1(n14781), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14727) );
  NAND2_X1 U16433 ( .A1(n14728), .A2(n14727), .ZN(n14759) );
  NAND2_X1 U16434 ( .A1(n14758), .A2(n14759), .ZN(n14729) );
  XNOR2_X1 U16435 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14732), .ZN(n14786) );
  NOR2_X1 U16436 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14756), .ZN(n14734) );
  NAND2_X1 U16437 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14756), .ZN(n14733) );
  NAND2_X1 U16438 ( .A1(n14793), .A2(n14794), .ZN(n14735) );
  XOR2_X1 U16439 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14795) );
  AND2_X1 U16440 ( .A1(n14740), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14739) );
  NOR2_X1 U16441 ( .A1(n14753), .A2(n14752), .ZN(n14741) );
  AOI21_X1 U16442 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14742), .A(n14741), 
        .ZN(n14798) );
  NAND2_X1 U16443 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14743), .ZN(n14744) );
  INV_X1 U16444 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14997) );
  AOI22_X1 U16445 ( .A1(n14798), .A2(n14744), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n14997), .ZN(n14802) );
  OR2_X1 U16446 ( .A1(n14746), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14745) );
  AOI22_X1 U16447 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14746), .B1(n14802), 
        .B2(n14745), .ZN(n14748) );
  INV_X1 U16448 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14747) );
  NAND2_X1 U16449 ( .A1(n14748), .A2(n14747), .ZN(n14750) );
  XNOR2_X1 U16450 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14748), .ZN(n14804) );
  NAND2_X1 U16451 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14804), .ZN(n14749) );
  NAND2_X1 U16452 ( .A1(n14750), .A2(n14749), .ZN(n14827) );
  NOR2_X1 U16453 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14830), .ZN(n14751) );
  AOI21_X1 U16454 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14830), .A(n14751), 
        .ZN(n14828) );
  XNOR2_X1 U16455 ( .A(n14827), .B(n14828), .ZN(n14825) );
  INV_X1 U16456 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14822) );
  INV_X1 U16457 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14969) );
  XOR2_X1 U16458 ( .A(n14753), .B(n14752), .Z(n14961) );
  INV_X1 U16459 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14959) );
  XOR2_X1 U16460 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14754) );
  XNOR2_X1 U16461 ( .A(n14755), .B(n14754), .ZN(n14957) );
  INV_X1 U16462 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14949) );
  XNOR2_X1 U16463 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n14757) );
  XOR2_X1 U16464 ( .A(n14757), .B(n14756), .Z(n14792) );
  XOR2_X1 U16465 ( .A(n14759), .B(n14758), .Z(n14785) );
  XNOR2_X1 U16466 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14760), .ZN(n14771) );
  NOR2_X1 U16467 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14771), .ZN(n14773) );
  INV_X1 U16468 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14812) );
  XNOR2_X1 U16469 ( .A(n14762), .B(n14761), .ZN(n14810) );
  NAND2_X1 U16470 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14765), .ZN(n14766) );
  AOI21_X1 U16471 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14764), .A(n14763), .ZN(
        n15466) );
  INV_X1 U16472 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15465) );
  NOR2_X1 U16473 ( .A1(n15466), .A2(n15465), .ZN(n15474) );
  NAND2_X1 U16474 ( .A1(n14810), .A2(n14811), .ZN(n14767) );
  NOR2_X1 U16475 ( .A1(n14810), .A2(n14811), .ZN(n14809) );
  AOI21_X1 U16476 ( .B1(n14812), .B2(n14767), .A(n14809), .ZN(n15470) );
  XNOR2_X1 U16477 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14768), .ZN(n15471) );
  NOR2_X1 U16478 ( .A1(n15470), .A2(n15471), .ZN(n14770) );
  INV_X1 U16479 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14769) );
  NAND2_X1 U16480 ( .A1(n15470), .A2(n15471), .ZN(n15469) );
  OAI21_X1 U16481 ( .B1(n14770), .B2(n14769), .A(n15469), .ZN(n15463) );
  XNOR2_X1 U16482 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14771), .ZN(n15462) );
  NOR2_X1 U16483 ( .A1(n15463), .A2(n15462), .ZN(n14772) );
  XNOR2_X1 U16484 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14774), .ZN(n14775) );
  NAND2_X1 U16485 ( .A1(n14777), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14780) );
  XNOR2_X1 U16486 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14779) );
  XNOR2_X1 U16487 ( .A(n14779), .B(n14778), .ZN(n14814) );
  NAND2_X1 U16488 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14782), .ZN(n14783) );
  XOR2_X1 U16489 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14781), .Z(n15468) );
  XNOR2_X1 U16490 ( .A(n14787), .B(n14786), .ZN(n14789) );
  NAND2_X1 U16491 ( .A1(n14788), .A2(n14789), .ZN(n14790) );
  XOR2_X1 U16492 ( .A(n14794), .B(n14793), .Z(n14948) );
  XNOR2_X1 U16493 ( .A(n14796), .B(n14795), .ZN(n14952) );
  XNOR2_X1 U16494 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14799) );
  XOR2_X1 U16495 ( .A(n14799), .B(n14798), .Z(n14800) );
  XOR2_X1 U16496 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .Z(n14801) );
  XNOR2_X1 U16497 ( .A(n14802), .B(n14801), .ZN(n14968) );
  NAND2_X1 U16498 ( .A1(n14967), .A2(n14968), .ZN(n14803) );
  NOR2_X1 U16499 ( .A1(n14967), .A2(n14968), .ZN(n14966) );
  XOR2_X1 U16500 ( .A(n14805), .B(n14804), .Z(n14820) );
  NAND2_X1 U16501 ( .A1(n14821), .A2(n14820), .ZN(n14806) );
  NOR2_X1 U16502 ( .A1(n14821), .A2(n14820), .ZN(n14819) );
  XNOR2_X1 U16503 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14824), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16504 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14807) );
  OAI21_X1 U16505 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14807), 
        .ZN(U28) );
  AOI21_X1 U16506 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14808) );
  OAI21_X1 U16507 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14808), 
        .ZN(U29) );
  AOI21_X1 U16508 ( .B1(n14811), .B2(n14810), .A(n14809), .ZN(n14813) );
  XNOR2_X1 U16509 ( .A(n14813), .B(n14812), .ZN(SUB_1596_U61) );
  XOR2_X1 U16510 ( .A(n14815), .B(n14814), .Z(SUB_1596_U57) );
  XNOR2_X1 U16511 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14816), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16512 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14817), .Z(SUB_1596_U54) );
  XNOR2_X1 U16513 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14818), .ZN(SUB_1596_U70)
         );
  AOI21_X1 U16514 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14823) );
  XNOR2_X1 U16515 ( .A(n14823), .B(n14822), .ZN(SUB_1596_U63) );
  NAND2_X1 U16516 ( .A1(n14828), .A2(n14827), .ZN(n14829) );
  OAI21_X1 U16517 ( .B1(n14830), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14829), 
        .ZN(n14833) );
  XNOR2_X1 U16518 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n14831) );
  XNOR2_X1 U16519 ( .A(n14831), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14832) );
  XNOR2_X1 U16520 ( .A(n14833), .B(n14832), .ZN(n14834) );
  XNOR2_X1 U16521 ( .A(n14835), .B(n14834), .ZN(SUB_1596_U4) );
  XNOR2_X1 U16522 ( .A(n14836), .B(n14844), .ZN(n14837) );
  NAND2_X1 U16523 ( .A1(n14837), .A2(n15218), .ZN(n14840) );
  AOI22_X1 U16524 ( .A1(n15212), .A2(n15197), .B1(n14838), .B2(n15215), .ZN(
        n14839) );
  NAND2_X1 U16525 ( .A1(n14840), .A2(n14839), .ZN(n14867) );
  AOI21_X1 U16526 ( .B1(n15244), .B2(n14841), .A(n14867), .ZN(n14849) );
  NAND2_X1 U16527 ( .A1(n14851), .A2(n14850), .ZN(n14843) );
  NAND2_X1 U16528 ( .A1(n14843), .A2(n14842), .ZN(n14845) );
  XNOR2_X1 U16529 ( .A(n14845), .B(n14844), .ZN(n14868) );
  NOR2_X1 U16530 ( .A1(n14846), .A2(n15281), .ZN(n14866) );
  AOI22_X1 U16531 ( .A1(n14868), .A2(n14847), .B1(n15228), .B2(n14866), .ZN(
        n14848) );
  OAI221_X1 U16532 ( .B1(n15250), .B2(n14849), .C1(n15248), .C2(n15329), .A(
        n14848), .ZN(P3_U3221) );
  XNOR2_X1 U16533 ( .A(n14851), .B(n14850), .ZN(n14875) );
  XNOR2_X1 U16534 ( .A(n14853), .B(n14852), .ZN(n14855) );
  OAI222_X1 U16535 ( .A1(n14859), .A2(n14858), .B1(n14857), .B2(n14856), .C1(
        n14855), .C2(n14854), .ZN(n14872) );
  AOI21_X1 U16536 ( .B1(n14875), .B2(n14860), .A(n14872), .ZN(n14865) );
  AND2_X1 U16537 ( .A1(n14861), .A2(n15287), .ZN(n14873) );
  NOR2_X1 U16538 ( .A1(n15234), .A2(n14862), .ZN(n14863) );
  AOI21_X1 U16539 ( .B1(n15228), .B2(n14873), .A(n14863), .ZN(n14864) );
  OAI221_X1 U16540 ( .B1(n15250), .B2(n14865), .C1(n15248), .C2(n7880), .A(
        n14864), .ZN(P3_U3222) );
  NOR2_X1 U16541 ( .A1(n14867), .A2(n14866), .ZN(n14870) );
  NAND2_X1 U16542 ( .A1(n14868), .A2(n14874), .ZN(n14869) );
  AND2_X1 U16543 ( .A1(n14870), .A2(n14869), .ZN(n14876) );
  AOI22_X1 U16544 ( .A1(n15308), .A2(n14876), .B1(n14871), .B2(n15306), .ZN(
        P3_U3471) );
  AOI211_X1 U16545 ( .C1(n14875), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14878) );
  AOI22_X1 U16546 ( .A1(n15308), .A2(n14878), .B1(n7879), .B2(n15306), .ZN(
        P3_U3470) );
  INV_X1 U16547 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14877) );
  AOI22_X1 U16548 ( .A1(n15295), .A2(n14877), .B1(n14876), .B2(n15293), .ZN(
        P3_U3426) );
  INV_X1 U16549 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14879) );
  AOI22_X1 U16550 ( .A1(n15295), .A2(n14879), .B1(n14878), .B2(n15293), .ZN(
        P3_U3423) );
  OAI21_X1 U16551 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14884) );
  AOI222_X1 U16552 ( .A1(n9631), .A2(n14887), .B1(n14886), .B2(n14885), .C1(
        n14884), .C2(n14883), .ZN(n14889) );
  OAI211_X1 U16553 ( .C1(n14891), .C2(n14890), .A(n14889), .B(n14888), .ZN(
        P2_U3187) );
  AND2_X1 U16554 ( .A1(n14893), .A2(n14892), .ZN(n14896) );
  OAI21_X1 U16555 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14901) );
  AOI22_X1 U16556 ( .A1(n14925), .A2(n14898), .B1(n14923), .B2(n14897), .ZN(
        n14899) );
  OAI21_X1 U16557 ( .B1(n14940), .B2(n14927), .A(n14899), .ZN(n14900) );
  AOI21_X1 U16558 ( .B1(n14901), .B2(n14930), .A(n14900), .ZN(n14903) );
  OAI211_X1 U16559 ( .C1(n14935), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        P1_U3215) );
  NAND2_X1 U16560 ( .A1(n14905), .A2(n15062), .ZN(n15103) );
  OAI211_X1 U16561 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14930), .ZN(
        n14912) );
  AOI22_X1 U16562 ( .A1(n14925), .A2(n14910), .B1(n14923), .B2(n14909), .ZN(
        n14911) );
  OAI211_X1 U16563 ( .C1(n14913), .C2(n15103), .A(n14912), .B(n14911), .ZN(
        n14914) );
  INV_X1 U16564 ( .A(n14914), .ZN(n14916) );
  OAI211_X1 U16565 ( .C1(n14935), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        P1_U3217) );
  AND2_X1 U16566 ( .A1(n14906), .A2(n14918), .ZN(n14921) );
  OAI21_X1 U16567 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14931) );
  AOI22_X1 U16568 ( .A1(n14925), .A2(n14924), .B1(n14923), .B2(n14922), .ZN(
        n14926) );
  OAI21_X1 U16569 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n14929) );
  AOI21_X1 U16570 ( .B1(n14931), .B2(n14930), .A(n14929), .ZN(n14933) );
  OAI211_X1 U16571 ( .C1(n14935), .C2(n14934), .A(n14933), .B(n14932), .ZN(
        P1_U3236) );
  NOR2_X1 U16572 ( .A1(n14937), .A2(n14936), .ZN(n14942) );
  OAI211_X1 U16573 ( .C1(n14940), .C2(n15072), .A(n14939), .B(n14938), .ZN(
        n14941) );
  AOI211_X1 U16574 ( .C1(n14943), .C2(n15108), .A(n14942), .B(n14941), .ZN(
        n14945) );
  AOI22_X1 U16575 ( .A1(n15123), .A2(n14945), .B1(n10148), .B2(n15120), .ZN(
        P1_U3542) );
  INV_X1 U16576 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U16577 ( .A1(n15111), .A2(n14945), .B1(n14944), .B2(n15109), .ZN(
        P1_U3501) );
  AOI21_X1 U16578 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n14950) );
  XNOR2_X1 U16579 ( .A(n14950), .B(n14949), .ZN(SUB_1596_U69) );
  AOI21_X1 U16580 ( .B1(n14953), .B2(n14952), .A(n14951), .ZN(n14955) );
  XNOR2_X1 U16581 ( .A(n14955), .B(n14954), .ZN(SUB_1596_U68) );
  AOI21_X1 U16582 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n14960) );
  XNOR2_X1 U16583 ( .A(n14960), .B(n14959), .ZN(SUB_1596_U67) );
  AOI21_X1 U16584 ( .B1(n14962), .B2(n14961), .A(n6575), .ZN(n14963) );
  XOR2_X1 U16585 ( .A(n14963), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16586 ( .A1(n14964), .A2(n6567), .ZN(n14965) );
  XOR2_X1 U16587 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14965), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16588 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n14970) );
  XNOR2_X1 U16589 ( .A(n14970), .B(n14969), .ZN(SUB_1596_U64) );
  AND2_X1 U16590 ( .A1(n9491), .A2(n9735), .ZN(n14973) );
  NOR2_X1 U16591 ( .A1(n14971), .A2(n14973), .ZN(n14972) );
  MUX2_X1 U16592 ( .A(n14973), .B(n14972), .S(P1_IR_REG_0__SCAN_IN), .Z(n14976) );
  INV_X1 U16593 ( .A(n14974), .ZN(n14975) );
  OR2_X1 U16594 ( .A1(n14976), .A2(n14975), .ZN(n14979) );
  AOI22_X1 U16595 ( .A1(n14977), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14978) );
  OAI21_X1 U16596 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(P1_U3243) );
  AOI21_X1 U16597 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14982), .A(n14981), 
        .ZN(n14984) );
  OR2_X1 U16598 ( .A1(n14984), .A2(n14983), .ZN(n14990) );
  AOI21_X1 U16599 ( .B1(n14986), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14985), 
        .ZN(n14988) );
  OR2_X1 U16600 ( .A1(n14988), .A2(n14987), .ZN(n14989) );
  OAI211_X1 U16601 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n14989), .ZN(
        n14993) );
  INV_X1 U16602 ( .A(n14993), .ZN(n14995) );
  OAI211_X1 U16603 ( .C1(n14997), .C2(n14996), .A(n14995), .B(n14994), .ZN(
        P1_U3258) );
  XNOR2_X1 U16604 ( .A(n14998), .B(n15003), .ZN(n15057) );
  NOR2_X1 U16605 ( .A1(n14999), .A2(n15053), .ZN(n15000) );
  NOR2_X1 U16606 ( .A1(n15001), .A2(n15000), .ZN(n15017) );
  XNOR2_X1 U16607 ( .A(n15017), .B(n15002), .ZN(n15005) );
  NOR2_X1 U16608 ( .A1(n15003), .A2(n15007), .ZN(n15004) );
  MUX2_X1 U16609 ( .A(n15005), .B(n15004), .S(n15006), .Z(n15009) );
  AOI21_X1 U16610 ( .B1(n15007), .B2(n15006), .A(n15079), .ZN(n15008) );
  NOR2_X1 U16611 ( .A1(n15009), .A2(n15008), .ZN(n15010) );
  AOI211_X1 U16612 ( .C1(n15068), .C2(n15057), .A(n15011), .B(n15010), .ZN(
        n15054) );
  OR2_X1 U16613 ( .A1(n15012), .A2(n15053), .ZN(n15015) );
  AOI22_X1 U16614 ( .A1(n15022), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n15013), .ZN(n15014) );
  AND2_X1 U16615 ( .A1(n15015), .A2(n15014), .ZN(n15021) );
  AND2_X1 U16616 ( .A1(n15017), .A2(n15016), .ZN(n15051) );
  AOI22_X1 U16617 ( .A1(n15019), .A2(n15057), .B1(n15018), .B2(n15051), .ZN(
        n15020) );
  OAI211_X1 U16618 ( .C1(n15022), .C2(n15054), .A(n15021), .B(n15020), .ZN(
        P1_U3292) );
  INV_X1 U16619 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15317) );
  NOR2_X1 U16620 ( .A1(n15050), .A2(n15317), .ZN(P1_U3294) );
  INV_X1 U16621 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15023) );
  NOR2_X1 U16622 ( .A1(n15050), .A2(n15023), .ZN(P1_U3295) );
  INV_X1 U16623 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15024) );
  NOR2_X1 U16624 ( .A1(n15050), .A2(n15024), .ZN(P1_U3296) );
  INV_X1 U16625 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15025) );
  NOR2_X1 U16626 ( .A1(n15050), .A2(n15025), .ZN(P1_U3297) );
  INV_X1 U16627 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15026) );
  NOR2_X1 U16628 ( .A1(n15050), .A2(n15026), .ZN(P1_U3298) );
  INV_X1 U16629 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15027) );
  NOR2_X1 U16630 ( .A1(n15050), .A2(n15027), .ZN(P1_U3299) );
  INV_X1 U16631 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15028) );
  NOR2_X1 U16632 ( .A1(n15050), .A2(n15028), .ZN(P1_U3300) );
  INV_X1 U16633 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15029) );
  NOR2_X1 U16634 ( .A1(n15050), .A2(n15029), .ZN(P1_U3301) );
  INV_X1 U16635 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15030) );
  NOR2_X1 U16636 ( .A1(n15050), .A2(n15030), .ZN(P1_U3302) );
  INV_X1 U16637 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15031) );
  NOR2_X1 U16638 ( .A1(n15050), .A2(n15031), .ZN(P1_U3303) );
  INV_X1 U16639 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15032) );
  NOR2_X1 U16640 ( .A1(n15050), .A2(n15032), .ZN(P1_U3304) );
  INV_X1 U16641 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15033) );
  NOR2_X1 U16642 ( .A1(n15050), .A2(n15033), .ZN(P1_U3305) );
  INV_X1 U16643 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15034) );
  NOR2_X1 U16644 ( .A1(n15050), .A2(n15034), .ZN(P1_U3306) );
  INV_X1 U16645 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15035) );
  NOR2_X1 U16646 ( .A1(n15050), .A2(n15035), .ZN(P1_U3307) );
  INV_X1 U16647 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15036) );
  NOR2_X1 U16648 ( .A1(n15050), .A2(n15036), .ZN(P1_U3308) );
  INV_X1 U16649 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15037) );
  NOR2_X1 U16650 ( .A1(n15050), .A2(n15037), .ZN(P1_U3309) );
  INV_X1 U16651 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15038) );
  NOR2_X1 U16652 ( .A1(n15050), .A2(n15038), .ZN(P1_U3310) );
  INV_X1 U16653 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15039) );
  NOR2_X1 U16654 ( .A1(n15050), .A2(n15039), .ZN(P1_U3311) );
  INV_X1 U16655 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15352) );
  NOR2_X1 U16656 ( .A1(n15050), .A2(n15352), .ZN(P1_U3312) );
  INV_X1 U16657 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15370) );
  NOR2_X1 U16658 ( .A1(n15050), .A2(n15370), .ZN(P1_U3313) );
  INV_X1 U16659 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15040) );
  NOR2_X1 U16660 ( .A1(n15050), .A2(n15040), .ZN(P1_U3314) );
  INV_X1 U16661 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15041) );
  NOR2_X1 U16662 ( .A1(n15050), .A2(n15041), .ZN(P1_U3315) );
  INV_X1 U16663 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15042) );
  NOR2_X1 U16664 ( .A1(n15050), .A2(n15042), .ZN(P1_U3316) );
  INV_X1 U16665 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15043) );
  NOR2_X1 U16666 ( .A1(n15050), .A2(n15043), .ZN(P1_U3317) );
  INV_X1 U16667 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15044) );
  NOR2_X1 U16668 ( .A1(n15050), .A2(n15044), .ZN(P1_U3318) );
  INV_X1 U16669 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15045) );
  NOR2_X1 U16670 ( .A1(n15050), .A2(n15045), .ZN(P1_U3319) );
  INV_X1 U16671 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15046) );
  NOR2_X1 U16672 ( .A1(n15050), .A2(n15046), .ZN(P1_U3320) );
  INV_X1 U16673 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15047) );
  NOR2_X1 U16674 ( .A1(n15050), .A2(n15047), .ZN(P1_U3321) );
  INV_X1 U16675 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U16676 ( .A1(n15050), .A2(n15048), .ZN(P1_U3322) );
  INV_X1 U16677 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15049) );
  NOR2_X1 U16678 ( .A1(n15050), .A2(n15049), .ZN(P1_U3323) );
  INV_X1 U16679 ( .A(n15051), .ZN(n15052) );
  OAI21_X1 U16680 ( .B1(n15053), .B2(n15072), .A(n15052), .ZN(n15056) );
  INV_X1 U16681 ( .A(n15054), .ZN(n15055) );
  AOI211_X1 U16682 ( .C1(n15098), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15113) );
  INV_X1 U16683 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16684 ( .A1(n15111), .A2(n15113), .B1(n15058), .B2(n15109), .ZN(
        P1_U3462) );
  INV_X1 U16685 ( .A(n15065), .ZN(n15067) );
  AOI211_X1 U16686 ( .C1(n15062), .C2(n15061), .A(n15060), .B(n15059), .ZN(
        n15063) );
  OAI21_X1 U16687 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15066) );
  AOI21_X1 U16688 ( .B1(n15068), .B2(n15067), .A(n15066), .ZN(n15114) );
  INV_X1 U16689 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U16690 ( .A1(n15111), .A2(n15114), .B1(n15069), .B2(n15109), .ZN(
        P1_U3468) );
  OAI211_X1 U16691 ( .C1(n15073), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        n15077) );
  NOR2_X1 U16692 ( .A1(n15075), .A2(n15074), .ZN(n15076) );
  AOI211_X1 U16693 ( .C1(n15079), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15115) );
  INV_X1 U16694 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U16695 ( .A1(n15111), .A2(n15115), .B1(n15080), .B2(n15109), .ZN(
        P1_U3471) );
  INV_X1 U16696 ( .A(n15081), .ZN(n15083) );
  NAND3_X1 U16697 ( .A1(n15084), .A2(n15083), .A3(n15082), .ZN(n15086) );
  AOI211_X1 U16698 ( .C1(n15108), .C2(n15087), .A(n15086), .B(n15085), .ZN(
        n15116) );
  INV_X1 U16699 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U16700 ( .A1(n15111), .A2(n15116), .B1(n15088), .B2(n15109), .ZN(
        P1_U3480) );
  NAND2_X1 U16701 ( .A1(n15090), .A2(n15089), .ZN(n15092) );
  AOI211_X1 U16702 ( .C1(n15108), .C2(n15093), .A(n15092), .B(n15091), .ZN(
        n15117) );
  INV_X1 U16703 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U16704 ( .A1(n15111), .A2(n15117), .B1(n15094), .B2(n15109), .ZN(
        P1_U3483) );
  INV_X1 U16705 ( .A(n15095), .ZN(n15097) );
  AOI211_X1 U16706 ( .C1(n15099), .C2(n15098), .A(n15097), .B(n15096), .ZN(
        n15100) );
  AND2_X1 U16707 ( .A1(n15101), .A2(n15100), .ZN(n15119) );
  INV_X1 U16708 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U16709 ( .A1(n15111), .A2(n15119), .B1(n15102), .B2(n15109), .ZN(
        P1_U3486) );
  NAND3_X1 U16710 ( .A1(n15105), .A2(n15104), .A3(n15103), .ZN(n15106) );
  AOI21_X1 U16711 ( .B1(n15108), .B2(n15107), .A(n15106), .ZN(n15122) );
  INV_X1 U16712 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U16713 ( .A1(n15111), .A2(n15122), .B1(n15110), .B2(n15109), .ZN(
        P1_U3489) );
  AOI22_X1 U16714 ( .A1(n15123), .A2(n15113), .B1(n15112), .B2(n15120), .ZN(
        P1_U3529) );
  AOI22_X1 U16715 ( .A1(n15123), .A2(n15114), .B1(n9479), .B2(n15120), .ZN(
        P1_U3531) );
  AOI22_X1 U16716 ( .A1(n15123), .A2(n15115), .B1(n9482), .B2(n15120), .ZN(
        P1_U3532) );
  AOI22_X1 U16717 ( .A1(n15123), .A2(n15116), .B1(n9508), .B2(n15120), .ZN(
        P1_U3535) );
  AOI22_X1 U16718 ( .A1(n9971), .A2(n15117), .B1(n9512), .B2(n15120), .ZN(
        P1_U3536) );
  AOI22_X1 U16719 ( .A1(n9971), .A2(n15119), .B1(n15118), .B2(n15120), .ZN(
        P1_U3537) );
  AOI22_X1 U16720 ( .A1(n15123), .A2(n15122), .B1(n15121), .B2(n15120), .ZN(
        P1_U3538) );
  NOR2_X1 U16721 ( .A1(n15154), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16722 ( .A1(n15155), .A2(n15124), .ZN(n15126) );
  OAI211_X1 U16723 ( .C1(n15127), .C2(n7106), .A(n15126), .B(n15125), .ZN(
        n15128) );
  INV_X1 U16724 ( .A(n15128), .ZN(n15139) );
  AOI21_X1 U16725 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n15133) );
  NAND2_X1 U16726 ( .A1(n15133), .A2(n15132), .ZN(n15138) );
  OAI211_X1 U16727 ( .C1(n15136), .C2(n15135), .A(n15161), .B(n15134), .ZN(
        n15137) );
  NAND3_X1 U16728 ( .A1(n15139), .A2(n15138), .A3(n15137), .ZN(P2_U3221) );
  INV_X1 U16729 ( .A(n15140), .ZN(n15141) );
  OAI21_X1 U16730 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n15144) );
  AOI21_X1 U16731 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n15154), .A(n15144), 
        .ZN(n15153) );
  OAI211_X1 U16732 ( .C1(n15147), .C2(n15146), .A(n15145), .B(n15158), .ZN(
        n15152) );
  OAI211_X1 U16733 ( .C1(n15150), .C2(n15149), .A(n15148), .B(n15161), .ZN(
        n15151) );
  NAND3_X1 U16734 ( .A1(n15153), .A2(n15152), .A3(n15151), .ZN(P2_U3227) );
  AOI22_X1 U16735 ( .A1(n15154), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15166) );
  NAND2_X1 U16736 ( .A1(n15156), .A2(n15155), .ZN(n15165) );
  OAI211_X1 U16737 ( .C1(n15159), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15158), 
        .B(n15157), .ZN(n15164) );
  OAI211_X1 U16738 ( .C1(n15162), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15161), 
        .B(n15160), .ZN(n15163) );
  NAND4_X1 U16739 ( .A1(n15166), .A2(n15165), .A3(n15164), .A4(n15163), .ZN(
        P2_U3229) );
  INV_X1 U16740 ( .A(n15168), .ZN(n15169) );
  AND2_X1 U16741 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15169), .ZN(P2_U3266) );
  AND2_X1 U16742 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15169), .ZN(P2_U3267) );
  AND2_X1 U16743 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15169), .ZN(P2_U3268) );
  AND2_X1 U16744 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15169), .ZN(P2_U3269) );
  AND2_X1 U16745 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15169), .ZN(P2_U3270) );
  AND2_X1 U16746 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15169), .ZN(P2_U3271) );
  AND2_X1 U16747 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15169), .ZN(P2_U3272) );
  INV_X1 U16748 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15410) );
  NOR2_X1 U16749 ( .A1(n15168), .A2(n15410), .ZN(P2_U3273) );
  AND2_X1 U16750 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15169), .ZN(P2_U3274) );
  AND2_X1 U16751 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15169), .ZN(P2_U3275) );
  AND2_X1 U16752 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15169), .ZN(P2_U3276) );
  AND2_X1 U16753 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15169), .ZN(P2_U3277) );
  AND2_X1 U16754 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15169), .ZN(P2_U3278) );
  AND2_X1 U16755 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15169), .ZN(P2_U3279) );
  AND2_X1 U16756 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15169), .ZN(P2_U3280) );
  INV_X1 U16757 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15367) );
  NOR2_X1 U16758 ( .A1(n15168), .A2(n15367), .ZN(P2_U3281) );
  AND2_X1 U16759 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15169), .ZN(P2_U3282) );
  AND2_X1 U16760 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15169), .ZN(P2_U3283) );
  INV_X1 U16761 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15310) );
  NOR2_X1 U16762 ( .A1(n15168), .A2(n15310), .ZN(P2_U3284) );
  AND2_X1 U16763 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15169), .ZN(P2_U3285) );
  AND2_X1 U16764 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15169), .ZN(P2_U3286) );
  AND2_X1 U16765 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15169), .ZN(P2_U3287) );
  AND2_X1 U16766 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15169), .ZN(P2_U3288) );
  AND2_X1 U16767 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15169), .ZN(P2_U3289) );
  AND2_X1 U16768 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15169), .ZN(P2_U3290) );
  AND2_X1 U16769 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15169), .ZN(P2_U3291) );
  AND2_X1 U16770 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15169), .ZN(P2_U3292) );
  AND2_X1 U16771 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15169), .ZN(P2_U3293) );
  AND2_X1 U16772 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15169), .ZN(P2_U3294) );
  AND2_X1 U16773 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15169), .ZN(P2_U3295) );
  NOR2_X1 U16774 ( .A1(n15170), .A2(n15173), .ZN(n15171) );
  AOI21_X1 U16775 ( .B1(n15173), .B2(n15172), .A(n15171), .ZN(P2_U3416) );
  AOI22_X1 U16776 ( .A1(n15176), .A2(n15175), .B1(n15174), .B2(n15173), .ZN(
        P2_U3417) );
  AOI21_X1 U16777 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(n15180) );
  OAI211_X1 U16778 ( .C1(n15183), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15184) );
  INV_X1 U16779 ( .A(n15184), .ZN(n15189) );
  INV_X1 U16780 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U16781 ( .A1(n15187), .A2(n15189), .B1(n15186), .B2(n15185), .ZN(
        P2_U3451) );
  AOI22_X1 U16782 ( .A1(n15190), .A2(n15189), .B1(n9538), .B2(n15188), .ZN(
        P2_U3506) );
  NOR2_X1 U16783 ( .A1(P3_U3897), .A2(n15191), .ZN(P3_U3150) );
  XNOR2_X1 U16784 ( .A(n15192), .B(n15194), .ZN(n15290) );
  INV_X1 U16785 ( .A(n15290), .ZN(n15203) );
  OAI211_X1 U16786 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n15218), .ZN(
        n15199) );
  AOI22_X1 U16787 ( .A1(n15215), .A2(n15197), .B1(n15196), .B2(n15212), .ZN(
        n15198) );
  NAND2_X1 U16788 ( .A1(n15199), .A2(n15198), .ZN(n15200) );
  AOI21_X1 U16789 ( .B1(n15290), .B2(n15201), .A(n15200), .ZN(n15292) );
  OAI21_X1 U16790 ( .B1(n15203), .B2(n15202), .A(n15292), .ZN(n15208) );
  OAI22_X1 U16791 ( .A1(n15206), .A2(n15205), .B1(n15204), .B2(n15248), .ZN(
        n15207) );
  AOI21_X1 U16792 ( .B1(n15208), .B2(n15248), .A(n15207), .ZN(n15209) );
  OAI21_X1 U16793 ( .B1(n15210), .B2(n15234), .A(n15209), .ZN(P3_U3223) );
  XNOR2_X1 U16794 ( .A(n15211), .B(n11041), .ZN(n15224) );
  INV_X1 U16795 ( .A(n15224), .ZN(n15269) );
  AOI22_X1 U16796 ( .A1(n15215), .A2(n15214), .B1(n15213), .B2(n15212), .ZN(
        n15222) );
  AND2_X1 U16797 ( .A1(n15217), .A2(n15216), .ZN(n15220) );
  OAI211_X1 U16798 ( .C1(n15220), .C2(n11041), .A(n15219), .B(n15218), .ZN(
        n15221) );
  OAI211_X1 U16799 ( .C1(n15224), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15267) );
  AOI21_X1 U16800 ( .B1(n15238), .B2(n15269), .A(n15267), .ZN(n15231) );
  NOR2_X1 U16801 ( .A1(n15225), .A2(n15281), .ZN(n15268) );
  NOR2_X1 U16802 ( .A1(n15234), .A2(n15226), .ZN(n15227) );
  AOI21_X1 U16803 ( .B1(n15228), .B2(n15268), .A(n15227), .ZN(n15229) );
  OAI221_X1 U16804 ( .B1(n15250), .B2(n15231), .C1(n15248), .C2(n15230), .A(
        n15229), .ZN(P3_U3227) );
  OAI22_X1 U16805 ( .A1(n15234), .A2(n10585), .B1(n15233), .B2(n15232), .ZN(
        n15236) );
  AOI211_X1 U16806 ( .C1(n15238), .C2(n15237), .A(n15236), .B(n15235), .ZN(
        n15239) );
  AOI22_X1 U16807 ( .A1(n15250), .A2(n11119), .B1(n15239), .B2(n15248), .ZN(
        P3_U3231) );
  INV_X1 U16808 ( .A(n15240), .ZN(n15241) );
  AOI21_X1 U16809 ( .B1(n15243), .B2(n15242), .A(n15241), .ZN(n15249) );
  AOI22_X1 U16810 ( .A1(n15246), .A2(n15245), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15244), .ZN(n15247) );
  OAI221_X1 U16811 ( .B1(n15250), .B2(n15249), .C1(n15248), .C2(n11079), .A(
        n15247), .ZN(P3_U3232) );
  AOI22_X1 U16812 ( .A1(n15295), .A2(n7705), .B1(n15251), .B2(n15293), .ZN(
        P3_U3393) );
  AOI22_X1 U16813 ( .A1(n15295), .A2(n7716), .B1(n15252), .B2(n15293), .ZN(
        P3_U3396) );
  INV_X1 U16814 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15257) );
  INV_X1 U16815 ( .A(n15253), .ZN(n15255) );
  AOI211_X1 U16816 ( .C1(n15256), .C2(n15289), .A(n15255), .B(n15254), .ZN(
        n15296) );
  AOI22_X1 U16817 ( .A1(n15295), .A2(n15257), .B1(n15296), .B2(n15293), .ZN(
        P3_U3399) );
  INV_X1 U16818 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15262) );
  INV_X1 U16819 ( .A(n15258), .ZN(n15259) );
  AOI211_X1 U16820 ( .C1(n15261), .C2(n15289), .A(n15260), .B(n15259), .ZN(
        n15298) );
  AOI22_X1 U16821 ( .A1(n15295), .A2(n15262), .B1(n15298), .B2(n15293), .ZN(
        P3_U3402) );
  INV_X1 U16822 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15266) );
  AOI211_X1 U16823 ( .C1(n15265), .C2(n15289), .A(n15264), .B(n15263), .ZN(
        n15299) );
  AOI22_X1 U16824 ( .A1(n15295), .A2(n15266), .B1(n15299), .B2(n15293), .ZN(
        P3_U3405) );
  INV_X1 U16825 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15270) );
  AOI211_X1 U16826 ( .C1(n15269), .C2(n15289), .A(n15268), .B(n15267), .ZN(
        n15301) );
  AOI22_X1 U16827 ( .A1(n15295), .A2(n15270), .B1(n15301), .B2(n15293), .ZN(
        P3_U3408) );
  INV_X1 U16828 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15275) );
  AOI21_X1 U16829 ( .B1(n15272), .B2(n15289), .A(n15271), .ZN(n15273) );
  AOI22_X1 U16830 ( .A1(n15295), .A2(n15275), .B1(n15302), .B2(n15293), .ZN(
        P3_U3411) );
  AOI21_X1 U16831 ( .B1(n15277), .B2(n15289), .A(n15276), .ZN(n15278) );
  AND2_X1 U16832 ( .A1(n15279), .A2(n15278), .ZN(n15304) );
  AOI22_X1 U16833 ( .A1(n15295), .A2(n7820), .B1(n15304), .B2(n15293), .ZN(
        P3_U3414) );
  INV_X1 U16834 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15286) );
  INV_X1 U16835 ( .A(n15280), .ZN(n15285) );
  NOR2_X1 U16836 ( .A1(n15282), .A2(n15281), .ZN(n15284) );
  AOI211_X1 U16837 ( .C1(n15285), .C2(n15289), .A(n15284), .B(n15283), .ZN(
        n15305) );
  AOI22_X1 U16838 ( .A1(n15295), .A2(n15286), .B1(n15305), .B2(n15293), .ZN(
        P3_U3417) );
  INV_X1 U16839 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15294) );
  AOI22_X1 U16840 ( .A1(n15290), .A2(n15289), .B1(n15288), .B2(n15287), .ZN(
        n15291) );
  AND2_X1 U16841 ( .A1(n15292), .A2(n15291), .ZN(n15307) );
  AOI22_X1 U16842 ( .A1(n15295), .A2(n15294), .B1(n15307), .B2(n15293), .ZN(
        P3_U3420) );
  AOI22_X1 U16843 ( .A1(n15308), .A2(n15296), .B1(n11090), .B2(n15306), .ZN(
        P3_U3462) );
  AOI22_X1 U16844 ( .A1(n15308), .A2(n15298), .B1(n15297), .B2(n15306), .ZN(
        P3_U3463) );
  AOI22_X1 U16845 ( .A1(n15308), .A2(n15299), .B1(n11101), .B2(n15306), .ZN(
        P3_U3464) );
  AOI22_X1 U16846 ( .A1(n15308), .A2(n15301), .B1(n15300), .B2(n15306), .ZN(
        P3_U3465) );
  AOI22_X1 U16847 ( .A1(n15308), .A2(n15302), .B1(n11110), .B2(n15306), .ZN(
        P3_U3466) );
  AOI22_X1 U16848 ( .A1(n15308), .A2(n15304), .B1(n15303), .B2(n15306), .ZN(
        P3_U3467) );
  AOI22_X1 U16849 ( .A1(n15308), .A2(n15305), .B1(n11161), .B2(n15306), .ZN(
        P3_U3468) );
  AOI22_X1 U16850 ( .A1(n15308), .A2(n15307), .B1(n11186), .B2(n15306), .ZN(
        P3_U3469) );
  AOI22_X1 U16851 ( .A1(n15443), .A2(keyinput10), .B1(n15310), .B2(keyinput43), 
        .ZN(n15309) );
  OAI221_X1 U16852 ( .B1(n15443), .B2(keyinput10), .C1(n15310), .C2(keyinput43), .A(n15309), .ZN(n15321) );
  INV_X1 U16853 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15312) );
  AOI22_X1 U16854 ( .A1(n15313), .A2(keyinput45), .B1(n15312), .B2(keyinput61), 
        .ZN(n15311) );
  OAI221_X1 U16855 ( .B1(n15313), .B2(keyinput45), .C1(n15312), .C2(keyinput61), .A(n15311), .ZN(n15320) );
  AOI22_X1 U16856 ( .A1(n15315), .A2(keyinput41), .B1(n15447), .B2(keyinput42), 
        .ZN(n15314) );
  OAI221_X1 U16857 ( .B1(n15315), .B2(keyinput41), .C1(n15447), .C2(keyinput42), .A(n15314), .ZN(n15319) );
  AOI22_X1 U16858 ( .A1(n15317), .A2(keyinput25), .B1(keyinput33), .B2(n15445), 
        .ZN(n15316) );
  OAI221_X1 U16859 ( .B1(n15317), .B2(keyinput25), .C1(n15445), .C2(keyinput33), .A(n15316), .ZN(n15318) );
  NOR4_X1 U16860 ( .A1(n15321), .A2(n15320), .A3(n15319), .A4(n15318), .ZN(
        n15365) );
  INV_X1 U16861 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15324) );
  AOI22_X1 U16862 ( .A1(n15324), .A2(keyinput48), .B1(keyinput29), .B2(n15323), 
        .ZN(n15322) );
  OAI221_X1 U16863 ( .B1(n15324), .B2(keyinput48), .C1(n15323), .C2(keyinput29), .A(n15322), .ZN(n15335) );
  INV_X1 U16864 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U16865 ( .A1(n15327), .A2(keyinput2), .B1(keyinput4), .B2(n15326), 
        .ZN(n15325) );
  OAI221_X1 U16866 ( .B1(n15327), .B2(keyinput2), .C1(n15326), .C2(keyinput4), 
        .A(n15325), .ZN(n15334) );
  INV_X1 U16867 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U16868 ( .A1(n15448), .A2(keyinput1), .B1(keyinput37), .B2(n15329), 
        .ZN(n15328) );
  OAI221_X1 U16869 ( .B1(n15448), .B2(keyinput1), .C1(n15329), .C2(keyinput37), 
        .A(n15328), .ZN(n15333) );
  XOR2_X1 U16870 ( .A(n7880), .B(keyinput52), .Z(n15331) );
  XNOR2_X1 U16871 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput16), .ZN(n15330) );
  NAND2_X1 U16872 ( .A1(n15331), .A2(n15330), .ZN(n15332) );
  NOR4_X1 U16873 ( .A1(n15335), .A2(n15334), .A3(n15333), .A4(n15332), .ZN(
        n15364) );
  AOI22_X1 U16874 ( .A1(n9391), .A2(keyinput27), .B1(keyinput9), .B2(n15337), 
        .ZN(n15336) );
  OAI221_X1 U16875 ( .B1(n9391), .B2(keyinput27), .C1(n15337), .C2(keyinput9), 
        .A(n15336), .ZN(n15346) );
  AOI22_X1 U16876 ( .A1(n10674), .A2(keyinput12), .B1(keyinput18), .B2(n15339), 
        .ZN(n15338) );
  OAI221_X1 U16877 ( .B1(n10674), .B2(keyinput12), .C1(n15339), .C2(keyinput18), .A(n15338), .ZN(n15345) );
  XNOR2_X1 U16878 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput59), .ZN(n15343) );
  XNOR2_X1 U16879 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput3), .ZN(n15342) );
  XNOR2_X1 U16880 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput53), .ZN(n15341) );
  XNOR2_X1 U16881 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput6), .ZN(n15340) );
  NAND4_X1 U16882 ( .A1(n15343), .A2(n15342), .A3(n15341), .A4(n15340), .ZN(
        n15344) );
  NOR3_X1 U16883 ( .A1(n15346), .A2(n15345), .A3(n15344), .ZN(n15363) );
  AOI22_X1 U16884 ( .A1(n15349), .A2(keyinput20), .B1(n15348), .B2(keyinput0), 
        .ZN(n15347) );
  OAI221_X1 U16885 ( .B1(n15349), .B2(keyinput20), .C1(n15348), .C2(keyinput0), 
        .A(n15347), .ZN(n15361) );
  AOI22_X1 U16886 ( .A1(n15352), .A2(keyinput13), .B1(n15351), .B2(keyinput47), 
        .ZN(n15350) );
  OAI221_X1 U16887 ( .B1(n15352), .B2(keyinput13), .C1(n15351), .C2(keyinput47), .A(n15350), .ZN(n15360) );
  INV_X1 U16888 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U16889 ( .A1(n15355), .A2(keyinput17), .B1(n15354), .B2(keyinput14), 
        .ZN(n15353) );
  OAI221_X1 U16890 ( .B1(n15355), .B2(keyinput17), .C1(n15354), .C2(keyinput14), .A(n15353), .ZN(n15359) );
  XNOR2_X1 U16891 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput36), .ZN(n15357) );
  XNOR2_X1 U16892 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput55), .ZN(n15356)
         );
  NAND2_X1 U16893 ( .A1(n15357), .A2(n15356), .ZN(n15358) );
  NOR4_X1 U16894 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15362) );
  NAND4_X1 U16895 ( .A1(n15365), .A2(n15364), .A3(n15363), .A4(n15362), .ZN(
        n15424) );
  AOI22_X1 U16896 ( .A1(n15367), .A2(keyinput50), .B1(keyinput22), .B2(n7763), 
        .ZN(n15366) );
  OAI221_X1 U16897 ( .B1(n15367), .B2(keyinput50), .C1(n7763), .C2(keyinput22), 
        .A(n15366), .ZN(n15377) );
  INV_X1 U16898 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U16899 ( .A1(n15370), .A2(keyinput30), .B1(n15369), .B2(keyinput34), 
        .ZN(n15368) );
  OAI221_X1 U16900 ( .B1(n15370), .B2(keyinput30), .C1(n15369), .C2(keyinput34), .A(n15368), .ZN(n15376) );
  AOI22_X1 U16901 ( .A1(n11090), .A2(keyinput31), .B1(n15204), .B2(keyinput40), 
        .ZN(n15371) );
  OAI221_X1 U16902 ( .B1(n11090), .B2(keyinput31), .C1(n15204), .C2(keyinput40), .A(n15371), .ZN(n15375) );
  XOR2_X1 U16903 ( .A(n9735), .B(keyinput5), .Z(n15373) );
  XNOR2_X1 U16904 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput58), .ZN(n15372) );
  NAND2_X1 U16905 ( .A1(n15373), .A2(n15372), .ZN(n15374) );
  NOR4_X1 U16906 ( .A1(n15377), .A2(n15376), .A3(n15375), .A4(n15374), .ZN(
        n15422) );
  AOI22_X1 U16907 ( .A1(n15428), .A2(keyinput23), .B1(n15379), .B2(keyinput28), 
        .ZN(n15378) );
  OAI221_X1 U16908 ( .B1(n15428), .B2(keyinput23), .C1(n15379), .C2(keyinput28), .A(n15378), .ZN(n15388) );
  XNOR2_X1 U16909 ( .A(SI_8_), .B(keyinput46), .ZN(n15383) );
  XNOR2_X1 U16910 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput19), .ZN(n15382) );
  XNOR2_X1 U16911 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput8), .ZN(n15381) );
  XNOR2_X1 U16912 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput60), .ZN(n15380)
         );
  NAND4_X1 U16913 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15387) );
  XNOR2_X1 U16914 ( .A(n15451), .B(keyinput35), .ZN(n15386) );
  INV_X1 U16915 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15384) );
  XNOR2_X1 U16916 ( .A(keyinput38), .B(n15384), .ZN(n15385) );
  NOR4_X1 U16917 ( .A1(n15388), .A2(n15387), .A3(n15386), .A4(n15385), .ZN(
        n15421) );
  INV_X1 U16918 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U16919 ( .A1(n15391), .A2(keyinput15), .B1(keyinput56), .B2(n15390), 
        .ZN(n15389) );
  OAI221_X1 U16920 ( .B1(n15391), .B2(keyinput15), .C1(n15390), .C2(keyinput56), .A(n15389), .ZN(n15401) );
  INV_X1 U16921 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15393) );
  AOI22_X1 U16922 ( .A1(n15446), .A2(keyinput24), .B1(keyinput26), .B2(n15393), 
        .ZN(n15392) );
  OAI221_X1 U16923 ( .B1(n15446), .B2(keyinput24), .C1(n15393), .C2(keyinput26), .A(n15392), .ZN(n15400) );
  INV_X1 U16924 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U16925 ( .A1(n15396), .A2(keyinput21), .B1(keyinput63), .B2(n15395), 
        .ZN(n15394) );
  OAI221_X1 U16926 ( .B1(n15396), .B2(keyinput21), .C1(n15395), .C2(keyinput63), .A(n15394), .ZN(n15399) );
  AOI22_X1 U16927 ( .A1(n11111), .A2(keyinput57), .B1(keyinput62), .B2(n15442), 
        .ZN(n15397) );
  OAI221_X1 U16928 ( .B1(n11111), .B2(keyinput57), .C1(n15442), .C2(keyinput62), .A(n15397), .ZN(n15398) );
  NOR4_X1 U16929 ( .A1(n15401), .A2(n15400), .A3(n15399), .A4(n15398), .ZN(
        n15420) );
  INV_X1 U16930 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U16931 ( .A1(n7838), .A2(keyinput54), .B1(keyinput11), .B2(n15403), 
        .ZN(n15402) );
  OAI221_X1 U16932 ( .B1(n7838), .B2(keyinput54), .C1(n15403), .C2(keyinput11), 
        .A(n15402), .ZN(n15408) );
  INV_X1 U16933 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15405) );
  AOI22_X1 U16934 ( .A1(n15406), .A2(keyinput32), .B1(keyinput7), .B2(n15405), 
        .ZN(n15404) );
  OAI221_X1 U16935 ( .B1(n15406), .B2(keyinput32), .C1(n15405), .C2(keyinput7), 
        .A(n15404), .ZN(n15407) );
  NOR2_X1 U16936 ( .A1(n15408), .A2(n15407), .ZN(n15418) );
  INV_X1 U16937 ( .A(keyinput49), .ZN(n15409) );
  XNOR2_X1 U16938 ( .A(n15410), .B(n15409), .ZN(n15417) );
  XNOR2_X1 U16939 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput51), .ZN(n15416) );
  AOI22_X1 U16940 ( .A1(n15413), .A2(keyinput39), .B1(keyinput44), .B2(n15412), 
        .ZN(n15411) );
  OAI221_X1 U16941 ( .B1(n15413), .B2(keyinput39), .C1(n15412), .C2(keyinput44), .A(n15411), .ZN(n15414) );
  INV_X1 U16942 ( .A(n15414), .ZN(n15415) );
  AND4_X1 U16943 ( .A1(n15418), .A2(n15417), .A3(n15416), .A4(n15415), .ZN(
        n15419) );
  NAND4_X1 U16944 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15423) );
  NOR2_X1 U16945 ( .A1(n15424), .A2(n15423), .ZN(n15427) );
  NAND2_X1 U16946 ( .A1(n15425), .A2(P3_D_REG_16__SCAN_IN), .ZN(n15426) );
  XNOR2_X1 U16947 ( .A(n15427), .B(n15426), .ZN(n15461) );
  NOR4_X1 U16948 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(P3_REG2_REG_11__SCAN_IN), 
        .A3(P2_DATAO_REG_30__SCAN_IN), .A4(P2_U3088), .ZN(n15459) );
  NAND3_X1 U16949 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(n15429), .A3(n15428), 
        .ZN(n15432) );
  NAND4_X1 U16950 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .A3(P3_DATAO_REG_10__SCAN_IN), .A4(P3_DATAO_REG_21__SCAN_IN), .ZN(
        n15431) );
  NAND4_X1 U16951 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), 
        .A3(P3_REG2_REG_7__SCAN_IN), .A4(P1_REG3_REG_8__SCAN_IN), .ZN(n15430)
         );
  NOR4_X1 U16952 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n15432), .A3(n15431), .A4(
        n15430), .ZN(n15458) );
  NAND4_X1 U16953 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_REG0_REG_19__SCAN_IN), 
        .A3(P3_REG3_REG_4__SCAN_IN), .A4(P3_REG2_REG_4__SCAN_IN), .ZN(n15436)
         );
  NAND4_X1 U16954 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_REG0_REG_2__SCAN_IN), .A4(P1_REG1_REG_25__SCAN_IN), .ZN(n15435) );
  NAND4_X1 U16955 ( .A1(SI_21_), .A2(SI_14_), .A3(P1_REG3_REG_10__SCAN_IN), 
        .A4(P1_REG1_REG_15__SCAN_IN), .ZN(n15434) );
  NAND4_X1 U16956 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(
        P2_DATAO_REG_22__SCAN_IN), .A3(P1_DATAO_REG_22__SCAN_IN), .A4(
        P2_REG2_REG_25__SCAN_IN), .ZN(n15433) );
  NOR4_X1 U16957 ( .A1(n15436), .A2(n15435), .A3(n15434), .A4(n15433), .ZN(
        n15457) );
  NOR4_X1 U16958 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .A3(P2_D_REG_24__SCAN_IN), .A4(SI_8_), .ZN(n15440) );
  NOR4_X1 U16959 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG0_REG_27__SCAN_IN), 
        .A3(P1_REG0_REG_26__SCAN_IN), .A4(P1_REG0_REG_31__SCAN_IN), .ZN(n15439) );
  NOR4_X1 U16960 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_REG0_REG_24__SCAN_IN), .ZN(n15438) );
  NOR4_X1 U16961 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .A3(P1_REG2_REG_24__SCAN_IN), .A4(P1_REG1_REG_0__SCAN_IN), .ZN(n15437)
         );
  NAND4_X1 U16962 ( .A1(n15440), .A2(n15439), .A3(n15438), .A4(n15437), .ZN(
        n15455) );
  INV_X1 U16963 ( .A(n15441), .ZN(n15454) );
  NAND4_X1 U16964 ( .A1(n15444), .A2(n15443), .A3(n7763), .A4(n15442), .ZN(
        n15453) );
  NOR4_X1 U16965 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .A3(P3_REG2_REG_10__SCAN_IN), .A4(P3_REG1_REG_3__SCAN_IN), .ZN(n15450)
         );
  AND4_X1 U16966 ( .A1(n15448), .A2(n15447), .A3(n15446), .A4(n15445), .ZN(
        n15449) );
  NAND4_X1 U16967 ( .A1(n15451), .A2(P3_ADDR_REG_2__SCAN_IN), .A3(n15450), 
        .A4(n15449), .ZN(n15452) );
  NOR4_X1 U16968 ( .A1(n15455), .A2(n15454), .A3(n15453), .A4(n15452), .ZN(
        n15456) );
  NAND4_X1 U16969 ( .A1(n15459), .A2(n15458), .A3(n15457), .A4(n15456), .ZN(
        n15460) );
  XNOR2_X1 U16970 ( .A(n15461), .B(n15460), .ZN(P3_U3249) );
  XNOR2_X1 U16971 ( .A(n15463), .B(n15462), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16972 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15464), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16973 ( .B1(n15466), .B2(n15465), .A(n15474), .ZN(SUB_1596_U53) );
  XOR2_X1 U16974 ( .A(n15468), .B(n15467), .Z(SUB_1596_U56) );
  OAI21_X1 U16975 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(n15472) );
  XNOR2_X1 U16976 ( .A(n15472), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16977 ( .A(n15474), .B(n15473), .Z(SUB_1596_U5) );
  CLKBUF_X1 U8484 ( .A(n8511), .Z(n9155) );
endmodule

