

module b15_C_gen_AntiSAT_k_128_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814;

  INV_X2 U3432 ( .A(n6050), .ZN(n6014) );
  OR2_X1 U3433 ( .A1(n5470), .A2(n4364), .ZN(n5460) );
  CLKBUF_X2 U3434 ( .A(n4024), .Z(n5484) );
  CLKBUF_X2 U3435 ( .A(n3199), .Z(n3852) );
  CLKBUF_X2 U3436 ( .A(n3279), .Z(n2986) );
  INV_X1 U3437 ( .A(n4339), .ZN(n4240) );
  INV_X1 U3438 ( .A(n3635), .ZN(n3280) );
  BUF_X1 U3439 ( .A(n3250), .Z(n3009) );
  NAND2_X1 U3440 ( .A1(n3235), .A2(n3251), .ZN(n4017) );
  OR2_X1 U3441 ( .A1(n3166), .A2(n3167), .ZN(n3252) );
  AND2_X1 U3442 ( .A1(n3118), .A2(n4523), .ZN(n3179) );
  AND2_X2 U3443 ( .A1(n4403), .A2(n4536), .ZN(n3177) );
  AND2_X2 U3444 ( .A1(n4536), .A2(n4414), .ZN(n3006) );
  AND2_X1 U34450 ( .A1(n3244), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3003) );
  INV_X1 U34480 ( .A(n3945), .ZN(n3980) );
  NAND2_X1 U3449 ( .A1(n4010), .A2(n4339), .ZN(n4118) );
  NAND2_X1 U3450 ( .A1(n4045), .A2(n4102), .ZN(n4315) );
  AND2_X2 U34510 ( .A1(n5375), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4404) );
  AND2_X1 U34520 ( .A1(n6020), .A2(n4358), .ZN(n6054) );
  NAND2_X1 U34530 ( .A1(n5434), .A2(n5435), .ZN(n5422) );
  INV_X1 U3454 ( .A(n6054), .ZN(n6024) );
  OR2_X1 U34550 ( .A1(n5434), .A2(n5450), .ZN(n5550) );
  OR2_X1 U34560 ( .A1(n4437), .A2(n4293), .ZN(n6134) );
  OAI222_X1 U3457 ( .A1(n4586), .A2(n5773), .B1(n5772), .B2(n5771), .C1(n6390), 
        .C2(n5770), .ZN(n5774) );
  AND2_X1 U3458 ( .A1(n3368), .A2(n3367), .ZN(n2984) );
  AND2_X1 U34590 ( .A1(n5280), .A2(n3041), .ZN(n5310) );
  AND2_X2 U34600 ( .A1(n3406), .A2(n3405), .ZN(n3945) );
  OAI21_X2 U34610 ( .B1(n4586), .B2(n4160), .A(n4159), .ZN(n4161) );
  AND2_X4 U34620 ( .A1(n3112), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4403) );
  AND2_X2 U34630 ( .A1(n4536), .A2(n4414), .ZN(n3007) );
  AND2_X4 U34640 ( .A1(n4404), .A2(n4522), .ZN(n3022) );
  OR2_X1 U34650 ( .A1(n5588), .A2(n5589), .ZN(n3005) );
  XNOR2_X1 U3466 ( .A(n4323), .B(n4322), .ZN(n5384) );
  INV_X4 U3467 ( .A(n3035), .ZN(n2985) );
  NAND2_X1 U34680 ( .A1(n4316), .A2(n5400), .ZN(n4318) );
  CLKBUF_X2 U34690 ( .A(n6118), .Z(n6122) );
  NAND2_X1 U34700 ( .A1(n5616), .A2(n4301), .ZN(n6162) );
  OR2_X1 U34710 ( .A1(n3027), .A2(n5314), .ZN(n5313) );
  AND3_X1 U34720 ( .A1(n3054), .A2(n3056), .A3(n3055), .ZN(n4726) );
  CLKBUF_X1 U34730 ( .A(n3003), .Z(n3399) );
  AND3_X2 U34740 ( .A1(n3247), .A2(n3280), .A3(n3246), .ZN(n4245) );
  CLKBUF_X2 U3475 ( .A(n3010), .Z(n3004) );
  CLKBUF_X1 U3476 ( .A(n3251), .Z(n4621) );
  CLKBUF_X2 U3477 ( .A(n3273), .Z(n3010) );
  CLKBUF_X3 U3478 ( .A(n3252), .Z(n3015) );
  NAND2_X2 U3479 ( .A1(n3176), .A2(n3028), .ZN(n3249) );
  AND4_X1 U3480 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3124)
         );
  BUF_X2 U3481 ( .A(n3304), .Z(n3021) );
  CLKBUF_X2 U3482 ( .A(n3869), .Z(n3851) );
  BUF_X2 U3483 ( .A(n3348), .Z(n3874) );
  BUF_X2 U3484 ( .A(n3185), .Z(n3018) );
  CLKBUF_X2 U3485 ( .A(n6106), .Z(n6603) );
  BUF_X2 U3486 ( .A(n3178), .Z(n3909) );
  AND2_X2 U3487 ( .A1(n3117), .A2(n3118), .ZN(n3150) );
  AOI21_X1 U3488 ( .B1(n5533), .B2(n5541), .A(n5532), .ZN(n5534) );
  OAI22_X1 U3489 ( .A1(n5572), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5582), .B2(n5563), .ZN(n5564) );
  AOI211_X1 U3490 ( .C1(n6130), .C2(n5547), .A(n5546), .B(n5545), .ZN(n5548)
         );
  NOR2_X1 U3491 ( .A1(n5588), .A2(n5589), .ZN(n5587) );
  CLKBUF_X1 U3492 ( .A(n2998), .Z(n5604) );
  NAND2_X1 U3493 ( .A1(n5612), .A2(n3068), .ZN(n5570) );
  AND2_X1 U3494 ( .A1(n2989), .A2(n2990), .ZN(n5603) );
  AND2_X1 U3495 ( .A1(n5489), .A2(n5503), .ZN(n6067) );
  NAND2_X1 U3496 ( .A1(n5049), .A2(n4207), .ZN(n5181) );
  NAND4_X1 U3497 ( .A1(n3501), .A2(n4834), .A3(n3093), .A4(n3579), .ZN(n3587)
         );
  OR2_X1 U3498 ( .A1(n2995), .A2(n6137), .ZN(n2994) );
  AND2_X1 U3499 ( .A1(n3063), .A2(n3034), .ZN(n4330) );
  NOR2_X1 U3500 ( .A1(n4212), .A2(n3086), .ZN(n3085) );
  OR2_X1 U3501 ( .A1(n5384), .A2(n6185), .ZN(n3063) );
  NAND2_X1 U3502 ( .A1(n3500), .A2(n3499), .ZN(n4834) );
  NAND2_X1 U3503 ( .A1(n4321), .A2(n4320), .ZN(n4323) );
  NAND2_X1 U3504 ( .A1(n4177), .A2(n4176), .ZN(n4178) );
  NAND2_X1 U3505 ( .A1(n3397), .A2(n3396), .ZN(n4508) );
  NOR2_X1 U3506 ( .A1(n6386), .A2(n4844), .ZN(n6374) );
  AND2_X1 U3507 ( .A1(n3447), .A2(n3446), .ZN(n4635) );
  NOR2_X1 U3508 ( .A1(n6555), .A2(n5961), .ZN(n5319) );
  NAND2_X1 U3509 ( .A1(n3450), .A2(n3421), .ZN(n4586) );
  NAND2_X1 U3510 ( .A1(n2984), .A2(n3420), .ZN(n3450) );
  AND2_X1 U3511 ( .A1(n6020), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5381) );
  AOI21_X1 U3512 ( .B1(n4498), .B2(n4499), .A(n4152), .ZN(n6155) );
  NAND2_X1 U3513 ( .A1(n5512), .A2(n4002), .ZN(n5848) );
  NAND2_X1 U3514 ( .A1(n4454), .A2(n4371), .ZN(n6601) );
  CLKBUF_X1 U3515 ( .A(n4521), .Z(n5119) );
  AND2_X2 U3516 ( .A1(n3982), .A2(n3981), .ZN(n6480) );
  NAND2_X1 U3517 ( .A1(n3329), .A2(n3328), .ZN(n3331) );
  AND2_X1 U3518 ( .A1(n4519), .A2(n3057), .ZN(n3056) );
  OR2_X1 U3519 ( .A1(n3059), .A2(n5060), .ZN(n3058) );
  INV_X1 U3520 ( .A(n4030), .ZN(n4519) );
  OR2_X1 U3521 ( .A1(n4837), .A2(n3060), .ZN(n3059) );
  NAND2_X1 U3522 ( .A1(n3243), .A2(n3242), .ZN(n3244) );
  NOR2_X1 U3523 ( .A1(n3036), .A2(n4037), .ZN(n4038) );
  INV_X1 U3524 ( .A(n4315), .ZN(n4110) );
  AND2_X1 U3525 ( .A1(n3281), .A2(n3229), .ZN(n3231) );
  NAND2_X1 U3526 ( .A1(n4118), .A2(n5484), .ZN(n4446) );
  NAND2_X1 U3527 ( .A1(n3228), .A2(n3269), .ZN(n3281) );
  AND2_X1 U3528 ( .A1(n3270), .A2(n4017), .ZN(n3067) );
  AND2_X1 U3529 ( .A1(n4609), .A2(n3275), .ZN(n3269) );
  AND2_X1 U3530 ( .A1(n3270), .A2(n4009), .ZN(n3228) );
  OR2_X1 U3531 ( .A1(n3343), .A2(n3342), .ZN(n4202) );
  NAND2_X2 U3532 ( .A1(n3124), .A2(n3123), .ZN(n3251) );
  NAND4_X1 U3533 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3273)
         );
  OR2_X1 U3534 ( .A1(n3354), .A2(n3353), .ZN(n4145) );
  AND2_X1 U3535 ( .A1(n3141), .A2(n3140), .ZN(n3157) );
  AND4_X1 U3536 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n3028)
         );
  AND4_X1 U3537 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3156)
         );
  AND4_X1 U3538 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3212)
         );
  AND4_X1 U3539 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3227)
         );
  AND4_X1 U3540 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3134)
         );
  AND4_X1 U3541 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3214)
         );
  AND4_X1 U3542 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3215)
         );
  AND4_X1 U3543 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3213)
         );
  AND4_X1 U3544 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3176)
         );
  AND4_X1 U3545 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3140)
         );
  AND3_X1 U3546 ( .A1(n3131), .A2(n3130), .A3(n3129), .ZN(n3133) );
  AND4_X1 U3547 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3155)
         );
  AND3_X1 U3548 ( .A1(n3153), .A2(n3152), .A3(n3151), .ZN(n3154) );
  AND4_X1 U3549 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3123)
         );
  BUF_X2 U3550 ( .A(n3193), .Z(n3332) );
  BUF_X2 U3551 ( .A(n3222), .Z(n3333) );
  AND2_X2 U3552 ( .A1(n3118), .A2(n4523), .ZN(n3019) );
  AND2_X2 U3553 ( .A1(n4404), .A2(n4536), .ZN(n3222) );
  CLKBUF_X1 U3554 ( .A(n3304), .Z(n2987) );
  AND2_X2 U3555 ( .A1(n3110), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4522)
         );
  INV_X1 U3556 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3110) );
  NOR2_X2 U3557 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3118) );
  NOR2_X2 U3558 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U3559 ( .A1(n4570), .A2(n4170), .ZN(n4730) );
  NAND2_X2 U3560 ( .A1(n4226), .A2(n3106), .ZN(n5528) );
  NOR4_X2 U3561 ( .A1(n3023), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4309), .ZN(n4310) );
  AND2_X1 U3562 ( .A1(n5312), .A2(n3041), .ZN(n2988) );
  INV_X2 U3563 ( .A(n3217), .ZN(n3235) );
  OR2_X1 U3564 ( .A1(n5448), .A2(n5458), .ZN(n5852) );
  NAND2_X1 U3565 ( .A1(n3102), .A2(n3100), .ZN(n4295) );
  AND2_X2 U3566 ( .A1(n5448), .A2(n5449), .ZN(n5434) );
  NAND2_X1 U3567 ( .A1(n4217), .A2(n2992), .ZN(n2989) );
  OR2_X1 U3568 ( .A1(n2991), .A2(n3068), .ZN(n2990) );
  INV_X1 U3569 ( .A(n4222), .ZN(n2991) );
  AND2_X1 U3570 ( .A1(n4216), .A2(n4222), .ZN(n2992) );
  NAND2_X1 U3571 ( .A1(n4731), .A2(n2996), .ZN(n2993) );
  AND2_X2 U3572 ( .A1(n2993), .A2(n2994), .ZN(n4955) );
  INV_X1 U3573 ( .A(n4189), .ZN(n2995) );
  AND2_X1 U3574 ( .A1(n4179), .A2(n4189), .ZN(n2996) );
  NOR2_X2 U3575 ( .A1(n5313), .A2(n5494), .ZN(n5481) );
  XNOR2_X1 U3577 ( .A(n4314), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5365)
         );
  INV_X2 U3578 ( .A(n4833), .ZN(n3501) );
  NAND2_X1 U3579 ( .A1(n4214), .A2(n4213), .ZN(n5342) );
  XNOR2_X1 U3580 ( .A(n4295), .B(n3927), .ZN(n5353) );
  OAI21_X1 U3581 ( .B1(n4585), .B2(n4160), .A(n4135), .ZN(n6154) );
  NAND2_X1 U3582 ( .A1(n5570), .A2(n4222), .ZN(n2998) );
  INV_X1 U3583 ( .A(n4007), .ZN(n2999) );
  NAND2_X1 U3585 ( .A1(n4217), .A2(n4216), .ZN(n5612) );
  NAND2_X2 U3586 ( .A1(n5273), .A2(n3600), .ZN(n5280) );
  CLKBUF_X1 U3587 ( .A(n4955), .Z(n3001) );
  NAND2_X1 U3588 ( .A1(n3368), .A2(n3367), .ZN(n3002) );
  BUF_X2 U3589 ( .A(n3217), .Z(n4609) );
  NAND3_X2 U3590 ( .A1(n3134), .A2(n3133), .A3(n3132), .ZN(n3217) );
  AND2_X2 U3591 ( .A1(n4403), .A2(n4522), .ZN(n3185) );
  NAND2_X2 U3592 ( .A1(n3233), .A2(n3252), .ZN(n3635) );
  AND2_X1 U3593 ( .A1(n3117), .A2(n4414), .ZN(n3008) );
  AND2_X1 U3594 ( .A1(n3117), .A2(n4414), .ZN(n3178) );
  INV_X2 U3595 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3111) );
  INV_X2 U3596 ( .A(n3249), .ZN(n4391) );
  AND2_X2 U3597 ( .A1(n4403), .A2(n4536), .ZN(n3011) );
  XNOR2_X2 U3598 ( .A(n3313), .B(n3312), .ZN(n3368) );
  XNOR2_X1 U3599 ( .A(n3450), .B(n3451), .ZN(n4163) );
  NAND2_X1 U3600 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  NAND2_X1 U3601 ( .A1(n3377), .A2(n3381), .ZN(n5009) );
  AND3_X1 U3602 ( .A1(n3004), .A2(n4339), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3972) );
  OR2_X1 U3603 ( .A1(n3004), .A2(n6504), .ZN(n3406) );
  OR2_X2 U3604 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  NAND2_X2 U3605 ( .A1(n3294), .A2(n3293), .ZN(n3398) );
  INV_X2 U3606 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5375) );
  AND2_X1 U3607 ( .A1(n4523), .A2(n4414), .ZN(n3012) );
  AND2_X1 U3608 ( .A1(n4523), .A2(n4414), .ZN(n3013) );
  NAND2_X2 U3609 ( .A1(n3135), .A2(n3217), .ZN(n3239) );
  INV_X2 U3610 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3112) );
  AND2_X1 U3611 ( .A1(n4246), .A2(n4339), .ZN(n3279) );
  BUF_X8 U3612 ( .A(n3298), .Z(n3017) );
  AND2_X2 U3613 ( .A1(n4523), .A2(n4403), .ZN(n3298) );
  NOR2_X2 U3614 ( .A1(n3277), .A2(n3248), .ZN(n4239) );
  AND2_X4 U3615 ( .A1(n3111), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4523)
         );
  AND2_X2 U3616 ( .A1(n4361), .A2(n5457), .ZN(n5448) );
  NOR2_X2 U3617 ( .A1(n4359), .A2(n4362), .ZN(n4361) );
  OAI21_X2 U3618 ( .B1(n5265), .B2(n3083), .A(n3081), .ZN(n5872) );
  NAND2_X2 U3619 ( .A1(n4208), .A2(n5180), .ZN(n5265) );
  OAI22_X2 U3620 ( .A1(n5603), .A2(n5605), .B1(n3035), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5597) );
  NOR2_X2 U3621 ( .A1(n5311), .A2(n3097), .ZN(n5478) );
  NAND2_X2 U3622 ( .A1(n2988), .A2(n5280), .ZN(n5311) );
  NOR2_X2 U3623 ( .A1(n4632), .A2(n4724), .ZN(n4723) );
  AND2_X4 U3624 ( .A1(n3331), .A2(n3330), .ZN(n3383) );
  AND2_X2 U3625 ( .A1(n3118), .A2(n4523), .ZN(n3020) );
  AND2_X1 U3626 ( .A1(n4523), .A2(n4414), .ZN(n3304) );
  AND2_X4 U3627 ( .A1(n4404), .A2(n4522), .ZN(n3194) );
  AND2_X4 U3628 ( .A1(n4523), .A2(n4404), .ZN(n3411) );
  NAND2_X1 U3629 ( .A1(n3452), .A2(n3451), .ZN(n3470) );
  INV_X1 U3630 ( .A(n3450), .ZN(n3452) );
  AND2_X1 U3631 ( .A1(n3239), .A2(n4339), .ZN(n3216) );
  NAND2_X1 U3632 ( .A1(n3439), .A2(n3438), .ZN(n3451) );
  NOR2_X1 U3633 ( .A1(n3983), .A2(n3984), .ZN(n4255) );
  INV_X1 U3634 ( .A(n5472), .ZN(n3089) );
  NOR2_X1 U3635 ( .A1(n4965), .A2(n3094), .ZN(n3093) );
  INV_X1 U3636 ( .A(n5058), .ZN(n3094) );
  NAND2_X1 U3637 ( .A1(n3233), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3614) );
  INV_X1 U3638 ( .A(n3614), .ZN(n3623) );
  AND2_X1 U3639 ( .A1(n4091), .A2(n3049), .ZN(n3048) );
  INV_X1 U3640 ( .A(n5711), .ZN(n3049) );
  INV_X1 U3641 ( .A(n4728), .ZN(n3055) );
  NOR2_X1 U3642 ( .A1(n4009), .A2(n3249), .ZN(n4019) );
  INV_X1 U3643 ( .A(n3801), .ZN(n5357) );
  NAND2_X1 U3644 ( .A1(n6480), .A2(n6501), .ZN(n4437) );
  INV_X1 U3645 ( .A(n5009), .ZN(n4912) );
  NAND2_X1 U3646 ( .A1(n4240), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3405) );
  NOR2_X2 U3647 ( .A1(n3470), .A2(n3469), .ZN(n3493) );
  OR2_X1 U3648 ( .A1(n3324), .A2(n3323), .ZN(n4137) );
  OR2_X1 U3649 ( .A1(n3310), .A2(n3309), .ZN(n3311) );
  AND2_X1 U3650 ( .A1(n4006), .A2(n4008), .ZN(n4238) );
  AOI22_X1 U3651 ( .A1(n3020), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3011), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U3652 ( .A1(n3016), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U3653 ( .A1(n3348), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U3654 ( .A1(n3869), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3131) );
  AOI21_X1 U3655 ( .B1(n6252), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3938), 
        .ZN(n3976) );
  INV_X1 U3656 ( .A(n5474), .ZN(n3754) );
  INV_X1 U3657 ( .A(n3924), .ZN(n3898) );
  AND2_X1 U3658 ( .A1(n3631), .A2(n5282), .ZN(n3096) );
  INV_X1 U3659 ( .A(n3311), .ZN(n4156) );
  OR3_X1 U3660 ( .A1(n2985), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5653), 
        .ZN(n4309) );
  OR2_X1 U3661 ( .A1(n5459), .A2(n5452), .ZN(n3064) );
  INV_X1 U3662 ( .A(n5475), .ZN(n3047) );
  OR2_X1 U3663 ( .A1(n3053), .A2(n5321), .ZN(n3052) );
  INV_X1 U3664 ( .A(n5288), .ZN(n3084) );
  NAND2_X1 U3665 ( .A1(n4102), .A2(n5484), .ZN(n4109) );
  AND2_X1 U3666 ( .A1(n4518), .A2(n4574), .ZN(n3057) );
  OR2_X1 U3667 ( .A1(n6480), .A2(n4418), .ZN(n4395) );
  OR2_X1 U3668 ( .A1(n3985), .A2(n3992), .ZN(n3993) );
  INV_X1 U3669 ( .A(n6108), .ZN(n4438) );
  NAND2_X1 U3670 ( .A1(n3904), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4354)
         );
  NOR2_X1 U3671 ( .A1(n5423), .A2(n3101), .ZN(n3100) );
  INV_X1 U3672 ( .A(n4296), .ZN(n3101) );
  AND2_X1 U3673 ( .A1(n3734), .A2(n3733), .ZN(n5591) );
  NAND2_X1 U3674 ( .A1(n5479), .A2(n3098), .ZN(n3097) );
  INV_X1 U3675 ( .A(n3099), .ZN(n3098) );
  NAND2_X1 U3676 ( .A1(n3584), .A2(n3585), .ZN(n3600) );
  AND4_X1 U3677 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n4965)
         );
  INV_X1 U3678 ( .A(n3077), .ZN(n3076) );
  AOI21_X1 U3679 ( .B1(n3075), .B2(n3077), .A(n3040), .ZN(n3074) );
  AND2_X1 U3680 ( .A1(n4090), .A2(n5493), .ZN(n4091) );
  NAND2_X1 U3681 ( .A1(n5481), .A2(n3048), .ZN(n5714) );
  INV_X1 U3682 ( .A(n5266), .ZN(n3086) );
  AND2_X1 U3683 ( .A1(n5892), .A2(n5302), .ZN(n5184) );
  INV_X1 U3684 ( .A(n6202), .ZN(n5725) );
  NAND2_X1 U3685 ( .A1(n4275), .A2(n6479), .ZN(n6211) );
  INV_X1 U3686 ( .A(n3420), .ZN(n4795) );
  NOR2_X1 U3687 ( .A1(n6475), .A2(n4246), .ZN(n4527) );
  AND2_X1 U3688 ( .A1(n4794), .A2(n4586), .ZN(n5010) );
  AND2_X1 U3689 ( .A1(n4585), .A2(n3070), .ZN(n4794) );
  OR2_X1 U3690 ( .A1(n4586), .A2(n5765), .ZN(n6386) );
  AND2_X1 U3691 ( .A1(n5012), .A2(n5119), .ZN(n6387) );
  NAND2_X1 U3692 ( .A1(n3404), .A2(n3403), .ZN(n5084) );
  INV_X1 U3693 ( .A(n4738), .ZN(n4849) );
  AOI22_X1 U3694 ( .A1(n3011), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3008), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U3695 ( .A1(n4600), .A2(n3070), .ZN(n4710) );
  INV_X1 U3696 ( .A(n4739), .ZN(n4712) );
  INV_X1 U3697 ( .A(n6389), .ZN(n4879) );
  AND2_X1 U3698 ( .A1(n6493), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3997) );
  INV_X2 U3699 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6503) );
  AND2_X1 U3700 ( .A1(n5800), .A2(n5378), .ZN(n5782) );
  NOR2_X1 U3701 ( .A1(n5362), .A2(n6493), .ZN(n4363) );
  OR2_X1 U3702 ( .A1(n5417), .A2(n5843), .ZN(n4132) );
  INV_X1 U3703 ( .A(n6066), .ZN(n5495) );
  NAND2_X1 U3704 ( .A1(n6066), .A2(n5513), .ZN(n5843) );
  AND2_X1 U3705 ( .A1(n5512), .A2(n4003), .ZN(n6074) );
  NAND2_X1 U3706 ( .A1(n6134), .A2(n4298), .ZN(n5616) );
  NOR2_X1 U3707 ( .A1(n5882), .A2(n4278), .ZN(n5736) );
  INV_X1 U3708 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6455) );
  OAI21_X1 U3709 ( .B1(n3070), .B2(STATEBS16_REG_SCAN_IN), .A(n6384), .ZN(
        n3072) );
  CLKBUF_X1 U3710 ( .A(n4399), .Z(n4400) );
  INV_X1 U3711 ( .A(n4585), .ZN(n5765) );
  AND2_X1 U3712 ( .A1(n3070), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6254) );
  NAND2_X1 U3713 ( .A1(n3398), .A2(n3297), .ZN(n4415) );
  INV_X1 U3714 ( .A(n5119), .ZN(n5771) );
  NAND2_X1 U3715 ( .A1(n5081), .A2(n3070), .ZN(n6445) );
  AND2_X1 U3716 ( .A1(n3635), .A2(n3249), .ZN(n3234) );
  AND2_X1 U3717 ( .A1(n2985), .A2(n5683), .ZN(n4228) );
  OR2_X1 U3718 ( .A1(n3462), .A2(n3461), .ZN(n4183) );
  OR2_X1 U3719 ( .A1(n3437), .A2(n3436), .ZN(n4172) );
  OAI211_X1 U3720 ( .C1(n4202), .C2(n3406), .A(n3362), .B(n3361), .ZN(n3370)
         );
  AND2_X1 U3721 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U3722 ( .A1(n3016), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3114) );
  NAND2_X1 U3723 ( .A1(n3972), .A2(n4190), .ZN(n3956) );
  OR2_X1 U3724 ( .A1(n3940), .A2(n3939), .ZN(n3973) );
  INV_X1 U3725 ( .A(n3973), .ZN(n3987) );
  AND4_X1 U3726 ( .A1(n4531), .A2(n3281), .A3(n6502), .A4(n3282), .ZN(n3283)
         );
  OR2_X1 U3727 ( .A1(n5502), .A2(n5490), .ZN(n3099) );
  INV_X1 U3728 ( .A(n5506), .ZN(n3095) );
  INV_X1 U3729 ( .A(n3493), .ZN(n3481) );
  INV_X1 U3730 ( .A(n3078), .ZN(n3075) );
  NOR2_X1 U3731 ( .A1(n4228), .A2(n3079), .ZN(n3078) );
  INV_X1 U3732 ( .A(n4227), .ZN(n3079) );
  OR2_X1 U3733 ( .A1(n5558), .A2(n4228), .ZN(n3077) );
  INV_X1 U3734 ( .A(n4967), .ZN(n3060) );
  NOR2_X1 U3735 ( .A1(n4109), .A2(EBX_REG_3__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U3736 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  OR2_X1 U3737 ( .A1(n3635), .A2(n3634), .ZN(n4016) );
  AND3_X1 U3738 ( .A1(n4015), .A2(n4238), .A3(n4014), .ZN(n4402) );
  INV_X1 U3739 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6461) );
  AOI22_X1 U3740 ( .A1(n3012), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U3741 ( .A1(n3348), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3225) );
  AOI22_X1 U3742 ( .A1(n3184), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3132) );
  AND2_X2 U3743 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4536) );
  INV_X1 U3744 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6466) );
  INV_X1 U3745 ( .A(n3956), .ZN(n3977) );
  AND2_X1 U3746 ( .A1(n4255), .A2(n3009), .ZN(n6473) );
  NOR2_X1 U3747 ( .A1(n3633), .A2(n3632), .ZN(n3649) );
  INV_X1 U3748 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3632) );
  XNOR2_X1 U3749 ( .A(n3398), .B(n5084), .ZN(n4521) );
  OAI21_X1 U3750 ( .B1(n4495), .B2(n4496), .A(n4029), .ZN(n4030) );
  AOI22_X1 U3751 ( .A1(n3903), .A2(n3902), .B1(n3920), .B2(n5404), .ZN(n4296)
         );
  OR2_X1 U3752 ( .A1(n3863), .A2(n5543), .ZN(n3865) );
  AOI22_X1 U3753 ( .A1(n3862), .A2(n3861), .B1(n3920), .B2(n5547), .ZN(n5435)
         );
  NAND2_X1 U3754 ( .A1(n3839), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3863)
         );
  OR2_X1 U3755 ( .A1(n3796), .A2(n5806), .ZN(n3797) );
  NOR2_X1 U3756 ( .A1(n3797), .A2(n4342), .ZN(n3838) );
  NAND2_X1 U3757 ( .A1(n3750), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3796)
         );
  AND2_X1 U3758 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n3716), .ZN(n3717)
         );
  NAND2_X1 U3759 ( .A1(n3717), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3749)
         );
  NOR2_X1 U3760 ( .A1(n3666), .A2(n3665), .ZN(n3667) );
  NAND2_X1 U3761 ( .A1(n3667), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3715)
         );
  AND3_X1 U3762 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n5318) );
  AND2_X1 U3763 ( .A1(n3580), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3581)
         );
  NAND2_X1 U3764 ( .A1(n3581), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3626)
         );
  NOR2_X1 U3765 ( .A1(n3562), .A2(n3547), .ZN(n3580) );
  INV_X1 U3766 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3547) );
  AND2_X1 U3767 ( .A1(n4834), .A2(n3093), .ZN(n3090) );
  AND2_X1 U3768 ( .A1(n3512), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3518)
         );
  AND2_X1 U3769 ( .A1(n4834), .A2(n3092), .ZN(n3091) );
  INV_X1 U3770 ( .A(n4965), .ZN(n3092) );
  AND2_X1 U3771 ( .A1(n3485), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3512)
         );
  INV_X1 U3772 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3483) );
  INV_X1 U3773 ( .A(n4635), .ZN(n3448) );
  OAI211_X1 U3774 ( .C1(n3444), .C2(n3110), .A(n3392), .B(n3391), .ZN(n4510)
         );
  NAND2_X1 U3775 ( .A1(n4493), .A2(n4494), .ZN(n4492) );
  NOR2_X1 U3776 ( .A1(n4229), .A2(n4309), .ZN(n4291) );
  AND2_X1 U3777 ( .A1(n4120), .A2(n4119), .ZN(n5437) );
  AND2_X1 U3778 ( .A1(n4115), .A2(n4114), .ZN(n5452) );
  NOR2_X1 U3779 ( .A1(n5460), .A2(n3064), .ZN(n5451) );
  NAND2_X1 U3780 ( .A1(n5481), .A2(n3026), .ZN(n5470) );
  NOR2_X1 U3781 ( .A1(n3069), .A2(n3039), .ZN(n3068) );
  INV_X1 U3782 ( .A(n4219), .ZN(n3069) );
  AND2_X1 U3783 ( .A1(n4097), .A2(n4096), .ZN(n5475) );
  AND2_X1 U3784 ( .A1(n4088), .A2(n4087), .ZN(n5482) );
  OR2_X1 U3785 ( .A1(n5278), .A2(n3051), .ZN(n3050) );
  INV_X1 U3786 ( .A(n5507), .ZN(n3051) );
  NOR2_X1 U3787 ( .A1(n3105), .A2(n4200), .ZN(n4201) );
  AOI21_X1 U3788 ( .B1(n3082), .B2(n4211), .A(n3046), .ZN(n3081) );
  NAND2_X1 U3789 ( .A1(n4211), .A2(n3084), .ZN(n3083) );
  NOR2_X1 U3790 ( .A1(n3085), .A2(n5288), .ZN(n3082) );
  NAND2_X1 U3791 ( .A1(n5066), .A2(n5065), .ZN(n5987) );
  OR2_X1 U3792 ( .A1(n5777), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4297) );
  NOR2_X1 U3793 ( .A1(n4836), .A2(n4837), .ZN(n4966) );
  CLKBUF_X1 U3794 ( .A(n4726), .Z(n4841) );
  NAND2_X1 U3795 ( .A1(n3054), .A2(n3056), .ZN(n4727) );
  NOR2_X1 U3796 ( .A1(n4516), .A2(n4515), .ZN(n4573) );
  INV_X1 U3797 ( .A(n4102), .ZN(n4496) );
  OAI21_X1 U3798 ( .B1(n5009), .B2(n4160), .A(n4147), .ZN(n4381) );
  INV_X1 U3799 ( .A(n4016), .ZN(n5367) );
  NAND4_X1 U3800 ( .A1(n4019), .A2(n4240), .A3(n3280), .A4(n3010), .ZN(n4531)
         );
  OR2_X1 U3801 ( .A1(n5119), .A2(n4846), .ZN(n4643) );
  OR2_X1 U3802 ( .A1(n5769), .A2(n4136), .ZN(n4911) );
  INV_X1 U3803 ( .A(n3070), .ZN(n4874) );
  NOR2_X1 U3804 ( .A1(n3070), .A2(n5923), .ZN(n4875) );
  AND2_X1 U3805 ( .A1(n3070), .A2(n5009), .ZN(n5193) );
  AND2_X1 U3806 ( .A1(n4600), .A2(n4874), .ZN(n4605) );
  NOR2_X1 U3807 ( .A1(n4415), .A2(n4400), .ZN(n6308) );
  NOR2_X1 U3808 ( .A1(n6587), .A2(n4595), .ZN(n4624) );
  NOR2_X2 U3809 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6384) );
  NAND2_X1 U3810 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4545) );
  AND2_X1 U3811 ( .A1(n5816), .A2(n4353), .ZN(n5800) );
  AND2_X1 U3812 ( .A1(n6020), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6051) );
  AND2_X1 U3813 ( .A1(n4102), .A2(n4367), .ZN(n6050) );
  INV_X1 U3814 ( .A(n6051), .ZN(n6036) );
  INV_X1 U3815 ( .A(n6047), .ZN(n5949) );
  INV_X1 U3816 ( .A(n5843), .ZN(n6062) );
  AND2_X1 U3817 ( .A1(n4022), .A2(n6501), .ZN(n6066) );
  INV_X1 U3818 ( .A(n3015), .ZN(n5513) );
  INV_X1 U3819 ( .A(n5848), .ZN(n6071) );
  OR2_X1 U3820 ( .A1(n6070), .A2(n6074), .ZN(n5338) );
  NAND2_X1 U3821 ( .A1(n4001), .A2(n6124), .ZN(n5512) );
  OAI21_X1 U3822 ( .B1(n4396), .B2(n3998), .A(n6501), .ZN(n4001) );
  INV_X1 U3823 ( .A(n5338), .ZN(n4953) );
  NOR2_X1 U3824 ( .A1(n4527), .A2(n4435), .ZN(n4436) );
  NOR2_X1 U3825 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4545), .ZN(n6106) );
  INV_X1 U3826 ( .A(n6110), .ZN(n6121) );
  INV_X1 U3827 ( .A(n6124), .ZN(n4489) );
  OR2_X1 U3828 ( .A1(n4454), .A2(n3275), .ZN(n6110) );
  XNOR2_X1 U3829 ( .A(n4357), .B(n4356), .ZN(n5362) );
  XNOR2_X1 U3830 ( .A(n5359), .B(n5358), .ZN(n5514) );
  INV_X1 U3831 ( .A(n5356), .ZN(n3927) );
  INV_X1 U3832 ( .A(n5550), .ZN(n5849) );
  INV_X1 U3833 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5590) );
  CLKBUF_X1 U3834 ( .A(n5273), .Z(n5274) );
  INV_X1 U3835 ( .A(n6162), .ZN(n6130) );
  CLKBUF_X1 U3836 ( .A(n5049), .Z(n5050) );
  CLKBUF_X1 U3837 ( .A(n4956), .Z(n4957) );
  CLKBUF_X1 U3838 ( .A(n4731), .Z(n4732) );
  INV_X1 U3839 ( .A(n5616), .ZN(n6153) );
  OR2_X1 U3840 ( .A1(n6511), .A2(n6390), .ZN(n5622) );
  INV_X1 U3841 ( .A(n6134), .ZN(n6158) );
  NAND2_X1 U3842 ( .A1(n4329), .A2(n3062), .ZN(n3061) );
  INV_X1 U3843 ( .A(n5360), .ZN(n3062) );
  INV_X1 U3844 ( .A(n4313), .ZN(n4314) );
  NAND2_X1 U3845 ( .A1(n5481), .A2(n4091), .ZN(n5712) );
  OR2_X1 U3846 ( .A1(n6242), .A2(n4264), .ZN(n4269) );
  NAND2_X1 U3847 ( .A1(n5265), .A2(n3085), .ZN(n3080) );
  CLKBUF_X1 U3848 ( .A(n4570), .Z(n4571) );
  INV_X1 U3849 ( .A(n6169), .ZN(n6241) );
  INV_X1 U3850 ( .A(n6384), .ZN(n6390) );
  CLKBUF_X1 U3851 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n4529) );
  NAND2_X1 U3852 ( .A1(n6589), .A2(n6493), .ZN(n5777) );
  OAI221_X1 U3853 ( .B1(n5016), .B2(n6589), .C1(n5016), .C2(n5015), .A(n5014), 
        .ZN(n5041) );
  AND2_X1 U3854 ( .A1(n4798), .A2(n4797), .ZN(n6298) );
  INV_X1 U3855 ( .A(n5232), .ZN(n6352) );
  NAND2_X1 U3856 ( .A1(n3070), .A2(n4912), .ZN(n4845) );
  INV_X1 U3857 ( .A(n6374), .ZN(n4873) );
  AND2_X1 U3858 ( .A1(n4857), .A2(n4856), .ZN(n6371) );
  INV_X1 U3859 ( .A(n6379), .ZN(n6353) );
  OR2_X1 U3860 ( .A1(n3070), .A2(n4912), .ZN(n4844) );
  OAI211_X1 U3861 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6503), .A(n5014), .B(n4979), .ZN(n5002) );
  AOI22_X1 U3862 ( .A1(n4978), .A2(n6387), .B1(n5196), .B2(n4975), .ZN(n5008)
         );
  OR2_X1 U3863 ( .A1(n5090), .A2(n5089), .ZN(n5141) );
  NOR2_X1 U3864 ( .A1(n6747), .A2(n4849), .ZN(n6396) );
  INV_X1 U3865 ( .A(n6381), .ZN(n4933) );
  NOR2_X1 U3866 ( .A1(n6737), .A2(n4849), .ZN(n6403) );
  NOR2_X1 U3867 ( .A1(n6719), .A2(n4849), .ZN(n6410) );
  NOR2_X1 U3868 ( .A1(n6786), .A2(n4849), .ZN(n6417) );
  NOR2_X1 U3869 ( .A1(n4718), .A2(n4849), .ZN(n6424) );
  INV_X1 U3870 ( .A(n6421), .ZN(n6333) );
  NOR2_X1 U3871 ( .A1(n6725), .A2(n4849), .ZN(n6431) );
  INV_X1 U3872 ( .A(n6428), .ZN(n6337) );
  AND2_X1 U3873 ( .A1(n4605), .A2(n5009), .ZN(n5145) );
  NAND2_X1 U3874 ( .A1(n4605), .A2(n4912), .ZN(n4821) );
  NOR2_X1 U3875 ( .A1(n6782), .A2(n4849), .ZN(n6438) );
  INV_X1 U3876 ( .A(n6435), .ZN(n4923) );
  INV_X1 U3877 ( .A(n4792), .ZN(n4827) );
  INV_X1 U3878 ( .A(n6443), .ZN(n6350) );
  INV_X1 U3879 ( .A(n6403), .ZN(n6360) );
  INV_X1 U3880 ( .A(n6410), .ZN(n6328) );
  INV_X1 U3881 ( .A(n6417), .ZN(n6365) );
  NOR2_X1 U3882 ( .A1(n5622), .A2(n6679), .ZN(n6367) );
  INV_X1 U3883 ( .A(n6424), .ZN(n6370) );
  NOR2_X1 U3884 ( .A1(n5622), .A2(n6682), .ZN(n6375) );
  INV_X1 U3885 ( .A(n4719), .ZN(n4789) );
  INV_X1 U3886 ( .A(n6438), .ZN(n6348) );
  INV_X1 U3887 ( .A(n6448), .ZN(n6358) );
  AND2_X1 U3888 ( .A1(n4714), .A2(n4713), .ZN(n4786) );
  OAI211_X1 U3889 ( .C1(n6384), .C2(n4712), .A(n4709), .B(n4879), .ZN(n4785)
         );
  AND2_X1 U3890 ( .A1(n6480), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6491) );
  AND2_X1 U3891 ( .A1(n3997), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U3892 ( .A1(n4235), .A2(n6523), .ZN(n6518) );
  INV_X1 U3893 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U3894 ( .A1(n6385), .A2(n3071), .ZN(n5763) );
  INV_X1 U3895 ( .A(n3072), .ZN(n3071) );
  NAND2_X1 U3896 ( .A1(n5557), .A2(n5558), .ZN(n3023) );
  NAND2_X1 U3897 ( .A1(n3000), .A2(n4219), .ZN(n5610) );
  AND2_X1 U3898 ( .A1(n3090), .A2(n3501), .ZN(n5057) );
  NAND2_X1 U3899 ( .A1(n5280), .A2(n5282), .ZN(n5281) );
  AND2_X1 U3900 ( .A1(n3091), .A2(n3501), .ZN(n4964) );
  INV_X1 U3901 ( .A(n3275), .ZN(n4246) );
  NOR2_X1 U3902 ( .A1(n4339), .A2(n3275), .ZN(n3250) );
  OAI211_X1 U3903 ( .C1(n3239), .C2(n3010), .A(n3015), .B(n4017), .ZN(n3272)
         );
  OR3_X1 U3904 ( .A1(n5252), .A2(n5278), .A3(n3053), .ZN(n3024) );
  AND2_X1 U3905 ( .A1(n3048), .A2(n3047), .ZN(n3025) );
  AND2_X1 U3906 ( .A1(n3025), .A2(n5468), .ZN(n3026) );
  AND2_X1 U3907 ( .A1(n3275), .A2(n4339), .ZN(n4102) );
  OR3_X1 U3908 ( .A1(n5252), .A2(n3050), .A3(n3052), .ZN(n3027) );
  NAND2_X1 U3909 ( .A1(n3089), .A2(n3754), .ZN(n5465) );
  AND4_X1 U3910 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3029)
         );
  NOR2_X1 U3911 ( .A1(n5311), .A2(n3099), .ZN(n3030) );
  OAI21_X1 U3912 ( .B1(n4315), .B2(EBX_REG_1__SCAN_IN), .A(n4026), .ZN(n4029)
         );
  OR2_X1 U3913 ( .A1(n5311), .A2(n5502), .ZN(n5489) );
  NAND2_X1 U3914 ( .A1(n3383), .A2(n6504), .ZN(n3377) );
  NAND2_X1 U3915 ( .A1(n3073), .A2(n3077), .ZN(n4229) );
  OAI21_X1 U3916 ( .B1(n5434), .B2(n5435), .A(n5422), .ZN(n5544) );
  INV_X1 U3917 ( .A(n3065), .ZN(n4316) );
  INV_X1 U3918 ( .A(n3273), .ZN(n3270) );
  NOR2_X1 U3919 ( .A1(n5540), .A2(n5652), .ZN(n4312) );
  NAND2_X1 U3920 ( .A1(n3493), .A2(n3492), .ZN(n4180) );
  AND3_X1 U3921 ( .A1(n3188), .A2(n3187), .A3(n3186), .ZN(n3031) );
  AND3_X1 U3922 ( .A1(n3285), .A2(n3284), .A3(n3283), .ZN(n3032) );
  OR2_X2 U3923 ( .A1(n3191), .A2(n3190), .ZN(n4009) );
  AND2_X1 U3924 ( .A1(n2985), .A2(n5343), .ZN(n3033) );
  NOR2_X1 U3926 ( .A1(n3061), .A2(n4326), .ZN(n3034) );
  INV_X1 U3928 ( .A(n3682), .ZN(n3921) );
  NOR2_X1 U3929 ( .A1(n3015), .A2(n6503), .ZN(n3385) );
  NAND2_X1 U3930 ( .A1(n5280), .A2(n3096), .ZN(n5316) );
  NOR2_X1 U3931 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3036)
         );
  NAND2_X1 U3932 ( .A1(n4245), .A2(n4339), .ZN(n3999) );
  INV_X1 U3933 ( .A(n3251), .ZN(n3233) );
  AND2_X1 U3934 ( .A1(n5481), .A2(n3025), .ZN(n3037) );
  NAND2_X1 U3935 ( .A1(n3080), .A2(n4211), .ZN(n5287) );
  NAND2_X1 U3936 ( .A1(n3501), .A2(n4834), .ZN(n4963) );
  OR2_X1 U3937 ( .A1(n5460), .A2(n5459), .ZN(n3038) );
  NAND2_X1 U3938 ( .A1(n5265), .A2(n5266), .ZN(n6125) );
  AND2_X1 U3939 ( .A1(n2985), .A2(n4278), .ZN(n3039) );
  NOR3_X1 U3940 ( .A1(n5460), .A2(n3066), .A3(n3064), .ZN(n5425) );
  NAND2_X1 U3941 ( .A1(n2985), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3040) );
  AND2_X1 U3942 ( .A1(n3719), .A2(n3718), .ZN(n5479) );
  AND2_X1 U3943 ( .A1(n3096), .A2(n3095), .ZN(n3041) );
  AND2_X1 U3944 ( .A1(n3600), .A2(n3588), .ZN(n3042) );
  AND2_X1 U3945 ( .A1(n3782), .A2(n3754), .ZN(n3043) );
  OR2_X1 U3946 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3044) );
  AND2_X1 U3947 ( .A1(n4275), .A2(n4262), .ZN(n6238) );
  INV_X1 U3948 ( .A(n6238), .ZN(n6185) );
  NOR2_X1 U3949 ( .A1(n5987), .A2(n5988), .ZN(n5250) );
  OR2_X1 U3950 ( .A1(n4836), .A2(n3059), .ZN(n3045) );
  AND2_X1 U3951 ( .A1(n2985), .A2(n5303), .ZN(n3046) );
  AND3_X1 U3952 ( .A1(n4101), .A2(n4100), .A3(n4099), .ZN(n5468) );
  NOR3_X1 U3953 ( .A1(n5252), .A2(n3052), .A3(n5278), .ZN(n5320) );
  INV_X1 U3954 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6504) );
  INV_X2 U3955 ( .A(n5622), .ZN(n6149) );
  AND2_X2 U3956 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U3957 ( .A1(n4519), .A2(n4518), .ZN(n4515) );
  XNOR2_X1 U3958 ( .A(n4029), .B(n4448), .ZN(n4495) );
  NAND2_X1 U3959 ( .A1(n4039), .A2(n4038), .ZN(n4516) );
  INV_X1 U3960 ( .A(n4516), .ZN(n3054) );
  INV_X1 U3961 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5643) );
  NOR2_X1 U3962 ( .A1(n5252), .A2(n5278), .ZN(n5277) );
  INV_X1 U3963 ( .A(n5284), .ZN(n3053) );
  NOR2_X2 U3964 ( .A1(n4836), .A2(n3058), .ZN(n5066) );
  NAND2_X1 U3965 ( .A1(n5425), .A2(n5424), .ZN(n3065) );
  INV_X1 U3966 ( .A(n5437), .ZN(n3066) );
  NAND2_X2 U3967 ( .A1(n3067), .A2(n3015), .ZN(n3277) );
  NAND2_X1 U3968 ( .A1(n3234), .A2(n3067), .ZN(n3238) );
  OAI21_X2 U3969 ( .B1(n5342), .B2(n3033), .A(n4215), .ZN(n5634) );
  NAND2_X1 U3970 ( .A1(n4136), .A2(n3275), .ZN(n4142) );
  CLKBUF_X1 U3971 ( .A(n4136), .Z(n3070) );
  NAND2_X1 U3972 ( .A1(n5528), .A2(n3078), .ZN(n3073) );
  NAND2_X1 U3973 ( .A1(n5528), .A2(n4227), .ZN(n5557) );
  OAI21_X1 U3974 ( .B1(n5528), .B2(n3076), .A(n3074), .ZN(n5540) );
  NAND2_X1 U3975 ( .A1(n3364), .A2(n3087), .ZN(n3365) );
  XNOR2_X2 U3976 ( .A(n3363), .B(n3087), .ZN(n3372) );
  OAI21_X2 U3977 ( .B1(n4399), .B2(STATE2_REG_0__SCAN_IN), .A(n3325), .ZN(
        n3087) );
  OAI21_X1 U3978 ( .B1(n4156), .B2(n3406), .A(n3088), .ZN(n3313) );
  NAND3_X1 U3979 ( .A1(n3398), .A2(n6504), .A3(n3297), .ZN(n3088) );
  NAND3_X1 U3980 ( .A1(n3600), .A2(n3588), .A3(n5275), .ZN(n5273) );
  NAND2_X1 U3981 ( .A1(n3089), .A2(n3043), .ZN(n4359) );
  NOR2_X1 U3982 ( .A1(n5422), .A2(n5423), .ZN(n4294) );
  INV_X1 U3983 ( .A(n5422), .ZN(n3102) );
  XNOR2_X1 U3984 ( .A(n4233), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5355)
         );
  NAND2_X1 U3985 ( .A1(n4232), .A2(n4231), .ZN(n4233) );
  XNOR2_X1 U3986 ( .A(n3372), .B(n3371), .ZN(n4136) );
  NAND2_X1 U3987 ( .A1(n3372), .A2(n3370), .ZN(n3366) );
  CLKBUF_X1 U3988 ( .A(n3393), .Z(n3395) );
  NAND2_X2 U3989 ( .A1(n4341), .A2(n4340), .ZN(n6047) );
  INV_X1 U3990 ( .A(READY_N), .ZN(n6708) );
  AND2_X1 U3991 ( .A1(n4255), .A2(n4254), .ZN(n6474) );
  INV_X1 U3992 ( .A(n6474), .ZN(n4293) );
  OR2_X1 U3993 ( .A1(n4297), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6183) );
  OR2_X1 U3994 ( .A1(n6066), .A2(n4131), .ZN(n3103) );
  AND2_X1 U3995 ( .A1(n4132), .A2(n3103), .ZN(n3104) );
  NAND2_X1 U3996 ( .A1(n4190), .A2(n3270), .ZN(n3105) );
  OR2_X1 U3997 ( .A1(n2985), .A2(n4225), .ZN(n3106) );
  OR2_X1 U3998 ( .A1(n3259), .A2(n4529), .ZN(n3107) );
  AND2_X1 U3999 ( .A1(n4005), .A2(n4004), .ZN(n3108) );
  INV_X1 U4000 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3665) );
  NOR2_X1 U4001 ( .A1(n5196), .A2(n4589), .ZN(n3109) );
  AND2_X2 U4002 ( .A1(n4404), .A2(n3117), .ZN(n3193) );
  OR2_X1 U4003 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6811), .ZN(n6579) );
  INV_X1 U4004 ( .A(n3009), .ZN(n3942) );
  AND2_X1 U4005 ( .A1(n3942), .A2(n3941), .ZN(n3962) );
  INV_X1 U4006 ( .A(n3962), .ZN(n3967) );
  OR2_X1 U4007 ( .A1(n4158), .A2(n6605), .ZN(n4159) );
  INV_X1 U4008 ( .A(n4247), .ZN(n3253) );
  AND2_X1 U4009 ( .A1(n3936), .A2(n3935), .ZN(n3938) );
  INV_X1 U4010 ( .A(n5467), .ZN(n3782) );
  INV_X1 U4011 ( .A(n5318), .ZN(n3631) );
  OR2_X1 U4012 ( .A1(n3480), .A2(n3479), .ZN(n4193) );
  INV_X1 U4013 ( .A(n5633), .ZN(n4216) );
  OR2_X1 U4014 ( .A1(n2985), .A2(n6164), .ZN(n4210) );
  OR2_X1 U4015 ( .A1(n3417), .A2(n3416), .ZN(n4164) );
  INV_X1 U4016 ( .A(n3901), .ZN(n3904) );
  INV_X1 U4017 ( .A(n3715), .ZN(n3716) );
  NAND2_X1 U4018 ( .A1(n5367), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3924) );
  INV_X1 U4019 ( .A(n3385), .ZN(n3682) );
  INV_X1 U4020 ( .A(n3498), .ZN(n3499) );
  INV_X1 U4021 ( .A(n3384), .ZN(n3444) );
  AND2_X1 U4022 ( .A1(n6126), .A2(n4210), .ZN(n4211) );
  INV_X1 U4023 ( .A(n4109), .ZN(n4116) );
  INV_X1 U4024 ( .A(n3972), .ZN(n3965) );
  AND2_X1 U4025 ( .A1(n6251), .A2(n3291), .ZN(n4593) );
  NOR2_X1 U4026 ( .A1(n3749), .A2(n5590), .ZN(n3750) );
  OR2_X1 U4027 ( .A1(n3626), .A2(n5959), .ZN(n3633) );
  OR2_X1 U4028 ( .A1(n3865), .A2(n3864), .ZN(n3901) );
  NOR2_X1 U4029 ( .A1(n3542), .A2(n5993), .ZN(n3546) );
  AND2_X1 U4030 ( .A1(n2985), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5527)
         );
  OR2_X1 U4031 ( .A1(n2985), .A2(n4221), .ZN(n4222) );
  OAI211_X1 U4032 ( .C1(n3965), .C2(n4692), .A(n3357), .B(n3356), .ZN(n3380)
         );
  AOI21_X1 U4033 ( .B1(n4543), .B2(n4545), .A(n6491), .ZN(n4595) );
  INV_X1 U4034 ( .A(n3370), .ZN(n3371) );
  NOR2_X1 U4035 ( .A1(n4593), .A2(n6503), .ZN(n5197) );
  NAND2_X1 U4036 ( .A1(n3979), .A2(n3978), .ZN(n3982) );
  AND2_X1 U4037 ( .A1(n5782), .A2(n5380), .ZN(n5429) );
  AND2_X1 U4038 ( .A1(n3838), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3839)
         );
  NAND2_X1 U4039 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5335), .ZN(n5838) );
  INV_X1 U4040 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5959) );
  INV_X1 U4041 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5993) );
  AND2_X1 U4042 ( .A1(n5362), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4358) );
  OR2_X1 U4043 ( .A1(n5239), .A2(n5240), .ZN(n5248) );
  NAND2_X1 U4044 ( .A1(n4291), .A2(n5643), .ZN(n4231) );
  NAND2_X1 U4045 ( .A1(n4229), .A2(n5527), .ZN(n5533) );
  OR2_X1 U4046 ( .A1(n5184), .A2(n4500), .ZN(n6242) );
  OR2_X1 U4047 ( .A1(n4437), .A2(n4250), .ZN(n4251) );
  INV_X1 U4048 ( .A(n6254), .ZN(n6385) );
  OR2_X1 U4049 ( .A1(n4397), .A2(n4396), .ZN(n6458) );
  AND2_X1 U4050 ( .A1(n5019), .A2(n5018), .ZN(n5043) );
  OR2_X1 U4051 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4908), .ZN(n6299)
         );
  NOR2_X1 U4052 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4595), .ZN(n4738) );
  OR2_X1 U4053 ( .A1(n5769), .A2(n5194), .ZN(n5232) );
  INV_X1 U4054 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6252) );
  AND2_X1 U4055 ( .A1(n5094), .A2(n5093), .ZN(n5142) );
  INV_X1 U4056 ( .A(DATAI_23_), .ZN(n6717) );
  INV_X1 U4057 ( .A(DATAI_19_), .ZN(n6679) );
  OR2_X1 U4058 ( .A1(n4710), .A2(n5009), .ZN(n4719) );
  INV_X1 U4059 ( .A(n2986), .ZN(n6605) );
  OAI211_X1 U4060 ( .C1(n6688), .C2(n5391), .A(n5390), .B(n5389), .ZN(n5392)
         );
  NOR2_X1 U4061 ( .A1(n5780), .A2(n5376), .ZN(n5441) );
  INV_X1 U4062 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4342) );
  AND2_X1 U4063 ( .A1(n4086), .A2(n4085), .ZN(n5494) );
  INV_X1 U4064 ( .A(n6038), .ZN(n5989) );
  OR3_X1 U4065 ( .A1(n6601), .A2(n6221), .A3(n4333), .ZN(n6020) );
  INV_X1 U4066 ( .A(n5313), .ZN(n5500) );
  INV_X1 U4067 ( .A(n5498), .ZN(n6063) );
  INV_X1 U4068 ( .A(n5512), .ZN(n6073) );
  OAI21_X1 U4069 ( .B1(n2986), .B2(n6708), .A(n4455), .ZN(n6118) );
  OR2_X1 U4070 ( .A1(n3999), .A2(n4000), .ZN(n4389) );
  INV_X1 U4071 ( .A(n5598), .ZN(n5863) );
  INV_X1 U4072 ( .A(n4382), .ZN(n4301) );
  OR2_X1 U4073 ( .A1(n5699), .A2(n4286), .ZN(n5691) );
  NAND2_X1 U4074 ( .A1(n5184), .A2(n6211), .ZN(n6202) );
  NAND2_X1 U4075 ( .A1(n4252), .A2(n4251), .ZN(n4275) );
  INV_X1 U4076 ( .A(n4671), .ZN(n4701) );
  OAI21_X1 U4077 ( .B1(n6264), .B2(n6261), .A(n6260), .ZN(n6289) );
  NAND2_X1 U4078 ( .A1(n4806), .A2(n4805), .ZN(n6302) );
  OAI21_X1 U4079 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6589), .A(n4738), 
        .ZN(n6389) );
  OAI21_X1 U4080 ( .B1(n6315), .B2(n6314), .A(n6313), .ZN(n6355) );
  OR2_X1 U4081 ( .A1(n4852), .A2(n4851), .ZN(n6376) );
  INV_X1 U4082 ( .A(n4980), .ZN(n5005) );
  NOR2_X1 U4083 ( .A1(n6386), .A2(n5009), .ZN(n5081) );
  INV_X1 U4084 ( .A(n6414), .ZN(n6329) );
  AND2_X1 U4085 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5086), .ZN(n4629)
         );
  NOR2_X1 U4086 ( .A1(n5622), .A2(n4620), .ZN(n6345) );
  NOR2_X1 U4087 ( .A1(n6648), .A2(n4849), .ZN(n6448) );
  NOR2_X1 U4088 ( .A1(n5622), .A2(n4612), .ZN(n6325) );
  INV_X1 U4089 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6493) );
  INV_X1 U4090 ( .A(n6575), .ZN(n6577) );
  OR2_X1 U4091 ( .A1(n4437), .A2(n3999), .ZN(n4454) );
  INV_X1 U4092 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5923) );
  INV_X1 U4093 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U4094 ( .A1(n6020), .A2(n4363), .ZN(n6038) );
  AND2_X1 U4095 ( .A1(n5100), .A2(n6038), .ZN(n6052) );
  NAND2_X1 U4096 ( .A1(n5353), .A2(n6063), .ZN(n4133) );
  NAND2_X1 U4097 ( .A1(n6066), .A2(n3015), .ZN(n5498) );
  INV_X1 U4098 ( .A(n6063), .ZN(n5844) );
  OR2_X1 U4099 ( .A1(n5057), .A2(n5059), .ZN(n5999) );
  INV_X1 U4100 ( .A(n6139), .ZN(n6039) );
  NAND2_X1 U4101 ( .A1(n4438), .A2(n4339), .ZN(n4562) );
  OR3_X1 U4102 ( .A1(n4437), .A2(n4436), .A3(n6518), .ZN(n6108) );
  INV_X1 U4103 ( .A(DATAI_6_), .ZN(n6782) );
  OR2_X1 U4104 ( .A1(n4437), .A2(n4389), .ZN(n6124) );
  AND2_X1 U4105 ( .A1(n4269), .A2(n4268), .ZN(n5882) );
  INV_X1 U4106 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U4107 ( .A1(n4275), .A2(n4261), .ZN(n6169) );
  OAI21_X1 U4108 ( .B1(n4544), .B2(n6586), .A(n4849), .ZN(n6249) );
  INV_X1 U4109 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5913) );
  INV_X1 U4110 ( .A(n4672), .ZN(n4704) );
  OR2_X1 U4111 ( .A1(n4651), .A2(n4912), .ZN(n4671) );
  NAND2_X1 U4112 ( .A1(n5010), .A2(n5009), .ZN(n6286) );
  NAND2_X1 U4113 ( .A1(n5010), .A2(n4912), .ZN(n6305) );
  AOI211_X2 U4114 ( .C1(n4908), .C2(n6390), .A(n6389), .B(n4906), .ZN(n4952)
         );
  NAND2_X1 U4115 ( .A1(n4913), .A2(n4912), .ZN(n5237) );
  AOI22_X1 U4116 ( .A1(n6311), .A2(n6314), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3400), .ZN(n6359) );
  OR2_X1 U4117 ( .A1(n5769), .A2(n4845), .ZN(n6379) );
  NAND2_X1 U4118 ( .A1(n5081), .A2(n4874), .ZN(n4980) );
  INV_X1 U4119 ( .A(n6396), .ZN(n6319) );
  INV_X1 U4120 ( .A(n6431), .ZN(n6342) );
  NAND2_X1 U4121 ( .A1(n4972), .A2(n5193), .ZN(n6452) );
  INV_X1 U4122 ( .A(n6345), .ZN(n6441) );
  NAND2_X1 U4123 ( .A1(n6149), .A2(DATAI_18_), .ZN(n6413) );
  INV_X1 U4124 ( .A(n6339), .ZN(n6429) );
  INV_X1 U4125 ( .A(n6321), .ZN(n6401) );
  OR2_X1 U4126 ( .A1(n4710), .A2(n4912), .ZN(n4792) );
  INV_X1 U4127 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6589) );
  NOR2_X1 U4128 ( .A1(n6812), .A2(n5921), .ZN(n6585) );
  INV_X1 U4129 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6555) );
  INV_X1 U4130 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U4131 ( .A1(n4133), .A2(n3104), .ZN(U2829) );
  AND2_X2 U4132 ( .A1(n4522), .A2(n3118), .ZN(n3869) );
  AOI22_X1 U4133 ( .A1(n3194), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4134 ( .A1(n3179), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4135 ( .A1(n3177), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3113) );
  AND2_X4 U4136 ( .A1(n4403), .A2(n3117), .ZN(n3184) );
  AOI22_X1 U4137 ( .A1(n3184), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3122) );
  AND2_X2 U4138 ( .A1(n4522), .A2(n4414), .ZN(n3348) );
  AOI22_X1 U4139 ( .A1(n3348), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4140 ( .A1(n3411), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3120) );
  AND2_X2 U4141 ( .A1(n3118), .A2(n4536), .ZN(n3199) );
  AOI22_X1 U4142 ( .A1(n3013), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3119) );
  INV_X1 U4143 ( .A(n3251), .ZN(n3135) );
  AOI22_X1 U4144 ( .A1(n3411), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4145 ( .A1(n3013), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4146 ( .A1(n3194), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U4147 ( .A1(n3304), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4148 ( .A1(n3411), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4149 ( .A1(n3348), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3138)
         );
  NAND2_X1 U4150 ( .A1(n3185), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U4151 ( .A1(n3222), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3136)
         );
  NAND2_X1 U4152 ( .A1(n3194), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3145)
         );
  NAND2_X1 U4153 ( .A1(n3017), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U4154 ( .A1(n3869), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U4155 ( .A1(n3006), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3142)
         );
  NAND2_X1 U4156 ( .A1(n3177), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3149)
         );
  NAND2_X1 U4157 ( .A1(n3019), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4158 ( .A1(n3193), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U4159 ( .A1(n3008), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4160 ( .A1(n3199), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3153)
         );
  NAND2_X1 U4161 ( .A1(n3150), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4162 ( .A1(n3184), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4163 ( .A1(n3020), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4164 ( .A1(n3022), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4165 ( .A1(n3177), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4166 ( .A1(n3016), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3158) );
  NAND4_X1 U4167 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3167)
         );
  AOI22_X1 U4168 ( .A1(n3411), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4169 ( .A1(n3348), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4170 ( .A1(n3184), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4171 ( .A1(n3304), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3162) );
  NAND4_X1 U4172 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3166)
         );
  INV_X1 U4173 ( .A(n3272), .ZN(n3192) );
  AOI22_X1 U4174 ( .A1(n3411), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4175 ( .A1(n3019), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4176 ( .A1(n3194), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4177 ( .A1(n3177), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3008), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4178 ( .A1(n3013), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4179 ( .A1(n3017), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4180 ( .A1(n3185), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4181 ( .A1(n3199), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4182 ( .A1(n3022), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4183 ( .A1(n3179), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4184 ( .A1(n3017), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3180) );
  NAND4_X1 U4185 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3191)
         );
  AOI22_X1 U4186 ( .A1(n3184), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4187 ( .A1(n3411), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4188 ( .A1(n3013), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4189 ( .A1(n3348), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4190 ( .A1(n3189), .A2(n3031), .ZN(n3190) );
  NAND2_X1 U4192 ( .A1(n3192), .A2(n3247), .ZN(n3983) );
  INV_X1 U4193 ( .A(n3983), .ZN(n3232) );
  NAND2_X1 U4194 ( .A1(n3193), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4195 ( .A1(n3020), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4196 ( .A1(n3194), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4197 ( .A1(n3869), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4198 ( .A1(n3013), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4199 ( .A1(n3411), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4200 ( .A1(n3185), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4201 ( .A1(n3199), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3200)
         );
  NAND2_X1 U4202 ( .A1(n3184), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4203 ( .A1(n3348), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3206)
         );
  NAND2_X1 U4204 ( .A1(n3222), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4205 ( .A1(n3006), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3204)
         );
  NAND2_X1 U4206 ( .A1(n3017), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4207 ( .A1(n3177), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3210)
         );
  NAND2_X1 U4208 ( .A1(n3150), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4209 ( .A1(n3008), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3208) );
  NAND4_X4 U4210 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n4339)
         );
  NAND2_X1 U4211 ( .A1(n3277), .A2(n3216), .ZN(n4006) );
  AOI22_X1 U4212 ( .A1(n3022), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4213 ( .A1(n3179), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4214 ( .A1(n3177), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4215 ( .A1(n3016), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4216 ( .A1(n3411), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4217 ( .A1(n3184), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3224) );
  NAND2_X4 U4218 ( .A1(n3227), .A2(n3029), .ZN(n3275) );
  XNOR2_X1 U4219 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3255) );
  INV_X1 U4220 ( .A(n3255), .ZN(n4235) );
  OAI21_X1 U4221 ( .B1(n4235), .B2(n3275), .A(n3235), .ZN(n3229) );
  NAND2_X1 U4222 ( .A1(n3277), .A2(n3279), .ZN(n3230) );
  AND4_X2 U4223 ( .A1(n3232), .A2(n4006), .A3(n3231), .A4(n3230), .ZN(n3243)
         );
  MUX2_X1 U4224 ( .A(n3010), .B(n3235), .S(n3251), .Z(n3236) );
  NAND2_X1 U4225 ( .A1(n3236), .A2(n4391), .ZN(n3237) );
  NAND2_X1 U4226 ( .A1(n3238), .A2(n3237), .ZN(n3241) );
  NAND2_X1 U4227 ( .A1(n3239), .A2(n4009), .ZN(n3278) );
  AND3_X1 U4228 ( .A1(n3278), .A2(n4246), .A3(n3015), .ZN(n3240) );
  NAND2_X1 U4229 ( .A1(n3241), .A2(n3240), .ZN(n3268) );
  NAND2_X1 U4230 ( .A1(n3268), .A2(n4240), .ZN(n3242) );
  NAND2_X1 U4231 ( .A1(n3244), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3262) );
  INV_X1 U4232 ( .A(n4297), .ZN(n3263) );
  XNOR2_X1 U4233 ( .A(n6455), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5196)
         );
  INV_X1 U4234 ( .A(n3997), .ZN(n3264) );
  AND2_X1 U4235 ( .A1(n3264), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3245)
         );
  AOI21_X1 U4236 ( .B1(n3263), .B2(n5196), .A(n3245), .ZN(n3258) );
  NOR2_X1 U4237 ( .A1(n4609), .A2(n3010), .ZN(n3246) );
  NAND3_X1 U4238 ( .A1(n3278), .A2(n3635), .A3(n3249), .ZN(n3248) );
  NAND2_X1 U4239 ( .A1(n4239), .A2(n3009), .ZN(n3985) );
  OAI21_X1 U4240 ( .B1(n3999), .B2(n4246), .A(n3985), .ZN(n4256) );
  NAND3_X1 U4241 ( .A1(n3009), .A2(n3235), .A3(n4019), .ZN(n3995) );
  INV_X1 U4242 ( .A(n3995), .ZN(n3254) );
  NAND2_X1 U4243 ( .A1(n4621), .A2(n3015), .ZN(n4247) );
  NAND2_X1 U4244 ( .A1(n3254), .A2(n3253), .ZN(n4257) );
  OAI21_X1 U4245 ( .B1(n3999), .B2(n3255), .A(n4257), .ZN(n3256) );
  OAI21_X1 U4246 ( .B1(n4256), .B2(n3256), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3257) );
  OAI211_X1 U4247 ( .C1(n3262), .C2(n3112), .A(n3258), .B(n3257), .ZN(n3287)
         );
  INV_X1 U4248 ( .A(n3257), .ZN(n3260) );
  INV_X1 U4249 ( .A(n3258), .ZN(n3259) );
  NAND2_X1 U4250 ( .A1(n3260), .A2(n3107), .ZN(n3261) );
  NAND2_X1 U4251 ( .A1(n3287), .A2(n3261), .ZN(n3314) );
  INV_X1 U4252 ( .A(n3314), .ZN(n3286) );
  NAND2_X1 U4253 ( .A1(n3003), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3267) );
  MUX2_X1 U4254 ( .A(n3264), .B(n3263), .S(n6455), .Z(n3265) );
  INV_X1 U4255 ( .A(n3265), .ZN(n3266) );
  NAND2_X1 U4256 ( .A1(n3267), .A2(n3266), .ZN(n3326) );
  AND2_X1 U4257 ( .A1(n3105), .A2(n4240), .ZN(n3271) );
  NAND2_X1 U4258 ( .A1(n3268), .A2(n3271), .ZN(n4015) );
  NAND2_X1 U4259 ( .A1(n2999), .A2(n3004), .ZN(n3274) );
  NAND2_X1 U4260 ( .A1(n3274), .A2(n4009), .ZN(n3276) );
  OAI21_X1 U4261 ( .B1(n3272), .B2(n3276), .A(n3275), .ZN(n3285) );
  OAI21_X1 U4262 ( .B1(n3277), .B2(n3278), .A(n2986), .ZN(n3284) );
  NOR2_X1 U4263 ( .A1(n5777), .A2(n6504), .ZN(n6502) );
  NAND2_X1 U4264 ( .A1(n3249), .A2(n4339), .ZN(n3282) );
  NAND2_X1 U4265 ( .A1(n4015), .A2(n3032), .ZN(n3327) );
  NAND2_X2 U4266 ( .A1(n3326), .A2(n3327), .ZN(n3330) );
  NAND2_X1 U4267 ( .A1(n3286), .A2(n3330), .ZN(n3288) );
  NAND2_X1 U4268 ( .A1(n3288), .A2(n3287), .ZN(n3296) );
  INV_X1 U4269 ( .A(n3296), .ZN(n3294) );
  NAND2_X1 U4270 ( .A1(n3289), .A2(n6466), .ZN(n6251) );
  INV_X1 U4271 ( .A(n3289), .ZN(n3290) );
  NAND2_X1 U4272 ( .A1(n3290), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3291) );
  OAI22_X1 U4273 ( .A1(n4593), .A2(n4297), .B1(n3997), .B2(n6466), .ZN(n3292)
         );
  AOI21_X1 U4274 ( .B1(n3399), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3292), 
        .ZN(n3295) );
  INV_X1 U4275 ( .A(n3295), .ZN(n3293) );
  NAND2_X1 U4276 ( .A1(n3296), .A2(n3295), .ZN(n3297) );
  AOI22_X1 U4277 ( .A1(n3179), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4278 ( .A1(n3022), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4279 ( .A1(n3177), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4280 ( .A1(n3017), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3299) );
  NAND4_X1 U4281 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3310)
         );
  BUF_X1 U4282 ( .A(n3411), .Z(n3303) );
  AOI22_X1 U4283 ( .A1(n3303), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4284 ( .A1(n3874), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4285 ( .A1(n3184), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4286 ( .A1(n3021), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3305) );
  NAND4_X1 U4287 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3309)
         );
  INV_X1 U4288 ( .A(n3405), .ZN(n3360) );
  AOI22_X1 U4289 ( .A1(n3972), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3360), 
        .B2(n3311), .ZN(n3312) );
  XNOR2_X1 U4290 ( .A(n3314), .B(n3330), .ZN(n4399) );
  INV_X1 U4291 ( .A(n3406), .ZN(n3358) );
  AOI22_X1 U4292 ( .A1(n3020), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4293 ( .A1(n3021), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4294 ( .A1(n3018), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4295 ( .A1(n3177), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3315) );
  NAND4_X1 U4296 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3324)
         );
  AOI22_X1 U4297 ( .A1(n3017), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4298 ( .A1(n3411), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4299 ( .A1(n3150), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4300 ( .A1(n3184), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3319) );
  NAND4_X1 U4301 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3323)
         );
  NAND2_X1 U4302 ( .A1(n3358), .A2(n4137), .ZN(n3325) );
  INV_X1 U4303 ( .A(n3326), .ZN(n3329) );
  INV_X1 U4304 ( .A(n3327), .ZN(n3328) );
  AOI22_X1 U4305 ( .A1(n3177), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4306 ( .A1(n3017), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4307 ( .A1(n3303), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4308 ( .A1(n3150), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3334) );
  NAND4_X1 U4309 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3343)
         );
  AOI22_X1 U4310 ( .A1(n2987), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4311 ( .A1(n3185), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4312 ( .A1(n3020), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4313 ( .A1(n3194), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4314 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3342)
         );
  AOI22_X1 U4315 ( .A1(n3179), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4316 ( .A1(n3022), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4317 ( .A1(n3011), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4318 ( .A1(n3017), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3344) );
  NAND4_X1 U4319 ( .A1(n3347), .A2(n3346), .A3(n3345), .A4(n3344), .ZN(n3354)
         );
  AOI22_X1 U4320 ( .A1(n3303), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4321 ( .A1(n3874), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4322 ( .A1(n3184), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4323 ( .A1(n2987), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3349) );
  NAND4_X1 U4324 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3353)
         );
  XNOR2_X1 U4325 ( .A(n4202), .B(n4145), .ZN(n3355) );
  NOR2_X1 U4326 ( .A1(n3355), .A2(n3406), .ZN(n3378) );
  INV_X1 U4327 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4692) );
  AOI21_X1 U4328 ( .B1(n3270), .B2(n4202), .A(n6504), .ZN(n3357) );
  NAND2_X1 U4329 ( .A1(n4240), .A2(n4145), .ZN(n3356) );
  AOI22_X1 U4330 ( .A1(n3378), .A2(n3380), .B1(n3358), .B2(n4202), .ZN(n3359)
         );
  AND2_X2 U4331 ( .A1(n3377), .A2(n3359), .ZN(n3363) );
  NAND2_X1 U4332 ( .A1(n3972), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U4333 ( .A1(n3360), .A2(n4137), .ZN(n3361) );
  INV_X1 U4334 ( .A(n3363), .ZN(n3364) );
  NAND2_X2 U4335 ( .A1(n3369), .A2(n3002), .ZN(n4585) );
  NAND2_X1 U4336 ( .A1(n6503), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3801) );
  OAI21_X2 U4337 ( .B1(n4585), .B2(n3614), .A(n3801), .ZN(n3393) );
  INV_X1 U4338 ( .A(n3393), .ZN(n3390) );
  NAND2_X1 U4339 ( .A1(n4136), .A2(n3623), .ZN(n3376) );
  AOI22_X1 U4340 ( .A1(n3921), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6503), .ZN(n3374) );
  AND2_X1 U4341 ( .A1(n3253), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4342 ( .A1(n3384), .A2(n4529), .ZN(n3373) );
  AND2_X1 U4343 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  NAND2_X1 U4344 ( .A1(n3376), .A2(n3375), .ZN(n4493) );
  INV_X1 U4345 ( .A(n3378), .ZN(n3379) );
  XNOR2_X1 U4346 ( .A(n3380), .B(n3379), .ZN(n3381) );
  NAND2_X1 U4347 ( .A1(n5009), .A2(n3280), .ZN(n3382) );
  NAND2_X1 U4348 ( .A1(n3382), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U4349 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6503), .ZN(n3387)
         );
  NAND2_X1 U4350 ( .A1(n3385), .A2(EAX_REG_0__SCAN_IN), .ZN(n3386) );
  OAI211_X1 U4351 ( .C1(n3444), .C2(n5375), .A(n3387), .B(n3386), .ZN(n3388)
         );
  AOI21_X1 U4352 ( .B1(n3383), .B2(n3623), .A(n3388), .ZN(n4377) );
  OR2_X1 U4353 ( .A1(n4378), .A2(n4377), .ZN(n4380) );
  NAND2_X1 U4354 ( .A1(n4377), .A2(n3920), .ZN(n3389) );
  NAND2_X1 U4355 ( .A1(n4380), .A2(n3389), .ZN(n4494) );
  NAND2_X1 U4356 ( .A1(n3390), .A2(n4492), .ZN(n4509) );
  INV_X2 U4357 ( .A(n3044), .ZN(n3920) );
  NAND2_X1 U4358 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3422) );
  OAI21_X1 U4359 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3422), .ZN(n6161) );
  AOI22_X1 U4360 ( .A1(n5357), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3920), 
        .B2(n6161), .ZN(n3392) );
  NAND2_X1 U4361 ( .A1(n3921), .A2(EAX_REG_2__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4362 ( .A1(n4509), .A2(n4510), .ZN(n3397) );
  INV_X1 U4363 ( .A(n4492), .ZN(n3394) );
  NAND2_X1 U4364 ( .A1(n3395), .A2(n3394), .ZN(n3396) );
  NAND2_X1 U4365 ( .A1(n3399), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3404) );
  NAND3_X1 U4366 ( .A1(n6252), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6312) );
  INV_X1 U4367 ( .A(n6312), .ZN(n3400) );
  NAND2_X1 U4368 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3400), .ZN(n6343) );
  NAND2_X1 U4369 ( .A1(n6252), .A2(n6343), .ZN(n3401) );
  NAND3_X1 U4370 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4739) );
  NAND2_X1 U4371 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4712), .ZN(n4787) );
  NAND2_X1 U4372 ( .A1(n3401), .A2(n4787), .ZN(n4848) );
  OAI22_X1 U4373 ( .A1(n4297), .A2(n4848), .B1(n3997), .B2(n6252), .ZN(n3402)
         );
  INV_X1 U4374 ( .A(n3402), .ZN(n3403) );
  NAND2_X1 U4375 ( .A1(n4521), .A2(n6504), .ZN(n3419) );
  AOI22_X1 U4376 ( .A1(n3020), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4377 ( .A1(n3194), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4378 ( .A1(n3177), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4379 ( .A1(n3017), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3407) );
  NAND4_X1 U4380 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3417)
         );
  AOI22_X1 U4381 ( .A1(n3303), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4382 ( .A1(n3874), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4383 ( .A1(n3184), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4384 ( .A1(n3021), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3412) );
  NAND4_X1 U4385 ( .A1(n3415), .A2(n3414), .A3(n3413), .A4(n3412), .ZN(n3416)
         );
  AOI22_X1 U4386 ( .A1(n3980), .A2(n4164), .B1(n3972), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4387 ( .A1(n3002), .A2(n4795), .ZN(n3421) );
  INV_X1 U4388 ( .A(n3422), .ZN(n3423) );
  NAND2_X1 U4389 ( .A1(n3423), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3440)
         );
  OAI21_X1 U4390 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3423), .A(n3440), 
        .ZN(n6152) );
  AOI22_X1 U4391 ( .A1(n3920), .A2(n6152), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4392 ( .A1(n3921), .A2(EAX_REG_3__SCAN_IN), .ZN(n3424) );
  OAI211_X1 U4393 ( .C1(n3444), .C2(n3111), .A(n3425), .B(n3424), .ZN(n3426)
         );
  INV_X1 U4394 ( .A(n3426), .ZN(n3427) );
  OAI21_X1 U4395 ( .B1(n4586), .B2(n3614), .A(n3427), .ZN(n4513) );
  NAND2_X1 U4396 ( .A1(n4508), .A2(n4513), .ZN(n4512) );
  INV_X1 U4397 ( .A(n4512), .ZN(n3449) );
  AOI22_X1 U4398 ( .A1(n3179), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4399 ( .A1(n3022), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4400 ( .A1(n3177), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4401 ( .A1(n3017), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4402 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3437)
         );
  AOI22_X1 U4403 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3411), .B1(n3018), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4404 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3333), .B1(n3874), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4405 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3184), .B1(n3875), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4406 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3021), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4407 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3436)
         );
  NAND2_X1 U4408 ( .A1(n3980), .A2(n4172), .ZN(n3439) );
  NAND2_X1 U4409 ( .A1(n3972), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3438) );
  NAND2_X1 U4410 ( .A1(n4163), .A2(n3623), .ZN(n3447) );
  INV_X1 U4411 ( .A(n3440), .ZN(n3441) );
  NAND2_X1 U4412 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3441), .ZN(n3484)
         );
  OAI21_X1 U4413 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3441), .A(n3484), 
        .ZN(n5166) );
  OAI21_X1 U4414 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n5923), .A(n6503), 
        .ZN(n3443) );
  NAND2_X1 U4415 ( .A1(n3921), .A2(EAX_REG_4__SCAN_IN), .ZN(n3442) );
  OAI211_X1 U4416 ( .C1(n3444), .C2(n5913), .A(n3443), .B(n3442), .ZN(n3445)
         );
  OAI21_X1 U4417 ( .B1(n3044), .B2(n5166), .A(n3445), .ZN(n3446) );
  NAND2_X1 U4418 ( .A1(n3449), .A2(n3448), .ZN(n4632) );
  AOI22_X1 U4419 ( .A1(n3019), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4420 ( .A1(n3022), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4421 ( .A1(n3011), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4422 ( .A1(n3017), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4423 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3462)
         );
  AOI22_X1 U4424 ( .A1(n3303), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4425 ( .A1(n3874), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4426 ( .A1(n3184), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4427 ( .A1(n3021), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3457) );
  NAND4_X1 U4428 ( .A1(n3460), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(n3461)
         );
  NAND2_X1 U4429 ( .A1(n3980), .A2(n4183), .ZN(n3464) );
  NAND2_X1 U4430 ( .A1(n3972), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3463) );
  NAND2_X1 U4431 ( .A1(n3464), .A2(n3463), .ZN(n3468) );
  XNOR2_X1 U4432 ( .A(n3470), .B(n3468), .ZN(n4171) );
  INV_X1 U4433 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3466) );
  XNOR2_X1 U4434 ( .A(n3483), .B(n3484), .ZN(n6053) );
  AOI22_X1 U4435 ( .A1(n6053), .A2(n3920), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3465) );
  OAI21_X1 U4436 ( .B1(n3682), .B2(n3466), .A(n3465), .ZN(n3467) );
  AOI21_X1 U4437 ( .B1(n4171), .B2(n3623), .A(n3467), .ZN(n4724) );
  INV_X1 U4438 ( .A(n3468), .ZN(n3469) );
  AOI22_X1 U4439 ( .A1(n3020), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4440 ( .A1(n3194), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4441 ( .A1(n3177), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4442 ( .A1(n3017), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3471) );
  NAND4_X1 U4443 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3480)
         );
  AOI22_X1 U4444 ( .A1(n3411), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4445 ( .A1(n3874), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4446 ( .A1(n3184), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4447 ( .A1(n3021), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3475) );
  NAND4_X1 U4448 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3479)
         );
  AOI22_X1 U4449 ( .A1(n3980), .A2(n4193), .B1(n3972), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U4450 ( .A1(n3481), .A2(n3491), .ZN(n4181) );
  NAND2_X1 U4451 ( .A1(n4181), .A2(n3623), .ZN(n3490) );
  INV_X1 U4452 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6037) );
  AOI21_X1 U4453 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6037), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3482) );
  AOI21_X1 U4454 ( .B1(n3921), .B2(EAX_REG_6__SCAN_IN), .A(n3482), .ZN(n3488)
         );
  NOR2_X1 U4455 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  NOR2_X1 U4456 ( .A1(n3485), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3486)
         );
  OR2_X1 U4457 ( .A1(n3512), .A2(n3486), .ZN(n6142) );
  NOR2_X1 U4458 ( .A1(n6142), .A2(n3044), .ZN(n3487) );
  OR2_X1 U4459 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  NAND2_X1 U4460 ( .A1(n3490), .A2(n3489), .ZN(n4839) );
  NAND2_X1 U4461 ( .A1(n4723), .A2(n4839), .ZN(n4833) );
  INV_X1 U4462 ( .A(n3491), .ZN(n3492) );
  INV_X1 U4463 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3495) );
  NAND2_X1 U4464 ( .A1(n3980), .A2(n4202), .ZN(n3494) );
  OAI21_X1 U4465 ( .B1(n3495), .B2(n3965), .A(n3494), .ZN(n3496) );
  XNOR2_X1 U4466 ( .A(n4180), .B(n3496), .ZN(n4191) );
  NAND2_X1 U4467 ( .A1(n4191), .A2(n3623), .ZN(n3500) );
  INV_X1 U4468 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4954) );
  XNOR2_X1 U4469 ( .A(n3512), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6025) );
  AOI22_X1 U4470 ( .A1(n6025), .A2(n3920), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3497) );
  OAI21_X1 U4471 ( .B1(n3682), .B2(n4954), .A(n3497), .ZN(n3498) );
  AOI22_X1 U4472 ( .A1(n3874), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4473 ( .A1(n3332), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4474 ( .A1(n3184), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4475 ( .A1(n3851), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3502) );
  NAND4_X1 U4476 ( .A1(n3505), .A2(n3504), .A3(n3503), .A4(n3502), .ZN(n3511)
         );
  AOI22_X1 U4477 ( .A1(n3017), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4478 ( .A1(n3411), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4479 ( .A1(n3019), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4480 ( .A1(n3021), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3506) );
  NAND4_X1 U4481 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n3510)
         );
  OAI21_X1 U4482 ( .B1(n3511), .B2(n3510), .A(n3623), .ZN(n3517) );
  NAND2_X1 U4483 ( .A1(n3921), .A2(EAX_REG_8__SCAN_IN), .ZN(n3516) );
  INV_X1 U4484 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3513) );
  XNOR2_X1 U4485 ( .A(n3518), .B(n3513), .ZN(n6008) );
  OR2_X1 U4486 ( .A1(n6008), .A2(n3044), .ZN(n3515) );
  NAND2_X1 U4487 ( .A1(n5357), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3514)
         );
  NAND2_X1 U4488 ( .A1(n3518), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3542)
         );
  XNOR2_X1 U4489 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3542), .ZN(n5997) );
  AOI22_X1 U4490 ( .A1(n3017), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4491 ( .A1(n3018), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4492 ( .A1(n3020), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4493 ( .A1(n3021), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4494 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3528)
         );
  AOI22_X1 U4495 ( .A1(n3011), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4496 ( .A1(n3411), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4497 ( .A1(n3022), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4498 ( .A1(n3184), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3523) );
  NAND4_X1 U4499 ( .A1(n3526), .A2(n3525), .A3(n3524), .A4(n3523), .ZN(n3527)
         );
  OR2_X1 U4500 ( .A1(n3528), .A2(n3527), .ZN(n3529) );
  AOI22_X1 U4501 ( .A1(n3623), .A2(n3529), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4502 ( .A1(n3921), .A2(EAX_REG_9__SCAN_IN), .ZN(n3530) );
  OAI211_X1 U4503 ( .C1(n5997), .C2(n3044), .A(n3531), .B(n3530), .ZN(n5058)
         );
  AOI22_X1 U4504 ( .A1(n3179), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3011), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4505 ( .A1(n3021), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4506 ( .A1(n3018), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4507 ( .A1(n3332), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3532) );
  NAND4_X1 U4508 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3541)
         );
  AOI22_X1 U4509 ( .A1(n3017), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4510 ( .A1(n3303), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4511 ( .A1(n3194), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4512 ( .A1(n3150), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4513 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3540)
         );
  NOR2_X1 U4514 ( .A1(n3541), .A2(n3540), .ZN(n3545) );
  XNOR2_X1 U4515 ( .A(n3546), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5268)
         );
  NAND2_X1 U4516 ( .A1(n5268), .A2(n3920), .ZN(n3544) );
  AOI22_X1 U4517 ( .A1(n3921), .A2(EAX_REG_10__SCAN_IN), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3543) );
  OAI211_X1 U4518 ( .C1(n3545), .C2(n3614), .A(n3544), .B(n3543), .ZN(n5063)
         );
  NAND2_X1 U4519 ( .A1(n3546), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3562)
         );
  XNOR2_X1 U4520 ( .A(n3580), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5291)
         );
  AOI22_X1 U4521 ( .A1(n3017), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4522 ( .A1(n3021), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4523 ( .A1(n3177), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4524 ( .A1(n3150), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4525 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3557)
         );
  AOI22_X1 U4526 ( .A1(n3019), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4527 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3303), .B1(n3018), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4528 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3874), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4529 ( .A1(n3851), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4530 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3556)
         );
  OAI21_X1 U4531 ( .B1(n3557), .B2(n3556), .A(n3623), .ZN(n3560) );
  NAND2_X1 U4532 ( .A1(n3921), .A2(EAX_REG_12__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4533 ( .A1(n5357), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3558)
         );
  NAND3_X1 U4534 ( .A1(n3560), .A2(n3559), .A3(n3558), .ZN(n3561) );
  AOI21_X1 U4535 ( .B1(n5291), .B2(n3920), .A(n3561), .ZN(n5249) );
  XNOR2_X1 U4536 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3562), .ZN(n6129)
         );
  INV_X1 U4537 ( .A(n6129), .ZN(n3577) );
  AOI22_X1 U4538 ( .A1(n3011), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4539 ( .A1(n3303), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4540 ( .A1(n3021), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4541 ( .A1(n3184), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4542 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3572)
         );
  AOI22_X1 U4543 ( .A1(n3022), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4544 ( .A1(n3179), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4545 ( .A1(n3017), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4546 ( .A1(n3333), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4547 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  OAI21_X1 U4548 ( .B1(n3572), .B2(n3571), .A(n3623), .ZN(n3575) );
  NAND2_X1 U4549 ( .A1(n3921), .A2(EAX_REG_11__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4550 ( .A1(n5357), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3573)
         );
  NAND3_X1 U4551 ( .A1(n3575), .A2(n3574), .A3(n3573), .ZN(n3576) );
  AOI21_X1 U4552 ( .B1(n3577), .B2(n3920), .A(n3576), .ZN(n5240) );
  NOR2_X1 U4553 ( .A1(n5249), .A2(n5240), .ZN(n3578) );
  AND2_X1 U4554 ( .A1(n5063), .A2(n3578), .ZN(n3579) );
  INV_X1 U4555 ( .A(n3587), .ZN(n3584) );
  NAND2_X1 U4556 ( .A1(n3921), .A2(EAX_REG_13__SCAN_IN), .ZN(n3583) );
  OAI21_X1 U4557 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3581), .A(n3626), 
        .ZN(n5975) );
  AOI22_X1 U4558 ( .A1(n3920), .A2(n5975), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4559 ( .A1(n3583), .A2(n3582), .ZN(n3585) );
  INV_X1 U4560 ( .A(n3585), .ZN(n3586) );
  NAND2_X1 U4561 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  AOI22_X1 U4562 ( .A1(n3019), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4563 ( .A1(n3021), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4564 ( .A1(n3194), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4565 ( .A1(n3184), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4566 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3598)
         );
  AOI22_X1 U4567 ( .A1(n3018), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4568 ( .A1(n3332), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4569 ( .A1(n3017), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4570 ( .A1(n3333), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3593) );
  NAND4_X1 U4571 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3597)
         );
  OR2_X1 U4572 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  AND2_X1 U4573 ( .A1(n3623), .A2(n3599), .ZN(n5275) );
  AOI22_X1 U4574 ( .A1(n3177), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4575 ( .A1(n3303), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4576 ( .A1(n3022), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4577 ( .A1(n3184), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3601) );
  NAND4_X1 U4578 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3610)
         );
  AOI22_X1 U4579 ( .A1(n3874), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4580 ( .A1(n3020), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4581 ( .A1(n3021), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4582 ( .A1(n3017), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3605) );
  NAND4_X1 U4583 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3609)
         );
  NOR2_X1 U4584 ( .A1(n3610), .A2(n3609), .ZN(n3613) );
  XNOR2_X1 U4585 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3626), .ZN(n5964)
         );
  INV_X1 U4586 ( .A(n5964), .ZN(n5347) );
  AOI22_X1 U4587 ( .A1(n5357), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3920), 
        .B2(n5347), .ZN(n3612) );
  NAND2_X1 U4588 ( .A1(n3921), .A2(EAX_REG_14__SCAN_IN), .ZN(n3611) );
  OAI211_X1 U4589 ( .C1(n3614), .C2(n3613), .A(n3612), .B(n3611), .ZN(n5282)
         );
  AOI22_X1 U4590 ( .A1(n3019), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4591 ( .A1(n3018), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4592 ( .A1(n3011), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4593 ( .A1(n3333), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4594 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3625)
         );
  AOI22_X1 U4595 ( .A1(n3021), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4596 ( .A1(n3022), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4597 ( .A1(n3184), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4598 ( .A1(n3017), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4599 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3624)
         );
  OAI21_X1 U4600 ( .B1(n3625), .B2(n3624), .A(n3623), .ZN(n3630) );
  NAND2_X1 U4601 ( .A1(n3921), .A2(EAX_REG_15__SCAN_IN), .ZN(n3629) );
  INV_X1 U4602 ( .A(n3633), .ZN(n3627) );
  XNOR2_X1 U4603 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3627), .ZN(n5638)
         );
  AOI22_X1 U4604 ( .A1(n3920), .A2(n5638), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3628) );
  XOR2_X1 U4605 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3649), .Z(n5955) );
  INV_X1 U4606 ( .A(n5955), .ZN(n5628) );
  NAND2_X1 U4607 ( .A1(n4609), .A2(n3004), .ZN(n3634) );
  AOI22_X1 U4608 ( .A1(n3011), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4609 ( .A1(n3021), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4610 ( .A1(n3018), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4611 ( .A1(n3017), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3636) );
  NAND4_X1 U4612 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3645)
         );
  AOI22_X1 U4613 ( .A1(n3022), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4614 ( .A1(n3020), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4615 ( .A1(n3184), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4616 ( .A1(n3411), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3640) );
  NAND4_X1 U4617 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3644)
         );
  NOR2_X1 U4618 ( .A1(n3645), .A2(n3644), .ZN(n3647) );
  AOI22_X1 U4619 ( .A1(n3921), .A2(EAX_REG_16__SCAN_IN), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3646) );
  OAI21_X1 U4620 ( .B1(n3924), .B2(n3647), .A(n3646), .ZN(n3648) );
  AOI21_X1 U4621 ( .B1(n5628), .B2(n3920), .A(n3648), .ZN(n5506) );
  NAND2_X1 U4622 ( .A1(n3649), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3666)
         );
  XNOR2_X1 U4623 ( .A(n3666), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5618)
         );
  AOI22_X1 U4624 ( .A1(n3179), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4625 ( .A1(n3022), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4626 ( .A1(n3177), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4627 ( .A1(n3017), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3650) );
  NAND4_X1 U4628 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3659)
         );
  AOI22_X1 U4629 ( .A1(n3303), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4630 ( .A1(n3874), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4631 ( .A1(n3184), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4632 ( .A1(n3021), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3654) );
  NAND4_X1 U4633 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n3658)
         );
  OR2_X1 U4634 ( .A1(n3659), .A2(n3658), .ZN(n3663) );
  INV_X1 U4635 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3661) );
  OAI21_X1 U4636 ( .B1(n5923), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6503), 
        .ZN(n3660) );
  OAI21_X1 U4637 ( .B1(n3682), .B2(n3661), .A(n3660), .ZN(n3662) );
  AOI21_X1 U4638 ( .B1(n3898), .B2(n3663), .A(n3662), .ZN(n3664) );
  AOI21_X1 U4639 ( .B1(n5618), .B2(n3920), .A(n3664), .ZN(n5312) );
  OR2_X1 U4640 ( .A1(n3667), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3668)
         );
  NAND2_X1 U4641 ( .A1(n3668), .A2(n3715), .ZN(n5948) );
  AOI22_X1 U4642 ( .A1(n3179), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4643 ( .A1(n3017), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4644 ( .A1(n3021), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4645 ( .A1(n3411), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4646 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3678)
         );
  AOI22_X1 U4647 ( .A1(n3011), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4648 ( .A1(n3184), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4649 ( .A1(n3018), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4650 ( .A1(n3851), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4651 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3677)
         );
  NOR2_X1 U4652 ( .A1(n3678), .A2(n3677), .ZN(n3679) );
  NOR2_X1 U4653 ( .A1(n3924), .A2(n3679), .ZN(n3684) );
  INV_X1 U4654 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3681) );
  NAND2_X1 U4655 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3680)
         );
  OAI211_X1 U4656 ( .C1(n3682), .C2(n3681), .A(n3044), .B(n3680), .ZN(n3683)
         );
  OAI22_X1 U4657 ( .A1(n5948), .A2(n3044), .B1(n3684), .B2(n3683), .ZN(n5502)
         );
  AOI22_X1 U4658 ( .A1(n3019), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3011), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4659 ( .A1(n3184), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4660 ( .A1(n3303), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4661 ( .A1(n3194), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4662 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3694)
         );
  AOI22_X1 U4663 ( .A1(n3021), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4664 ( .A1(n3017), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4665 ( .A1(n3332), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4666 ( .A1(n3875), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4667 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3693)
         );
  NOR2_X1 U4668 ( .A1(n3694), .A2(n3693), .ZN(n3698) );
  NAND2_X1 U4669 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3695)
         );
  NAND2_X1 U4670 ( .A1(n3044), .A2(n3695), .ZN(n3696) );
  AOI21_X1 U4671 ( .B1(n3921), .B2(EAX_REG_19__SCAN_IN), .A(n3696), .ZN(n3697)
         );
  OAI21_X1 U4672 ( .B1(n3924), .B2(n3698), .A(n3697), .ZN(n3700) );
  XNOR2_X1 U4673 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3715), .ZN(n5832)
         );
  NAND2_X1 U4674 ( .A1(n3920), .A2(n5832), .ZN(n3699) );
  NAND2_X1 U4675 ( .A1(n3700), .A2(n3699), .ZN(n5490) );
  AOI22_X1 U4676 ( .A1(n3177), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4677 ( .A1(n3411), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4678 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3194), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4679 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3017), .B1(n3875), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4680 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3710)
         );
  AOI22_X1 U4681 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3333), .B1(n3874), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4682 ( .A1(n3020), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4683 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3021), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4684 ( .A1(n3184), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4685 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  NOR2_X1 U4686 ( .A1(n3710), .A2(n3709), .ZN(n3714) );
  NAND2_X1 U4687 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3711)
         );
  NAND2_X1 U4688 ( .A1(n3044), .A2(n3711), .ZN(n3712) );
  AOI21_X1 U4689 ( .B1(n3921), .B2(EAX_REG_20__SCAN_IN), .A(n3712), .ZN(n3713)
         );
  OAI21_X1 U4690 ( .B1(n3924), .B2(n3714), .A(n3713), .ZN(n3719) );
  OAI21_X1 U4691 ( .B1(n3717), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3749), 
        .ZN(n5823) );
  OR2_X1 U4692 ( .A1(n5823), .A2(n3044), .ZN(n3718) );
  AOI22_X1 U4693 ( .A1(n3019), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4694 ( .A1(n3194), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4695 ( .A1(n3177), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4696 ( .A1(n3017), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3720) );
  NAND4_X1 U4697 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3729)
         );
  AOI22_X1 U4698 ( .A1(n3303), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4699 ( .A1(n3874), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4700 ( .A1(n3184), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4701 ( .A1(n3021), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3724) );
  NAND4_X1 U4702 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3728)
         );
  NOR2_X1 U4703 ( .A1(n3729), .A2(n3728), .ZN(n3732) );
  AOI21_X1 U4704 ( .B1(n5590), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3730) );
  AOI21_X1 U4705 ( .B1(n3921), .B2(EAX_REG_21__SCAN_IN), .A(n3730), .ZN(n3731)
         );
  OAI21_X1 U4706 ( .B1(n3924), .B2(n3732), .A(n3731), .ZN(n3734) );
  XNOR2_X1 U4707 ( .A(n3749), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5817)
         );
  NAND2_X1 U4708 ( .A1(n5817), .A2(n3920), .ZN(n3733) );
  NAND2_X1 U4709 ( .A1(n5478), .A2(n5591), .ZN(n5472) );
  AOI22_X1 U4710 ( .A1(n3332), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4711 ( .A1(n3411), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4712 ( .A1(n3021), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4713 ( .A1(n3011), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3735) );
  NAND4_X1 U4714 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3744)
         );
  AOI22_X1 U4715 ( .A1(n3019), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4716 ( .A1(n3874), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4717 ( .A1(n3017), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4718 ( .A1(n3150), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3739) );
  NAND4_X1 U4719 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3743)
         );
  NOR2_X1 U4720 ( .A1(n3744), .A2(n3743), .ZN(n3748) );
  NAND2_X1 U4721 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3745)
         );
  NAND2_X1 U4722 ( .A1(n3044), .A2(n3745), .ZN(n3746) );
  AOI21_X1 U4723 ( .B1(n3921), .B2(EAX_REG_22__SCAN_IN), .A(n3746), .ZN(n3747)
         );
  OAI21_X1 U4724 ( .B1(n3924), .B2(n3748), .A(n3747), .ZN(n3753) );
  OR2_X1 U4725 ( .A1(n3750), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3751)
         );
  AND2_X1 U4726 ( .A1(n3796), .A2(n3751), .ZN(n5810) );
  NAND2_X1 U4727 ( .A1(n5810), .A2(n3920), .ZN(n3752) );
  NAND2_X1 U4728 ( .A1(n3753), .A2(n3752), .ZN(n5474) );
  AOI22_X1 U4729 ( .A1(n3011), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4730 ( .A1(n3017), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4731 ( .A1(n3303), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4732 ( .A1(n3184), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3755) );
  NAND4_X1 U4733 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3764)
         );
  AOI22_X1 U4734 ( .A1(n3021), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4735 ( .A1(n3019), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4736 ( .A1(n3150), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4737 ( .A1(n3851), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4738 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3763)
         );
  NOR2_X1 U4739 ( .A1(n3764), .A2(n3763), .ZN(n3783) );
  AOI22_X1 U4740 ( .A1(n3021), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4741 ( .A1(n3179), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4742 ( .A1(n3332), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4743 ( .A1(n3184), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4744 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3774)
         );
  AOI22_X1 U4745 ( .A1(n3017), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4746 ( .A1(n3411), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4747 ( .A1(n3022), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4748 ( .A1(n3333), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4749 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  NOR2_X1 U4750 ( .A1(n3774), .A2(n3773), .ZN(n3784) );
  XOR2_X1 U4751 ( .A(n3783), .B(n3784), .Z(n3775) );
  NAND2_X1 U4752 ( .A1(n3775), .A2(n3898), .ZN(n3779) );
  NAND2_X1 U4753 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3776)
         );
  NAND2_X1 U4754 ( .A1(n3044), .A2(n3776), .ZN(n3777) );
  AOI21_X1 U4755 ( .B1(n3921), .B2(EAX_REG_23__SCAN_IN), .A(n3777), .ZN(n3778)
         );
  NAND2_X1 U4756 ( .A1(n3779), .A2(n3778), .ZN(n3781) );
  XNOR2_X1 U4757 ( .A(n3796), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5798)
         );
  NAND2_X1 U4758 ( .A1(n5798), .A2(n3920), .ZN(n3780) );
  NAND2_X1 U4759 ( .A1(n3781), .A2(n3780), .ZN(n5467) );
  NOR2_X1 U4760 ( .A1(n3784), .A2(n3783), .ZN(n3815) );
  AOI22_X1 U4761 ( .A1(n3019), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4762 ( .A1(n3022), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4763 ( .A1(n3011), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4764 ( .A1(n3017), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4765 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4766 ( .A1(n3303), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4767 ( .A1(n3874), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4768 ( .A1(n3184), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4769 ( .A1(n3021), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4770 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  OR2_X1 U4771 ( .A1(n3794), .A2(n3793), .ZN(n3814) );
  INV_X1 U4772 ( .A(n3814), .ZN(n3795) );
  XNOR2_X1 U4773 ( .A(n3815), .B(n3795), .ZN(n3803) );
  NAND2_X1 U4774 ( .A1(n3921), .A2(EAX_REG_24__SCAN_IN), .ZN(n3800) );
  AND2_X1 U4775 ( .A1(n3797), .A2(n4342), .ZN(n3798) );
  OR2_X1 U4776 ( .A1(n3798), .A2(n3838), .ZN(n5566) );
  NAND2_X1 U4777 ( .A1(n5566), .A2(n3920), .ZN(n3799) );
  OAI211_X1 U4778 ( .C1(n4342), .C2(n3801), .A(n3800), .B(n3799), .ZN(n3802)
         );
  AOI21_X1 U4779 ( .B1(n3803), .B2(n3898), .A(n3802), .ZN(n4362) );
  AOI22_X1 U4780 ( .A1(n3019), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4781 ( .A1(n3194), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4782 ( .A1(n3177), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4783 ( .A1(n3017), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4784 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4785 ( .A1(n3303), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4786 ( .A1(n3874), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4787 ( .A1(n3184), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4788 ( .A1(n3021), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4789 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  NOR2_X1 U4790 ( .A1(n3813), .A2(n3812), .ZN(n3823) );
  NAND2_X1 U4791 ( .A1(n3815), .A2(n3814), .ZN(n3822) );
  XOR2_X1 U4792 ( .A(n3823), .B(n3822), .Z(n3816) );
  NAND2_X1 U4793 ( .A1(n3816), .A2(n3898), .ZN(n3821) );
  NAND2_X1 U4794 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3817)
         );
  NAND2_X1 U4795 ( .A1(n3044), .A2(n3817), .ZN(n3818) );
  AOI21_X1 U4796 ( .B1(n3385), .B2(EAX_REG_25__SCAN_IN), .A(n3818), .ZN(n3820)
         );
  INV_X1 U4797 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5555) );
  XNOR2_X1 U4798 ( .A(n3838), .B(n5555), .ZN(n5789) );
  AND2_X1 U4799 ( .A1(n5789), .A2(n3920), .ZN(n3819) );
  AOI21_X1 U4800 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n5457) );
  NOR2_X1 U4801 ( .A1(n3823), .A2(n3822), .ZN(n3846) );
  AOI22_X1 U4802 ( .A1(n3179), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4803 ( .A1(n3022), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4804 ( .A1(n3011), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4805 ( .A1(n3017), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4806 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3833)
         );
  AOI22_X1 U4807 ( .A1(n3303), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4808 ( .A1(n3874), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4809 ( .A1(n3184), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4810 ( .A1(n3021), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4811 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3832)
         );
  OR2_X1 U4812 ( .A1(n3833), .A2(n3832), .ZN(n3845) );
  INV_X1 U4813 ( .A(n3845), .ZN(n3834) );
  XNOR2_X1 U4814 ( .A(n3846), .B(n3834), .ZN(n3835) );
  NAND2_X1 U4815 ( .A1(n3835), .A2(n3898), .ZN(n3844) );
  NAND2_X1 U4816 ( .A1(n6503), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3836)
         );
  NAND2_X1 U4817 ( .A1(n3044), .A2(n3836), .ZN(n3837) );
  AOI21_X1 U4818 ( .B1(n3921), .B2(EAX_REG_26__SCAN_IN), .A(n3837), .ZN(n3843)
         );
  INV_X1 U4819 ( .A(n3839), .ZN(n3840) );
  INV_X1 U4820 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U4821 ( .A1(n3840), .A2(n5551), .ZN(n3841) );
  NAND2_X1 U4822 ( .A1(n3863), .A2(n3841), .ZN(n5787) );
  NOR2_X1 U4823 ( .A1(n5787), .A2(n3044), .ZN(n3842) );
  AOI21_X1 U4824 ( .B1(n3844), .B2(n3843), .A(n3842), .ZN(n5449) );
  NAND2_X1 U4825 ( .A1(n3846), .A2(n3845), .ZN(n3867) );
  AOI22_X1 U4826 ( .A1(n3177), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4827 ( .A1(n3021), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4828 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3333), .B1(n3874), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4829 ( .A1(n3017), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4830 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3858)
         );
  AOI22_X1 U4831 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3303), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4832 ( .A1(n3194), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4833 ( .A1(n3020), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4834 ( .A1(n3852), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4835 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  NOR2_X1 U4836 ( .A1(n3858), .A2(n3857), .ZN(n3868) );
  XOR2_X1 U4837 ( .A(n3867), .B(n3868), .Z(n3859) );
  NAND2_X1 U4838 ( .A1(n3859), .A2(n3898), .ZN(n3862) );
  INV_X1 U4839 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5543) );
  NOR2_X1 U4840 ( .A1(n5543), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3860) );
  AOI211_X1 U4841 ( .C1(n3921), .C2(EAX_REG_27__SCAN_IN), .A(n3920), .B(n3860), 
        .ZN(n3861) );
  XNOR2_X1 U4842 ( .A(n3863), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5547)
         );
  INV_X1 U4843 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4844 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  NAND2_X1 U4845 ( .A1(n3901), .A2(n3866), .ZN(n5536) );
  NOR2_X1 U4846 ( .A1(n3868), .A2(n3867), .ZN(n3887) );
  AOI22_X1 U4847 ( .A1(n3019), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4848 ( .A1(n3022), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4849 ( .A1(n3011), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4850 ( .A1(n3017), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4851 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3881)
         );
  AOI22_X1 U4852 ( .A1(n3303), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4853 ( .A1(n3874), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4854 ( .A1(n3184), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4855 ( .A1(n3021), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4856 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3880)
         );
  OR2_X1 U4857 ( .A1(n3881), .A2(n3880), .ZN(n3886) );
  XNOR2_X1 U4858 ( .A(n3887), .B(n3886), .ZN(n3884) );
  AOI21_X1 U4859 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6503), .A(n3920), 
        .ZN(n3883) );
  NAND2_X1 U4860 ( .A1(n3921), .A2(EAX_REG_28__SCAN_IN), .ZN(n3882) );
  OAI211_X1 U4861 ( .C1(n3884), .C2(n3924), .A(n3883), .B(n3882), .ZN(n3885)
         );
  OAI21_X1 U4862 ( .B1(n3044), .B2(n5536), .A(n3885), .ZN(n5423) );
  NAND2_X1 U4863 ( .A1(n3887), .A2(n3886), .ZN(n3916) );
  AOI22_X1 U4864 ( .A1(n3411), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4865 ( .A1(n3021), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4866 ( .A1(n3184), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4867 ( .A1(n3909), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4868 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3897)
         );
  AOI22_X1 U4869 ( .A1(n3019), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4870 ( .A1(n3194), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4871 ( .A1(n3017), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4872 ( .A1(n3333), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4873 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  NOR2_X1 U4874 ( .A1(n3897), .A2(n3896), .ZN(n3917) );
  XOR2_X1 U4875 ( .A(n3916), .B(n3917), .Z(n3899) );
  NAND2_X1 U4876 ( .A1(n3899), .A2(n3898), .ZN(n3903) );
  INV_X1 U4877 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4302) );
  NOR2_X1 U4878 ( .A1(n4302), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3900) );
  AOI211_X1 U4879 ( .C1(n3385), .C2(EAX_REG_29__SCAN_IN), .A(n3920), .B(n3900), 
        .ZN(n3902) );
  XOR2_X1 U4880 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n3904), .Z(n5404) );
  XOR2_X1 U4881 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4354), .Z(n5412) );
  AOI22_X1 U4882 ( .A1(n3019), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3011), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4883 ( .A1(n3303), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4884 ( .A1(n3851), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4885 ( .A1(n3333), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4886 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3915)
         );
  AOI22_X1 U4887 ( .A1(n3017), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4888 ( .A1(n3021), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3874), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4889 ( .A1(n3332), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4890 ( .A1(n3150), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3006), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4891 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  NOR2_X1 U4892 ( .A1(n3915), .A2(n3914), .ZN(n3919) );
  NOR2_X1 U4893 ( .A1(n3917), .A2(n3916), .ZN(n3918) );
  XOR2_X1 U4894 ( .A(n3919), .B(n3918), .Z(n3925) );
  AOI21_X1 U4895 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6503), .A(n3920), 
        .ZN(n3923) );
  NAND2_X1 U4896 ( .A1(n3921), .A2(EAX_REG_30__SCAN_IN), .ZN(n3922) );
  OAI211_X1 U4897 ( .C1(n3925), .C2(n3924), .A(n3923), .B(n3922), .ZN(n3926)
         );
  OAI21_X1 U4898 ( .B1(n3044), .B2(n5412), .A(n3926), .ZN(n5356) );
  INV_X1 U4899 ( .A(n5353), .ZN(n5421) );
  NAND2_X1 U4900 ( .A1(n6455), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3947) );
  INV_X1 U4901 ( .A(n3947), .ZN(n3928) );
  XNOR2_X1 U4902 ( .A(n4529), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3948)
         );
  NAND2_X1 U4903 ( .A1(n3928), .A2(n3948), .ZN(n3930) );
  NAND2_X1 U4904 ( .A1(n6461), .A2(n4529), .ZN(n3929) );
  NAND2_X1 U4905 ( .A1(n3930), .A2(n3929), .ZN(n3964) );
  XNOR2_X1 U4906 ( .A(n3110), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3963)
         );
  INV_X1 U4907 ( .A(n3963), .ZN(n3931) );
  NAND2_X1 U4908 ( .A1(n3964), .A2(n3931), .ZN(n3933) );
  NAND2_X1 U4909 ( .A1(n6466), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U4910 ( .A1(n3933), .A2(n3932), .ZN(n3936) );
  XNOR2_X1 U4911 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4912 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3976), .ZN(n3934) );
  NOR2_X1 U4913 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3934), .ZN(n3940)
         );
  NOR2_X1 U4914 ( .A1(n3936), .A2(n3935), .ZN(n3937) );
  OR2_X1 U4915 ( .A1(n3938), .A2(n3937), .ZN(n3939) );
  NAND2_X1 U4916 ( .A1(n4246), .A2(n4609), .ZN(n3941) );
  NAND2_X1 U4917 ( .A1(n3270), .A2(n4609), .ZN(n4253) );
  NAND2_X1 U4918 ( .A1(n5375), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3943) );
  AND2_X1 U4919 ( .A1(n3947), .A2(n3943), .ZN(n3949) );
  NAND2_X1 U4920 ( .A1(n4253), .A2(n3949), .ZN(n3944) );
  NAND2_X1 U4921 ( .A1(n3944), .A2(n4339), .ZN(n3946) );
  AOI22_X1 U4922 ( .A1(n3962), .A2(n3946), .B1(n3945), .B2(n3956), .ZN(n3953)
         );
  AOI21_X1 U4923 ( .B1(n3980), .B2(n3275), .A(n3235), .ZN(n3954) );
  XNOR2_X1 U4924 ( .A(n3948), .B(n3947), .ZN(n3989) );
  NAND2_X1 U4925 ( .A1(n3989), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3955) );
  NAND2_X1 U4926 ( .A1(n3954), .A2(n3955), .ZN(n3952) );
  INV_X1 U4927 ( .A(n3949), .ZN(n3950) );
  NAND2_X1 U4928 ( .A1(n3956), .A2(n3950), .ZN(n3951) );
  NAND3_X1 U4929 ( .A1(n3953), .A2(n3952), .A3(n3951), .ZN(n3961) );
  INV_X1 U4930 ( .A(n3954), .ZN(n3959) );
  INV_X1 U4931 ( .A(n3955), .ZN(n3958) );
  INV_X1 U4932 ( .A(n3989), .ZN(n3957) );
  AOI22_X1 U4933 ( .A1(n3959), .A2(n3958), .B1(n3957), .B2(n3977), .ZN(n3960)
         );
  NAND2_X1 U4934 ( .A1(n3961), .A2(n3960), .ZN(n3966) );
  XNOR2_X1 U4935 ( .A(n3964), .B(n3963), .ZN(n3988) );
  OAI211_X1 U4936 ( .C1(n3966), .C2(n3967), .A(n3988), .B(n3980), .ZN(n3970)
         );
  NOR2_X1 U4937 ( .A1(n3965), .A2(n3988), .ZN(n3968) );
  OAI21_X1 U4938 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n3969) );
  NAND2_X1 U4939 ( .A1(n3970), .A2(n3969), .ZN(n3971) );
  OAI21_X1 U4940 ( .B1(n3972), .B2(n3987), .A(n3971), .ZN(n3975) );
  AOI22_X1 U4941 ( .A1(n3973), .A2(n3977), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6504), .ZN(n3974) );
  NAND2_X1 U4942 ( .A1(n3975), .A2(n3974), .ZN(n3979) );
  OAI222_X1 U4943 ( .A1(n5913), .A2(n3976), .B1(n5913), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3976), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U4944 ( .A1(n3986), .A2(n3977), .ZN(n3978) );
  NAND2_X1 U4945 ( .A1(n3986), .A2(n3980), .ZN(n3981) );
  AND2_X1 U4946 ( .A1(n4016), .A2(n4240), .ZN(n3984) );
  NAND2_X1 U4947 ( .A1(n6480), .A2(n6473), .ZN(n3994) );
  INV_X1 U4948 ( .A(n3986), .ZN(n3991) );
  NAND3_X1 U4949 ( .A1(n3989), .A2(n3988), .A3(n3987), .ZN(n3990) );
  NAND2_X1 U4950 ( .A1(n3991), .A2(n3990), .ZN(n5916) );
  NOR2_X1 U4951 ( .A1(READY_N), .A2(n5916), .ZN(n4236) );
  INV_X1 U4952 ( .A(n4236), .ZN(n3992) );
  NAND2_X1 U4953 ( .A1(n3994), .A2(n3993), .ZN(n4396) );
  NOR2_X1 U4954 ( .A1(n3015), .A2(n3004), .ZN(n4018) );
  NAND2_X1 U4955 ( .A1(n4018), .A2(n4621), .ZN(n3996) );
  NOR2_X1 U4956 ( .A1(n3995), .A2(n3996), .ZN(n3998) );
  NAND2_X1 U4957 ( .A1(n3275), .A2(n6708), .ZN(n4000) );
  NAND2_X1 U4958 ( .A1(n2999), .A2(n3015), .ZN(n4002) );
  AND2_X1 U4959 ( .A1(n5512), .A2(n3253), .ZN(n6070) );
  AOI22_X1 U4960 ( .A1(n6070), .A2(DATAI_30_), .B1(n6073), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4005) );
  NOR2_X1 U4961 ( .A1(n5513), .A2(n4609), .ZN(n4003) );
  NAND2_X1 U4962 ( .A1(n6074), .A2(DATAI_14_), .ZN(n4004) );
  OAI21_X1 U4963 ( .B1(n5421), .B2(n5848), .A(n3108), .ZN(U2861) );
  INV_X1 U4964 ( .A(n3239), .ZN(n4007) );
  NAND2_X1 U4965 ( .A1(n4007), .A2(n2986), .ZN(n4008) );
  INV_X1 U4966 ( .A(n4009), .ZN(n4010) );
  NAND2_X1 U4967 ( .A1(n4009), .A2(n3275), .ZN(n4024) );
  AND2_X1 U4968 ( .A1(n4240), .A2(n3275), .ZN(n5104) );
  NAND2_X1 U4969 ( .A1(n5104), .A2(n4019), .ZN(n4012) );
  OAI21_X1 U4970 ( .B1(n4247), .B2(n4339), .A(n3249), .ZN(n4011) );
  NAND2_X1 U4971 ( .A1(n4012), .A2(n4011), .ZN(n4013) );
  AOI21_X1 U4972 ( .B1(n3983), .B2(n4446), .A(n4013), .ZN(n4014) );
  NOR2_X1 U4973 ( .A1(n4016), .A2(n4246), .ZN(n4234) );
  NAND2_X1 U4974 ( .A1(n4402), .A2(n4234), .ZN(n4418) );
  INV_X1 U4975 ( .A(n4017), .ZN(n4020) );
  NAND4_X1 U4976 ( .A1(n4020), .A2(n4019), .A3(n4102), .A4(n4018), .ZN(n4021)
         );
  NAND2_X1 U4977 ( .A1(n4395), .A2(n4021), .ZN(n4022) );
  INV_X1 U4978 ( .A(n4024), .ZN(n4045) );
  INV_X1 U4979 ( .A(n4118), .ZN(n4058) );
  INV_X1 U4980 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U4981 ( .A1(n4102), .A2(n4023), .ZN(n4025) );
  OAI211_X1 U4982 ( .C1(n4058), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4025), 
        .B(n5484), .ZN(n4026) );
  NAND2_X1 U4983 ( .A1(n4118), .A2(EBX_REG_0__SCAN_IN), .ZN(n4028) );
  INV_X1 U4984 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U4985 ( .A1(n5484), .A2(n5178), .ZN(n4027) );
  AND2_X1 U4986 ( .A1(n4028), .A2(n4027), .ZN(n4448) );
  INV_X1 U4987 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4988 ( .A1(n4110), .A2(n4032), .ZN(n4036) );
  NAND2_X1 U4989 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4031)
         );
  NAND2_X1 U4990 ( .A1(n4118), .A2(n4031), .ZN(n4034) );
  NAND2_X1 U4991 ( .A1(n4102), .A2(n4032), .ZN(n4033) );
  NAND2_X1 U4992 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  NAND2_X1 U4993 ( .A1(n4036), .A2(n4035), .ZN(n4518) );
  NAND2_X1 U4994 ( .A1(n4045), .A2(EBX_REG_3__SCAN_IN), .ZN(n4039) );
  INV_X1 U4995 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U4996 ( .A1(n4102), .A2(n4040), .ZN(n4041) );
  OAI211_X1 U4997 ( .C1(n4058), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4041), 
        .B(n5484), .ZN(n4042) );
  OAI21_X1 U4998 ( .B1(n4315), .B2(EBX_REG_4__SCAN_IN), .A(n4042), .ZN(n4574)
         );
  INV_X1 U4999 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4044) );
  INV_X1 U5000 ( .A(n4446), .ZN(n4125) );
  INV_X1 U5001 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6204) );
  AOI22_X1 U5002 ( .A1(n4125), .A2(n6204), .B1(n4116), .B2(n4044), .ZN(n4043)
         );
  OAI21_X1 U5003 ( .B1(n5484), .B2(n4044), .A(n4043), .ZN(n4728) );
  INV_X1 U5004 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6209) );
  AOI21_X1 U5005 ( .B1(n6209), .B2(n4118), .A(n4045), .ZN(n4046) );
  OAI21_X1 U5006 ( .B1(EBX_REG_6__SCAN_IN), .B2(n4496), .A(n4046), .ZN(n4047)
         );
  OAI21_X1 U5007 ( .B1(n4315), .B2(EBX_REG_6__SCAN_IN), .A(n4047), .ZN(n4840)
         );
  NAND2_X1 U5008 ( .A1(n4726), .A2(n4840), .ZN(n4836) );
  INV_X1 U5009 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4049) );
  INV_X1 U5010 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6182) );
  AOI22_X1 U5011 ( .A1(n4125), .A2(n6182), .B1(n4116), .B2(n4049), .ZN(n4048)
         );
  OAI21_X1 U5012 ( .B1(n5484), .B2(n4049), .A(n4048), .ZN(n4837) );
  INV_X1 U5013 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4050) );
  NAND2_X1 U5014 ( .A1(n4110), .A2(n4050), .ZN(n4054) );
  INV_X1 U5015 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U5016 ( .A1(n4118), .A2(n6190), .ZN(n4052) );
  NAND2_X1 U5017 ( .A1(n4102), .A2(n4050), .ZN(n4051) );
  NAND3_X1 U5018 ( .A1(n4052), .A2(n5484), .A3(n4051), .ZN(n4053) );
  NAND2_X1 U5019 ( .A1(n4054), .A2(n4053), .ZN(n4967) );
  INV_X1 U5020 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4056) );
  INV_X1 U5021 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5189) );
  AOI22_X1 U5022 ( .A1(n4125), .A2(n5189), .B1(n4116), .B2(n4056), .ZN(n4055)
         );
  OAI21_X1 U5023 ( .B1(n5484), .B2(n4056), .A(n4055), .ZN(n5060) );
  INV_X1 U5024 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U5025 ( .A1(n4102), .A2(n5077), .ZN(n4057) );
  OAI211_X1 U5026 ( .C1(n4058), .C2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4057), .B(n5484), .ZN(n4059) );
  OAI21_X1 U5027 ( .B1(n4315), .B2(EBX_REG_10__SCAN_IN), .A(n4059), .ZN(n5065)
         );
  INV_X1 U5028 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6164) );
  INV_X1 U5029 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U5030 ( .A1(n4102), .A2(n6065), .ZN(n4060) );
  OAI211_X1 U5031 ( .C1(n4045), .C2(n6164), .A(n4060), .B(n4118), .ZN(n4061)
         );
  OAI21_X1 U5032 ( .B1(n4109), .B2(EBX_REG_11__SCAN_IN), .A(n4061), .ZN(n5988)
         );
  INV_X1 U5033 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5034 ( .A1(n4110), .A2(n4062), .ZN(n4066) );
  INV_X1 U5035 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U5036 ( .A1(n4118), .A2(n5303), .ZN(n4064) );
  NAND2_X1 U5037 ( .A1(n4102), .A2(n4062), .ZN(n4063) );
  NAND3_X1 U5038 ( .A1(n4064), .A2(n5484), .A3(n4063), .ZN(n4065) );
  NAND2_X1 U5039 ( .A1(n4066), .A2(n4065), .ZN(n5251) );
  NAND2_X1 U5040 ( .A1(n5250), .A2(n5251), .ZN(n5252) );
  INV_X1 U5041 ( .A(EBX_REG_13__SCAN_IN), .ZN(n4068) );
  INV_X1 U5042 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5908) );
  AOI22_X1 U5043 ( .A1(n4125), .A2(n5908), .B1(n4116), .B2(n4068), .ZN(n4067)
         );
  OAI21_X1 U5044 ( .B1(n5484), .B2(n4068), .A(n4067), .ZN(n5278) );
  INV_X1 U5045 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U5046 ( .A1(n4110), .A2(n5286), .ZN(n4073) );
  NAND2_X1 U5047 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4069) );
  NAND2_X1 U5048 ( .A1(n4118), .A2(n4069), .ZN(n4071) );
  NAND2_X1 U5049 ( .A1(n4102), .A2(n5286), .ZN(n4070) );
  NAND2_X1 U5050 ( .A1(n4071), .A2(n4070), .ZN(n4072) );
  NAND2_X1 U5051 ( .A1(n4073), .A2(n4072), .ZN(n5284) );
  NAND2_X1 U5052 ( .A1(n4045), .A2(EBX_REG_15__SCAN_IN), .ZN(n4075) );
  OR2_X1 U5053 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4074)
         );
  OAI211_X1 U5054 ( .C1(n4109), .C2(EBX_REG_15__SCAN_IN), .A(n4075), .B(n4074), 
        .ZN(n5321) );
  INV_X1 U5055 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U5056 ( .A1(n4110), .A2(n5509), .ZN(n4079) );
  INV_X1 U5057 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U5058 ( .A1(n4118), .A2(n5758), .ZN(n4077) );
  NAND2_X1 U5059 ( .A1(n4102), .A2(n5509), .ZN(n4076) );
  NAND3_X1 U5060 ( .A1(n4077), .A2(n5484), .A3(n4076), .ZN(n4078) );
  NAND2_X1 U5061 ( .A1(n4079), .A2(n4078), .ZN(n5507) );
  NAND2_X1 U5062 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4080) );
  OAI211_X1 U5063 ( .C1(n4496), .C2(EBX_REG_17__SCAN_IN), .A(n4118), .B(n4080), 
        .ZN(n4081) );
  OAI21_X1 U5064 ( .B1(n4109), .B2(EBX_REG_17__SCAN_IN), .A(n4081), .ZN(n5314)
         );
  INV_X1 U5065 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4082) );
  NAND2_X1 U5066 ( .A1(n4110), .A2(n4082), .ZN(n4086) );
  INV_X1 U5067 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U5068 ( .A1(n4118), .A2(n5735), .ZN(n4084) );
  NAND2_X1 U5069 ( .A1(n4102), .A2(n4082), .ZN(n4083) );
  NAND3_X1 U5070 ( .A1(n4084), .A2(n5484), .A3(n4083), .ZN(n4085) );
  OR2_X1 U5071 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4088)
         );
  INV_X1 U5072 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U5073 ( .A1(n4102), .A2(n5505), .ZN(n4087) );
  OAI22_X1 U5074 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4496), .ZN(n5485) );
  AOI22_X1 U5075 ( .A1(n5482), .A2(n5485), .B1(n4045), .B2(EBX_REG_20__SCAN_IN), .ZN(n4090) );
  INV_X1 U5076 ( .A(n5482), .ZN(n4089) );
  NAND2_X1 U5077 ( .A1(n4089), .A2(n5484), .ZN(n5493) );
  NAND2_X1 U5078 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4092) );
  OAI211_X1 U5079 ( .C1(n4496), .C2(EBX_REG_21__SCAN_IN), .A(n4118), .B(n4092), 
        .ZN(n4093) );
  OAI21_X1 U5080 ( .B1(n4109), .B2(EBX_REG_21__SCAN_IN), .A(n4093), .ZN(n5711)
         );
  INV_X1 U5081 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U5082 ( .A1(n4110), .A2(n5813), .ZN(n4097) );
  NAND2_X1 U5083 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4094) );
  NAND2_X1 U5084 ( .A1(n4118), .A2(n4094), .ZN(n4095) );
  OAI21_X1 U5085 ( .B1(EBX_REG_22__SCAN_IN), .B2(n4496), .A(n4095), .ZN(n4096)
         );
  NAND2_X1 U5086 ( .A1(n4045), .A2(EBX_REG_23__SCAN_IN), .ZN(n4101) );
  OR2_X1 U5087 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4100)
         );
  INV_X1 U5088 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U5089 ( .A1(n4116), .A2(n4098), .ZN(n4099) );
  INV_X1 U5090 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5091 ( .A1(n4110), .A2(n4343), .ZN(n4106) );
  INV_X1 U5092 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U5093 ( .A1(n4118), .A2(n5685), .ZN(n4104) );
  NAND2_X1 U5094 ( .A1(n4102), .A2(n4343), .ZN(n4103) );
  NAND3_X1 U5095 ( .A1(n4104), .A2(n5484), .A3(n4103), .ZN(n4105) );
  AND2_X1 U5096 ( .A1(n4106), .A2(n4105), .ZN(n4364) );
  OR2_X1 U5097 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4108)
         );
  NAND2_X1 U5098 ( .A1(n4045), .A2(EBX_REG_25__SCAN_IN), .ZN(n4107) );
  OAI211_X1 U5099 ( .C1(n4109), .C2(EBX_REG_25__SCAN_IN), .A(n4108), .B(n4107), 
        .ZN(n5459) );
  INV_X1 U5100 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4111) );
  NAND2_X1 U5101 ( .A1(n4110), .A2(n4111), .ZN(n4115) );
  INV_X1 U5102 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U5103 ( .A1(n4118), .A2(n5531), .ZN(n4113) );
  NAND2_X1 U5104 ( .A1(n4102), .A2(n4111), .ZN(n4112) );
  NAND3_X1 U5105 ( .A1(n4113), .A2(n5484), .A3(n4112), .ZN(n4114) );
  INV_X1 U5106 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U5107 ( .A1(n4116), .A2(n5445), .ZN(n4120) );
  NAND2_X1 U5108 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4117) );
  OAI211_X1 U5109 ( .C1(n4496), .C2(EBX_REG_27__SCAN_IN), .A(n4118), .B(n4117), 
        .ZN(n4119) );
  NAND2_X1 U5110 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4121) );
  NAND2_X1 U5111 ( .A1(n4118), .A2(n4121), .ZN(n4122) );
  OAI21_X1 U5112 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4496), .A(n4122), .ZN(n4123)
         );
  OAI21_X1 U5113 ( .B1(n4315), .B2(EBX_REG_28__SCAN_IN), .A(n4123), .ZN(n5424)
         );
  NOR2_X1 U5114 ( .A1(n4496), .A2(EBX_REG_29__SCAN_IN), .ZN(n4124) );
  AOI21_X1 U5115 ( .B1(n4125), .B2(n5643), .A(n4124), .ZN(n5400) );
  INV_X1 U5116 ( .A(n4318), .ZN(n4128) );
  NAND2_X1 U5117 ( .A1(n4318), .A2(n5484), .ZN(n4320) );
  AND2_X1 U5118 ( .A1(n4496), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4126)
         );
  AOI21_X1 U5119 ( .B1(n4446), .B2(EBX_REG_30__SCAN_IN), .A(n4126), .ZN(n4319)
         );
  INV_X1 U5120 ( .A(n4319), .ZN(n4127) );
  OAI211_X1 U5121 ( .C1(n4128), .C2(n3065), .A(n4320), .B(n4127), .ZN(n4130)
         );
  OAI211_X1 U5122 ( .C1(n4316), .C2(n5484), .A(n4318), .B(n4319), .ZN(n4129)
         );
  NAND2_X1 U5123 ( .A1(n4130), .A2(n4129), .ZN(n5417) );
  INV_X1 U5124 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4131) );
  INV_X1 U5125 ( .A(n4190), .ZN(n4160) );
  NAND2_X1 U5126 ( .A1(n4137), .A2(n4145), .ZN(n4157) );
  XNOR2_X1 U5127 ( .A(n4157), .B(n4156), .ZN(n4134) );
  AND2_X1 U5128 ( .A1(n4240), .A2(n4009), .ZN(n4143) );
  AOI21_X1 U5129 ( .B1(n4134), .B2(n2986), .A(n4143), .ZN(n4135) );
  OR2_X1 U5130 ( .A1(n6154), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4155)
         );
  NAND2_X1 U5131 ( .A1(n6154), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4153)
         );
  INV_X1 U5132 ( .A(n4145), .ZN(n4138) );
  XNOR2_X1 U5133 ( .A(n4138), .B(n4137), .ZN(n4140) );
  NAND3_X1 U5134 ( .A1(n4391), .A2(n4609), .A3(n4009), .ZN(n4139) );
  AOI21_X1 U5135 ( .B1(n4140), .B2(n2986), .A(n4139), .ZN(n4141) );
  NAND2_X1 U5136 ( .A1(n4142), .A2(n4141), .ZN(n4498) );
  INV_X1 U5137 ( .A(n4143), .ZN(n4144) );
  OAI21_X1 U5138 ( .B1(n6605), .B2(n4145), .A(n4144), .ZN(n4146) );
  INV_X1 U5139 ( .A(n4146), .ZN(n4147) );
  NAND2_X1 U5140 ( .A1(n4381), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4148)
         );
  INV_X1 U5141 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5142 ( .A1(n4148), .A2(n4576), .ZN(n4150) );
  AND2_X1 U5143 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4149) );
  NAND2_X1 U5144 ( .A1(n4381), .A2(n4149), .ZN(n4151) );
  AND2_X1 U5145 ( .A1(n4150), .A2(n4151), .ZN(n4499) );
  INV_X1 U5146 ( .A(n4151), .ZN(n4152) );
  NAND2_X1 U5147 ( .A1(n4153), .A2(n6155), .ZN(n4154) );
  AND2_X2 U5148 ( .A1(n4155), .A2(n4154), .ZN(n6145) );
  NAND2_X1 U5149 ( .A1(n4157), .A2(n4156), .ZN(n4165) );
  XNOR2_X1 U5150 ( .A(n4165), .B(n4164), .ZN(n4158) );
  INV_X1 U5151 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U5152 ( .A(n4161), .B(n6230), .ZN(n6143) );
  NAND2_X1 U5153 ( .A1(n6145), .A2(n6143), .ZN(n6144) );
  NAND2_X1 U5154 ( .A1(n4161), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4162)
         );
  NAND2_X1 U5155 ( .A1(n6144), .A2(n4162), .ZN(n4569) );
  NAND2_X1 U5156 ( .A1(n4163), .A2(n4190), .ZN(n4168) );
  NAND2_X1 U5157 ( .A1(n4165), .A2(n4164), .ZN(n4174) );
  XNOR2_X1 U5158 ( .A(n4174), .B(n4172), .ZN(n4166) );
  NAND2_X1 U5159 ( .A1(n4166), .A2(n2986), .ZN(n4167) );
  NAND2_X1 U5160 ( .A1(n4168), .A2(n4167), .ZN(n4169) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4580) );
  XNOR2_X1 U5162 ( .A(n4169), .B(n4580), .ZN(n4572) );
  NAND2_X1 U5163 ( .A1(n4569), .A2(n4572), .ZN(n4570) );
  NAND2_X1 U5164 ( .A1(n4169), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4170)
         );
  NAND2_X1 U5165 ( .A1(n4171), .A2(n4190), .ZN(n4177) );
  INV_X1 U5166 ( .A(n4172), .ZN(n4173) );
  OR2_X1 U5167 ( .A1(n4174), .A2(n4173), .ZN(n4182) );
  XNOR2_X1 U5168 ( .A(n4182), .B(n4183), .ZN(n4175) );
  NAND2_X1 U5169 ( .A1(n4175), .A2(n2986), .ZN(n4176) );
  XNOR2_X1 U5170 ( .A(n4178), .B(n6204), .ZN(n4733) );
  NAND2_X1 U5171 ( .A1(n4730), .A2(n4733), .ZN(n4731) );
  NAND2_X1 U5172 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4179)
         );
  NAND2_X1 U5173 ( .A1(n4731), .A2(n4179), .ZN(n6135) );
  NAND3_X1 U5174 ( .A1(n4180), .A2(n4190), .A3(n4181), .ZN(n4187) );
  INV_X1 U5175 ( .A(n4182), .ZN(n4184) );
  NAND2_X1 U5176 ( .A1(n4184), .A2(n4183), .ZN(n4192) );
  XNOR2_X1 U5177 ( .A(n4192), .B(n4193), .ZN(n4185) );
  NAND2_X1 U5178 ( .A1(n4185), .A2(n2986), .ZN(n4186) );
  NAND2_X1 U5179 ( .A1(n4187), .A2(n4186), .ZN(n4188) );
  XNOR2_X1 U5180 ( .A(n4188), .B(n6209), .ZN(n6137) );
  NAND2_X1 U5181 ( .A1(n6135), .A2(n6137), .ZN(n6136) );
  NAND2_X1 U5182 ( .A1(n4188), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4189)
         );
  NAND2_X1 U5183 ( .A1(n4191), .A2(n4190), .ZN(n4197) );
  INV_X1 U5184 ( .A(n4192), .ZN(n4194) );
  NAND2_X1 U5185 ( .A1(n4194), .A2(n4193), .ZN(n4204) );
  XNOR2_X1 U5186 ( .A(n4204), .B(n4202), .ZN(n4195) );
  NAND2_X1 U5187 ( .A1(n4195), .A2(n2986), .ZN(n4196) );
  NAND2_X1 U5188 ( .A1(n4197), .A2(n4196), .ZN(n4198) );
  XNOR2_X1 U5189 ( .A(n4198), .B(n6182), .ZN(n4958) );
  NAND2_X1 U5190 ( .A1(n4955), .A2(n4958), .ZN(n4956) );
  NAND2_X1 U5191 ( .A1(n4198), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4199)
         );
  NAND2_X1 U5192 ( .A1(n4956), .A2(n4199), .ZN(n5048) );
  NAND2_X1 U5193 ( .A1(n4202), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4200) );
  NAND2_X1 U5194 ( .A1(n2986), .A2(n4202), .ZN(n4203) );
  OR2_X1 U5195 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  NAND2_X1 U5196 ( .A1(n2985), .A2(n4205), .ZN(n4206) );
  XNOR2_X1 U5197 ( .A(n4206), .B(n6190), .ZN(n5051) );
  NAND2_X1 U5198 ( .A1(n5048), .A2(n5051), .ZN(n5049) );
  NAND2_X1 U5199 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4207)
         );
  NAND2_X1 U5200 ( .A1(n2985), .A2(n5189), .ZN(n5179) );
  NAND2_X1 U5201 ( .A1(n5181), .A2(n5179), .ZN(n4208) );
  OR2_X1 U5202 ( .A1(n2985), .A2(n5189), .ZN(n5180) );
  INV_X1 U5203 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4209) );
  NAND2_X1 U5204 ( .A1(n2985), .A2(n4209), .ZN(n5266) );
  AND2_X1 U5205 ( .A1(n2985), .A2(n6164), .ZN(n4212) );
  OR2_X1 U5206 ( .A1(n2985), .A2(n4209), .ZN(n6126) );
  NOR2_X1 U5207 ( .A1(n2985), .A2(n5303), .ZN(n5288) );
  XNOR2_X1 U5208 ( .A(n2985), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5873)
         );
  NAND2_X1 U5209 ( .A1(n5872), .A2(n5873), .ZN(n4214) );
  NAND2_X1 U5210 ( .A1(n2985), .A2(n5908), .ZN(n4213) );
  INV_X1 U5211 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5343) );
  OR2_X1 U5212 ( .A1(n2985), .A2(n5343), .ZN(n4215) );
  INV_X1 U5213 ( .A(n5634), .ZN(n4217) );
  NOR2_X1 U5214 ( .A1(n2985), .A2(n5890), .ZN(n5633) );
  NAND2_X1 U5215 ( .A1(n2985), .A2(n5890), .ZN(n5631) );
  NAND2_X1 U5216 ( .A1(n2985), .A2(n5758), .ZN(n4218) );
  AND2_X1 U5217 ( .A1(n5631), .A2(n4218), .ZN(n4219) );
  NAND2_X1 U5218 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4278) );
  INV_X1 U5219 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5747) );
  INV_X1 U5220 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4220) );
  AND3_X1 U5221 ( .A1(n5747), .A2(n4220), .A3(n5758), .ZN(n4221) );
  INV_X1 U5222 ( .A(n2998), .ZN(n4226) );
  INV_X1 U5223 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5686) );
  INV_X1 U5224 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4223) );
  INV_X1 U5225 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5703) );
  NAND4_X1 U5226 ( .A1(n5685), .A2(n5686), .A3(n4223), .A4(n5703), .ZN(n4224)
         );
  INV_X1 U5227 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U5228 ( .A1(n5595), .A2(n5735), .ZN(n5729) );
  NOR2_X1 U5229 ( .A1(n4224), .A2(n5729), .ZN(n4225) );
  AND2_X1 U5230 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5727) );
  AND2_X1 U5231 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U5232 ( .A1(n5727), .A2(n4281), .ZN(n4270) );
  NAND2_X1 U5233 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4284) );
  OAI21_X1 U5234 ( .B1(n4270), .B2(n4284), .A(n2985), .ZN(n4227) );
  XNOR2_X1 U5235 ( .A(n2985), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5558)
         );
  INV_X1 U5236 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U5237 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U5238 ( .A1(n4312), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4232) );
  INV_X1 U5239 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5666) );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U5241 ( .A1(n5666), .A2(n4230), .ZN(n5653) );
  INV_X1 U5242 ( .A(n4234), .ZN(n4243) );
  INV_X1 U5243 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U5244 ( .A1(n3275), .A2(n6518), .ZN(n4237) );
  NAND3_X1 U5245 ( .A1(n4237), .A2(n4236), .A3(n3249), .ZN(n4242) );
  NAND2_X1 U5246 ( .A1(n4255), .A2(n4238), .ZN(n4241) );
  NAND2_X1 U5247 ( .A1(n4239), .A2(n4240), .ZN(n6475) );
  NAND2_X1 U5248 ( .A1(n4241), .A2(n6475), .ZN(n4393) );
  OAI211_X1 U5249 ( .C1(n6480), .C2(n4243), .A(n4242), .B(n4393), .ZN(n4244)
         );
  NAND2_X1 U5250 ( .A1(n4244), .A2(n6501), .ZN(n4252) );
  NAND2_X1 U5251 ( .A1(n4246), .A2(n6518), .ZN(n4335) );
  NAND3_X1 U5252 ( .A1(n4245), .A2(n4335), .A3(n6708), .ZN(n4248) );
  NAND3_X1 U5253 ( .A1(n4248), .A2(n4339), .A3(n4247), .ZN(n4249) );
  NAND2_X1 U5254 ( .A1(n4249), .A2(n4391), .ZN(n4250) );
  INV_X1 U5255 ( .A(n4253), .ZN(n4254) );
  INV_X1 U5256 ( .A(n6473), .ZN(n4417) );
  INV_X1 U5257 ( .A(n4256), .ZN(n4260) );
  INV_X1 U5258 ( .A(n4257), .ZN(n4258) );
  NAND2_X1 U5259 ( .A1(n4258), .A2(n3004), .ZN(n4259) );
  NAND4_X1 U5260 ( .A1(n4293), .A2(n4417), .A3(n4260), .A4(n4259), .ZN(n4261)
         );
  INV_X1 U5261 ( .A(n5417), .ZN(n4274) );
  NAND2_X1 U5262 ( .A1(n4245), .A2(n2986), .ZN(n4434) );
  OAI21_X1 U5263 ( .B1(n4257), .B2(n3004), .A(n4434), .ZN(n4262) );
  NAND2_X1 U5264 ( .A1(n6221), .A2(REIP_REG_30__SCAN_IN), .ZN(n5351) );
  INV_X1 U5265 ( .A(n5351), .ZN(n4273) );
  OAI211_X1 U5266 ( .C1(n3281), .C2(n4339), .A(n4402), .B(n4531), .ZN(n4263)
         );
  NAND2_X1 U5267 ( .A1(n4275), .A2(n4263), .ZN(n5892) );
  NAND2_X1 U5268 ( .A1(n4275), .A2(n4527), .ZN(n5302) );
  AND2_X1 U5269 ( .A1(n5302), .A2(n5369), .ZN(n4500) );
  NAND4_X1 U5270 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U5271 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4265) );
  NOR2_X1 U5272 ( .A1(n6212), .A2(n4265), .ZN(n5183) );
  NAND2_X1 U5273 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U5274 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6175) );
  NOR2_X1 U5275 ( .A1(n5188), .A2(n6175), .ZN(n5296) );
  NAND2_X1 U5276 ( .A1(n5183), .A2(n5296), .ZN(n5301) );
  NAND3_X1 U5277 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5902) );
  NOR2_X1 U5278 ( .A1(n5343), .A2(n5902), .ZN(n5757) );
  NAND3_X1 U5279 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5757), .ZN(n4266) );
  NOR2_X1 U5280 ( .A1(n5301), .A2(n4266), .ZN(n4277) );
  INV_X1 U5281 ( .A(n4277), .ZN(n4264) );
  INV_X1 U5282 ( .A(n4418), .ZN(n6479) );
  INV_X1 U5283 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U5284 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U5285 ( .A1(n6243), .A2(n6234), .ZN(n6233) );
  NAND3_X1 U5286 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6233), .ZN(n6210) );
  NOR2_X1 U5287 ( .A1(n4265), .A2(n6210), .ZN(n5187) );
  NAND2_X1 U5288 ( .A1(n5296), .A2(n5187), .ZN(n5299) );
  NOR2_X1 U5289 ( .A1(n4266), .A2(n5299), .ZN(n5721) );
  INV_X1 U5290 ( .A(n5721), .ZN(n4267) );
  OR2_X1 U5291 ( .A1(n6211), .A2(n4267), .ZN(n4268) );
  INV_X1 U5292 ( .A(n4270), .ZN(n5571) );
  NAND2_X1 U5293 ( .A1(n5736), .A2(n5571), .ZN(n5697) );
  NOR2_X1 U5294 ( .A1(n5697), .A2(n4284), .ZN(n5680) );
  NAND2_X1 U5295 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5671) );
  INV_X1 U5296 ( .A(n5671), .ZN(n4271) );
  NAND2_X1 U5297 ( .A1(n5680), .A2(n4271), .ZN(n5651) );
  NOR4_X1 U5298 ( .A1(n5651), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5652), 
        .A4(n5643), .ZN(n4272) );
  AOI211_X1 U5299 ( .C1(n4274), .C2(n6238), .A(n4273), .B(n4272), .ZN(n4289)
         );
  INV_X1 U5300 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5369) );
  INV_X1 U5301 ( .A(n5892), .ZN(n4276) );
  NOR2_X1 U5302 ( .A1(n4275), .A2(n6221), .ZN(n4503) );
  AOI21_X1 U5303 ( .B1(n5369), .B2(n4276), .A(n4503), .ZN(n5295) );
  OAI21_X1 U5304 ( .B1(n5184), .B2(n4277), .A(n5295), .ZN(n5723) );
  INV_X1 U5305 ( .A(n4278), .ZN(n5726) );
  AND2_X1 U5306 ( .A1(n5726), .A2(n5727), .ZN(n5702) );
  NAND2_X1 U5307 ( .A1(n5721), .A2(n5702), .ZN(n4279) );
  AND2_X1 U5308 ( .A1(n6202), .A2(n4279), .ZN(n4280) );
  NOR2_X1 U5309 ( .A1(n5723), .A2(n4280), .ZN(n5706) );
  INV_X1 U5310 ( .A(n4281), .ZN(n4282) );
  NAND2_X1 U5311 ( .A1(n6202), .A2(n4282), .ZN(n4283) );
  NAND2_X1 U5312 ( .A1(n5706), .A2(n4283), .ZN(n5699) );
  INV_X1 U5313 ( .A(n4284), .ZN(n4285) );
  AOI21_X1 U5314 ( .B1(n6242), .B2(n6211), .A(n4285), .ZN(n4286) );
  INV_X1 U5315 ( .A(n5652), .ZN(n4287) );
  AOI21_X1 U5316 ( .B1(n6202), .B2(n5671), .A(n5691), .ZN(n5663) );
  OAI211_X1 U5317 ( .C1(n4287), .C2(n5725), .A(n5663), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U5318 ( .C1(n6202), .C2(n5691), .A(n5648), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4288) );
  AND2_X1 U5319 ( .A1(n4289), .A2(n4288), .ZN(n4290) );
  OAI21_X1 U5320 ( .B1(n5355), .B2(n6169), .A(n4290), .ZN(U2988) );
  NOR2_X1 U5321 ( .A1(n4312), .A2(n4291), .ZN(n4292) );
  XNOR2_X1 U5322 ( .A(n4292), .B(n5643), .ZN(n5650) );
  OAI21_X1 U5323 ( .B1(n4294), .B2(n4296), .A(n4295), .ZN(n5395) );
  AND2_X1 U5324 ( .A1(n6504), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U5325 ( .A1(n4332), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6511) );
  NOR2_X1 U5326 ( .A1(n5395), .A2(n5622), .ZN(n4307) );
  NAND2_X1 U5327 ( .A1(n6390), .A2(n4297), .ZN(n6602) );
  NAND2_X1 U5328 ( .A1(n6602), .A2(n6504), .ZN(n4298) );
  NAND2_X1 U5329 ( .A1(n6504), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U5330 ( .A1(n5923), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4299) );
  AND2_X1 U5331 ( .A1(n4300), .A2(n4299), .ZN(n4382) );
  NAND2_X1 U5332 ( .A1(n5404), .A2(n6130), .ZN(n4305) );
  NAND2_X1 U5333 ( .A1(n6221), .A2(REIP_REG_29__SCAN_IN), .ZN(n5644) );
  OAI21_X1 U5334 ( .B1(n5616), .B2(n4302), .A(n5644), .ZN(n4303) );
  INV_X1 U5335 ( .A(n4303), .ZN(n4304) );
  NAND2_X1 U5336 ( .A1(n4305), .A2(n4304), .ZN(n4306) );
  NOR2_X1 U5337 ( .A1(n4307), .A2(n4306), .ZN(n4308) );
  OAI21_X1 U5338 ( .B1(n5650), .B2(n6134), .A(n4308), .ZN(U2957) );
  INV_X1 U5339 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4324) );
  NOR2_X1 U5340 ( .A1(n5643), .A2(n4324), .ZN(n4311) );
  AOI21_X1 U5341 ( .B1(n4312), .B2(n4311), .A(n4310), .ZN(n4313) );
  NOR2_X1 U5342 ( .A1(n4315), .A2(EBX_REG_29__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U5343 ( .A1(n4316), .A2(n5399), .ZN(n4317) );
  OAI21_X2 U5344 ( .B1(n4318), .B2(n4045), .A(n4317), .ZN(n5398) );
  NAND2_X1 U5345 ( .A1(n5398), .A2(n4319), .ZN(n4321) );
  OAI22_X1 U5346 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4496), .ZN(n4322) );
  INV_X1 U5347 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6688) );
  NOR2_X1 U5348 ( .A1(n6183), .A2(n6688), .ZN(n5360) );
  NOR3_X1 U5349 ( .A1(n5652), .A2(n5643), .A3(n4324), .ZN(n4327) );
  INV_X1 U5350 ( .A(n4327), .ZN(n4325) );
  NOR3_X1 U5351 ( .A1(n5651), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4325), 
        .ZN(n4326) );
  OAI21_X1 U5352 ( .B1(n5725), .B2(n4327), .A(n5663), .ZN(n4328) );
  NAND2_X1 U5353 ( .A1(n4328), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4329) );
  OAI21_X1 U5354 ( .B1(n5365), .B2(n6169), .A(n4330), .ZN(U2987) );
  NAND3_X1 U5355 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4350) );
  INV_X1 U5356 ( .A(n5916), .ZN(n6476) );
  INV_X1 U5357 ( .A(n6501), .ZN(n6499) );
  NOR2_X1 U5358 ( .A1(n6475), .A2(n6499), .ZN(n4331) );
  NAND2_X1 U5359 ( .A1(n6476), .A2(n4331), .ZN(n4371) );
  NAND2_X1 U5360 ( .A1(n4332), .A2(n3920), .ZN(n6507) );
  NAND2_X1 U5361 ( .A1(n6493), .A2(n6503), .ZN(n4543) );
  INV_X1 U5362 ( .A(n4543), .ZN(n6606) );
  NAND3_X1 U5363 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6606), .ZN(n6497) );
  NAND2_X1 U5364 ( .A1(n6507), .A2(n6497), .ZN(n4333) );
  AND2_X1 U5365 ( .A1(n6708), .A2(n5923), .ZN(n4334) );
  AND3_X1 U5366 ( .A1(n4335), .A2(n4339), .A3(n4334), .ZN(n4336) );
  NAND2_X2 U5367 ( .A1(n5381), .A2(n4336), .ZN(n6046) );
  INV_X2 U5368 ( .A(n6046), .ZN(n6023) );
  INV_X1 U5369 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6553) );
  INV_X1 U5370 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6549) );
  INV_X1 U5371 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6545) );
  INV_X1 U5372 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6541) );
  INV_X1 U5373 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6537) );
  INV_X1 U5374 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6590) );
  INV_X1 U5375 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6533) );
  INV_X1 U5376 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6531) );
  NOR3_X1 U5377 ( .A1(n6590), .A2(n6533), .A3(n6531), .ZN(n5156) );
  NAND2_X1 U5378 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5156), .ZN(n6045) );
  NOR2_X1 U5379 ( .A1(n6537), .A2(n6045), .ZN(n6022) );
  NAND2_X1 U5380 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6022), .ZN(n6015) );
  NOR2_X1 U5381 ( .A1(n6541), .A2(n6015), .ZN(n6009) );
  NAND2_X1 U5382 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6009), .ZN(n5072) );
  NOR2_X1 U5383 ( .A1(n6545), .A2(n5072), .ZN(n5069) );
  NAND2_X1 U5384 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5069), .ZN(n5984) );
  NOR2_X1 U5385 ( .A1(n6549), .A2(n5984), .ZN(n5258) );
  NAND2_X1 U5386 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5258), .ZN(n5969) );
  NOR2_X1 U5387 ( .A1(n6553), .A2(n5969), .ZN(n4344) );
  NAND2_X1 U5388 ( .A1(n6023), .A2(n4344), .ZN(n5961) );
  NAND2_X1 U5389 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5319), .ZN(n5950) );
  NOR2_X2 U5390 ( .A1(n6559), .A2(n5950), .ZN(n5335) );
  NOR2_X2 U5391 ( .A1(n4350), .A2(n5838), .ZN(n5807) );
  NAND4_X1 U5392 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5807), .ZN(n5780) );
  NOR2_X1 U5393 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5780), .ZN(n5793) );
  OR3_X1 U5394 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6518), .ZN(
        n6487) );
  AND2_X1 U5395 ( .A1(n2986), .A2(n6487), .ZN(n4337) );
  NAND2_X1 U5396 ( .A1(n5381), .A2(n4337), .ZN(n4341) );
  INV_X1 U5397 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5366) );
  OAI21_X1 U5398 ( .B1(READY_N), .B2(STATEBS16_REG_SCAN_IN), .A(n5381), .ZN(
        n4338) );
  INV_X1 U5399 ( .A(n4338), .ZN(n4366) );
  NAND3_X1 U5400 ( .A1(n4339), .A2(n5366), .A3(n4366), .ZN(n4340) );
  OAI22_X1 U5401 ( .A1(n5949), .A2(n4343), .B1(n6036), .B2(n4342), .ZN(n4370)
         );
  NAND2_X1 U5402 ( .A1(n6046), .A2(n6020), .ZN(n5377) );
  INV_X1 U5403 ( .A(n4344), .ZN(n4345) );
  NOR2_X1 U5404 ( .A1(n4345), .A2(n6555), .ZN(n4346) );
  NAND2_X1 U5405 ( .A1(n6020), .A2(n4346), .ZN(n4347) );
  NAND2_X1 U5406 ( .A1(n5377), .A2(n4347), .ZN(n5960) );
  INV_X1 U5407 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6561) );
  INV_X1 U5408 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6557) );
  NOR3_X1 U5409 ( .A1(n6561), .A2(n6559), .A3(n6557), .ZN(n4348) );
  OR2_X1 U5410 ( .A1(n6046), .A2(n4348), .ZN(n4349) );
  NAND2_X1 U5411 ( .A1(n5960), .A2(n4349), .ZN(n5942) );
  AND2_X1 U5412 ( .A1(n5377), .A2(n4350), .ZN(n4351) );
  NOR2_X1 U5413 ( .A1(n5942), .A2(n4351), .ZN(n5816) );
  INV_X1 U5414 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6723) );
  INV_X1 U5415 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6750) );
  INV_X1 U5416 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6751) );
  NOR3_X1 U5417 ( .A1(n6723), .A2(n6750), .A3(n6751), .ZN(n4352) );
  OR2_X1 U5418 ( .A1(n6046), .A2(n4352), .ZN(n4353) );
  INV_X1 U5419 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6628) );
  INV_X1 U5420 ( .A(n4354), .ZN(n4355) );
  NAND2_X1 U5421 ( .A1(n4355), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4357)
         );
  INV_X1 U5422 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4356) );
  OAI22_X1 U5423 ( .A1(n5800), .A2(n6628), .B1(n5566), .B2(n6024), .ZN(n4369)
         );
  BUF_X1 U5424 ( .A(n4359), .Z(n4360) );
  AOI21_X1 U5425 ( .B1(n4362), .B2(n4360), .A(n4361), .ZN(n5568) );
  INV_X1 U5426 ( .A(n5568), .ZN(n5524) );
  NAND2_X1 U5427 ( .A1(n5470), .A2(n4364), .ZN(n4365) );
  NAND2_X1 U5428 ( .A1(n5460), .A2(n4365), .ZN(n5688) );
  AND2_X1 U5429 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4366), .ZN(n4367) );
  OAI22_X1 U5430 ( .A1(n5524), .A2(n6038), .B1(n5688), .B2(n6014), .ZN(n4368)
         );
  OR4_X1 U5431 ( .A1(n5793), .A2(n4370), .A3(n4369), .A4(n4368), .ZN(U2803) );
  INV_X1 U5432 ( .A(n4371), .ZN(n4373) );
  INV_X1 U5433 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6707) );
  AND2_X1 U5434 ( .A1(n6384), .A2(n6493), .ZN(n5068) );
  INV_X1 U5435 ( .A(n5068), .ZN(n4372) );
  OAI211_X1 U5436 ( .C1(n4373), .C2(n6707), .A(n4454), .B(n4372), .ZN(U2788)
         );
  INV_X1 U5437 ( .A(n6601), .ZN(n4376) );
  INV_X1 U5438 ( .A(n5104), .ZN(n4374) );
  NAND2_X1 U5439 ( .A1(n6605), .A2(n4374), .ZN(n5924) );
  OAI21_X1 U5440 ( .B1(n5068), .B2(READREQUEST_REG_SCAN_IN), .A(n4376), .ZN(
        n4375) );
  OAI21_X1 U5441 ( .B1(n4376), .B2(n5924), .A(n4375), .ZN(U3474) );
  NAND2_X1 U5442 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  NAND2_X1 U5443 ( .A1(n4380), .A2(n4379), .ZN(n5172) );
  XNOR2_X1 U5444 ( .A(n4381), .B(n5369), .ZN(n4452) );
  NAND2_X1 U5445 ( .A1(n4452), .A2(n6158), .ZN(n4386) );
  NAND2_X1 U5446 ( .A1(n4382), .A2(n5616), .ZN(n4384) );
  NAND2_X1 U5447 ( .A1(n6221), .A2(REIP_REG_0__SCAN_IN), .ZN(n4449) );
  INV_X1 U5448 ( .A(n4449), .ZN(n4383) );
  AOI21_X1 U5449 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4384), .A(n4383), 
        .ZN(n4385) );
  OAI211_X1 U5450 ( .C1(n5622), .C2(n5172), .A(n4386), .B(n4385), .ZN(U2986)
         );
  NAND2_X1 U5451 ( .A1(n6504), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6587) );
  INV_X1 U5452 ( .A(n6518), .ZN(n4387) );
  NAND2_X1 U5453 ( .A1(n4387), .A2(n6708), .ZN(n4388) );
  NAND2_X1 U5454 ( .A1(n4389), .A2(n4388), .ZN(n4390) );
  OAI211_X1 U5455 ( .C1(n4245), .C2(n4527), .A(n6480), .B(n4390), .ZN(n4394)
         );
  NAND2_X1 U5456 ( .A1(n5104), .A2(n4391), .ZN(n4392) );
  NAND4_X1 U5457 ( .A1(n4395), .A2(n4394), .A3(n4393), .A4(n4392), .ZN(n4397)
         );
  OR2_X1 U5458 ( .A1(n6504), .A2(n4545), .ZN(n6586) );
  INV_X1 U5459 ( .A(n6586), .ZN(n4398) );
  AOI22_X1 U5460 ( .A1(n6458), .A2(n6501), .B1(n4398), .B2(FLUSH_REG_SCAN_IN), 
        .ZN(n5910) );
  NAND2_X1 U5461 ( .A1(n6587), .A2(n5910), .ZN(n5914) );
  INV_X1 U5462 ( .A(n5914), .ZN(n4413) );
  INV_X1 U5463 ( .A(n4245), .ZN(n6488) );
  AND4_X1 U5464 ( .A1(n3985), .A2(n3281), .A3(n6488), .A4(n3995), .ZN(n4401)
         );
  NAND2_X1 U5465 ( .A1(n4402), .A2(n4401), .ZN(n5368) );
  INV_X1 U5466 ( .A(n5368), .ZN(n4416) );
  INV_X1 U5467 ( .A(n4403), .ZN(n4406) );
  INV_X1 U5468 ( .A(n4404), .ZN(n4405) );
  NAND2_X1 U5469 ( .A1(n4406), .A2(n4405), .ZN(n4409) );
  AOI22_X1 U5470 ( .A1(n4527), .A2(n3112), .B1(n5367), .B2(n4409), .ZN(n4407)
         );
  OAI21_X1 U5471 ( .B1(n4400), .B2(n4416), .A(n4407), .ZN(n6459) );
  INV_X1 U5472 ( .A(n5777), .ZN(n5372) );
  NOR2_X1 U5473 ( .A1(n6493), .A2(n5369), .ZN(n4427) );
  INV_X1 U5474 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4408) );
  AOI22_X1 U5475 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4408), .B2(n4576), .ZN(n4428)
         );
  INV_X1 U5476 ( .A(n4428), .ZN(n4410) );
  AOI222_X1 U5477 ( .A1(n6459), .A2(n5372), .B1(n4427), .B2(n4410), .C1(n4409), 
        .C2(n6491), .ZN(n4412) );
  NAND2_X1 U5478 ( .A1(n4413), .A2(n4529), .ZN(n4411) );
  OAI21_X1 U5479 ( .B1(n4413), .B2(n4412), .A(n4411), .ZN(U3460) );
  INV_X1 U5480 ( .A(n6491), .ZN(n5775) );
  OAI21_X1 U5481 ( .B1(n4414), .B2(n5775), .A(n5914), .ZN(n4432) );
  OR2_X1 U5482 ( .A1(n4415), .A2(n4416), .ZN(n4425) );
  AND2_X1 U5483 ( .A1(n4418), .A2(n4417), .ZN(n4526) );
  INV_X1 U5484 ( .A(n4526), .ZN(n4423) );
  XNOR2_X1 U5485 ( .A(n4414), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4422)
         );
  XNOR2_X1 U5486 ( .A(n3112), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4419)
         );
  NAND2_X1 U5487 ( .A1(n4527), .A2(n4419), .ZN(n4420) );
  OAI21_X1 U5488 ( .B1(n4422), .B2(n4531), .A(n4420), .ZN(n4421) );
  AOI21_X1 U5489 ( .B1(n4423), .B2(n4422), .A(n4421), .ZN(n4424) );
  NAND2_X1 U5490 ( .A1(n4425), .A2(n4424), .ZN(n4535) );
  INV_X1 U5491 ( .A(n4535), .ZN(n4430) );
  INV_X1 U5492 ( .A(n4414), .ZN(n4524) );
  NOR3_X1 U5493 ( .A1(n5775), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4524), 
        .ZN(n4426) );
  AOI21_X1 U5494 ( .B1(n4428), .B2(n4427), .A(n4426), .ZN(n4429) );
  OAI21_X1 U5495 ( .B1(n4430), .B2(n5777), .A(n4429), .ZN(n4431) );
  AOI22_X1 U5496 ( .A1(n4432), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n5914), .B2(n4431), .ZN(n4433) );
  INV_X1 U5497 ( .A(n4433), .ZN(U3459) );
  INV_X1 U5498 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4487) );
  INV_X1 U5499 ( .A(n4434), .ZN(n4435) );
  NOR2_X4 U5500 ( .A1(n4438), .A2(n6603), .ZN(n6105) );
  AOI22_X1 U5501 ( .A1(n6603), .A2(UWORD_REG_9__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4439) );
  OAI21_X1 U5502 ( .B1(n4487), .B2(n4562), .A(n4439), .ZN(U2898) );
  INV_X1 U5503 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5504 ( .A1(n6603), .A2(UWORD_REG_10__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4440) );
  OAI21_X1 U5505 ( .B1(n4491), .B2(n4562), .A(n4440), .ZN(U2897) );
  INV_X1 U5506 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U5507 ( .A1(n6603), .A2(UWORD_REG_8__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4441) );
  OAI21_X1 U5508 ( .B1(n4482), .B2(n4562), .A(n4441), .ZN(U2899) );
  INV_X1 U5509 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4459) );
  AOI22_X1 U5510 ( .A1(n6603), .A2(UWORD_REG_12__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4442) );
  OAI21_X1 U5511 ( .B1(n4459), .B2(n4562), .A(n4442), .ZN(U2895) );
  INV_X1 U5512 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U5513 ( .A1(n6603), .A2(UWORD_REG_13__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U5514 ( .B1(n4457), .B2(n4562), .A(n4443), .ZN(U2894) );
  INV_X1 U5515 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5516 ( .A1(n6603), .A2(UWORD_REG_11__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4444) );
  OAI21_X1 U5517 ( .B1(n4484), .B2(n4562), .A(n4444), .ZN(U2896) );
  INV_X1 U5518 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U5519 ( .A1(n6603), .A2(UWORD_REG_14__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4445) );
  OAI21_X1 U5520 ( .B1(n4461), .B2(n4562), .A(n4445), .ZN(U2893) );
  AOI21_X1 U5521 ( .B1(n5892), .B2(n6211), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4504) );
  NOR2_X1 U5522 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4447)
         );
  OR2_X1 U5523 ( .A1(n4448), .A2(n4447), .ZN(n5171) );
  INV_X1 U5524 ( .A(n5302), .ZN(n5894) );
  OAI21_X1 U5525 ( .B1(n4503), .B2(n5894), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4450) );
  OAI211_X1 U5526 ( .C1(n6185), .C2(n5171), .A(n4450), .B(n4449), .ZN(n4451)
         );
  AOI211_X1 U5527 ( .C1(n6241), .C2(n4452), .A(n4504), .B(n4451), .ZN(n4453)
         );
  INV_X1 U5528 ( .A(n4453), .ZN(U3018) );
  INV_X1 U5529 ( .A(n4454), .ZN(n4455) );
  AOI22_X1 U5530 ( .A1(n6122), .A2(UWORD_REG_13__SCAN_IN), .B1(n4489), .B2(
        DATAI_13_), .ZN(n4456) );
  OAI21_X1 U5531 ( .B1(n4457), .B2(n6110), .A(n4456), .ZN(U2937) );
  AOI22_X1 U5532 ( .A1(n6122), .A2(UWORD_REG_12__SCAN_IN), .B1(n4489), .B2(
        DATAI_12_), .ZN(n4458) );
  OAI21_X1 U5533 ( .B1(n4459), .B2(n6110), .A(n4458), .ZN(U2936) );
  AOI22_X1 U5534 ( .A1(n6122), .A2(UWORD_REG_14__SCAN_IN), .B1(n4489), .B2(
        DATAI_14_), .ZN(n4460) );
  OAI21_X1 U5535 ( .B1(n4461), .B2(n6110), .A(n4460), .ZN(U2938) );
  INV_X1 U5536 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U5537 ( .A1(n6122), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4462) );
  NAND2_X1 U5538 ( .A1(n4489), .A2(DATAI_0_), .ZN(n4470) );
  OAI211_X1 U5539 ( .C1(n6109), .C2(n6110), .A(n4462), .B(n4470), .ZN(U2939)
         );
  INV_X1 U5540 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U5541 ( .A1(n6122), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5542 ( .A1(n4489), .A2(DATAI_1_), .ZN(n4472) );
  OAI211_X1 U5543 ( .C1(n6104), .C2(n6110), .A(n4463), .B(n4472), .ZN(U2940)
         );
  NAND2_X1 U5544 ( .A1(n6122), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U5545 ( .A1(n4489), .A2(DATAI_5_), .ZN(n4474) );
  OAI211_X1 U5546 ( .C1(n3466), .C2(n6110), .A(n4464), .B(n4474), .ZN(U2944)
         );
  INV_X1 U5547 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U5548 ( .A1(n6122), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U5549 ( .A1(n4489), .A2(DATAI_2_), .ZN(n4476) );
  OAI211_X1 U5550 ( .C1(n6102), .C2(n6110), .A(n4465), .B(n4476), .ZN(U2941)
         );
  INV_X1 U5551 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U5552 ( .A1(n6122), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5553 ( .A1(n4489), .A2(DATAI_3_), .ZN(n4478) );
  OAI211_X1 U5554 ( .C1(n6100), .C2(n6110), .A(n4466), .B(n4478), .ZN(U2942)
         );
  INV_X1 U5555 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U5556 ( .A1(n6122), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5557 ( .A1(n4489), .A2(DATAI_4_), .ZN(n4468) );
  OAI211_X1 U5558 ( .C1(n6098), .C2(n6110), .A(n4467), .B(n4468), .ZN(U2943)
         );
  INV_X1 U5559 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U5560 ( .A1(n6122), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4469) );
  OAI211_X1 U5561 ( .C1(n4563), .C2(n6110), .A(n4469), .B(n4468), .ZN(U2928)
         );
  INV_X1 U5562 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5563 ( .A1(n6122), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4471) );
  OAI211_X1 U5564 ( .C1(n4551), .C2(n6110), .A(n4471), .B(n4470), .ZN(U2924)
         );
  NAND2_X1 U5565 ( .A1(n6122), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4473) );
  OAI211_X1 U5566 ( .C1(n3661), .C2(n6110), .A(n4473), .B(n4472), .ZN(U2925)
         );
  INV_X1 U5567 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U5568 ( .A1(n6122), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4475) );
  OAI211_X1 U5569 ( .C1(n4554), .C2(n6110), .A(n4475), .B(n4474), .ZN(U2929)
         );
  NAND2_X1 U5570 ( .A1(n6122), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4477) );
  OAI211_X1 U5571 ( .C1(n3681), .C2(n6110), .A(n4477), .B(n4476), .ZN(U2926)
         );
  INV_X1 U5572 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5573 ( .A1(n6122), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4479) );
  OAI211_X1 U5574 ( .C1(n4556), .C2(n6110), .A(n4479), .B(n4478), .ZN(U2927)
         );
  INV_X1 U5575 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4558) );
  AOI22_X1 U5576 ( .A1(n6122), .A2(UWORD_REG_7__SCAN_IN), .B1(n4489), .B2(
        DATAI_7_), .ZN(n4480) );
  OAI21_X1 U5577 ( .B1(n4558), .B2(n6110), .A(n4480), .ZN(U2931) );
  AOI22_X1 U5578 ( .A1(n6122), .A2(UWORD_REG_8__SCAN_IN), .B1(n4489), .B2(
        DATAI_8_), .ZN(n4481) );
  OAI21_X1 U5579 ( .B1(n4482), .B2(n6110), .A(n4481), .ZN(U2932) );
  AOI22_X1 U5580 ( .A1(n6122), .A2(UWORD_REG_11__SCAN_IN), .B1(n4489), .B2(
        DATAI_11_), .ZN(n4483) );
  OAI21_X1 U5581 ( .B1(n4484), .B2(n6110), .A(n4483), .ZN(U2935) );
  INV_X1 U5582 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6078) );
  AOI22_X1 U5583 ( .A1(n6122), .A2(LWORD_REG_15__SCAN_IN), .B1(n4489), .B2(
        DATAI_15_), .ZN(n4485) );
  OAI21_X1 U5584 ( .B1(n6078), .B2(n6110), .A(n4485), .ZN(U2954) );
  AOI22_X1 U5585 ( .A1(n6122), .A2(UWORD_REG_9__SCAN_IN), .B1(n4489), .B2(
        DATAI_9_), .ZN(n4486) );
  OAI21_X1 U5586 ( .B1(n4487), .B2(n6110), .A(n4486), .ZN(U2933) );
  INV_X1 U5587 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5588 ( .A1(n6122), .A2(UWORD_REG_6__SCAN_IN), .B1(n4489), .B2(
        DATAI_6_), .ZN(n4488) );
  OAI21_X1 U5589 ( .B1(n4560), .B2(n6110), .A(n4488), .ZN(U2930) );
  AOI22_X1 U5590 ( .A1(n6122), .A2(UWORD_REG_10__SCAN_IN), .B1(n4489), .B2(
        DATAI_10_), .ZN(n4490) );
  OAI21_X1 U5591 ( .B1(n4491), .B2(n6110), .A(n4490), .ZN(U2934) );
  OAI21_X1 U5592 ( .B1(n4494), .B2(n4493), .A(n4492), .ZN(n5108) );
  XNOR2_X1 U5593 ( .A(n4495), .B(n4496), .ZN(n4502) );
  AOI22_X1 U5594 ( .A1(n6062), .A2(n4502), .B1(n5495), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4497) );
  OAI21_X1 U5595 ( .B1(n5108), .B2(n5844), .A(n4497), .ZN(U2858) );
  XOR2_X1 U5596 ( .A(n4499), .B(n4498), .Z(n4564) );
  INV_X1 U5597 ( .A(n4564), .ZN(n4507) );
  INV_X2 U5598 ( .A(n6183), .ZN(n6221) );
  AND2_X1 U5599 ( .A1(n6221), .A2(REIP_REG_1__SCAN_IN), .ZN(n4566) );
  NOR3_X1 U5600 ( .A1(n5725), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4500), 
        .ZN(n4501) );
  AOI211_X1 U5601 ( .C1(n6238), .C2(n4502), .A(n4566), .B(n4501), .ZN(n4506)
         );
  OAI21_X1 U5602 ( .B1(n4504), .B2(n4503), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4505) );
  OAI211_X1 U5603 ( .C1(n4507), .C2(n6169), .A(n4506), .B(n4505), .ZN(U3017)
         );
  OAI222_X1 U5604 ( .A1(n5171), .A2(n5843), .B1(n6066), .B2(n5178), .C1(n5172), 
        .C2(n5844), .ZN(U2859) );
  INV_X1 U5605 ( .A(DATAI_1_), .ZN(n6737) );
  OAI222_X1 U5606 ( .A1(n5108), .A2(n5848), .B1(n4953), .B2(n6737), .C1(n5512), 
        .C2(n6104), .ZN(U2890) );
  NOR2_X1 U5607 ( .A1(n4509), .A2(n4510), .ZN(n4511) );
  NOR2_X1 U5608 ( .A1(n4508), .A2(n4511), .ZN(n6157) );
  INV_X1 U5609 ( .A(n6157), .ZN(n5155) );
  INV_X1 U5610 ( .A(DATAI_2_), .ZN(n6719) );
  OAI222_X1 U5611 ( .A1(n5155), .A2(n5848), .B1(n4953), .B2(n6719), .C1(n5512), 
        .C2(n6102), .ZN(U2889) );
  CLKBUF_X1 U5612 ( .A(n4512), .Z(n4634) );
  OR2_X1 U5613 ( .A1(n4508), .A2(n4513), .ZN(n4514) );
  NAND2_X1 U5614 ( .A1(n4634), .A2(n4514), .ZN(n6147) );
  AOI21_X1 U5615 ( .B1(n4516), .B2(n4515), .A(n4573), .ZN(n6222) );
  AOI22_X1 U5616 ( .A1(n6062), .A2(n6222), .B1(EBX_REG_3__SCAN_IN), .B2(n5495), 
        .ZN(n4517) );
  OAI21_X1 U5617 ( .B1(n6147), .B2(n5844), .A(n4517), .ZN(U2856) );
  INV_X1 U5618 ( .A(DATAI_0_), .ZN(n6747) );
  OAI222_X1 U5619 ( .A1(n5172), .A2(n5848), .B1(n4953), .B2(n6747), .C1(n5512), 
        .C2(n6109), .ZN(U2891) );
  OR2_X1 U5620 ( .A1(n4519), .A2(n4518), .ZN(n4520) );
  NAND2_X1 U5621 ( .A1(n4520), .A2(n4515), .ZN(n6232) );
  OAI222_X1 U5622 ( .A1(n6232), .A2(n5843), .B1(n6066), .B2(n4032), .C1(n5155), 
        .C2(n5844), .ZN(U2857) );
  INV_X1 U5623 ( .A(DATAI_3_), .ZN(n6786) );
  OAI222_X1 U5624 ( .A1(n6147), .A2(n5848), .B1(n4953), .B2(n6786), .C1(n5512), 
        .C2(n6100), .ZN(U2888) );
  AOI211_X1 U5625 ( .C1(n4522), .C2(n4524), .A(n4523), .B(n3909), .ZN(n4525)
         );
  NOR2_X1 U5626 ( .A1(n4526), .A2(n4525), .ZN(n4534) );
  INV_X1 U5627 ( .A(n4527), .ZN(n5371) );
  INV_X1 U5628 ( .A(n4522), .ZN(n4528) );
  OAI21_X1 U5629 ( .B1(n4529), .B2(n3111), .A(n4528), .ZN(n4530) );
  AOI21_X1 U5630 ( .B1(n4529), .B2(n4523), .A(n4530), .ZN(n4532) );
  NOR3_X1 U5631 ( .A1(n4530), .A2(n3021), .A3(n3333), .ZN(n5776) );
  OAI22_X1 U5632 ( .A1(n5371), .A2(n4532), .B1(n5776), .B2(n4531), .ZN(n4533)
         );
  AOI211_X1 U5633 ( .C1(n5119), .C2(n5368), .A(n4534), .B(n4533), .ZN(n5778)
         );
  MUX2_X1 U5634 ( .A(n3111), .B(n5778), .S(n6458), .Z(n6469) );
  MUX2_X1 U5635 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4535), .S(n6458), 
        .Z(n6464) );
  NAND2_X1 U5636 ( .A1(n6464), .A2(n6493), .ZN(n4539) );
  INV_X1 U5637 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6741) );
  NAND2_X1 U5638 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6741), .ZN(n4538) );
  INV_X1 U5639 ( .A(n4536), .ZN(n4537) );
  OAI22_X1 U5640 ( .A1(n6469), .A2(n4539), .B1(n4538), .B2(n4537), .ZN(n6483)
         );
  INV_X1 U5641 ( .A(n6483), .ZN(n4540) );
  NOR2_X1 U5642 ( .A1(n4540), .A2(n3118), .ZN(n4546) );
  MUX2_X1 U5643 ( .A(n6458), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4542) );
  INV_X1 U5644 ( .A(n5084), .ZN(n6307) );
  NOR2_X1 U5645 ( .A1(n3398), .A2(n6307), .ZN(n4541) );
  XNOR2_X1 U5646 ( .A(n4541), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5160)
         );
  OR3_X1 U5647 ( .A1(n5160), .A2(STATE2_REG_1__SCAN_IN), .A3(n3985), .ZN(n5911) );
  OAI21_X1 U5648 ( .B1(n4542), .B2(n5913), .A(n5911), .ZN(n6470) );
  NOR3_X1 U5649 ( .A1(n4546), .A2(n6470), .A3(FLUSH_REG_SCAN_IN), .ZN(n4544)
         );
  NOR3_X1 U5650 ( .A1(n4546), .A2(n4545), .A3(n6470), .ZN(n6494) );
  INV_X1 U5651 ( .A(n3383), .ZN(n6257) );
  AND2_X1 U5652 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6589), .ZN(n5772) );
  OAI22_X1 U5653 ( .A1(n5009), .A2(n6390), .B1(n6257), .B2(n5772), .ZN(n4547)
         );
  OAI21_X1 U5654 ( .B1(n6494), .B2(n4547), .A(n6249), .ZN(n4548) );
  OAI21_X1 U5655 ( .B1(n6249), .B2(n6455), .A(n4548), .ZN(U3465) );
  AOI22_X1 U5656 ( .A1(n6106), .A2(UWORD_REG_1__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4549) );
  OAI21_X1 U5657 ( .B1(n3661), .B2(n4562), .A(n4549), .ZN(U2906) );
  AOI22_X1 U5658 ( .A1(n6106), .A2(UWORD_REG_0__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4550) );
  OAI21_X1 U5659 ( .B1(n4551), .B2(n4562), .A(n4550), .ZN(U2907) );
  AOI22_X1 U5660 ( .A1(n6603), .A2(UWORD_REG_2__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4552) );
  OAI21_X1 U5661 ( .B1(n3681), .B2(n4562), .A(n4552), .ZN(U2905) );
  AOI22_X1 U5662 ( .A1(n6603), .A2(UWORD_REG_5__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4553) );
  OAI21_X1 U5663 ( .B1(n4554), .B2(n4562), .A(n4553), .ZN(U2902) );
  AOI22_X1 U5664 ( .A1(n6603), .A2(UWORD_REG_3__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4555) );
  OAI21_X1 U5665 ( .B1(n4556), .B2(n4562), .A(n4555), .ZN(U2904) );
  AOI22_X1 U5666 ( .A1(n6603), .A2(UWORD_REG_7__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4557) );
  OAI21_X1 U5667 ( .B1(n4558), .B2(n4562), .A(n4557), .ZN(U2900) );
  AOI22_X1 U5668 ( .A1(n6603), .A2(UWORD_REG_6__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4559) );
  OAI21_X1 U5669 ( .B1(n4560), .B2(n4562), .A(n4559), .ZN(U2901) );
  AOI22_X1 U5670 ( .A1(n6603), .A2(UWORD_REG_4__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4561) );
  OAI21_X1 U5671 ( .B1(n4563), .B2(n4562), .A(n4561), .ZN(U2903) );
  NAND2_X1 U5672 ( .A1(n4564), .A2(n6158), .ZN(n4568) );
  NOR2_X1 U5673 ( .A1(n6162), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4565)
         );
  AOI211_X1 U5674 ( .C1(n6153), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4566), 
        .B(n4565), .ZN(n4567) );
  OAI211_X1 U5675 ( .C1(n5622), .C2(n5108), .A(n4568), .B(n4567), .ZN(U2985)
         );
  OAI21_X1 U5676 ( .B1(n4569), .B2(n4572), .A(n4571), .ZN(n4640) );
  OAI21_X1 U5677 ( .B1(n4574), .B2(n4573), .A(n4727), .ZN(n4575) );
  INV_X1 U5678 ( .A(n4575), .ZN(n5164) );
  AND2_X1 U5679 ( .A1(n6221), .A2(REIP_REG_4__SCAN_IN), .ZN(n4636) );
  NOR2_X1 U5680 ( .A1(n6230), .A2(n4580), .ZN(n4582) );
  NOR2_X1 U5681 ( .A1(n6243), .A2(n4576), .ZN(n4579) );
  INV_X1 U5682 ( .A(n4579), .ZN(n4577) );
  OR2_X1 U5683 ( .A1(n6242), .A2(n4577), .ZN(n4578) );
  NAND2_X1 U5684 ( .A1(n4578), .A2(n6211), .ZN(n6223) );
  OAI211_X1 U5685 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6223), .B(n6233), .ZN(n4581) );
  INV_X1 U5686 ( .A(n6211), .ZN(n6236) );
  INV_X1 U5687 ( .A(n6233), .ZN(n6225) );
  OAI21_X1 U5688 ( .B1(n5184), .B2(n4579), .A(n5295), .ZN(n6239) );
  AOI21_X1 U5689 ( .B1(n6236), .B2(n6225), .A(n6239), .ZN(n6231) );
  OAI22_X1 U5690 ( .A1(n4582), .A2(n4581), .B1(n6231), .B2(n4580), .ZN(n4583)
         );
  AOI211_X1 U5691 ( .C1(n6238), .C2(n5164), .A(n4636), .B(n4583), .ZN(n4584)
         );
  OAI21_X1 U5692 ( .B1(n6169), .B2(n4640), .A(n4584), .ZN(U3014) );
  NOR2_X1 U5693 ( .A1(n4585), .A2(n4795), .ZN(n4600) );
  AND2_X1 U5694 ( .A1(n4585), .A2(n4874), .ZN(n4587) );
  NAND2_X1 U5695 ( .A1(n4587), .A2(n4586), .ZN(n4651) );
  NOR3_X1 U5696 ( .A1(n4789), .A2(n4701), .A3(n6390), .ZN(n4588) );
  NAND2_X1 U5697 ( .A1(n6384), .A2(n5923), .ZN(n5773) );
  INV_X1 U5698 ( .A(n5773), .ZN(n4802) );
  NAND2_X1 U5699 ( .A1(n4415), .A2(n4400), .ZN(n4846) );
  OAI21_X1 U5700 ( .B1(n4588), .B2(n4802), .A(n4643), .ZN(n4592) );
  NAND3_X1 U5701 ( .A1(n6252), .A2(n6466), .A3(n6461), .ZN(n4648) );
  NOR2_X1 U5702 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4648), .ZN(n4698)
         );
  INV_X1 U5703 ( .A(n4698), .ZN(n4590) );
  INV_X1 U5704 ( .A(n4848), .ZN(n4589) );
  OAI21_X1 U5705 ( .B1(n3109), .B2(n6503), .A(n4738), .ZN(n4804) );
  AOI211_X1 U5706 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4590), .A(n5197), .B(
        n4804), .ZN(n4591) );
  NAND2_X1 U5707 ( .A1(n4592), .A2(n4591), .ZN(n4672) );
  NAND2_X1 U5708 ( .A1(n6149), .A2(DATAI_31_), .ZN(n6453) );
  INV_X1 U5709 ( .A(DATAI_7_), .ZN(n6648) );
  AND2_X1 U5710 ( .A1(n4593), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5711 ( .A1(n3109), .A2(n5017), .ZN(n4594) );
  OAI21_X1 U5712 ( .B1(n4643), .B2(n6390), .A(n4594), .ZN(n4697) );
  NAND2_X1 U5713 ( .A1(n4624), .A2(n3015), .ZN(n6443) );
  AOI22_X1 U5714 ( .A1(n6448), .A2(n4697), .B1(n6350), .B2(n4698), .ZN(n4597)
         );
  NOR2_X1 U5715 ( .A1(n5622), .A2(n6717), .ZN(n6354) );
  NAND2_X1 U5716 ( .A1(n4701), .A2(n6354), .ZN(n4596) );
  OAI211_X1 U5717 ( .C1(n4719), .C2(n6453), .A(n4597), .B(n4596), .ZN(n4598)
         );
  AOI21_X1 U5718 ( .B1(n4672), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n4598), 
        .ZN(n4599) );
  INV_X1 U5719 ( .A(n4599), .ZN(U3027) );
  NAND2_X1 U5720 ( .A1(n6149), .A2(DATAI_17_), .ZN(n6406) );
  NAND2_X1 U5721 ( .A1(n6461), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4799) );
  NOR2_X1 U5722 ( .A1(n6252), .A2(n4799), .ZN(n5086) );
  AND2_X1 U5723 ( .A1(n5119), .A2(n3383), .ZN(n4877) );
  INV_X1 U5724 ( .A(n4400), .ZN(n4974) );
  NOR2_X1 U5725 ( .A1(n4415), .A2(n4974), .ZN(n5085) );
  AOI21_X1 U5726 ( .B1(n4877), .B2(n5085), .A(n4629), .ZN(n4604) );
  NAND2_X1 U5727 ( .A1(n4605), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5768) );
  NAND3_X1 U5728 ( .A1(n6384), .A2(n4604), .A3(n5768), .ZN(n4601) );
  OAI211_X1 U5729 ( .C1(n6384), .C2(n5086), .A(n4879), .B(n4601), .ZN(n4628)
         );
  NAND2_X1 U5730 ( .A1(n6384), .A2(n5768), .ZN(n4603) );
  NAND2_X1 U5731 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4602) );
  OAI22_X1 U5732 ( .A1(n4604), .A2(n4603), .B1(n4799), .B2(n4602), .ZN(n4627)
         );
  AOI22_X1 U5733 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4628), .B1(n6403), 
        .B2(n4627), .ZN(n4608) );
  INV_X1 U5734 ( .A(DATAI_25_), .ZN(n4606) );
  NOR2_X1 U5735 ( .A1(n5622), .A2(n4606), .ZN(n6321) );
  NAND2_X1 U5736 ( .A1(n4624), .A2(n3275), .ZN(n6400) );
  INV_X1 U5737 ( .A(n6400), .ZN(n4928) );
  AOI22_X1 U5738 ( .A1(n5145), .A2(n6321), .B1(n4928), .B2(n4629), .ZN(n4607)
         );
  OAI211_X1 U5739 ( .C1(n6406), .C2(n4821), .A(n4608), .B(n4607), .ZN(U3125)
         );
  INV_X1 U5740 ( .A(DATAI_21_), .ZN(n6788) );
  NOR2_X1 U5741 ( .A1(n5622), .A2(n6788), .ZN(n6339) );
  INV_X1 U5742 ( .A(DATAI_5_), .ZN(n6725) );
  AOI22_X1 U5743 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4628), .B1(n6431), 
        .B2(n4627), .ZN(n4611) );
  NAND2_X1 U5744 ( .A1(n6149), .A2(DATAI_29_), .ZN(n6434) );
  INV_X1 U5745 ( .A(n6434), .ZN(n6338) );
  NAND2_X1 U5746 ( .A1(n4624), .A2(n4609), .ZN(n6428) );
  AOI22_X1 U5747 ( .A1(n5145), .A2(n6338), .B1(n6337), .B2(n4629), .ZN(n4610)
         );
  OAI211_X1 U5748 ( .C1(n6429), .C2(n4821), .A(n4611), .B(n4610), .ZN(U3129)
         );
  AOI22_X1 U5749 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4628), .B1(n6410), 
        .B2(n4627), .ZN(n4614) );
  INV_X1 U5750 ( .A(DATAI_26_), .ZN(n4612) );
  NAND2_X1 U5751 ( .A1(n4624), .A2(n3249), .ZN(n6407) );
  INV_X1 U5752 ( .A(n6407), .ZN(n4914) );
  AOI22_X1 U5753 ( .A1(n5145), .A2(n6325), .B1(n4914), .B2(n4629), .ZN(n4613)
         );
  OAI211_X1 U5754 ( .C1(n6413), .C2(n4821), .A(n4614), .B(n4613), .ZN(U3126)
         );
  INV_X1 U5755 ( .A(n6367), .ZN(n6415) );
  AOI22_X1 U5756 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4628), .B1(n6417), 
        .B2(n4627), .ZN(n4616) );
  NAND2_X1 U5757 ( .A1(n6149), .A2(DATAI_27_), .ZN(n6420) );
  INV_X1 U5758 ( .A(n6420), .ZN(n6330) );
  NAND2_X1 U5759 ( .A1(n4624), .A2(n4009), .ZN(n6414) );
  AOI22_X1 U5760 ( .A1(n5145), .A2(n6330), .B1(n6329), .B2(n4629), .ZN(n4615)
         );
  OAI211_X1 U5761 ( .C1(n6415), .C2(n4821), .A(n4616), .B(n4615), .ZN(U3127)
         );
  NAND2_X1 U5762 ( .A1(n6149), .A2(DATAI_16_), .ZN(n6382) );
  AOI22_X1 U5763 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4628), .B1(n6396), 
        .B2(n4627), .ZN(n4619) );
  INV_X1 U5764 ( .A(DATAI_24_), .ZN(n4617) );
  NOR2_X1 U5765 ( .A1(n5622), .A2(n4617), .ZN(n6316) );
  NAND2_X1 U5766 ( .A1(n4624), .A2(n4339), .ZN(n6381) );
  AOI22_X1 U5767 ( .A1(n5145), .A2(n6316), .B1(n4933), .B2(n4629), .ZN(n4618)
         );
  OAI211_X1 U5768 ( .C1(n6382), .C2(n4821), .A(n4619), .B(n4618), .ZN(U3124)
         );
  NAND2_X1 U5769 ( .A1(n6149), .A2(DATAI_22_), .ZN(n6436) );
  AOI22_X1 U5770 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4628), .B1(n6438), 
        .B2(n4627), .ZN(n4623) );
  INV_X1 U5771 ( .A(DATAI_30_), .ZN(n4620) );
  NAND2_X1 U5772 ( .A1(n4624), .A2(n4621), .ZN(n6435) );
  AOI22_X1 U5773 ( .A1(n5145), .A2(n6345), .B1(n4923), .B2(n4629), .ZN(n4622)
         );
  OAI211_X1 U5774 ( .C1(n6436), .C2(n4821), .A(n4623), .B(n4622), .ZN(U3130)
         );
  INV_X1 U5775 ( .A(DATAI_20_), .ZN(n6682) );
  INV_X1 U5776 ( .A(n6375), .ZN(n6427) );
  INV_X1 U5777 ( .A(DATAI_4_), .ZN(n4718) );
  AOI22_X1 U5778 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4628), .B1(n6424), 
        .B2(n4627), .ZN(n4626) );
  NAND2_X1 U5779 ( .A1(n6149), .A2(DATAI_28_), .ZN(n6422) );
  INV_X1 U5780 ( .A(n6422), .ZN(n6334) );
  NAND2_X1 U5781 ( .A1(n4624), .A2(n3004), .ZN(n6421) );
  AOI22_X1 U5782 ( .A1(n5145), .A2(n6334), .B1(n6333), .B2(n4629), .ZN(n4625)
         );
  OAI211_X1 U5783 ( .C1(n6427), .C2(n4821), .A(n4626), .B(n4625), .ZN(U3128)
         );
  INV_X1 U5784 ( .A(n6354), .ZN(n6444) );
  AOI22_X1 U5785 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4628), .B1(n6448), 
        .B2(n4627), .ZN(n4631) );
  INV_X1 U5786 ( .A(n6453), .ZN(n6351) );
  AOI22_X1 U5787 ( .A1(n5145), .A2(n6351), .B1(n6350), .B2(n4629), .ZN(n4630)
         );
  OAI211_X1 U5788 ( .C1(n6444), .C2(n4821), .A(n4631), .B(n4630), .ZN(U3131)
         );
  INV_X1 U5789 ( .A(n4632), .ZN(n4633) );
  AOI21_X1 U5790 ( .B1(n4635), .B2(n4634), .A(n4633), .ZN(n4641) );
  AOI21_X1 U5791 ( .B1(n6153), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4636), 
        .ZN(n4637) );
  OAI21_X1 U5792 ( .B1(n5166), .B2(n6162), .A(n4637), .ZN(n4638) );
  AOI21_X1 U5793 ( .B1(n4641), .B2(n6149), .A(n4638), .ZN(n4639) );
  OAI21_X1 U5794 ( .B1(n6134), .B2(n4640), .A(n4639), .ZN(U2982) );
  INV_X1 U5795 ( .A(n4641), .ZN(n5169) );
  AOI22_X1 U5796 ( .A1(n6062), .A2(n5164), .B1(n5495), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4642) );
  OAI21_X1 U5797 ( .B1(n5169), .B2(n5844), .A(n4642), .ZN(U2855) );
  INV_X1 U5798 ( .A(n6316), .ZN(n6399) );
  INV_X1 U5799 ( .A(n4643), .ZN(n4644) );
  NOR2_X1 U5800 ( .A1(n6455), .A2(n4648), .ZN(n4668) );
  AOI21_X1 U5801 ( .B1(n4644), .B2(n3383), .A(n4668), .ZN(n4649) );
  OR2_X1 U5802 ( .A1(n4651), .A2(n5923), .ZN(n4645) );
  NAND2_X1 U5803 ( .A1(n4645), .A2(n6384), .ZN(n4650) );
  INV_X1 U5804 ( .A(n4650), .ZN(n4646) );
  AOI22_X1 U5805 ( .A1(n4649), .A2(n4646), .B1(n6390), .B2(n4648), .ZN(n4647)
         );
  NAND2_X1 U5806 ( .A1(n4879), .A2(n4647), .ZN(n4667) );
  OAI22_X1 U5807 ( .A1(n4650), .A2(n4649), .B1(n6503), .B2(n4648), .ZN(n4666)
         );
  AOI22_X1 U5808 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4667), .B1(n6396), 
        .B2(n4666), .ZN(n4653) );
  NOR2_X2 U5809 ( .A1(n4651), .A2(n5009), .ZN(n5045) );
  INV_X1 U5810 ( .A(n6382), .ZN(n5219) );
  AOI22_X1 U5811 ( .A1(n5045), .A2(n5219), .B1(n4933), .B2(n4668), .ZN(n4652)
         );
  OAI211_X1 U5812 ( .C1(n6399), .C2(n4671), .A(n4653), .B(n4652), .ZN(U3028)
         );
  AOI22_X1 U5813 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4667), .B1(n6438), 
        .B2(n4666), .ZN(n4655) );
  INV_X1 U5814 ( .A(n6436), .ZN(n5138) );
  AOI22_X1 U5815 ( .A1(n5045), .A2(n5138), .B1(n4923), .B2(n4668), .ZN(n4654)
         );
  OAI211_X1 U5816 ( .C1(n6441), .C2(n4671), .A(n4655), .B(n4654), .ZN(U3034)
         );
  AOI22_X1 U5817 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4667), .B1(n6431), 
        .B2(n4666), .ZN(n4657) );
  AOI22_X1 U5818 ( .A1(n5045), .A2(n6339), .B1(n6337), .B2(n4668), .ZN(n4656)
         );
  OAI211_X1 U5819 ( .C1(n6434), .C2(n4671), .A(n4657), .B(n4656), .ZN(U3033)
         );
  AOI22_X1 U5820 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4667), .B1(n6424), 
        .B2(n4666), .ZN(n4659) );
  AOI22_X1 U5821 ( .A1(n5045), .A2(n6375), .B1(n6333), .B2(n4668), .ZN(n4658)
         );
  OAI211_X1 U5822 ( .C1(n6422), .C2(n4671), .A(n4659), .B(n4658), .ZN(U3032)
         );
  AOI22_X1 U5823 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4667), .B1(n6417), 
        .B2(n4666), .ZN(n4661) );
  AOI22_X1 U5824 ( .A1(n5045), .A2(n6367), .B1(n6329), .B2(n4668), .ZN(n4660)
         );
  OAI211_X1 U5825 ( .C1(n6420), .C2(n4671), .A(n4661), .B(n4660), .ZN(U3031)
         );
  AOI22_X1 U5826 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4667), .B1(n6448), 
        .B2(n4666), .ZN(n4663) );
  AOI22_X1 U5827 ( .A1(n5045), .A2(n6354), .B1(n6350), .B2(n4668), .ZN(n4662)
         );
  OAI211_X1 U5828 ( .C1(n6453), .C2(n4671), .A(n4663), .B(n4662), .ZN(U3035)
         );
  AOI22_X1 U5829 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4667), .B1(n6403), 
        .B2(n4666), .ZN(n4665) );
  INV_X1 U5830 ( .A(n6406), .ZN(n6362) );
  AOI22_X1 U5831 ( .A1(n5045), .A2(n6362), .B1(n4928), .B2(n4668), .ZN(n4664)
         );
  OAI211_X1 U5832 ( .C1(n6401), .C2(n4671), .A(n4665), .B(n4664), .ZN(U3029)
         );
  INV_X1 U5833 ( .A(n6325), .ZN(n6408) );
  AOI22_X1 U5834 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4667), .B1(n6410), 
        .B2(n4666), .ZN(n4670) );
  INV_X1 U5835 ( .A(n6413), .ZN(n5212) );
  AOI22_X1 U5836 ( .A1(n5045), .A2(n5212), .B1(n4914), .B2(n4668), .ZN(n4669)
         );
  OAI211_X1 U5837 ( .C1(n6408), .C2(n4671), .A(n4670), .B(n4669), .ZN(U3030)
         );
  INV_X1 U5838 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5839 ( .A1(n6337), .A2(n4698), .B1(n6431), .B2(n4697), .ZN(n4673)
         );
  OAI21_X1 U5840 ( .B1(n6434), .B2(n4719), .A(n4673), .ZN(n4674) );
  AOI21_X1 U5841 ( .B1(n6339), .B2(n4701), .A(n4674), .ZN(n4675) );
  OAI21_X1 U5842 ( .B1(n4704), .B2(n4676), .A(n4675), .ZN(U3025) );
  INV_X1 U5843 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5844 ( .A1(n6438), .A2(n4697), .B1(n4923), .B2(n4698), .ZN(n4677)
         );
  OAI21_X1 U5845 ( .B1(n6441), .B2(n4719), .A(n4677), .ZN(n4678) );
  AOI21_X1 U5846 ( .B1(n5138), .B2(n4701), .A(n4678), .ZN(n4679) );
  OAI21_X1 U5847 ( .B1(n4704), .B2(n4680), .A(n4679), .ZN(U3026) );
  INV_X1 U5848 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5849 ( .A1(n4914), .A2(n4698), .B1(n6410), .B2(n4697), .ZN(n4681)
         );
  OAI21_X1 U5850 ( .B1(n6408), .B2(n4719), .A(n4681), .ZN(n4682) );
  AOI21_X1 U5851 ( .B1(n5212), .B2(n4701), .A(n4682), .ZN(n4683) );
  OAI21_X1 U5852 ( .B1(n4704), .B2(n4684), .A(n4683), .ZN(U3022) );
  INV_X1 U5853 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4688) );
  AOI22_X1 U5854 ( .A1(n6329), .A2(n4698), .B1(n6417), .B2(n4697), .ZN(n4685)
         );
  OAI21_X1 U5855 ( .B1(n6420), .B2(n4719), .A(n4685), .ZN(n4686) );
  AOI21_X1 U5856 ( .B1(n6367), .B2(n4701), .A(n4686), .ZN(n4687) );
  OAI21_X1 U5857 ( .B1(n4704), .B2(n4688), .A(n4687), .ZN(U3023) );
  AOI22_X1 U5858 ( .A1(n4933), .A2(n4698), .B1(n6396), .B2(n4697), .ZN(n4689)
         );
  OAI21_X1 U5859 ( .B1(n6399), .B2(n4719), .A(n4689), .ZN(n4690) );
  AOI21_X1 U5860 ( .B1(n5219), .B2(n4701), .A(n4690), .ZN(n4691) );
  OAI21_X1 U5861 ( .B1(n4704), .B2(n4692), .A(n4691), .ZN(U3020) );
  INV_X1 U5862 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5863 ( .A1(n4928), .A2(n4698), .B1(n6403), .B2(n4697), .ZN(n4693)
         );
  OAI21_X1 U5864 ( .B1(n6401), .B2(n4719), .A(n4693), .ZN(n4694) );
  AOI21_X1 U5865 ( .B1(n6362), .B2(n4701), .A(n4694), .ZN(n4695) );
  OAI21_X1 U5866 ( .B1(n4704), .B2(n4696), .A(n4695), .ZN(U3021) );
  INV_X1 U5867 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5868 ( .A1(n6333), .A2(n4698), .B1(n6424), .B2(n4697), .ZN(n4699)
         );
  OAI21_X1 U5869 ( .B1(n6422), .B2(n4719), .A(n4699), .ZN(n4700) );
  AOI21_X1 U5870 ( .B1(n6375), .B2(n4701), .A(n4700), .ZN(n4702) );
  OAI21_X1 U5871 ( .B1(n4704), .B2(n4703), .A(n4702), .ZN(U3024) );
  INV_X1 U5872 ( .A(n4710), .ZN(n4705) );
  OAI21_X1 U5873 ( .B1(n4705), .B2(n5622), .A(n5773), .ZN(n4708) );
  NAND2_X1 U5874 ( .A1(n4877), .A2(n6308), .ZN(n4706) );
  NAND2_X1 U5875 ( .A1(n4706), .A2(n4787), .ZN(n4711) );
  INV_X1 U5876 ( .A(n4711), .ZN(n4707) );
  NAND2_X1 U5877 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  OAI22_X1 U5878 ( .A1(n6441), .A2(n4792), .B1(n4719), .B2(n6436), .ZN(n4716)
         );
  NAND2_X1 U5879 ( .A1(n4711), .A2(n6384), .ZN(n4714) );
  NAND2_X1 U5880 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4712), .ZN(n4713) );
  OAI22_X1 U5881 ( .A1(n6348), .A2(n4786), .B1(n4787), .B2(n6435), .ZN(n4715)
         );
  AOI211_X1 U5882 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n4785), .A(n4716), 
        .B(n4715), .ZN(n4717) );
  INV_X1 U5883 ( .A(n4717), .ZN(U3146) );
  OAI222_X1 U5884 ( .A1(n5169), .A2(n5848), .B1(n4953), .B2(n4718), .C1(n5512), 
        .C2(n6098), .ZN(U2887) );
  OAI22_X1 U5885 ( .A1(n6453), .A2(n4792), .B1(n4719), .B2(n6444), .ZN(n4721)
         );
  OAI22_X1 U5886 ( .A1(n6358), .A2(n4786), .B1(n4787), .B2(n6443), .ZN(n4720)
         );
  AOI211_X1 U5887 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n4785), .A(n4721), 
        .B(n4720), .ZN(n4722) );
  INV_X1 U5888 ( .A(n4722), .ZN(U3147) );
  AND2_X1 U5889 ( .A1(n4724), .A2(n4632), .ZN(n4725) );
  NOR2_X1 U5890 ( .A1(n4723), .A2(n4725), .ZN(n6057) );
  INV_X1 U5891 ( .A(n6057), .ZN(n4793) );
  AOI21_X1 U5892 ( .B1(n4728), .B2(n4727), .A(n4841), .ZN(n6215) );
  AOI22_X1 U5893 ( .A1(n6062), .A2(n6215), .B1(EBX_REG_5__SCAN_IN), .B2(n5495), 
        .ZN(n4729) );
  OAI21_X1 U5894 ( .B1(n4793), .B2(n5844), .A(n4729), .ZN(U2854) );
  OAI21_X1 U5895 ( .B1(n4730), .B2(n4733), .A(n4732), .ZN(n6214) );
  AOI22_X1 U5896 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4734) );
  OAI21_X1 U5897 ( .B1(n6053), .B2(n6162), .A(n4734), .ZN(n4735) );
  AOI21_X1 U5898 ( .B1(n6057), .B2(n6149), .A(n4735), .ZN(n4736) );
  OAI21_X1 U5899 ( .B1(n6214), .B2(n6134), .A(n4736), .ZN(U2981) );
  NAND3_X1 U5900 ( .A1(n4821), .A2(n6384), .A3(n4792), .ZN(n4737) );
  AOI21_X1 U5901 ( .B1(n5773), .B2(n4737), .A(n6308), .ZN(n4742) );
  OAI21_X1 U5902 ( .B1(n5196), .B2(n6503), .A(n4738), .ZN(n4976) );
  NOR2_X1 U5903 ( .A1(n5017), .A2(n4976), .ZN(n5202) );
  INV_X1 U5904 ( .A(n5202), .ZN(n4741) );
  NOR2_X1 U5905 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4739), .ZN(n4825)
         );
  OAI21_X1 U5906 ( .B1(n6589), .B2(n4825), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n4740) );
  NOR3_X2 U5907 ( .A1(n4742), .A2(n4741), .A3(n4740), .ZN(n4832) );
  INV_X1 U5908 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4749) );
  INV_X1 U5909 ( .A(n6308), .ZN(n4743) );
  NOR2_X1 U5910 ( .A1(n4743), .A2(n6390), .ZN(n5195) );
  NAND2_X1 U5911 ( .A1(n5195), .A2(n5119), .ZN(n4745) );
  NAND3_X1 U5912 ( .A1(n5197), .A2(n5196), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U5913 ( .A1(n4745), .A2(n4744), .ZN(n4826) );
  AOI22_X1 U5914 ( .A1(n6329), .A2(n4825), .B1(n6417), .B2(n4826), .ZN(n4746)
         );
  OAI21_X1 U5915 ( .B1(n6420), .B2(n4821), .A(n4746), .ZN(n4747) );
  AOI21_X1 U5916 ( .B1(n6367), .B2(n4827), .A(n4747), .ZN(n4748) );
  OAI21_X1 U5917 ( .B1(n4832), .B2(n4749), .A(n4748), .ZN(U3135) );
  INV_X1 U5918 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U5919 ( .A1(n6337), .A2(n4825), .B1(n6431), .B2(n4826), .ZN(n4750)
         );
  OAI21_X1 U5920 ( .B1(n6434), .B2(n4821), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5921 ( .B1(n6339), .B2(n4827), .A(n4751), .ZN(n4752) );
  OAI21_X1 U5922 ( .B1(n4832), .B2(n4753), .A(n4752), .ZN(U3137) );
  INV_X1 U5923 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4757) );
  AOI22_X1 U5924 ( .A1(n4914), .A2(n4825), .B1(n6410), .B2(n4826), .ZN(n4754)
         );
  OAI21_X1 U5925 ( .B1(n6408), .B2(n4821), .A(n4754), .ZN(n4755) );
  AOI21_X1 U5926 ( .B1(n5212), .B2(n4827), .A(n4755), .ZN(n4756) );
  OAI21_X1 U5927 ( .B1(n4832), .B2(n4757), .A(n4756), .ZN(U3134) );
  INV_X1 U5928 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5929 ( .A1(n4933), .A2(n4825), .B1(n6396), .B2(n4826), .ZN(n4758)
         );
  OAI21_X1 U5930 ( .B1(n6399), .B2(n4821), .A(n4758), .ZN(n4759) );
  AOI21_X1 U5931 ( .B1(n5219), .B2(n4827), .A(n4759), .ZN(n4760) );
  OAI21_X1 U5932 ( .B1(n4832), .B2(n4761), .A(n4760), .ZN(U3132) );
  INV_X1 U5933 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5934 ( .A1(n4928), .A2(n4825), .B1(n6403), .B2(n4826), .ZN(n4762)
         );
  OAI21_X1 U5935 ( .B1(n6401), .B2(n4821), .A(n4762), .ZN(n4763) );
  AOI21_X1 U5936 ( .B1(n6362), .B2(n4827), .A(n4763), .ZN(n4764) );
  OAI21_X1 U5937 ( .B1(n4832), .B2(n4765), .A(n4764), .ZN(U3133) );
  INV_X1 U5938 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4769) );
  AOI22_X1 U5939 ( .A1(n6333), .A2(n4825), .B1(n6424), .B2(n4826), .ZN(n4766)
         );
  OAI21_X1 U5940 ( .B1(n6422), .B2(n4821), .A(n4766), .ZN(n4767) );
  AOI21_X1 U5941 ( .B1(n6375), .B2(n4827), .A(n4767), .ZN(n4768) );
  OAI21_X1 U5942 ( .B1(n4832), .B2(n4769), .A(n4768), .ZN(U3136) );
  NAND2_X1 U5943 ( .A1(n4785), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4772)
         );
  OAI22_X1 U5944 ( .A1(n6407), .A2(n4787), .B1(n4786), .B2(n6328), .ZN(n4770)
         );
  AOI21_X1 U5945 ( .B1(n4789), .B2(n5212), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5946 ( .C1(n4792), .C2(n6408), .A(n4772), .B(n4771), .ZN(U3142)
         );
  NAND2_X1 U5947 ( .A1(n4785), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4775)
         );
  OAI22_X1 U5948 ( .A1(n6381), .A2(n4787), .B1(n4786), .B2(n6319), .ZN(n4773)
         );
  AOI21_X1 U5949 ( .B1(n4789), .B2(n5219), .A(n4773), .ZN(n4774) );
  OAI211_X1 U5950 ( .C1(n4792), .C2(n6399), .A(n4775), .B(n4774), .ZN(U3140)
         );
  NAND2_X1 U5951 ( .A1(n4785), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4778)
         );
  OAI22_X1 U5952 ( .A1(n6400), .A2(n4787), .B1(n4786), .B2(n6360), .ZN(n4776)
         );
  AOI21_X1 U5953 ( .B1(n4789), .B2(n6362), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5954 ( .C1(n4792), .C2(n6401), .A(n4778), .B(n4777), .ZN(U3141)
         );
  NAND2_X1 U5955 ( .A1(n4785), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4781)
         );
  OAI22_X1 U5956 ( .A1(n6428), .A2(n4787), .B1(n4786), .B2(n6342), .ZN(n4779)
         );
  AOI21_X1 U5957 ( .B1(n4789), .B2(n6339), .A(n4779), .ZN(n4780) );
  OAI211_X1 U5958 ( .C1(n4792), .C2(n6434), .A(n4781), .B(n4780), .ZN(U3145)
         );
  NAND2_X1 U5959 ( .A1(n4785), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4784)
         );
  OAI22_X1 U5960 ( .A1(n6414), .A2(n4787), .B1(n4786), .B2(n6365), .ZN(n4782)
         );
  AOI21_X1 U5961 ( .B1(n4789), .B2(n6367), .A(n4782), .ZN(n4783) );
  OAI211_X1 U5962 ( .C1(n4792), .C2(n6420), .A(n4784), .B(n4783), .ZN(U3143)
         );
  NAND2_X1 U5963 ( .A1(n4785), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4791)
         );
  OAI22_X1 U5964 ( .A1(n6421), .A2(n4787), .B1(n4786), .B2(n6370), .ZN(n4788)
         );
  AOI21_X1 U5965 ( .B1(n4789), .B2(n6375), .A(n4788), .ZN(n4790) );
  OAI211_X1 U5966 ( .C1(n4792), .C2(n6422), .A(n4791), .B(n4790), .ZN(U3144)
         );
  OAI222_X1 U5967 ( .A1(n4793), .A2(n5848), .B1(n4953), .B2(n6725), .C1(n5512), 
        .C2(n3466), .ZN(U2886) );
  NAND2_X1 U5968 ( .A1(n5765), .A2(n4795), .ZN(n5769) );
  NOR2_X2 U5969 ( .A1(n4911), .A2(n4912), .ZN(n6301) );
  INV_X1 U5970 ( .A(n5085), .ZN(n4796) );
  NOR2_X1 U5971 ( .A1(n4796), .A2(n6390), .ZN(n5091) );
  NAND2_X1 U5972 ( .A1(n5091), .A2(n5771), .ZN(n4798) );
  NAND2_X1 U5973 ( .A1(n5197), .A2(n3109), .ZN(n4797) );
  OR2_X1 U5974 ( .A1(n4799), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4908)
         );
  OAI22_X1 U5975 ( .A1(n6348), .A2(n6298), .B1(n6435), .B2(n6299), .ZN(n4800)
         );
  AOI21_X1 U5976 ( .B1(n5138), .B2(n6301), .A(n4800), .ZN(n4808) );
  INV_X1 U5977 ( .A(n6305), .ZN(n4801) );
  NOR3_X1 U5978 ( .A1(n6301), .A2(n4801), .A3(n6390), .ZN(n4803) );
  NAND2_X1 U5979 ( .A1(n5085), .A2(n6307), .ZN(n4903) );
  OAI21_X1 U5980 ( .B1(n4803), .B2(n4802), .A(n4903), .ZN(n4806) );
  AOI211_X1 U5981 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6299), .A(n5017), .B(
        n4804), .ZN(n4805) );
  NAND2_X1 U5982 ( .A1(n6302), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4807) );
  OAI211_X1 U5983 ( .C1(n6305), .C2(n6441), .A(n4808), .B(n4807), .ZN(U3058)
         );
  OAI22_X1 U5984 ( .A1(n6358), .A2(n6298), .B1(n6443), .B2(n6299), .ZN(n4809)
         );
  AOI21_X1 U5985 ( .B1(n6354), .B2(n6301), .A(n4809), .ZN(n4811) );
  NAND2_X1 U5986 ( .A1(n6302), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4810) );
  OAI211_X1 U5987 ( .C1(n6305), .C2(n6453), .A(n4811), .B(n4810), .ZN(U3059)
         );
  NAND2_X1 U5988 ( .A1(n6302), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4814) );
  OAI22_X1 U5989 ( .A1(n6381), .A2(n6299), .B1(n6298), .B2(n6319), .ZN(n4812)
         );
  AOI21_X1 U5990 ( .B1(n6301), .B2(n5219), .A(n4812), .ZN(n4813) );
  OAI211_X1 U5991 ( .C1(n6305), .C2(n6399), .A(n4814), .B(n4813), .ZN(U3052)
         );
  NAND2_X1 U5992 ( .A1(n6302), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4817) );
  OAI22_X1 U5993 ( .A1(n6407), .A2(n6299), .B1(n6298), .B2(n6328), .ZN(n4815)
         );
  AOI21_X1 U5994 ( .B1(n6301), .B2(n5212), .A(n4815), .ZN(n4816) );
  OAI211_X1 U5995 ( .C1(n6305), .C2(n6408), .A(n4817), .B(n4816), .ZN(U3054)
         );
  NAND2_X1 U5996 ( .A1(n6302), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4820) );
  OAI22_X1 U5997 ( .A1(n6428), .A2(n6299), .B1(n6298), .B2(n6342), .ZN(n4818)
         );
  AOI21_X1 U5998 ( .B1(n6301), .B2(n6339), .A(n4818), .ZN(n4819) );
  OAI211_X1 U5999 ( .C1(n6305), .C2(n6434), .A(n4820), .B(n4819), .ZN(U3057)
         );
  INV_X1 U6000 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U6001 ( .A1(n6448), .A2(n4826), .B1(n6350), .B2(n4825), .ZN(n4823)
         );
  INV_X1 U6002 ( .A(n4821), .ZN(n4828) );
  AOI22_X1 U6003 ( .A1(n6351), .A2(n4828), .B1(n4827), .B2(n6354), .ZN(n4822)
         );
  OAI211_X1 U6004 ( .C1(n4832), .C2(n4824), .A(n4823), .B(n4822), .ZN(U3139)
         );
  INV_X1 U6005 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U6006 ( .A1(n6438), .A2(n4826), .B1(n4923), .B2(n4825), .ZN(n4830)
         );
  AOI22_X1 U6007 ( .A1(n6345), .A2(n4828), .B1(n4827), .B2(n5138), .ZN(n4829)
         );
  OAI211_X1 U6008 ( .C1(n4832), .C2(n4831), .A(n4830), .B(n4829), .ZN(U3138)
         );
  INV_X1 U6009 ( .A(n4834), .ZN(n4835) );
  XOR2_X1 U6010 ( .A(n4833), .B(n4835), .Z(n4961) );
  INV_X1 U6011 ( .A(n4961), .ZN(n6026) );
  AOI21_X1 U6012 ( .B1(n4837), .B2(n4836), .A(n4966), .ZN(n6194) );
  AOI22_X1 U6013 ( .A1(n6062), .A2(n6194), .B1(EBX_REG_7__SCAN_IN), .B2(n5495), 
        .ZN(n4838) );
  OAI21_X1 U6014 ( .B1(n6026), .B2(n5844), .A(n4838), .ZN(U2852) );
  XOR2_X1 U6015 ( .A(n4723), .B(n4839), .Z(n6139) );
  XOR2_X1 U6016 ( .A(n4841), .B(n4840), .Z(n6203) );
  AOI22_X1 U6017 ( .A1(n6062), .A2(n6203), .B1(EBX_REG_6__SCAN_IN), .B2(n5495), 
        .ZN(n4842) );
  OAI21_X1 U6018 ( .B1(n6039), .B2(n5498), .A(n4842), .ZN(U2853) );
  AOI22_X1 U6019 ( .A1(n5338), .A2(DATAI_6_), .B1(EAX_REG_6__SCAN_IN), .B2(
        n6073), .ZN(n4843) );
  OAI21_X1 U6020 ( .B1(n6039), .B2(n5848), .A(n4843), .ZN(U2885) );
  NAND3_X1 U6021 ( .A1(n4873), .A2(n6384), .A3(n6379), .ZN(n4847) );
  INV_X1 U6022 ( .A(n4846), .ZN(n4876) );
  AND2_X1 U6023 ( .A1(n4876), .A2(n5119), .ZN(n4854) );
  AOI21_X1 U6024 ( .B1(n4847), .B2(n5773), .A(n4854), .ZN(n4852) );
  NAND3_X1 U6025 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6466), .A3(n6461), .ZN(n4881) );
  NOR2_X1 U6026 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4881), .ZN(n4853)
         );
  INV_X1 U6027 ( .A(n5197), .ZN(n4850) );
  OR2_X1 U6028 ( .A1(n5196), .A2(n4848), .ZN(n4855) );
  AOI21_X1 U6029 ( .B1(n4855), .B2(STATE2_REG_2__SCAN_IN), .A(n4849), .ZN(
        n5087) );
  OAI211_X1 U6030 ( .C1(n6589), .C2(n4853), .A(n4850), .B(n5087), .ZN(n4851)
         );
  NAND2_X1 U6031 ( .A1(n6376), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4860) );
  INV_X1 U6032 ( .A(n4853), .ZN(n6372) );
  NAND2_X1 U6033 ( .A1(n4854), .A2(n6384), .ZN(n4857) );
  INV_X1 U6034 ( .A(n4855), .ZN(n5092) );
  NAND2_X1 U6035 ( .A1(n5092), .A2(n5017), .ZN(n4856) );
  OAI22_X1 U6036 ( .A1(n6381), .A2(n6372), .B1(n6371), .B2(n6319), .ZN(n4858)
         );
  AOI21_X1 U6037 ( .B1(n6316), .B2(n6353), .A(n4858), .ZN(n4859) );
  OAI211_X1 U6038 ( .C1(n4873), .C2(n6382), .A(n4860), .B(n4859), .ZN(U3084)
         );
  NAND2_X1 U6039 ( .A1(n6376), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4863) );
  OAI22_X1 U6040 ( .A1(n6407), .A2(n6372), .B1(n6371), .B2(n6328), .ZN(n4861)
         );
  AOI21_X1 U6041 ( .B1(n6325), .B2(n6353), .A(n4861), .ZN(n4862) );
  OAI211_X1 U6042 ( .C1(n4873), .C2(n6413), .A(n4863), .B(n4862), .ZN(U3086)
         );
  NAND2_X1 U6043 ( .A1(n6376), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4866) );
  OAI22_X1 U6044 ( .A1(n6428), .A2(n6372), .B1(n6371), .B2(n6342), .ZN(n4864)
         );
  AOI21_X1 U6045 ( .B1(n6338), .B2(n6353), .A(n4864), .ZN(n4865) );
  OAI211_X1 U6046 ( .C1(n4873), .C2(n6429), .A(n4866), .B(n4865), .ZN(U3089)
         );
  OAI22_X1 U6047 ( .A1(n6348), .A2(n6371), .B1(n6435), .B2(n6372), .ZN(n4867)
         );
  AOI21_X1 U6048 ( .B1(n6345), .B2(n6353), .A(n4867), .ZN(n4869) );
  NAND2_X1 U6049 ( .A1(n6376), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4868) );
  OAI211_X1 U6050 ( .C1(n4873), .C2(n6436), .A(n4869), .B(n4868), .ZN(U3090)
         );
  OAI22_X1 U6051 ( .A1(n6358), .A2(n6371), .B1(n6443), .B2(n6372), .ZN(n4870)
         );
  AOI21_X1 U6052 ( .B1(n6351), .B2(n6353), .A(n4870), .ZN(n4872) );
  NAND2_X1 U6053 ( .A1(n6376), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4871) );
  OAI211_X1 U6054 ( .C1(n4873), .C2(n6444), .A(n4872), .B(n4871), .ZN(U3091)
         );
  INV_X1 U6055 ( .A(n6386), .ZN(n4972) );
  AOI21_X1 U6056 ( .B1(n4972), .B2(n4875), .A(n6390), .ZN(n4880) );
  NOR2_X1 U6057 ( .A1(n6455), .A2(n4881), .ZN(n4900) );
  AOI21_X1 U6058 ( .B1(n4877), .B2(n4876), .A(n4900), .ZN(n4883) );
  AOI22_X1 U6059 ( .A1(n4880), .A2(n4883), .B1(n6390), .B2(n4881), .ZN(n4878)
         );
  NAND2_X1 U6060 ( .A1(n4879), .A2(n4878), .ZN(n4899) );
  INV_X1 U6061 ( .A(n4880), .ZN(n4882) );
  OAI22_X1 U6062 ( .A1(n4883), .A2(n4882), .B1(n6503), .B2(n4881), .ZN(n4898)
         );
  AOI22_X1 U6063 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4899), .B1(n6396), 
        .B2(n4898), .ZN(n4885) );
  AOI22_X1 U6064 ( .A1(n6374), .A2(n6316), .B1(n4933), .B2(n4900), .ZN(n4884)
         );
  OAI211_X1 U6065 ( .C1(n4980), .C2(n6382), .A(n4885), .B(n4884), .ZN(U3092)
         );
  AOI22_X1 U6066 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4899), .B1(n6417), 
        .B2(n4898), .ZN(n4887) );
  AOI22_X1 U6067 ( .A1(n6374), .A2(n6330), .B1(n6329), .B2(n4900), .ZN(n4886)
         );
  OAI211_X1 U6068 ( .C1(n4980), .C2(n6415), .A(n4887), .B(n4886), .ZN(U3095)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4899), .B1(n6410), 
        .B2(n4898), .ZN(n4889) );
  AOI22_X1 U6070 ( .A1(n6374), .A2(n6325), .B1(n4914), .B2(n4900), .ZN(n4888)
         );
  OAI211_X1 U6071 ( .C1(n4980), .C2(n6413), .A(n4889), .B(n4888), .ZN(U3094)
         );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4899), .B1(n6403), 
        .B2(n4898), .ZN(n4891) );
  AOI22_X1 U6073 ( .A1(n6374), .A2(n6321), .B1(n4928), .B2(n4900), .ZN(n4890)
         );
  OAI211_X1 U6074 ( .C1(n4980), .C2(n6406), .A(n4891), .B(n4890), .ZN(U3093)
         );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4899), .B1(n6431), 
        .B2(n4898), .ZN(n4893) );
  AOI22_X1 U6076 ( .A1(n6374), .A2(n6338), .B1(n6337), .B2(n4900), .ZN(n4892)
         );
  OAI211_X1 U6077 ( .C1(n4980), .C2(n6429), .A(n4893), .B(n4892), .ZN(U3097)
         );
  AOI22_X1 U6078 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4899), .B1(n6438), 
        .B2(n4898), .ZN(n4895) );
  AOI22_X1 U6079 ( .A1(n6374), .A2(n6345), .B1(n4923), .B2(n4900), .ZN(n4894)
         );
  OAI211_X1 U6080 ( .C1(n4980), .C2(n6436), .A(n4895), .B(n4894), .ZN(U3098)
         );
  AOI22_X1 U6081 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4899), .B1(n6424), 
        .B2(n4898), .ZN(n4897) );
  AOI22_X1 U6082 ( .A1(n6374), .A2(n6334), .B1(n6333), .B2(n4900), .ZN(n4896)
         );
  OAI211_X1 U6083 ( .C1(n4980), .C2(n6427), .A(n4897), .B(n4896), .ZN(U3096)
         );
  AOI22_X1 U6084 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4899), .B1(n6448), 
        .B2(n4898), .ZN(n4902) );
  AOI22_X1 U6085 ( .A1(n6374), .A2(n6351), .B1(n6350), .B2(n4900), .ZN(n4901)
         );
  OAI211_X1 U6086 ( .C1(n4980), .C2(n6444), .A(n4902), .B(n4901), .ZN(U3099)
         );
  OAI21_X1 U6087 ( .B1(n4911), .B2(n5923), .A(n6384), .ZN(n4910) );
  OR2_X1 U6088 ( .A1(n4903), .A2(n6257), .ZN(n4905) );
  NOR2_X1 U6089 ( .A1(n6455), .A2(n4908), .ZN(n4946) );
  INV_X1 U6090 ( .A(n4946), .ZN(n4904) );
  NAND2_X1 U6091 ( .A1(n4905), .A2(n4904), .ZN(n4907) );
  NOR2_X1 U6092 ( .A1(n4910), .A2(n4907), .ZN(n4906) );
  INV_X1 U6093 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4918) );
  INV_X1 U6094 ( .A(n4907), .ZN(n4909) );
  OAI22_X1 U6095 ( .A1(n4910), .A2(n4909), .B1(n4908), .B2(n6503), .ZN(n4949)
         );
  INV_X1 U6096 ( .A(n4911), .ZN(n4913) );
  AOI22_X1 U6097 ( .A1(n6301), .A2(n6325), .B1(n4914), .B2(n4946), .ZN(n4915)
         );
  OAI21_X1 U6098 ( .B1(n6413), .B2(n5237), .A(n4915), .ZN(n4916) );
  AOI21_X1 U6099 ( .B1(n6410), .B2(n4949), .A(n4916), .ZN(n4917) );
  OAI21_X1 U6100 ( .B1(n4952), .B2(n4918), .A(n4917), .ZN(U3062) );
  INV_X1 U6101 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4922) );
  AOI22_X1 U6102 ( .A1(n6301), .A2(n6334), .B1(n6333), .B2(n4946), .ZN(n4919)
         );
  OAI21_X1 U6103 ( .B1(n6427), .B2(n5237), .A(n4919), .ZN(n4920) );
  AOI21_X1 U6104 ( .B1(n6424), .B2(n4949), .A(n4920), .ZN(n4921) );
  OAI21_X1 U6105 ( .B1(n4952), .B2(n4922), .A(n4921), .ZN(U3064) );
  INV_X1 U6106 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4927) );
  AOI22_X1 U6107 ( .A1(n6301), .A2(n6345), .B1(n4923), .B2(n4946), .ZN(n4924)
         );
  OAI21_X1 U6108 ( .B1(n6436), .B2(n5237), .A(n4924), .ZN(n4925) );
  AOI21_X1 U6109 ( .B1(n6438), .B2(n4949), .A(n4925), .ZN(n4926) );
  OAI21_X1 U6110 ( .B1(n4952), .B2(n4927), .A(n4926), .ZN(U3066) );
  INV_X1 U6111 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4932) );
  AOI22_X1 U6112 ( .A1(n6301), .A2(n6321), .B1(n4928), .B2(n4946), .ZN(n4929)
         );
  OAI21_X1 U6113 ( .B1(n6406), .B2(n5237), .A(n4929), .ZN(n4930) );
  AOI21_X1 U6114 ( .B1(n6403), .B2(n4949), .A(n4930), .ZN(n4931) );
  OAI21_X1 U6115 ( .B1(n4952), .B2(n4932), .A(n4931), .ZN(U3061) );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U6117 ( .A1(n6301), .A2(n6316), .B1(n4933), .B2(n4946), .ZN(n4934)
         );
  OAI21_X1 U6118 ( .B1(n6382), .B2(n5237), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6119 ( .B1(n6396), .B2(n4949), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6120 ( .B1(n4952), .B2(n4937), .A(n4936), .ZN(U3060) );
  INV_X1 U6121 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U6122 ( .A1(n6301), .A2(n6338), .B1(n6337), .B2(n4946), .ZN(n4938)
         );
  OAI21_X1 U6123 ( .B1(n6429), .B2(n5237), .A(n4938), .ZN(n4939) );
  AOI21_X1 U6124 ( .B1(n6431), .B2(n4949), .A(n4939), .ZN(n4940) );
  OAI21_X1 U6125 ( .B1(n4952), .B2(n4941), .A(n4940), .ZN(U3065) );
  INV_X1 U6126 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6127 ( .A1(n6301), .A2(n6351), .B1(n6350), .B2(n4946), .ZN(n4942)
         );
  OAI21_X1 U6128 ( .B1(n6444), .B2(n5237), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6129 ( .B1(n6448), .B2(n4949), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6130 ( .B1(n4952), .B2(n4945), .A(n4944), .ZN(U3067) );
  INV_X1 U6131 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4951) );
  AOI22_X1 U6132 ( .A1(n6301), .A2(n6330), .B1(n6329), .B2(n4946), .ZN(n4947)
         );
  OAI21_X1 U6133 ( .B1(n6415), .B2(n5237), .A(n4947), .ZN(n4948) );
  AOI21_X1 U6134 ( .B1(n6417), .B2(n4949), .A(n4948), .ZN(n4950) );
  OAI21_X1 U6135 ( .B1(n4952), .B2(n4951), .A(n4950), .ZN(U3063) );
  OAI222_X1 U6136 ( .A1(n5512), .A2(n4954), .B1(n6648), .B2(n4953), .C1(n5848), 
        .C2(n6026), .ZN(U2884) );
  OAI21_X1 U6137 ( .B1(n3001), .B2(n4958), .A(n4957), .ZN(n6195) );
  NAND2_X1 U6138 ( .A1(n6221), .A2(REIP_REG_7__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U6139 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4959)
         );
  OAI211_X1 U6140 ( .C1(n6162), .C2(n6025), .A(n6192), .B(n4959), .ZN(n4960)
         );
  AOI21_X1 U6141 ( .B1(n4961), .B2(n6149), .A(n4960), .ZN(n4962) );
  OAI21_X1 U6142 ( .B1(n6195), .B2(n6134), .A(n4962), .ZN(U2979) );
  AOI21_X1 U6143 ( .B1(n4965), .B2(n4963), .A(n4964), .ZN(n5055) );
  INV_X1 U6144 ( .A(n5055), .ZN(n6006) );
  OR2_X1 U6145 ( .A1(n4967), .A2(n4966), .ZN(n4968) );
  NAND2_X1 U6146 ( .A1(n4968), .A2(n3045), .ZN(n6184) );
  INV_X1 U6147 ( .A(n6184), .ZN(n4969) );
  AOI22_X1 U6148 ( .A1(n6062), .A2(n4969), .B1(n5495), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4970) );
  OAI21_X1 U6149 ( .B1(n6006), .B2(n5844), .A(n4970), .ZN(U2851) );
  AOI22_X1 U6150 ( .A1(n5338), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6073), .ZN(n4971) );
  OAI21_X1 U6151 ( .B1(n6006), .B2(n5848), .A(n4971), .ZN(U2883) );
  NAND2_X1 U6152 ( .A1(n4980), .A2(n6452), .ZN(n4973) );
  AOI21_X1 U6153 ( .B1(n4973), .B2(STATEBS16_REG_SCAN_IN), .A(n6390), .ZN(
        n4978) );
  AND2_X1 U6154 ( .A1(n4415), .A2(n4974), .ZN(n5012) );
  INV_X1 U6155 ( .A(n5017), .ZN(n5088) );
  NOR2_X1 U6156 ( .A1(n5088), .A2(n6252), .ZN(n4975) );
  NOR2_X1 U6157 ( .A1(n5197), .A2(n4976), .ZN(n5014) );
  INV_X1 U6158 ( .A(n6387), .ZN(n4977) );
  NAND3_X1 U6159 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6466), .ZN(n6393) );
  OR2_X1 U6160 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6393), .ZN(n5003)
         );
  AOI22_X1 U6161 ( .A1(n4978), .A2(n4977), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5003), .ZN(n4979) );
  NAND2_X1 U6162 ( .A1(n5002), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4983)
         );
  OAI22_X1 U6163 ( .A1(n6452), .A2(n6382), .B1(n5003), .B2(n6381), .ZN(n4981)
         );
  AOI21_X1 U6164 ( .B1(n5005), .B2(n6316), .A(n4981), .ZN(n4982) );
  OAI211_X1 U6165 ( .C1(n5008), .C2(n6319), .A(n4983), .B(n4982), .ZN(U3100)
         );
  NAND2_X1 U6166 ( .A1(n5002), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4986)
         );
  OAI22_X1 U6167 ( .A1(n6452), .A2(n6429), .B1(n5003), .B2(n6428), .ZN(n4984)
         );
  AOI21_X1 U6168 ( .B1(n5005), .B2(n6338), .A(n4984), .ZN(n4985) );
  OAI211_X1 U6169 ( .C1(n5008), .C2(n6342), .A(n4986), .B(n4985), .ZN(U3105)
         );
  NAND2_X1 U6170 ( .A1(n5002), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4989)
         );
  OAI22_X1 U6171 ( .A1(n6452), .A2(n6444), .B1(n5003), .B2(n6443), .ZN(n4987)
         );
  AOI21_X1 U6172 ( .B1(n5005), .B2(n6351), .A(n4987), .ZN(n4988) );
  OAI211_X1 U6173 ( .C1(n5008), .C2(n6358), .A(n4989), .B(n4988), .ZN(U3107)
         );
  NAND2_X1 U6174 ( .A1(n5002), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4992)
         );
  OAI22_X1 U6175 ( .A1(n6452), .A2(n6436), .B1(n5003), .B2(n6435), .ZN(n4990)
         );
  AOI21_X1 U6176 ( .B1(n5005), .B2(n6345), .A(n4990), .ZN(n4991) );
  OAI211_X1 U6177 ( .C1(n5008), .C2(n6348), .A(n4992), .B(n4991), .ZN(U3106)
         );
  NAND2_X1 U6178 ( .A1(n5002), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4995)
         );
  OAI22_X1 U6179 ( .A1(n6452), .A2(n6406), .B1(n5003), .B2(n6400), .ZN(n4993)
         );
  AOI21_X1 U6180 ( .B1(n5005), .B2(n6321), .A(n4993), .ZN(n4994) );
  OAI211_X1 U6181 ( .C1(n5008), .C2(n6360), .A(n4995), .B(n4994), .ZN(U3101)
         );
  NAND2_X1 U6182 ( .A1(n5002), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4998)
         );
  OAI22_X1 U6183 ( .A1(n6452), .A2(n6413), .B1(n5003), .B2(n6407), .ZN(n4996)
         );
  AOI21_X1 U6184 ( .B1(n5005), .B2(n6325), .A(n4996), .ZN(n4997) );
  OAI211_X1 U6185 ( .C1(n5008), .C2(n6328), .A(n4998), .B(n4997), .ZN(U3102)
         );
  NAND2_X1 U6186 ( .A1(n5002), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5001)
         );
  OAI22_X1 U6187 ( .A1(n6452), .A2(n6427), .B1(n5003), .B2(n6421), .ZN(n4999)
         );
  AOI21_X1 U6188 ( .B1(n5005), .B2(n6334), .A(n4999), .ZN(n5000) );
  OAI211_X1 U6189 ( .C1(n5008), .C2(n6370), .A(n5001), .B(n5000), .ZN(U3104)
         );
  NAND2_X1 U6190 ( .A1(n5002), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5007)
         );
  OAI22_X1 U6191 ( .A1(n6452), .A2(n6415), .B1(n5003), .B2(n6414), .ZN(n5004)
         );
  AOI21_X1 U6192 ( .B1(n5005), .B2(n6330), .A(n5004), .ZN(n5006) );
  OAI211_X1 U6193 ( .C1(n5008), .C2(n6365), .A(n5007), .B(n5006), .ZN(U3103)
         );
  NAND3_X1 U6194 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6252), .A3(n6466), .ZN(n6262) );
  NOR2_X1 U6195 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6262), .ZN(n5016)
         );
  INV_X1 U6196 ( .A(n6286), .ZN(n5011) );
  OAI21_X1 U6197 ( .B1(n5011), .B2(n5045), .A(n5773), .ZN(n5013) );
  NAND2_X1 U6198 ( .A1(n5771), .A2(n5012), .ZN(n6258) );
  NAND2_X1 U6199 ( .A1(n5013), .A2(n6258), .ZN(n5015) );
  NAND2_X1 U6200 ( .A1(n5041), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5022) );
  INV_X1 U6201 ( .A(n5016), .ZN(n5042) );
  OR2_X1 U6202 ( .A1(n6258), .A2(n6390), .ZN(n5019) );
  NAND3_X1 U6203 ( .A1(n5017), .A2(n5196), .A3(n6252), .ZN(n5018) );
  OAI22_X1 U6204 ( .A1(n6400), .A2(n5042), .B1(n5043), .B2(n6360), .ZN(n5020)
         );
  AOI21_X1 U6205 ( .B1(n6321), .B2(n5045), .A(n5020), .ZN(n5021) );
  OAI211_X1 U6206 ( .C1(n6286), .C2(n6406), .A(n5022), .B(n5021), .ZN(U3037)
         );
  NAND2_X1 U6207 ( .A1(n5041), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5025) );
  OAI22_X1 U6208 ( .A1(n6407), .A2(n5042), .B1(n5043), .B2(n6328), .ZN(n5023)
         );
  AOI21_X1 U6209 ( .B1(n6325), .B2(n5045), .A(n5023), .ZN(n5024) );
  OAI211_X1 U6210 ( .C1(n6286), .C2(n6413), .A(n5025), .B(n5024), .ZN(U3038)
         );
  NAND2_X1 U6211 ( .A1(n5041), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5028) );
  OAI22_X1 U6212 ( .A1(n6421), .A2(n5042), .B1(n5043), .B2(n6370), .ZN(n5026)
         );
  AOI21_X1 U6213 ( .B1(n6334), .B2(n5045), .A(n5026), .ZN(n5027) );
  OAI211_X1 U6214 ( .C1(n6286), .C2(n6427), .A(n5028), .B(n5027), .ZN(U3040)
         );
  NAND2_X1 U6215 ( .A1(n5041), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5031) );
  OAI22_X1 U6216 ( .A1(n6381), .A2(n5042), .B1(n5043), .B2(n6319), .ZN(n5029)
         );
  AOI21_X1 U6217 ( .B1(n6316), .B2(n5045), .A(n5029), .ZN(n5030) );
  OAI211_X1 U6218 ( .C1(n6382), .C2(n6286), .A(n5031), .B(n5030), .ZN(U3036)
         );
  NAND2_X1 U6219 ( .A1(n5041), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5034) );
  OAI22_X1 U6220 ( .A1(n6348), .A2(n5043), .B1(n6435), .B2(n5042), .ZN(n5032)
         );
  AOI21_X1 U6221 ( .B1(n6345), .B2(n5045), .A(n5032), .ZN(n5033) );
  OAI211_X1 U6222 ( .C1(n6286), .C2(n6436), .A(n5034), .B(n5033), .ZN(U3042)
         );
  NAND2_X1 U6223 ( .A1(n5041), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5037) );
  OAI22_X1 U6224 ( .A1(n6428), .A2(n5042), .B1(n5043), .B2(n6342), .ZN(n5035)
         );
  AOI21_X1 U6225 ( .B1(n6338), .B2(n5045), .A(n5035), .ZN(n5036) );
  OAI211_X1 U6226 ( .C1(n6286), .C2(n6429), .A(n5037), .B(n5036), .ZN(U3041)
         );
  NAND2_X1 U6227 ( .A1(n5041), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5040) );
  OAI22_X1 U6228 ( .A1(n6414), .A2(n5042), .B1(n5043), .B2(n6365), .ZN(n5038)
         );
  AOI21_X1 U6229 ( .B1(n6330), .B2(n5045), .A(n5038), .ZN(n5039) );
  OAI211_X1 U6230 ( .C1(n6286), .C2(n6415), .A(n5040), .B(n5039), .ZN(U3039)
         );
  NAND2_X1 U6231 ( .A1(n5041), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5047) );
  OAI22_X1 U6232 ( .A1(n6358), .A2(n5043), .B1(n6443), .B2(n5042), .ZN(n5044)
         );
  AOI21_X1 U6233 ( .B1(n6351), .B2(n5045), .A(n5044), .ZN(n5046) );
  OAI211_X1 U6234 ( .C1(n6286), .C2(n6444), .A(n5047), .B(n5046), .ZN(U3043)
         );
  OAI21_X1 U6235 ( .B1(n5048), .B2(n5051), .A(n5050), .ZN(n6180) );
  INV_X1 U6236 ( .A(n6008), .ZN(n5053) );
  AOI22_X1 U6237 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5052) );
  OAI21_X1 U6238 ( .B1(n5053), .B2(n6162), .A(n5052), .ZN(n5054) );
  AOI21_X1 U6239 ( .B1(n5055), .B2(n6149), .A(n5054), .ZN(n5056) );
  OAI21_X1 U6240 ( .B1(n6180), .B2(n6134), .A(n5056), .ZN(U2978) );
  NOR2_X1 U6241 ( .A1(n4964), .A2(n5058), .ZN(n5059) );
  AOI21_X1 U6242 ( .B1(n5060), .B2(n3045), .A(n5066), .ZN(n5996) );
  AOI22_X1 U6243 ( .A1(n6062), .A2(n5996), .B1(EBX_REG_9__SCAN_IN), .B2(n5495), 
        .ZN(n5061) );
  OAI21_X1 U6244 ( .B1(n5999), .B2(n5844), .A(n5061), .ZN(U2850) );
  AOI22_X1 U6245 ( .A1(n5338), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6073), .ZN(n5062) );
  OAI21_X1 U6246 ( .B1(n5999), .B2(n5848), .A(n5062), .ZN(U2882) );
  NAND2_X1 U6247 ( .A1(n5057), .A2(n5063), .ZN(n5239) );
  OAI21_X1 U6248 ( .B1(n5057), .B2(n5063), .A(n5239), .ZN(n5272) );
  AOI22_X1 U6249 ( .A1(n5338), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6073), .ZN(n5064) );
  OAI21_X1 U6250 ( .B1(n5272), .B2(n5848), .A(n5064), .ZN(U2881) );
  XOR2_X1 U6251 ( .A(n5066), .B(n5065), .Z(n6172) );
  AOI22_X1 U6252 ( .A1(n6062), .A2(n6172), .B1(n5495), .B2(EBX_REG_10__SCAN_IN), .ZN(n5067) );
  OAI21_X1 U6253 ( .B1(n5272), .B2(n5844), .A(n5067), .ZN(U2849) );
  INV_X1 U6254 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6255 ( .A1(n6020), .A2(n5068), .ZN(n6058) );
  INV_X1 U6256 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6547) );
  NAND3_X1 U6257 ( .A1(n6023), .A2(n6547), .A3(n5069), .ZN(n5070) );
  OAI211_X1 U6258 ( .C1(n6036), .C2(n5071), .A(n6058), .B(n5070), .ZN(n5079)
         );
  NOR3_X1 U6259 ( .A1(n6046), .A2(REIP_REG_9__SCAN_IN), .A3(n5072), .ZN(n5995)
         );
  INV_X1 U6260 ( .A(n5072), .ZN(n5073) );
  OAI21_X1 U6261 ( .B1(n6046), .B2(n5073), .A(n6020), .ZN(n6010) );
  OAI21_X1 U6262 ( .B1(n5995), .B2(n6010), .A(REIP_REG_10__SCAN_IN), .ZN(n5076) );
  INV_X1 U6263 ( .A(n5268), .ZN(n5074) );
  AOI22_X1 U6264 ( .A1(n6054), .A2(n5074), .B1(n6050), .B2(n6172), .ZN(n5075)
         );
  OAI211_X1 U6265 ( .C1(n5949), .C2(n5077), .A(n5076), .B(n5075), .ZN(n5078)
         );
  NOR2_X1 U6266 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  OAI21_X1 U6267 ( .B1(n5272), .B2(n6038), .A(n5080), .ZN(U2817) );
  INV_X1 U6268 ( .A(n5145), .ZN(n5082) );
  AOI21_X1 U6269 ( .B1(n5082), .B2(n6445), .A(n5923), .ZN(n5083) );
  AOI211_X1 U6270 ( .C1(n5085), .C2(n5084), .A(n6390), .B(n5083), .ZN(n5090)
         );
  AND2_X1 U6271 ( .A1(n6455), .A2(n5086), .ZN(n5121) );
  OAI211_X1 U6272 ( .C1(n6589), .C2(n5121), .A(n5088), .B(n5087), .ZN(n5089)
         );
  NAND2_X1 U6273 ( .A1(n5091), .A2(n5119), .ZN(n5094) );
  NAND2_X1 U6274 ( .A1(n5197), .A2(n5092), .ZN(n5093) );
  INV_X1 U6275 ( .A(n5142), .ZN(n5095) );
  AOI22_X1 U6276 ( .A1(n6448), .A2(n5095), .B1(n6350), .B2(n5121), .ZN(n5097)
         );
  NAND2_X1 U6277 ( .A1(n5145), .A2(n6354), .ZN(n5096) );
  OAI211_X1 U6278 ( .C1(n6445), .C2(n6453), .A(n5097), .B(n5096), .ZN(n5098)
         );
  AOI21_X1 U6279 ( .B1(n5141), .B2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n5098), 
        .ZN(n5099) );
  INV_X1 U6280 ( .A(n5099), .ZN(U3123) );
  NAND2_X1 U6281 ( .A1(n5381), .A2(n3009), .ZN(n5100) );
  INV_X1 U6282 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5103) );
  OAI22_X1 U6283 ( .A1(n6020), .A2(n6590), .B1(n4495), .B2(n6014), .ZN(n5101)
         );
  AOI21_X1 U6284 ( .B1(n6054), .B2(n5103), .A(n5101), .ZN(n5102) );
  OAI21_X1 U6285 ( .B1(n5103), .B2(n6036), .A(n5102), .ZN(n5106) );
  NAND2_X1 U6286 ( .A1(n5381), .A2(n5104), .ZN(n5159) );
  NAND2_X1 U6287 ( .A1(n6023), .A2(n6590), .ZN(n5113) );
  OAI21_X1 U6288 ( .B1(n5159), .B2(n4400), .A(n5113), .ZN(n5105) );
  AOI211_X1 U6289 ( .C1(n6047), .C2(EBX_REG_1__SCAN_IN), .A(n5106), .B(n5105), 
        .ZN(n5107) );
  OAI21_X1 U6290 ( .B1(n5108), .B2(n6052), .A(n5107), .ZN(U2826) );
  INV_X1 U6291 ( .A(n5159), .ZN(n5175) );
  NAND2_X1 U6292 ( .A1(n6047), .A2(EBX_REG_3__SCAN_IN), .ZN(n5112) );
  INV_X1 U6293 ( .A(n6152), .ZN(n5109) );
  AOI22_X1 U6294 ( .A1(n6054), .A2(n5109), .B1(n6050), .B2(n6222), .ZN(n5111)
         );
  NAND2_X1 U6295 ( .A1(n6051), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5110)
         );
  NAND3_X1 U6296 ( .A1(n5112), .A2(n5111), .A3(n5110), .ZN(n5118) );
  NAND2_X1 U6297 ( .A1(n5113), .A2(n6020), .ZN(n5153) );
  OR2_X1 U6298 ( .A1(n5153), .A2(n6531), .ZN(n5116) );
  INV_X1 U6299 ( .A(n6020), .ZN(n5115) );
  INV_X1 U6300 ( .A(n5156), .ZN(n5114) );
  OAI21_X1 U6301 ( .B1(n5115), .B2(n5114), .A(n5377), .ZN(n5161) );
  AOI21_X1 U6302 ( .B1(n6533), .B2(n5116), .A(n5161), .ZN(n5117) );
  AOI211_X1 U6303 ( .C1(n5175), .C2(n5119), .A(n5118), .B(n5117), .ZN(n5120)
         );
  OAI21_X1 U6304 ( .B1(n6052), .B2(n6147), .A(n5120), .ZN(U2824) );
  NAND2_X1 U6305 ( .A1(n5141), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5124)
         );
  INV_X1 U6306 ( .A(n5121), .ZN(n5143) );
  OAI22_X1 U6307 ( .A1(n6400), .A2(n5143), .B1(n5142), .B2(n6360), .ZN(n5122)
         );
  AOI21_X1 U6308 ( .B1(n5145), .B2(n6362), .A(n5122), .ZN(n5123) );
  OAI211_X1 U6309 ( .C1(n6445), .C2(n6401), .A(n5124), .B(n5123), .ZN(U3117)
         );
  NAND2_X1 U6310 ( .A1(n5141), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5127)
         );
  OAI22_X1 U6311 ( .A1(n6407), .A2(n5143), .B1(n5142), .B2(n6328), .ZN(n5125)
         );
  AOI21_X1 U6312 ( .B1(n5145), .B2(n5212), .A(n5125), .ZN(n5126) );
  OAI211_X1 U6313 ( .C1(n6445), .C2(n6408), .A(n5127), .B(n5126), .ZN(U3118)
         );
  NAND2_X1 U6314 ( .A1(n5141), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5130)
         );
  OAI22_X1 U6315 ( .A1(n6421), .A2(n5143), .B1(n5142), .B2(n6370), .ZN(n5128)
         );
  AOI21_X1 U6316 ( .B1(n5145), .B2(n6375), .A(n5128), .ZN(n5129) );
  OAI211_X1 U6317 ( .C1(n6445), .C2(n6422), .A(n5130), .B(n5129), .ZN(U3120)
         );
  NAND2_X1 U6318 ( .A1(n5141), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5133)
         );
  OAI22_X1 U6319 ( .A1(n6428), .A2(n5143), .B1(n5142), .B2(n6342), .ZN(n5131)
         );
  AOI21_X1 U6320 ( .B1(n5145), .B2(n6339), .A(n5131), .ZN(n5132) );
  OAI211_X1 U6321 ( .C1(n6445), .C2(n6434), .A(n5133), .B(n5132), .ZN(U3121)
         );
  NAND2_X1 U6322 ( .A1(n5141), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5136)
         );
  OAI22_X1 U6323 ( .A1(n6414), .A2(n5143), .B1(n5142), .B2(n6365), .ZN(n5134)
         );
  AOI21_X1 U6324 ( .B1(n5145), .B2(n6367), .A(n5134), .ZN(n5135) );
  OAI211_X1 U6325 ( .C1(n6445), .C2(n6420), .A(n5136), .B(n5135), .ZN(U3119)
         );
  NAND2_X1 U6326 ( .A1(n5141), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5140)
         );
  OAI22_X1 U6327 ( .A1(n6348), .A2(n5142), .B1(n6435), .B2(n5143), .ZN(n5137)
         );
  AOI21_X1 U6328 ( .B1(n5138), .B2(n5145), .A(n5137), .ZN(n5139) );
  OAI211_X1 U6329 ( .C1(n6445), .C2(n6441), .A(n5140), .B(n5139), .ZN(U3122)
         );
  NAND2_X1 U6330 ( .A1(n5141), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5147)
         );
  OAI22_X1 U6331 ( .A1(n6381), .A2(n5143), .B1(n5142), .B2(n6319), .ZN(n5144)
         );
  AOI21_X1 U6332 ( .B1(n5145), .B2(n5219), .A(n5144), .ZN(n5146) );
  OAI211_X1 U6333 ( .C1(n6445), .C2(n6399), .A(n5147), .B(n5146), .ZN(U3116)
         );
  OAI22_X1 U6334 ( .A1(n5159), .A2(n4415), .B1(n6014), .B2(n6232), .ZN(n5152)
         );
  INV_X1 U6335 ( .A(n6161), .ZN(n5148) );
  AOI22_X1 U6336 ( .A1(n6051), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6054), 
        .B2(n5148), .ZN(n5150) );
  NAND3_X1 U6337 ( .A1(n6023), .A2(REIP_REG_1__SCAN_IN), .A3(n6531), .ZN(n5149) );
  OAI211_X1 U6338 ( .C1(n5949), .C2(n4032), .A(n5150), .B(n5149), .ZN(n5151)
         );
  AOI211_X1 U6339 ( .C1(REIP_REG_2__SCAN_IN), .C2(n5153), .A(n5152), .B(n5151), 
        .ZN(n5154) );
  OAI21_X1 U6340 ( .B1(n5155), .B2(n6052), .A(n5154), .ZN(U2825) );
  INV_X1 U6341 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5158) );
  INV_X1 U6342 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6535) );
  NAND3_X1 U6343 ( .A1(n6023), .A2(n6535), .A3(n5156), .ZN(n5157) );
  OAI211_X1 U6344 ( .C1(n6036), .C2(n5158), .A(n6058), .B(n5157), .ZN(n5163)
         );
  OAI22_X1 U6345 ( .A1(n5161), .A2(n6535), .B1(n5160), .B2(n5159), .ZN(n5162)
         );
  AOI211_X1 U6346 ( .C1(n5164), .C2(n6050), .A(n5163), .B(n5162), .ZN(n5165)
         );
  OAI21_X1 U6347 ( .B1(n6024), .B2(n5166), .A(n5165), .ZN(n5167) );
  AOI21_X1 U6348 ( .B1(EBX_REG_4__SCAN_IN), .B2(n6047), .A(n5167), .ZN(n5168)
         );
  OAI21_X1 U6349 ( .B1(n5169), .B2(n6052), .A(n5168), .ZN(U2823) );
  OAI21_X1 U6350 ( .B1(n6051), .B2(n6054), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5170) );
  OAI21_X1 U6351 ( .B1(n5171), .B2(n6014), .A(n5170), .ZN(n5174) );
  NOR2_X1 U6352 ( .A1(n6052), .A2(n5172), .ZN(n5173) );
  AOI211_X1 U6353 ( .C1(n5175), .C2(n3383), .A(n5174), .B(n5173), .ZN(n5177)
         );
  NAND2_X1 U6354 ( .A1(n5377), .A2(REIP_REG_0__SCAN_IN), .ZN(n5176) );
  OAI211_X1 U6355 ( .C1(n5949), .C2(n5178), .A(n5177), .B(n5176), .ZN(U2827)
         );
  NAND2_X1 U6356 ( .A1(n5180), .A2(n5179), .ZN(n5182) );
  XOR2_X1 U6357 ( .A(n5182), .B(n5181), .Z(n5247) );
  INV_X1 U6358 ( .A(n5188), .ZN(n6181) );
  OAI22_X1 U6359 ( .A1(n5184), .A2(n5183), .B1(n5187), .B2(n6211), .ZN(n5185)
         );
  INV_X1 U6360 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6361 ( .A1(n5295), .A2(n5186), .ZN(n6196) );
  INV_X1 U6362 ( .A(n6196), .ZN(n6191) );
  OAI21_X1 U6363 ( .B1(n5725), .B2(n6181), .A(n6191), .ZN(n6173) );
  NAND2_X1 U6364 ( .A1(n5187), .A2(n6223), .ZN(n6200) );
  NOR2_X1 U6365 ( .A1(n5188), .A2(n6200), .ZN(n6176) );
  AOI22_X1 U6366 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6173), .B1(n6176), 
        .B2(n5189), .ZN(n5192) );
  NAND2_X1 U6367 ( .A1(n6221), .A2(REIP_REG_9__SCAN_IN), .ZN(n5243) );
  INV_X1 U6368 ( .A(n5243), .ZN(n5190) );
  AOI21_X1 U6369 ( .B1(n6238), .B2(n5996), .A(n5190), .ZN(n5191) );
  OAI211_X1 U6370 ( .C1(n5247), .C2(n6169), .A(n5192), .B(n5191), .ZN(U3009)
         );
  INV_X1 U6371 ( .A(n5193), .ZN(n5194) );
  NAND2_X1 U6372 ( .A1(n6455), .A2(n3400), .ZN(n5231) );
  NAND2_X1 U6373 ( .A1(n5195), .A2(n5771), .ZN(n5199) );
  NAND3_X1 U6374 ( .A1(n5197), .A2(n5196), .A3(n6252), .ZN(n5198) );
  NAND2_X1 U6375 ( .A1(n5199), .A2(n5198), .ZN(n5235) );
  NAND3_X1 U6376 ( .A1(n6384), .A2(n5237), .A3(n5232), .ZN(n5200) );
  AOI21_X1 U6377 ( .B1(n5200), .B2(n5773), .A(n6308), .ZN(n5201) );
  AOI21_X1 U6378 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5231), .A(n5201), .ZN(
        n5203) );
  NAND3_X1 U6379 ( .A1(n6252), .A2(n5203), .A3(n5202), .ZN(n5224) );
  AOI22_X1 U6380 ( .A1(n5235), .A2(n6431), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n5224), .ZN(n5204) );
  OAI21_X1 U6381 ( .B1(n6428), .B2(n5231), .A(n5204), .ZN(n5205) );
  AOI21_X1 U6382 ( .B1(n6339), .B2(n6352), .A(n5205), .ZN(n5206) );
  OAI21_X1 U6383 ( .B1(n6434), .B2(n5237), .A(n5206), .ZN(U3073) );
  AOI22_X1 U6384 ( .A1(n5235), .A2(n6424), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n5224), .ZN(n5207) );
  OAI21_X1 U6385 ( .B1(n6421), .B2(n5231), .A(n5207), .ZN(n5208) );
  AOI21_X1 U6386 ( .B1(n6375), .B2(n6352), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6387 ( .B1(n6422), .B2(n5237), .A(n5209), .ZN(U3072) );
  AOI22_X1 U6388 ( .A1(n5235), .A2(n6410), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n5224), .ZN(n5210) );
  OAI21_X1 U6389 ( .B1(n6407), .B2(n5231), .A(n5210), .ZN(n5211) );
  AOI21_X1 U6390 ( .B1(n5212), .B2(n6352), .A(n5211), .ZN(n5213) );
  OAI21_X1 U6391 ( .B1(n6408), .B2(n5237), .A(n5213), .ZN(U3070) );
  AOI22_X1 U6392 ( .A1(n5235), .A2(n6403), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n5224), .ZN(n5214) );
  OAI21_X1 U6393 ( .B1(n6400), .B2(n5231), .A(n5214), .ZN(n5215) );
  AOI21_X1 U6394 ( .B1(n6362), .B2(n6352), .A(n5215), .ZN(n5216) );
  OAI21_X1 U6395 ( .B1(n6401), .B2(n5237), .A(n5216), .ZN(U3069) );
  AOI22_X1 U6396 ( .A1(n5235), .A2(n6396), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n5224), .ZN(n5217) );
  OAI21_X1 U6397 ( .B1(n6381), .B2(n5231), .A(n5217), .ZN(n5218) );
  AOI21_X1 U6398 ( .B1(n5219), .B2(n6352), .A(n5218), .ZN(n5220) );
  OAI21_X1 U6399 ( .B1(n6399), .B2(n5237), .A(n5220), .ZN(U3068) );
  AOI22_X1 U6400 ( .A1(n5235), .A2(n6417), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n5224), .ZN(n5221) );
  OAI21_X1 U6401 ( .B1(n6414), .B2(n5231), .A(n5221), .ZN(n5222) );
  AOI21_X1 U6402 ( .B1(n6367), .B2(n6352), .A(n5222), .ZN(n5223) );
  OAI21_X1 U6403 ( .B1(n6420), .B2(n5237), .A(n5223), .ZN(U3071) );
  INV_X1 U6404 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5225) );
  INV_X1 U6405 ( .A(n5224), .ZN(n5229) );
  OAI22_X1 U6406 ( .A1(n6435), .A2(n5231), .B1(n5225), .B2(n5229), .ZN(n5227)
         );
  NOR2_X1 U6407 ( .A1(n5232), .A2(n6436), .ZN(n5226) );
  AOI211_X1 U6408 ( .C1(n6438), .C2(n5235), .A(n5227), .B(n5226), .ZN(n5228)
         );
  OAI21_X1 U6409 ( .B1(n6441), .B2(n5237), .A(n5228), .ZN(U3074) );
  INV_X1 U6410 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5230) );
  OAI22_X1 U6411 ( .A1(n6443), .A2(n5231), .B1(n5230), .B2(n5229), .ZN(n5234)
         );
  NOR2_X1 U6412 ( .A1(n5232), .A2(n6444), .ZN(n5233) );
  AOI211_X1 U6413 ( .C1(n6448), .C2(n5235), .A(n5234), .B(n5233), .ZN(n5236)
         );
  OAI21_X1 U6414 ( .B1(n6453), .B2(n5237), .A(n5236), .ZN(U3075) );
  INV_X1 U6415 ( .A(n5248), .ZN(n5238) );
  AOI21_X1 U6416 ( .B1(n5240), .B2(n5239), .A(n5238), .ZN(n6131) );
  INV_X1 U6417 ( .A(n6131), .ZN(n5242) );
  AOI22_X1 U6418 ( .A1(n5338), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6073), .ZN(n5241) );
  OAI21_X1 U6419 ( .B1(n5242), .B2(n5848), .A(n5241), .ZN(U2880) );
  OAI21_X1 U6420 ( .B1(n5616), .B2(n5993), .A(n5243), .ZN(n5245) );
  NOR2_X1 U6421 ( .A1(n5999), .A2(n5622), .ZN(n5244) );
  AOI211_X1 U6422 ( .C1(n6130), .C2(n5997), .A(n5245), .B(n5244), .ZN(n5246)
         );
  OAI21_X1 U6423 ( .B1(n5247), .B2(n6134), .A(n5246), .ZN(U2977) );
  XOR2_X1 U6424 ( .A(n5249), .B(n5248), .Z(n5293) );
  INV_X1 U6425 ( .A(n5293), .ZN(n5264) );
  OR2_X1 U6426 ( .A1(n5251), .A2(n5250), .ZN(n5253) );
  NAND2_X1 U6427 ( .A1(n5253), .A2(n5252), .ZN(n5304) );
  INV_X1 U6428 ( .A(n5304), .ZN(n5254) );
  AOI22_X1 U6429 ( .A1(n6062), .A2(n5254), .B1(n5495), .B2(EBX_REG_12__SCAN_IN), .ZN(n5255) );
  OAI21_X1 U6430 ( .B1(n5264), .B2(n5844), .A(n5255), .ZN(U2847) );
  AOI22_X1 U6431 ( .A1(n5338), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6073), .ZN(n5256) );
  OAI21_X1 U6432 ( .B1(n5264), .B2(n5848), .A(n5256), .ZN(U2879) );
  INV_X1 U6433 ( .A(n5291), .ZN(n5262) );
  INV_X1 U6434 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6551) );
  OR2_X1 U6435 ( .A1(n6046), .A2(n5258), .ZN(n5257) );
  AND2_X1 U6436 ( .A1(n5257), .A2(n6020), .ZN(n5983) );
  OAI22_X1 U6437 ( .A1(n6551), .A2(n5983), .B1(n6014), .B2(n5304), .ZN(n5261)
         );
  AOI22_X1 U6438 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6051), .B1(
        EBX_REG_12__SCAN_IN), .B2(n6047), .ZN(n5259) );
  NAND3_X1 U6439 ( .A1(n6023), .A2(n6551), .A3(n5258), .ZN(n5974) );
  NAND3_X1 U6440 ( .A1(n5259), .A2(n6058), .A3(n5974), .ZN(n5260) );
  AOI211_X1 U6441 ( .C1(n6054), .C2(n5262), .A(n5261), .B(n5260), .ZN(n5263)
         );
  OAI21_X1 U6442 ( .B1(n5264), .B2(n6038), .A(n5263), .ZN(U2815) );
  NAND2_X1 U6443 ( .A1(n6126), .A2(n5266), .ZN(n5267) );
  XNOR2_X1 U6444 ( .A(n5265), .B(n5267), .ZN(n6174) );
  NAND2_X1 U6445 ( .A1(n6174), .A2(n6158), .ZN(n5271) );
  AND2_X1 U6446 ( .A1(n6221), .A2(REIP_REG_10__SCAN_IN), .ZN(n6171) );
  NOR2_X1 U6447 ( .A1(n6162), .A2(n5268), .ZN(n5269) );
  AOI211_X1 U6448 ( .C1(n6153), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6171), 
        .B(n5269), .ZN(n5270) );
  OAI211_X1 U6449 ( .C1(n5622), .C2(n5272), .A(n5271), .B(n5270), .ZN(U2976)
         );
  OAI21_X1 U6450 ( .B1(n3042), .B2(n5275), .A(n5274), .ZN(n5976) );
  AOI22_X1 U6451 ( .A1(n5338), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6073), .ZN(n5276) );
  OAI21_X1 U6452 ( .B1(n5976), .B2(n5848), .A(n5276), .ZN(U2878) );
  AOI21_X1 U6453 ( .B1(n5278), .B2(n5252), .A(n5277), .ZN(n5979) );
  AOI22_X1 U6454 ( .A1(n6062), .A2(n5979), .B1(EBX_REG_13__SCAN_IN), .B2(n5495), .ZN(n5279) );
  OAI21_X1 U6455 ( .B1(n5976), .B2(n5844), .A(n5279), .ZN(U2846) );
  OAI21_X1 U6456 ( .B1(n5280), .B2(n5282), .A(n5281), .ZN(n5345) );
  AOI22_X1 U6457 ( .A1(n5338), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6073), .ZN(n5283) );
  OAI21_X1 U6458 ( .B1(n5345), .B2(n5848), .A(n5283), .ZN(U2877) );
  OR2_X1 U6459 ( .A1(n5284), .A2(n5277), .ZN(n5285) );
  NAND2_X1 U6460 ( .A1(n5285), .A2(n3024), .ZN(n5968) );
  OAI222_X1 U6461 ( .A1(n5345), .A2(n5844), .B1(n5286), .B2(n6066), .C1(n5968), 
        .C2(n5843), .ZN(U2845) );
  NOR2_X1 U6462 ( .A1(n5288), .A2(n3046), .ZN(n5289) );
  XNOR2_X1 U6463 ( .A(n5287), .B(n5289), .ZN(n5309) );
  AOI22_X1 U6464 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5290) );
  OAI21_X1 U6465 ( .B1(n5291), .B2(n6162), .A(n5290), .ZN(n5292) );
  AOI21_X1 U6466 ( .B1(n5293), .B2(n6149), .A(n5292), .ZN(n5294) );
  OAI21_X1 U6467 ( .B1(n5309), .B2(n6134), .A(n5294), .ZN(U2974) );
  AOI22_X1 U6468 ( .A1(n5296), .A2(n6191), .B1(n5295), .B2(n5725), .ZN(n6166)
         );
  OR3_X1 U6469 ( .A1(n5892), .A2(n5369), .A3(n5301), .ZN(n5298) );
  NAND3_X1 U6470 ( .A1(n5302), .A2(n5298), .A3(n6211), .ZN(n5297) );
  OAI221_X1 U6471 ( .B1(n6166), .B2(n6164), .C1(n6166), .C2(n5297), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5308) );
  OAI21_X1 U6472 ( .B1(n5299), .B2(n6211), .A(n5298), .ZN(n5300) );
  INV_X1 U6473 ( .A(n5300), .ZN(n5895) );
  OAI21_X1 U6474 ( .B1(n5302), .B2(n5301), .A(n5895), .ZN(n6165) );
  AND3_X1 U6475 ( .A1(n5303), .A2(n6165), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5306) );
  OAI22_X1 U6476 ( .A1(n6185), .A2(n5304), .B1(n6551), .B2(n6183), .ZN(n5305)
         );
  NOR2_X1 U6477 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  OAI211_X1 U6478 ( .C1(n5309), .C2(n6169), .A(n5308), .B(n5307), .ZN(U3006)
         );
  OAI21_X1 U6479 ( .B1(n5310), .B2(n5312), .A(n5311), .ZN(n5621) );
  AOI21_X1 U6480 ( .B1(n3027), .B2(n5314), .A(n5500), .ZN(n5878) );
  AOI22_X1 U6481 ( .A1(n6062), .A2(n5878), .B1(EBX_REG_17__SCAN_IN), .B2(n5495), .ZN(n5315) );
  OAI21_X1 U6482 ( .B1(n5621), .B2(n5498), .A(n5315), .ZN(U2842) );
  INV_X1 U6483 ( .A(n5316), .ZN(n5317) );
  AOI21_X1 U6484 ( .B1(n5318), .B2(n5281), .A(n5317), .ZN(n5640) );
  NAND2_X1 U6485 ( .A1(n5319), .A2(n6557), .ZN(n5953) );
  AOI21_X1 U6486 ( .B1(n5321), .B2(n3024), .A(n5320), .ZN(n5886) );
  INV_X1 U6487 ( .A(n5886), .ZN(n5325) );
  INV_X1 U6488 ( .A(n5638), .ZN(n5322) );
  NAND2_X1 U6489 ( .A1(n6054), .A2(n5322), .ZN(n5324) );
  INV_X1 U6490 ( .A(n6058), .ZN(n6032) );
  AOI21_X1 U6491 ( .B1(n6051), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6032), 
        .ZN(n5323) );
  OAI211_X1 U6492 ( .C1(n5325), .C2(n6014), .A(n5324), .B(n5323), .ZN(n5326)
         );
  AOI21_X1 U6493 ( .B1(EBX_REG_15__SCAN_IN), .B2(n6047), .A(n5326), .ZN(n5327)
         );
  OAI211_X1 U6494 ( .C1(n6557), .C2(n5960), .A(n5953), .B(n5327), .ZN(n5328)
         );
  AOI21_X1 U6495 ( .B1(n5640), .B2(n5989), .A(n5328), .ZN(n5329) );
  INV_X1 U6496 ( .A(n5329), .ZN(U2812) );
  AOI22_X1 U6497 ( .A1(n6070), .A2(DATAI_17_), .B1(n6073), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6498 ( .A1(n6074), .A2(DATAI_1_), .ZN(n5330) );
  OAI211_X1 U6499 ( .C1(n5621), .C2(n5848), .A(n5331), .B(n5330), .ZN(U2874)
         );
  INV_X1 U6500 ( .A(n5878), .ZN(n5333) );
  AOI22_X1 U6501 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6051), .B1(n6054), 
        .B2(n5618), .ZN(n5332) );
  OAI211_X1 U6502 ( .C1(n5333), .C2(n6014), .A(n5332), .B(n6058), .ZN(n5334)
         );
  AOI21_X1 U6503 ( .B1(EBX_REG_17__SCAN_IN), .B2(n6047), .A(n5334), .ZN(n5337)
         );
  OAI21_X1 U6504 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5335), .A(n5942), .ZN(n5336) );
  OAI211_X1 U6505 ( .C1(n5621), .C2(n6038), .A(n5337), .B(n5336), .ZN(U2810)
         );
  INV_X1 U6506 ( .A(n5640), .ZN(n5341) );
  AOI22_X1 U6507 ( .A1(n5338), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6073), .ZN(n5339) );
  OAI21_X1 U6508 ( .B1(n5341), .B2(n5848), .A(n5339), .ZN(U2876) );
  AOI22_X1 U6509 ( .A1(n6062), .A2(n5886), .B1(EBX_REG_15__SCAN_IN), .B2(n5495), .ZN(n5340) );
  OAI21_X1 U6510 ( .B1(n5341), .B2(n5844), .A(n5340), .ZN(U2844) );
  XNOR2_X1 U6511 ( .A(n2985), .B(n5343), .ZN(n5344) );
  XNOR2_X1 U6512 ( .A(n2997), .B(n5344), .ZN(n5896) );
  INV_X1 U6513 ( .A(n5345), .ZN(n5965) );
  AOI22_X1 U6514 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5346) );
  OAI21_X1 U6515 ( .B1(n6162), .B2(n5347), .A(n5346), .ZN(n5348) );
  AOI21_X1 U6516 ( .B1(n5965), .B2(n6149), .A(n5348), .ZN(n5349) );
  OAI21_X1 U6517 ( .B1(n5896), .B2(n6134), .A(n5349), .ZN(U2972) );
  NAND2_X1 U6518 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5350)
         );
  OAI211_X1 U6519 ( .C1(n6162), .C2(n5412), .A(n5351), .B(n5350), .ZN(n5352)
         );
  AOI21_X1 U6520 ( .B1(n5353), .B2(n6149), .A(n5352), .ZN(n5354) );
  OAI21_X1 U6521 ( .B1(n5355), .B2(n6134), .A(n5354), .ZN(U2956) );
  NOR2_X2 U6522 ( .A1(n4295), .A2(n5356), .ZN(n5359) );
  AOI22_X1 U6523 ( .A1(n3385), .A2(EAX_REG_31__SCAN_IN), .B1(n5357), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5358) );
  AOI21_X1 U6524 ( .B1(n6153), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5360), 
        .ZN(n5361) );
  OAI21_X1 U6525 ( .B1(n6162), .B2(n5362), .A(n5361), .ZN(n5363) );
  AOI21_X1 U6526 ( .B1(n5514), .B2(n6149), .A(n5363), .ZN(n5364) );
  OAI21_X1 U6527 ( .B1(n5365), .B2(n6134), .A(n5364), .ZN(U2955) );
  OAI22_X1 U6528 ( .A1(n5384), .A2(n5843), .B1(n6066), .B2(n5366), .ZN(U2828)
         );
  AOI22_X1 U6529 ( .A1(n3383), .A2(n5368), .B1(n5367), .B2(n5375), .ZN(n6454)
         );
  AOI22_X1 U6530 ( .A1(n6491), .A2(n5375), .B1(n5369), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n5370) );
  OAI21_X1 U6531 ( .B1(n6454), .B2(n5777), .A(n5370), .ZN(n5373) );
  NOR2_X1 U6532 ( .A1(n5371), .A2(n5375), .ZN(n6457) );
  AOI22_X1 U6533 ( .A1(n5914), .A2(n5373), .B1(n5372), .B2(n6457), .ZN(n5374)
         );
  OAI21_X1 U6534 ( .B1(n5914), .B2(n5375), .A(n5374), .ZN(U3461) );
  INV_X1 U6535 ( .A(n5514), .ZN(n5394) );
  NAND3_X1 U6536 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5376) );
  NAND3_X1 U6537 ( .A1(n5441), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5386) );
  INV_X1 U6538 ( .A(n5386), .ZN(n5411) );
  INV_X1 U6539 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U6540 ( .A1(n5411), .A2(n6685), .ZN(n5408) );
  NAND2_X1 U6541 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  INV_X1 U6542 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U6543 ( .A1(n6733), .A2(n6726), .ZN(n5379) );
  OR2_X1 U6544 ( .A1(n6046), .A2(n5379), .ZN(n5380) );
  NAND2_X1 U6545 ( .A1(n5408), .A2(n5429), .ZN(n5419) );
  INV_X1 U6546 ( .A(n5419), .ZN(n5391) );
  NAND2_X1 U6547 ( .A1(n6051), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5383)
         );
  NAND4_X1 U6548 ( .A1(n5381), .A2(n2986), .A3(EBX_REG_31__SCAN_IN), .A4(n6487), .ZN(n5382) );
  OAI211_X1 U6549 ( .C1(n5384), .C2(n6014), .A(n5383), .B(n5382), .ZN(n5385)
         );
  INV_X1 U6550 ( .A(n5385), .ZN(n5390) );
  INV_X1 U6551 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6748) );
  AOI21_X1 U6552 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6688), .A(n6748), .ZN(n5387) );
  AOI211_X1 U6553 ( .C1(n6748), .C2(n6688), .A(n5387), .B(n5386), .ZN(n5388)
         );
  INV_X1 U6554 ( .A(n5388), .ZN(n5389) );
  INV_X1 U6555 ( .A(n5392), .ZN(n5393) );
  OAI21_X1 U6556 ( .B1(n5394), .B2(n6038), .A(n5393), .ZN(U2796) );
  AOI22_X1 U6557 ( .A1(n6070), .A2(DATAI_29_), .B1(n6073), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6558 ( .A1(n6074), .A2(DATAI_13_), .ZN(n5396) );
  OAI211_X1 U6559 ( .C1(n5395), .C2(n5848), .A(n5397), .B(n5396), .ZN(U2862)
         );
  INV_X1 U6560 ( .A(n5398), .ZN(n5403) );
  AOI21_X1 U6561 ( .B1(n5400), .B2(n5484), .A(n5399), .ZN(n5401) );
  NAND2_X1 U6562 ( .A1(n3065), .A2(n5401), .ZN(n5402) );
  NAND2_X1 U6563 ( .A1(n5403), .A2(n5402), .ZN(n5645) );
  AOI22_X1 U6564 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6051), .B1(n6054), 
        .B2(n5404), .ZN(n5405) );
  OAI21_X1 U6565 ( .B1(n5645), .B2(n6014), .A(n5405), .ZN(n5407) );
  NOR2_X1 U6566 ( .A1(n5429), .A2(n6685), .ZN(n5406) );
  AOI211_X1 U6567 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6047), .A(n5407), .B(n5406), 
        .ZN(n5409) );
  OAI211_X1 U6568 ( .C1(n5395), .C2(n6038), .A(n5409), .B(n5408), .ZN(U2798)
         );
  INV_X1 U6569 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5410) );
  OAI222_X1 U6570 ( .A1(n5498), .A2(n5395), .B1(n5410), .B2(n6066), .C1(n5645), 
        .C2(n5843), .ZN(U2830) );
  NAND3_X1 U6571 ( .A1(n5411), .A2(REIP_REG_29__SCAN_IN), .A3(n6748), .ZN(
        n5416) );
  INV_X1 U6572 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5413) );
  OAI22_X1 U6573 ( .A1(n5413), .A2(n6036), .B1(n6024), .B2(n5412), .ZN(n5414)
         );
  AOI21_X1 U6574 ( .B1(EBX_REG_30__SCAN_IN), .B2(n6047), .A(n5414), .ZN(n5415)
         );
  OAI211_X1 U6575 ( .C1(n6014), .C2(n5417), .A(n5416), .B(n5415), .ZN(n5418)
         );
  AOI21_X1 U6576 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5419), .A(n5418), .ZN(n5420) );
  OAI21_X1 U6577 ( .B1(n5421), .B2(n6038), .A(n5420), .ZN(U2797) );
  AOI21_X1 U6578 ( .B1(n5423), .B2(n5422), .A(n4294), .ZN(n5538) );
  INV_X1 U6579 ( .A(n5538), .ZN(n5519) );
  INV_X1 U6580 ( .A(n5424), .ZN(n5427) );
  INV_X1 U6581 ( .A(n5425), .ZN(n5426) );
  AOI21_X1 U6582 ( .B1(n5427), .B2(n5426), .A(n4316), .ZN(n5656) );
  AOI22_X1 U6583 ( .A1(n5656), .A2(n6050), .B1(PHYADDRPOINTER_REG_28__SCAN_IN), 
        .B2(n6051), .ZN(n5428) );
  OAI21_X1 U6584 ( .B1(n5536), .B2(n6024), .A(n5428), .ZN(n5431) );
  NOR2_X1 U6585 ( .A1(n5429), .A2(n6733), .ZN(n5430) );
  AOI211_X1 U6586 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6047), .A(n5431), .B(n5430), 
        .ZN(n5433) );
  NAND3_X1 U6587 ( .A1(n5441), .A2(REIP_REG_27__SCAN_IN), .A3(n6733), .ZN(
        n5432) );
  OAI211_X1 U6588 ( .C1(n5519), .C2(n6038), .A(n5433), .B(n5432), .ZN(U2799)
         );
  AOI22_X1 U6589 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6051), .B1(
        EBX_REG_27__SCAN_IN), .B2(n6047), .ZN(n5436) );
  OAI21_X1 U6590 ( .B1(n5782), .B2(n6726), .A(n5436), .ZN(n5440) );
  NOR2_X1 U6591 ( .A1(n5451), .A2(n5437), .ZN(n5438) );
  OR2_X1 U6592 ( .A1(n5425), .A2(n5438), .ZN(n5662) );
  NOR2_X1 U6593 ( .A1(n5662), .A2(n6014), .ZN(n5439) );
  AOI211_X1 U6594 ( .C1(n6054), .C2(n5547), .A(n5440), .B(n5439), .ZN(n5443)
         );
  NAND2_X1 U6595 ( .A1(n5441), .A2(n6726), .ZN(n5442) );
  OAI211_X1 U6596 ( .C1(n5544), .C2(n6038), .A(n5443), .B(n5442), .ZN(U2800)
         );
  AOI22_X1 U6597 ( .A1(n5656), .A2(n6062), .B1(EBX_REG_28__SCAN_IN), .B2(n5495), .ZN(n5444) );
  OAI21_X1 U6598 ( .B1(n5519), .B2(n5498), .A(n5444), .ZN(U2831) );
  OAI22_X1 U6599 ( .A1(n5662), .A2(n5843), .B1(n5445), .B2(n6066), .ZN(n5446)
         );
  INV_X1 U6600 ( .A(n5446), .ZN(n5447) );
  OAI21_X1 U6601 ( .B1(n5544), .B2(n5498), .A(n5447), .ZN(U2832) );
  NOR2_X1 U6602 ( .A1(n5448), .A2(n5449), .ZN(n5450) );
  INV_X1 U6603 ( .A(n5451), .ZN(n5454) );
  NAND2_X1 U6604 ( .A1(n3038), .A2(n5452), .ZN(n5453) );
  NAND2_X1 U6605 ( .A1(n5454), .A2(n5453), .ZN(n5781) );
  INV_X1 U6606 ( .A(n5781), .ZN(n5455) );
  AOI22_X1 U6607 ( .A1(n5455), .A2(n6062), .B1(EBX_REG_26__SCAN_IN), .B2(n5495), .ZN(n5456) );
  OAI21_X1 U6608 ( .B1(n5550), .B2(n5498), .A(n5456), .ZN(U2833) );
  NOR2_X1 U6609 ( .A1(n4361), .A2(n5457), .ZN(n5458) );
  INV_X1 U6610 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6611 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U6612 ( .A1(n3038), .A2(n5461), .ZN(n5790) );
  OAI222_X1 U6613 ( .A1(n5852), .A2(n5498), .B1(n5462), .B2(n6066), .C1(n5790), 
        .C2(n5843), .ZN(U2834) );
  INV_X1 U6614 ( .A(n5688), .ZN(n5463) );
  AOI22_X1 U6615 ( .A1(n6062), .A2(n5463), .B1(EBX_REG_24__SCAN_IN), .B2(n5495), .ZN(n5464) );
  OAI21_X1 U6616 ( .B1(n5524), .B2(n5498), .A(n5464), .ZN(U2835) );
  INV_X1 U6617 ( .A(n4360), .ZN(n5466) );
  AOI21_X1 U6618 ( .B1(n5467), .B2(n5465), .A(n5466), .ZN(n5578) );
  INV_X1 U6619 ( .A(n5578), .ZN(n5801) );
  OR2_X1 U6620 ( .A1(n3037), .A2(n5468), .ZN(n5469) );
  AND2_X1 U6621 ( .A1(n5470), .A2(n5469), .ZN(n5803) );
  AOI22_X1 U6622 ( .A1(n6062), .A2(n5803), .B1(EBX_REG_23__SCAN_IN), .B2(n5495), .ZN(n5471) );
  OAI21_X1 U6623 ( .B1(n5801), .B2(n5498), .A(n5471), .ZN(U2836) );
  INV_X1 U6624 ( .A(n5465), .ZN(n5473) );
  AOI21_X1 U6625 ( .B1(n5474), .B2(n5472), .A(n5473), .ZN(n5856) );
  INV_X1 U6626 ( .A(n5856), .ZN(n5477) );
  AOI21_X1 U6627 ( .B1(n5475), .B2(n5714), .A(n3037), .ZN(n5809) );
  INV_X1 U6628 ( .A(n5809), .ZN(n5476) );
  OAI222_X1 U6629 ( .A1(n5498), .A2(n5477), .B1(n6066), .B2(n5813), .C1(n5476), 
        .C2(n5843), .ZN(U2837) );
  NOR2_X1 U6630 ( .A1(n3030), .A2(n5479), .ZN(n5480) );
  OR2_X1 U6631 ( .A1(n5478), .A2(n5480), .ZN(n5598) );
  INV_X1 U6632 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6633 ( .A1(n5481), .A2(n5482), .ZN(n5483) );
  OAI21_X1 U6634 ( .B1(n5481), .B2(n5484), .A(n5483), .ZN(n5487) );
  INV_X1 U6635 ( .A(n5485), .ZN(n5486) );
  XNOR2_X1 U6636 ( .A(n5487), .B(n5486), .ZN(n5830) );
  OAI222_X1 U6637 ( .A1(n5598), .A2(n5498), .B1(n5488), .B2(n6066), .C1(n5843), 
        .C2(n5830), .ZN(U2839) );
  AND2_X1 U6638 ( .A1(n5489), .A2(n5490), .ZN(n5491) );
  OR2_X1 U6639 ( .A1(n5491), .A2(n3030), .ZN(n5831) );
  NAND2_X1 U6640 ( .A1(n4045), .A2(EBX_REG_18__SCAN_IN), .ZN(n5492) );
  AND2_X1 U6641 ( .A1(n5493), .A2(n5492), .ZN(n5501) );
  NAND2_X1 U6642 ( .A1(n5501), .A2(n5500), .ZN(n5499) );
  XNOR2_X1 U6643 ( .A(n5499), .B(n5494), .ZN(n5841) );
  INV_X1 U6644 ( .A(n5841), .ZN(n5496) );
  AOI22_X1 U6645 ( .A1(n6062), .A2(n5496), .B1(EBX_REG_19__SCAN_IN), .B2(n5495), .ZN(n5497) );
  OAI21_X1 U6646 ( .B1(n5831), .B2(n5498), .A(n5497), .ZN(U2840) );
  OAI21_X1 U6647 ( .B1(n5501), .B2(n5500), .A(n5499), .ZN(n5940) );
  NAND2_X1 U6648 ( .A1(n5311), .A2(n5502), .ZN(n5503) );
  INV_X1 U6649 ( .A(n6067), .ZN(n5504) );
  OAI222_X1 U6650 ( .A1(n5940), .A2(n5843), .B1(n5505), .B2(n6066), .C1(n5504), 
        .C2(n5844), .ZN(U2841) );
  AOI21_X1 U6651 ( .B1(n5506), .B2(n5316), .A(n5310), .ZN(n6072) );
  OR2_X1 U6652 ( .A1(n5507), .A2(n5320), .ZN(n5508) );
  NAND2_X1 U6653 ( .A1(n5508), .A2(n3027), .ZN(n5958) );
  OAI22_X1 U6654 ( .A1(n5843), .A2(n5958), .B1(n6066), .B2(n5509), .ZN(n5510)
         );
  AOI21_X1 U6655 ( .B1(n6072), .B2(n6063), .A(n5510), .ZN(n5511) );
  INV_X1 U6656 ( .A(n5511), .ZN(U2843) );
  NAND3_X1 U6657 ( .A1(n5514), .A2(n5513), .A3(n5512), .ZN(n5516) );
  AOI22_X1 U6658 ( .A1(n6070), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6073), .ZN(n5515) );
  NAND2_X1 U6659 ( .A1(n5516), .A2(n5515), .ZN(U2860) );
  AOI22_X1 U6660 ( .A1(n6070), .A2(DATAI_28_), .B1(n6073), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U6661 ( .A1(n6074), .A2(DATAI_12_), .ZN(n5517) );
  OAI211_X1 U6662 ( .C1(n5519), .C2(n5848), .A(n5518), .B(n5517), .ZN(U2863)
         );
  AOI22_X1 U6663 ( .A1(n6070), .A2(DATAI_27_), .B1(n6073), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U6664 ( .A1(n6074), .A2(DATAI_11_), .ZN(n5520) );
  OAI211_X1 U6665 ( .C1(n5544), .C2(n5848), .A(n5521), .B(n5520), .ZN(U2864)
         );
  AOI22_X1 U6666 ( .A1(n6074), .A2(DATAI_8_), .B1(n6073), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U6667 ( .A1(n6070), .A2(DATAI_24_), .ZN(n5522) );
  OAI211_X1 U6668 ( .C1(n5524), .C2(n5848), .A(n5523), .B(n5522), .ZN(U2867)
         );
  AOI22_X1 U6669 ( .A1(n6074), .A2(DATAI_7_), .B1(n6073), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6670 ( .A1(n6070), .A2(DATAI_23_), .ZN(n5525) );
  OAI211_X1 U6671 ( .C1(n5801), .C2(n5848), .A(n5526), .B(n5525), .ZN(U2868)
         );
  INV_X1 U6672 ( .A(n5528), .ZN(n5530) );
  NAND2_X1 U6673 ( .A1(n5683), .A2(n5531), .ZN(n5670) );
  NOR2_X1 U6674 ( .A1(n2985), .A2(n5670), .ZN(n5529) );
  NAND2_X1 U6675 ( .A1(n5530), .A2(n5529), .ZN(n5541) );
  AND2_X1 U6676 ( .A1(n5531), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5532)
         );
  XNOR2_X1 U6677 ( .A(n5534), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5660)
         );
  NOR2_X1 U6678 ( .A1(n6183), .A2(n6733), .ZN(n5655) );
  AOI21_X1 U6679 ( .B1(n6153), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5655), 
        .ZN(n5535) );
  OAI21_X1 U6680 ( .B1(n5536), .B2(n6162), .A(n5535), .ZN(n5537) );
  AOI21_X1 U6681 ( .B1(n5538), .B2(n6149), .A(n5537), .ZN(n5539) );
  OAI21_X1 U6682 ( .B1(n6134), .B2(n5660), .A(n5539), .ZN(U2958) );
  NAND2_X1 U6683 ( .A1(n5540), .A2(n5541), .ZN(n5542) );
  XNOR2_X1 U6684 ( .A(n5542), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5669)
         );
  NAND2_X1 U6685 ( .A1(n6221), .A2(REIP_REG_27__SCAN_IN), .ZN(n5661) );
  OAI21_X1 U6686 ( .B1(n5616), .B2(n5543), .A(n5661), .ZN(n5546) );
  NOR2_X1 U6687 ( .A1(n5544), .A2(n5622), .ZN(n5545) );
  OAI21_X1 U6688 ( .B1(n5669), .B2(n6134), .A(n5548), .ZN(U2959) );
  XNOR2_X1 U6689 ( .A(n2985), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5549)
         );
  XNOR2_X1 U6690 ( .A(n4229), .B(n5549), .ZN(n5676) );
  NOR2_X1 U6691 ( .A1(n6162), .A2(n5787), .ZN(n5553) );
  NAND2_X1 U6692 ( .A1(n6221), .A2(REIP_REG_26__SCAN_IN), .ZN(n5672) );
  OAI21_X1 U6693 ( .B1(n5616), .B2(n5551), .A(n5672), .ZN(n5552) );
  AOI211_X1 U6694 ( .C1(n5849), .C2(n6149), .A(n5553), .B(n5552), .ZN(n5554)
         );
  OAI21_X1 U6695 ( .B1(n6134), .B2(n5676), .A(n5554), .ZN(U2960) );
  NAND2_X1 U6696 ( .A1(n6221), .A2(REIP_REG_25__SCAN_IN), .ZN(n5678) );
  OAI21_X1 U6697 ( .B1(n5616), .B2(n5555), .A(n5678), .ZN(n5556) );
  AOI21_X1 U6698 ( .B1(n6130), .B2(n5789), .A(n5556), .ZN(n5560) );
  OAI21_X1 U6699 ( .B1(n5558), .B2(n5557), .A(n3023), .ZN(n5677) );
  NAND2_X1 U6700 ( .A1(n5677), .A2(n6158), .ZN(n5559) );
  OAI211_X1 U6701 ( .C1(n5852), .C2(n5622), .A(n5560), .B(n5559), .ZN(U2961)
         );
  XNOR2_X1 U6702 ( .A(n2985), .B(n5735), .ZN(n5605) );
  AND2_X1 U6703 ( .A1(n2985), .A2(n5595), .ZN(n5562) );
  OR2_X1 U6704 ( .A1(n2985), .A2(n5595), .ZN(n5561) );
  OAI21_X2 U6705 ( .B1(n5597), .B2(n5562), .A(n5561), .ZN(n5588) );
  XNOR2_X1 U6706 ( .A(n2985), .B(n5703), .ZN(n5589) );
  NOR2_X1 U6707 ( .A1(n2985), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5580)
         );
  NAND2_X1 U6708 ( .A1(n5587), .A2(n5580), .ZN(n5572) );
  OAI21_X1 U6709 ( .B1(n3035), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n3005), 
        .ZN(n5582) );
  NAND3_X1 U6710 ( .A1(n2985), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5563) );
  XNOR2_X1 U6711 ( .A(n5564), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5693)
         );
  NAND2_X1 U6712 ( .A1(n6221), .A2(REIP_REG_24__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U6713 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5565)
         );
  OAI211_X1 U6714 ( .C1(n6162), .C2(n5566), .A(n5687), .B(n5565), .ZN(n5567)
         );
  AOI21_X1 U6715 ( .B1(n5568), .B2(n6149), .A(n5567), .ZN(n5569) );
  OAI21_X1 U6716 ( .B1(n5693), .B2(n6134), .A(n5569), .ZN(U2962) );
  NAND2_X1 U6717 ( .A1(n2985), .A2(n5571), .ZN(n5573) );
  OAI21_X1 U6718 ( .B1(n5570), .B2(n5573), .A(n5572), .ZN(n5574) );
  XNOR2_X1 U6719 ( .A(n5574), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5701)
         );
  INV_X1 U6720 ( .A(n5798), .ZN(n5576) );
  NAND2_X1 U6721 ( .A1(n6221), .A2(REIP_REG_23__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6722 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5575)
         );
  OAI211_X1 U6723 ( .C1(n6162), .C2(n5576), .A(n5694), .B(n5575), .ZN(n5577)
         );
  AOI21_X1 U6724 ( .B1(n5578), .B2(n6149), .A(n5577), .ZN(n5579) );
  OAI21_X1 U6725 ( .B1(n5701), .B2(n6134), .A(n5579), .ZN(U2963) );
  AOI21_X1 U6726 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2985), .A(n5580), 
        .ZN(n5581) );
  XNOR2_X1 U6727 ( .A(n5582), .B(n5581), .ZN(n5710) );
  INV_X1 U6728 ( .A(n5810), .ZN(n5584) );
  AND2_X1 U6729 ( .A1(n6221), .A2(REIP_REG_22__SCAN_IN), .ZN(n5705) );
  AOI21_X1 U6730 ( .B1(n6153), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5705), 
        .ZN(n5583) );
  OAI21_X1 U6731 ( .B1(n5584), .B2(n6162), .A(n5583), .ZN(n5585) );
  AOI21_X1 U6732 ( .B1(n5856), .B2(n6149), .A(n5585), .ZN(n5586) );
  OAI21_X1 U6733 ( .B1(n5710), .B2(n6134), .A(n5586), .ZN(U2964) );
  AOI21_X1 U6734 ( .B1(n5589), .B2(n5588), .A(n5587), .ZN(n5720) );
  NAND2_X1 U6735 ( .A1(n6221), .A2(REIP_REG_21__SCAN_IN), .ZN(n5715) );
  OAI21_X1 U6736 ( .B1(n5616), .B2(n5590), .A(n5715), .ZN(n5593) );
  XNOR2_X1 U6737 ( .A(n5478), .B(n5591), .ZN(n5859) );
  NOR2_X1 U6738 ( .A1(n5859), .A2(n5622), .ZN(n5592) );
  AOI211_X1 U6739 ( .C1(n6130), .C2(n5817), .A(n5593), .B(n5592), .ZN(n5594)
         );
  OAI21_X1 U6740 ( .B1(n5720), .B2(n6134), .A(n5594), .ZN(U2965) );
  XNOR2_X1 U6741 ( .A(n2985), .B(n5595), .ZN(n5596) );
  XNOR2_X1 U6742 ( .A(n5597), .B(n5596), .ZN(n5734) );
  NAND2_X1 U6743 ( .A1(n6221), .A2(REIP_REG_20__SCAN_IN), .ZN(n5730) );
  INV_X1 U6744 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5599) );
  OR2_X1 U6745 ( .A1(n5616), .A2(n5599), .ZN(n5600) );
  OAI211_X1 U6746 ( .C1(n6162), .C2(n5823), .A(n5730), .B(n5600), .ZN(n5601)
         );
  AOI21_X1 U6747 ( .B1(n5863), .B2(n6149), .A(n5601), .ZN(n5602) );
  OAI21_X1 U6748 ( .B1(n5734), .B2(n6134), .A(n5602), .ZN(U2966) );
  XOR2_X1 U6749 ( .A(n5605), .B(n5604), .Z(n5742) );
  INV_X1 U6750 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6751 ( .A1(n6221), .A2(REIP_REG_19__SCAN_IN), .ZN(n5737) );
  OAI21_X1 U6752 ( .B1(n5616), .B2(n5606), .A(n5737), .ZN(n5608) );
  NOR2_X1 U6753 ( .A1(n5831), .A2(n5622), .ZN(n5607) );
  AOI211_X1 U6754 ( .C1(n6130), .C2(n5832), .A(n5608), .B(n5607), .ZN(n5609)
         );
  OAI21_X1 U6755 ( .B1(n5742), .B2(n6134), .A(n5609), .ZN(U2967) );
  OR2_X1 U6756 ( .A1(n2985), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5613)
         );
  AOI21_X1 U6757 ( .B1(n3035), .B2(n5747), .A(n5610), .ZN(n5611) );
  AOI21_X1 U6758 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5613), .A(n5611), 
        .ZN(n5615) );
  NOR3_X1 U6759 ( .A1(n5610), .A2(n3035), .A3(n5747), .ZN(n5744) );
  NOR3_X1 U6760 ( .A1(n3000), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5613), 
        .ZN(n5743) );
  INV_X1 U6761 ( .A(n5743), .ZN(n5614) );
  OAI21_X1 U6762 ( .B1(n5615), .B2(n5744), .A(n5614), .ZN(n5879) );
  NAND2_X1 U6763 ( .A1(n5879), .A2(n6158), .ZN(n5620) );
  OAI22_X1 U6764 ( .A1(n5616), .A2(n3665), .B1(n6183), .B2(n6561), .ZN(n5617)
         );
  AOI21_X1 U6765 ( .B1(n6130), .B2(n5618), .A(n5617), .ZN(n5619) );
  OAI211_X1 U6766 ( .C1(n5622), .C2(n5621), .A(n5620), .B(n5619), .ZN(U2969)
         );
  OAI211_X1 U6767 ( .C1(n3035), .C2(n3000), .A(n5610), .B(n5631), .ZN(n5623)
         );
  NAND2_X1 U6768 ( .A1(n5623), .A2(n5758), .ZN(n5626) );
  INV_X1 U6769 ( .A(n3000), .ZN(n5624) );
  NAND3_X1 U6770 ( .A1(n5624), .A2(n3035), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5625) );
  OAI211_X1 U6771 ( .C1(n3035), .C2(n5610), .A(n5626), .B(n5625), .ZN(n5762)
         );
  NAND2_X1 U6772 ( .A1(n6221), .A2(REIP_REG_16__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6773 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5627)
         );
  OAI211_X1 U6774 ( .C1(n6162), .C2(n5628), .A(n5756), .B(n5627), .ZN(n5629)
         );
  AOI21_X1 U6775 ( .B1(n6072), .B2(n6149), .A(n5629), .ZN(n5630) );
  OAI21_X1 U6776 ( .B1(n5762), .B2(n6134), .A(n5630), .ZN(U2970) );
  INV_X1 U6777 ( .A(n5631), .ZN(n5632) );
  NOR2_X1 U6778 ( .A1(n5633), .A2(n5632), .ZN(n5636) );
  BUF_X1 U6779 ( .A(n5634), .Z(n5635) );
  XOR2_X1 U6780 ( .A(n5636), .B(n5635), .Z(n5887) );
  INV_X1 U6781 ( .A(n5887), .ZN(n5642) );
  AOI22_X1 U6782 ( .A1(n6153), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5637) );
  OAI21_X1 U6783 ( .B1(n5638), .B2(n6162), .A(n5637), .ZN(n5639) );
  AOI21_X1 U6784 ( .B1(n5640), .B2(n6149), .A(n5639), .ZN(n5641) );
  OAI21_X1 U6785 ( .B1(n5642), .B2(n6134), .A(n5641), .ZN(U2971) );
  OAI21_X1 U6786 ( .B1(n5651), .B2(n5652), .A(n5643), .ZN(n5647) );
  OAI21_X1 U6787 ( .B1(n5645), .B2(n6185), .A(n5644), .ZN(n5646) );
  AOI21_X1 U6788 ( .B1(n5648), .B2(n5647), .A(n5646), .ZN(n5649) );
  OAI21_X1 U6789 ( .B1(n5650), .B2(n6169), .A(n5649), .ZN(U2989) );
  INV_X1 U6790 ( .A(n5651), .ZN(n5667) );
  AND3_X1 U6791 ( .A1(n5667), .A2(n5653), .A3(n5652), .ZN(n5654) );
  AOI211_X1 U6792 ( .C1(n6238), .C2(n5656), .A(n5655), .B(n5654), .ZN(n5659)
         );
  INV_X1 U6793 ( .A(n5663), .ZN(n5657) );
  NAND2_X1 U6794 ( .A1(n5657), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5658) );
  OAI211_X1 U6795 ( .C1(n5660), .C2(n6169), .A(n5659), .B(n5658), .ZN(U2990)
         );
  OAI21_X1 U6796 ( .B1(n5662), .B2(n6185), .A(n5661), .ZN(n5665) );
  NOR2_X1 U6797 ( .A1(n5663), .A2(n5666), .ZN(n5664) );
  AOI211_X1 U6798 ( .C1(n5667), .C2(n5666), .A(n5665), .B(n5664), .ZN(n5668)
         );
  OAI21_X1 U6799 ( .B1(n5669), .B2(n6169), .A(n5668), .ZN(U2991) );
  NAND3_X1 U6800 ( .A1(n5680), .A2(n5671), .A3(n5670), .ZN(n5673) );
  OAI211_X1 U6801 ( .C1(n6185), .C2(n5781), .A(n5673), .B(n5672), .ZN(n5674)
         );
  AOI21_X1 U6802 ( .B1(n5691), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5674), 
        .ZN(n5675) );
  OAI21_X1 U6803 ( .B1(n5676), .B2(n6169), .A(n5675), .ZN(U2992) );
  INV_X1 U6804 ( .A(n5691), .ZN(n5684) );
  NAND2_X1 U6805 ( .A1(n5677), .A2(n6241), .ZN(n5682) );
  OAI21_X1 U6806 ( .B1(n6185), .B2(n5790), .A(n5678), .ZN(n5679) );
  AOI21_X1 U6807 ( .B1(n5680), .B2(n5683), .A(n5679), .ZN(n5681) );
  OAI211_X1 U6808 ( .C1(n5684), .C2(n5683), .A(n5682), .B(n5681), .ZN(U2993)
         );
  OAI21_X1 U6809 ( .B1(n5697), .B2(n5686), .A(n5685), .ZN(n5690) );
  OAI21_X1 U6810 ( .B1(n6185), .B2(n5688), .A(n5687), .ZN(n5689) );
  AOI21_X1 U6811 ( .B1(n5691), .B2(n5690), .A(n5689), .ZN(n5692) );
  OAI21_X1 U6812 ( .B1(n5693), .B2(n6169), .A(n5692), .ZN(U2994) );
  INV_X1 U6813 ( .A(n5694), .ZN(n5695) );
  AOI21_X1 U6814 ( .B1(n6238), .B2(n5803), .A(n5695), .ZN(n5696) );
  OAI21_X1 U6815 ( .B1(n5697), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5696), 
        .ZN(n5698) );
  AOI21_X1 U6816 ( .B1(n5699), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5698), 
        .ZN(n5700) );
  OAI21_X1 U6817 ( .B1(n5701), .B2(n6169), .A(n5700), .ZN(U2995) );
  INV_X1 U6818 ( .A(n5702), .ZN(n5707) );
  NOR4_X1 U6819 ( .A1(n5882), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n5703), 
        .A4(n5707), .ZN(n5704) );
  AOI211_X1 U6820 ( .C1(n6238), .C2(n5809), .A(n5705), .B(n5704), .ZN(n5709)
         );
  INV_X1 U6821 ( .A(n5706), .ZN(n5718) );
  NOR3_X1 U6822 ( .A1(n5882), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5707), 
        .ZN(n5717) );
  OAI21_X1 U6823 ( .B1(n5718), .B2(n5717), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5708) );
  OAI211_X1 U6824 ( .C1(n5710), .C2(n6169), .A(n5709), .B(n5708), .ZN(U2996)
         );
  NAND2_X1 U6825 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  NAND2_X1 U6826 ( .A1(n5714), .A2(n5713), .ZN(n5842) );
  OAI21_X1 U6827 ( .B1(n6185), .B2(n5842), .A(n5715), .ZN(n5716) );
  AOI211_X1 U6828 ( .C1(n5718), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5717), .B(n5716), .ZN(n5719) );
  OAI21_X1 U6829 ( .B1(n5720), .B2(n6169), .A(n5719), .ZN(U2997) );
  NOR2_X1 U6830 ( .A1(n6211), .A2(n5721), .ZN(n5722) );
  OR2_X1 U6831 ( .A1(n5723), .A2(n5722), .ZN(n5877) );
  INV_X1 U6832 ( .A(n5877), .ZN(n5724) );
  OAI21_X1 U6833 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5740) );
  INV_X1 U6834 ( .A(n5727), .ZN(n5728) );
  NAND3_X1 U6835 ( .A1(n5736), .A2(n5729), .A3(n5728), .ZN(n5731) );
  OAI211_X1 U6836 ( .C1(n5830), .C2(n6185), .A(n5731), .B(n5730), .ZN(n5732)
         );
  AOI21_X1 U6837 ( .B1(n5740), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5732), 
        .ZN(n5733) );
  OAI21_X1 U6838 ( .B1(n5734), .B2(n6169), .A(n5733), .ZN(U2998) );
  NAND2_X1 U6839 ( .A1(n5736), .A2(n5735), .ZN(n5738) );
  OAI211_X1 U6840 ( .C1(n5841), .C2(n6185), .A(n5738), .B(n5737), .ZN(n5739)
         );
  AOI21_X1 U6841 ( .B1(n5740), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5739), 
        .ZN(n5741) );
  OAI21_X1 U6842 ( .B1(n5742), .B2(n6169), .A(n5741), .ZN(U2999) );
  NOR2_X1 U6843 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  XNOR2_X1 U6844 ( .A(n5745), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5869)
         );
  NOR2_X1 U6845 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5882), .ZN(n5746)
         );
  OAI21_X1 U6846 ( .B1(n5877), .B2(n5746), .A(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n5751) );
  INV_X1 U6847 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U6848 ( .A1(n6183), .A2(n6563), .ZN(n5749) );
  NOR3_X1 U6849 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5882), .A3(n5747), 
        .ZN(n5748) );
  NOR2_X1 U6850 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  OAI211_X1 U6851 ( .C1(n6185), .C2(n5940), .A(n5751), .B(n5750), .ZN(n5752)
         );
  AOI21_X1 U6852 ( .B1(n5869), .B2(n6241), .A(n5752), .ZN(n5753) );
  INV_X1 U6853 ( .A(n5753), .ZN(U3000) );
  INV_X1 U6854 ( .A(n5757), .ZN(n5754) );
  AND2_X1 U6855 ( .A1(n6202), .A2(n5754), .ZN(n5755) );
  OR2_X1 U6856 ( .A1(n6166), .A2(n5755), .ZN(n5883) );
  OAI21_X1 U6857 ( .B1(n6185), .B2(n5958), .A(n5756), .ZN(n5760) );
  NAND2_X1 U6858 ( .A1(n5757), .A2(n6165), .ZN(n5884) );
  AOI221_X1 U6859 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5890), .C2(n5758), .A(n5884), 
        .ZN(n5759) );
  AOI211_X1 U6860 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5883), .A(n5760), .B(n5759), .ZN(n5761) );
  OAI21_X1 U6861 ( .B1(n5762), .B2(n6169), .A(n5761), .ZN(U3002) );
  OAI21_X1 U6862 ( .B1(n5772), .B2(n4400), .A(n5763), .ZN(n5764) );
  MUX2_X1 U6863 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5764), .S(n6249), 
        .Z(U3464) );
  XNOR2_X1 U6864 ( .A(n5765), .B(n6254), .ZN(n5766) );
  OAI22_X1 U6865 ( .A1(n5766), .A2(n6390), .B1(n4415), .B2(n5772), .ZN(n5767)
         );
  MUX2_X1 U6866 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5767), .S(n6249), 
        .Z(U3463) );
  NAND2_X1 U6867 ( .A1(n5768), .A2(n6386), .ZN(n6256) );
  NOR2_X1 U6868 ( .A1(n5769), .A2(n6385), .ZN(n6306) );
  NOR2_X1 U6869 ( .A1(n6256), .A2(n6306), .ZN(n5770) );
  MUX2_X1 U6870 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5774), .S(n6249), 
        .Z(U3462) );
  OAI22_X1 U6871 ( .A1(n5778), .A2(n5777), .B1(n5776), .B2(n5775), .ZN(n5779)
         );
  MUX2_X1 U6872 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5779), .S(n5914), 
        .Z(U3456) );
  AND2_X1 U6873 ( .A1(n6105), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6874 ( .A1(n6047), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6051), .ZN(n5786) );
  NOR2_X1 U6875 ( .A1(n6628), .A2(n5780), .ZN(n5788) );
  AOI21_X1 U6876 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5788), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5783) );
  OAI22_X1 U6877 ( .A1(n5783), .A2(n5782), .B1(n5781), .B2(n6014), .ZN(n5784)
         );
  AOI21_X1 U6878 ( .B1(n5849), .B2(n5989), .A(n5784), .ZN(n5785) );
  OAI211_X1 U6879 ( .C1(n5787), .C2(n6024), .A(n5786), .B(n5785), .ZN(U2801)
         );
  AOI22_X1 U6880 ( .A1(n6047), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6051), .ZN(n5797) );
  INV_X1 U6881 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6785) );
  AOI22_X1 U6882 ( .A1(n5789), .A2(n6054), .B1(n5788), .B2(n6785), .ZN(n5796)
         );
  OAI22_X1 U6883 ( .A1(n5852), .A2(n6038), .B1(n6014), .B2(n5790), .ZN(n5791)
         );
  INV_X1 U6884 ( .A(n5791), .ZN(n5795) );
  INV_X1 U6885 ( .A(n5800), .ZN(n5792) );
  OAI21_X1 U6886 ( .B1(n5793), .B2(n5792), .A(REIP_REG_25__SCAN_IN), .ZN(n5794) );
  NAND4_X1 U6887 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(U2802)
         );
  AOI22_X1 U6888 ( .A1(n6047), .A2(EBX_REG_23__SCAN_IN), .B1(n5798), .B2(n6054), .ZN(n5805) );
  AND2_X1 U6889 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5807), .ZN(n5808) );
  AOI21_X1 U6890 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5808), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5799) );
  OAI22_X1 U6891 ( .A1(n5801), .A2(n6038), .B1(n5800), .B2(n5799), .ZN(n5802)
         );
  AOI21_X1 U6892 ( .B1(n5803), .B2(n6050), .A(n5802), .ZN(n5804) );
  OAI211_X1 U6893 ( .C1(n5806), .C2(n6036), .A(n5805), .B(n5804), .ZN(U2804)
         );
  NAND2_X1 U6894 ( .A1(n5807), .A2(n6751), .ZN(n5819) );
  AOI22_X1 U6895 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6051), .B1(n5808), 
        .B2(n6750), .ZN(n5812) );
  AOI22_X1 U6896 ( .A1(n6054), .A2(n5810), .B1(n5809), .B2(n6050), .ZN(n5811)
         );
  OAI211_X1 U6897 ( .C1(n5949), .C2(n5813), .A(n5812), .B(n5811), .ZN(n5814)
         );
  AOI21_X1 U6898 ( .B1(n5856), .B2(n5989), .A(n5814), .ZN(n5815) );
  OAI221_X1 U6899 ( .B1(n6750), .B2(n5816), .C1(n6750), .C2(n5819), .A(n5815), 
        .ZN(U2805) );
  AOI22_X1 U6900 ( .A1(n6047), .A2(EBX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6051), .ZN(n5822) );
  INV_X1 U6901 ( .A(n5816), .ZN(n5826) );
  AOI22_X1 U6902 ( .A1(n5817), .A2(n6054), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5826), .ZN(n5821) );
  OAI22_X1 U6903 ( .A1(n5859), .A2(n6038), .B1(n6014), .B2(n5842), .ZN(n5818)
         );
  INV_X1 U6904 ( .A(n5818), .ZN(n5820) );
  NAND4_X1 U6905 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(U2806)
         );
  OAI22_X1 U6906 ( .A1(n5599), .A2(n6036), .B1(n6024), .B2(n5823), .ZN(n5824)
         );
  AOI21_X1 U6907 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6047), .A(n5824), .ZN(n5829)
         );
  NAND2_X1 U6908 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5825) );
  INV_X1 U6909 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6705) );
  OAI21_X1 U6910 ( .B1(n5825), .B2(n5838), .A(n6705), .ZN(n5827) );
  AOI22_X1 U6911 ( .A1(n5863), .A2(n5989), .B1(n5827), .B2(n5826), .ZN(n5828)
         );
  OAI211_X1 U6912 ( .C1(n5830), .C2(n6014), .A(n5829), .B(n5828), .ZN(U2807)
         );
  INV_X1 U6913 ( .A(n5831), .ZN(n5866) );
  NOR3_X1 U6914 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6563), .A3(n5838), .ZN(n5837) );
  INV_X1 U6915 ( .A(n5832), .ZN(n5835) );
  AOI21_X1 U6916 ( .B1(n6051), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6032), 
        .ZN(n5834) );
  NAND2_X1 U6917 ( .A1(n6047), .A2(EBX_REG_19__SCAN_IN), .ZN(n5833) );
  OAI211_X1 U6918 ( .C1(n5835), .C2(n6024), .A(n5834), .B(n5833), .ZN(n5836)
         );
  AOI211_X1 U6919 ( .C1(n5866), .C2(n5989), .A(n5837), .B(n5836), .ZN(n5840)
         );
  NOR2_X1 U6920 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5838), .ZN(n5939) );
  OAI21_X1 U6921 ( .B1(n5939), .B2(n5942), .A(REIP_REG_19__SCAN_IN), .ZN(n5839) );
  OAI211_X1 U6922 ( .C1(n5841), .C2(n6014), .A(n5840), .B(n5839), .ZN(U2808)
         );
  INV_X1 U6923 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5847) );
  OAI22_X1 U6924 ( .A1(n5859), .A2(n5844), .B1(n5843), .B2(n5842), .ZN(n5845)
         );
  INV_X1 U6925 ( .A(n5845), .ZN(n5846) );
  OAI21_X1 U6926 ( .B1(n6066), .B2(n5847), .A(n5846), .ZN(U2838) );
  AOI22_X1 U6927 ( .A1(n5849), .A2(n6071), .B1(n6070), .B2(DATAI_26_), .ZN(
        n5851) );
  AOI22_X1 U6928 ( .A1(n6074), .A2(DATAI_10_), .B1(n6073), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6929 ( .A1(n5851), .A2(n5850), .ZN(U2865) );
  INV_X1 U6930 ( .A(n5852), .ZN(n5853) );
  AOI22_X1 U6931 ( .A1(n5853), .A2(n6071), .B1(n6070), .B2(DATAI_25_), .ZN(
        n5855) );
  AOI22_X1 U6932 ( .A1(n6074), .A2(DATAI_9_), .B1(n6073), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6933 ( .A1(n5855), .A2(n5854), .ZN(U2866) );
  AOI22_X1 U6934 ( .A1(n5856), .A2(n6071), .B1(n6070), .B2(DATAI_22_), .ZN(
        n5858) );
  AOI22_X1 U6935 ( .A1(n6074), .A2(DATAI_6_), .B1(n6073), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6936 ( .A1(n5858), .A2(n5857), .ZN(U2869) );
  INV_X1 U6937 ( .A(n5859), .ZN(n5860) );
  AOI22_X1 U6938 ( .A1(n5860), .A2(n6071), .B1(n6070), .B2(DATAI_21_), .ZN(
        n5862) );
  AOI22_X1 U6939 ( .A1(n6074), .A2(DATAI_5_), .B1(n6073), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U6940 ( .A1(n5862), .A2(n5861), .ZN(U2870) );
  AOI22_X1 U6941 ( .A1(n5863), .A2(n6071), .B1(n6070), .B2(DATAI_20_), .ZN(
        n5865) );
  AOI22_X1 U6942 ( .A1(n6074), .A2(DATAI_4_), .B1(n6073), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U6943 ( .A1(n5865), .A2(n5864), .ZN(U2871) );
  AOI22_X1 U6944 ( .A1(n5866), .A2(n6071), .B1(n6070), .B2(DATAI_19_), .ZN(
        n5868) );
  AOI22_X1 U6945 ( .A1(n6074), .A2(DATAI_3_), .B1(n6073), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6946 ( .A1(n5868), .A2(n5867), .ZN(U2872) );
  AOI22_X1 U6947 ( .A1(n6221), .A2(REIP_REG_18__SCAN_IN), .B1(n6153), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5871) );
  AOI22_X1 U6948 ( .A1(n5869), .A2(n6158), .B1(n6149), .B2(n6067), .ZN(n5870)
         );
  OAI211_X1 U6949 ( .C1(n6162), .C2(n5948), .A(n5871), .B(n5870), .ZN(U2968)
         );
  AOI22_X1 U6950 ( .A1(n6221), .A2(REIP_REG_13__SCAN_IN), .B1(n6153), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U6951 ( .A(n5872), .B(n5873), .ZN(n5905) );
  INV_X1 U6952 ( .A(n5976), .ZN(n5874) );
  AOI22_X1 U6953 ( .A1(n5905), .A2(n6158), .B1(n6149), .B2(n5874), .ZN(n5875)
         );
  OAI211_X1 U6954 ( .C1(n6162), .C2(n5975), .A(n5876), .B(n5875), .ZN(U2973)
         );
  AOI22_X1 U6955 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5877), .B1(n6221), .B2(REIP_REG_17__SCAN_IN), .ZN(n5881) );
  AOI22_X1 U6956 ( .A1(n5879), .A2(n6241), .B1(n6238), .B2(n5878), .ZN(n5880)
         );
  OAI211_X1 U6957 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5882), .A(n5881), .B(n5880), .ZN(U3001) );
  INV_X1 U6958 ( .A(n5883), .ZN(n5891) );
  INV_X1 U6959 ( .A(n5884), .ZN(n5885) );
  AOI22_X1 U6960 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6221), .B1(n5885), .B2(
        n5890), .ZN(n5889) );
  AOI22_X1 U6961 ( .A1(n5887), .A2(n6241), .B1(n6238), .B2(n5886), .ZN(n5888)
         );
  OAI211_X1 U6962 ( .C1(n5891), .C2(n5890), .A(n5889), .B(n5888), .ZN(U3003)
         );
  NAND2_X1 U6963 ( .A1(n5343), .A2(n6165), .ZN(n5901) );
  NAND3_X1 U6964 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n5908), .ZN(n5903) );
  AOI22_X1 U6965 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .B1(n5892), .B2(n6211), .ZN(n5893)
         );
  AOI211_X1 U6966 ( .C1(n5894), .C2(n5902), .A(n6166), .B(n5893), .ZN(n5909)
         );
  OAI21_X1 U6967 ( .B1(n5895), .B2(n5903), .A(n5909), .ZN(n5898) );
  OAI22_X1 U6968 ( .A1(n5896), .A2(n6169), .B1(n6185), .B2(n5968), .ZN(n5897)
         );
  AOI21_X1 U6969 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5898), .A(n5897), 
        .ZN(n5900) );
  NAND2_X1 U6970 ( .A1(n6221), .A2(REIP_REG_14__SCAN_IN), .ZN(n5899) );
  OAI211_X1 U6971 ( .C1(n5902), .C2(n5901), .A(n5900), .B(n5899), .ZN(U3004)
         );
  INV_X1 U6972 ( .A(n5903), .ZN(n5904) );
  AOI22_X1 U6973 ( .A1(n6221), .A2(REIP_REG_13__SCAN_IN), .B1(n5904), .B2(
        n6165), .ZN(n5907) );
  AOI22_X1 U6974 ( .A1(n5905), .A2(n6241), .B1(n6238), .B2(n5979), .ZN(n5906)
         );
  OAI211_X1 U6975 ( .C1(n5909), .C2(n5908), .A(n5907), .B(n5906), .ZN(U3005)
         );
  OR3_X1 U6976 ( .A1(n5911), .A2(STATE2_REG_3__SCAN_IN), .A3(n5910), .ZN(n5912) );
  OAI21_X1 U6977 ( .B1(n5914), .B2(n5913), .A(n5912), .ZN(U3455) );
  INV_X1 U6978 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6513) );
  AOI21_X1 U6979 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6513), .A(n6523), .ZN(n5921) );
  INV_X1 U6980 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5915) );
  INV_X1 U6981 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6519) );
  NOR2_X2 U6982 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6519), .ZN(n6812) );
  AOI21_X1 U6983 ( .B1(n5921), .B2(n5915), .A(n6812), .ZN(U2789) );
  NAND2_X1 U6984 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6606), .ZN(n5919) );
  OAI21_X1 U6985 ( .B1(n5916), .B2(n6475), .A(n3999), .ZN(n5917) );
  OAI21_X1 U6986 ( .B1(n6480), .B2(n3009), .A(n5917), .ZN(n5925) );
  OAI21_X1 U6987 ( .B1(n5925), .B2(n6499), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5918) );
  OAI21_X1 U6988 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5919), .A(n5918), .ZN(
        U2790) );
  INV_X1 U6989 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6678) );
  NOR2_X1 U6990 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5922) );
  NOR2_X1 U6991 ( .A1(n6812), .A2(n5922), .ZN(n5920) );
  AOI22_X1 U6992 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6812), .B1(n6678), .B2(
        n5920), .ZN(U2791) );
  OAI21_X1 U6993 ( .B1(BS16_N), .B2(n5922), .A(n6585), .ZN(n6583) );
  OAI21_X1 U6994 ( .B1(n6585), .B2(n5923), .A(n6583), .ZN(U2792) );
  AOI21_X1 U6995 ( .B1(n5924), .B2(n6518), .A(READY_N), .ZN(n6604) );
  NOR2_X1 U6996 ( .A1(n5925), .A2(n6604), .ZN(n6471) );
  NOR2_X1 U6997 ( .A1(n6471), .A2(n6499), .ZN(n6600) );
  OAI21_X1 U6998 ( .B1(n6600), .B2(n6741), .A(n6134), .ZN(U2793) );
  NOR4_X1 U6999 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5929) );
  NOR4_X1 U7000 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5928) );
  NOR4_X1 U7001 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5927) );
  NOR4_X1 U7002 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5926) );
  NAND4_X1 U7003 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(n5935)
         );
  NOR4_X1 U7004 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5933) );
  AOI211_X1 U7005 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5932) );
  NOR4_X1 U7006 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5931) );
  NOR4_X1 U7007 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5930) );
  NAND4_X1 U7008 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n5934)
         );
  NOR2_X1 U7009 ( .A1(n5935), .A2(n5934), .ZN(n6597) );
  INV_X1 U7010 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6710) );
  NOR3_X1 U7011 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5937) );
  OAI21_X1 U7012 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5937), .A(n6597), .ZN(n5936)
         );
  OAI21_X1 U7013 ( .B1(n6597), .B2(n6710), .A(n5936), .ZN(U2794) );
  INV_X1 U7014 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6584) );
  AOI21_X1 U7015 ( .B1(n6590), .B2(n6584), .A(n5937), .ZN(n5938) );
  INV_X1 U7016 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6755) );
  INV_X1 U7017 ( .A(n6597), .ZN(n6592) );
  AOI22_X1 U7018 ( .A1(n6597), .A2(n5938), .B1(n6755), .B2(n6592), .ZN(U2795)
         );
  AOI211_X1 U7019 ( .C1(n6051), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5939), 
        .B(n6032), .ZN(n5945) );
  NOR2_X1 U7020 ( .A1(n5940), .A2(n6014), .ZN(n5941) );
  AOI21_X1 U7021 ( .B1(n6047), .B2(EBX_REG_18__SCAN_IN), .A(n5941), .ZN(n5944)
         );
  NAND2_X1 U7022 ( .A1(n5942), .A2(REIP_REG_18__SCAN_IN), .ZN(n5943) );
  NAND3_X1 U7023 ( .A1(n5945), .A2(n5944), .A3(n5943), .ZN(n5946) );
  AOI21_X1 U7024 ( .B1(n6067), .B2(n5989), .A(n5946), .ZN(n5947) );
  OAI21_X1 U7025 ( .B1(n5948), .B2(n6024), .A(n5947), .ZN(U2809) );
  OAI22_X1 U7026 ( .A1(n5950), .A2(REIP_REG_16__SCAN_IN), .B1(n5949), .B2(
        n5509), .ZN(n5951) );
  INV_X1 U7027 ( .A(n5951), .ZN(n5952) );
  OAI221_X1 U7028 ( .B1(n6559), .B2(n5960), .C1(n6559), .C2(n5953), .A(n5952), 
        .ZN(n5954) );
  AOI211_X1 U7029 ( .C1(n6051), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6032), 
        .B(n5954), .ZN(n5957) );
  AOI22_X1 U7030 ( .A1(n6072), .A2(n5989), .B1(n6054), .B2(n5955), .ZN(n5956)
         );
  OAI211_X1 U7031 ( .C1(n6014), .C2(n5958), .A(n5957), .B(n5956), .ZN(U2811)
         );
  OAI21_X1 U7032 ( .B1(n6036), .B2(n5959), .A(n6058), .ZN(n5963) );
  AOI21_X1 U7033 ( .B1(n6555), .B2(n5961), .A(n5960), .ZN(n5962) );
  AOI211_X1 U7034 ( .C1(EBX_REG_14__SCAN_IN), .C2(n6047), .A(n5963), .B(n5962), 
        .ZN(n5967) );
  AOI22_X1 U7035 ( .A1(n5965), .A2(n5989), .B1(n6054), .B2(n5964), .ZN(n5966)
         );
  OAI211_X1 U7036 ( .C1(n6014), .C2(n5968), .A(n5967), .B(n5966), .ZN(U2813)
         );
  INV_X1 U7037 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5982) );
  INV_X1 U7038 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U7039 ( .A1(n6553), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7040 ( .A1(n6047), .A2(EBX_REG_13__SCAN_IN), .ZN(n5971) );
  OAI211_X1 U7041 ( .C1(n6046), .C2(n5972), .A(n5971), .B(n6058), .ZN(n5973)
         );
  INV_X1 U7042 ( .A(n5973), .ZN(n5981) );
  AOI21_X1 U7043 ( .B1(n5983), .B2(n5974), .A(n6553), .ZN(n5978) );
  OAI22_X1 U7044 ( .A1(n5976), .A2(n6038), .B1(n5975), .B2(n6024), .ZN(n5977)
         );
  AOI211_X1 U7045 ( .C1(n5979), .C2(n6050), .A(n5978), .B(n5977), .ZN(n5980)
         );
  OAI211_X1 U7046 ( .C1(n5982), .C2(n6036), .A(n5981), .B(n5980), .ZN(U2814)
         );
  INV_X1 U7047 ( .A(n5983), .ZN(n5986) );
  OAI21_X1 U7048 ( .B1(n6046), .B2(n5984), .A(n6549), .ZN(n5985) );
  AOI22_X1 U7049 ( .A1(n5986), .A2(n5985), .B1(EBX_REG_11__SCAN_IN), .B2(n6047), .ZN(n5992) );
  AOI21_X1 U7050 ( .B1(n5988), .B2(n5987), .A(n5250), .ZN(n6163) );
  AOI22_X1 U7051 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6051), .B1(n6050), 
        .B2(n6163), .ZN(n5991) );
  AOI22_X1 U7052 ( .A1(n6131), .A2(n5989), .B1(n6054), .B2(n6129), .ZN(n5990)
         );
  NAND4_X1 U7053 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n6058), .ZN(U2816)
         );
  AOI22_X1 U7054 ( .A1(n6010), .A2(REIP_REG_9__SCAN_IN), .B1(
        EBX_REG_9__SCAN_IN), .B2(n6047), .ZN(n6003) );
  OAI21_X1 U7055 ( .B1(n6036), .B2(n5993), .A(n6058), .ZN(n5994) );
  AOI211_X1 U7056 ( .C1(n5996), .C2(n6050), .A(n5995), .B(n5994), .ZN(n6002)
         );
  INV_X1 U7057 ( .A(n5997), .ZN(n5998) );
  OAI22_X1 U7058 ( .A1(n5999), .A2(n6038), .B1(n6024), .B2(n5998), .ZN(n6000)
         );
  INV_X1 U7059 ( .A(n6000), .ZN(n6001) );
  NAND3_X1 U7060 ( .A1(n6003), .A2(n6002), .A3(n6001), .ZN(U2818) );
  AOI21_X1 U7061 ( .B1(n6051), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6032), 
        .ZN(n6005) );
  NAND2_X1 U7062 ( .A1(n6047), .A2(EBX_REG_8__SCAN_IN), .ZN(n6004) );
  OAI211_X1 U7063 ( .C1(n6006), .C2(n6038), .A(n6005), .B(n6004), .ZN(n6007)
         );
  AOI21_X1 U7064 ( .B1(n6008), .B2(n6054), .A(n6007), .ZN(n6013) );
  AND2_X1 U7065 ( .A1(n6023), .A2(n6009), .ZN(n6011) );
  OAI21_X1 U7066 ( .B1(n6011), .B2(REIP_REG_8__SCAN_IN), .A(n6010), .ZN(n6012)
         );
  OAI211_X1 U7067 ( .C1(n6184), .C2(n6014), .A(n6013), .B(n6012), .ZN(U2819)
         );
  INV_X1 U7068 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6031) );
  INV_X1 U7069 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7070 ( .A1(n6541), .A2(n6016), .ZN(n6018) );
  NAND2_X1 U7071 ( .A1(n6047), .A2(EBX_REG_7__SCAN_IN), .ZN(n6017) );
  OAI211_X1 U7072 ( .C1(n6046), .C2(n6018), .A(n6017), .B(n6058), .ZN(n6019)
         );
  INV_X1 U7073 ( .A(n6019), .ZN(n6030) );
  OR2_X1 U7074 ( .A1(n6046), .A2(n6022), .ZN(n6021) );
  AND2_X1 U7075 ( .A1(n6021), .A2(n6020), .ZN(n6044) );
  INV_X1 U7076 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6539) );
  NAND3_X1 U7077 ( .A1(n6023), .A2(n6022), .A3(n6539), .ZN(n6035) );
  AOI21_X1 U7078 ( .B1(n6044), .B2(n6035), .A(n6541), .ZN(n6028) );
  OAI22_X1 U7079 ( .A1(n6026), .A2(n6038), .B1(n6025), .B2(n6024), .ZN(n6027)
         );
  AOI211_X1 U7080 ( .C1(n6194), .C2(n6050), .A(n6028), .B(n6027), .ZN(n6029)
         );
  OAI211_X1 U7081 ( .C1(n6031), .C2(n6036), .A(n6030), .B(n6029), .ZN(U2820)
         );
  INV_X1 U7082 ( .A(n6142), .ZN(n6033) );
  AOI21_X1 U7083 ( .B1(n6054), .B2(n6033), .A(n6032), .ZN(n6034) );
  OAI211_X1 U7084 ( .C1(n6037), .C2(n6036), .A(n6035), .B(n6034), .ZN(n6041)
         );
  NOR2_X1 U7085 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  AOI211_X1 U7086 ( .C1(EBX_REG_6__SCAN_IN), .C2(n6047), .A(n6041), .B(n6040), 
        .ZN(n6043) );
  NAND2_X1 U7087 ( .A1(n6050), .A2(n6203), .ZN(n6042) );
  OAI211_X1 U7088 ( .C1(n6044), .C2(n6539), .A(n6043), .B(n6042), .ZN(U2821)
         );
  INV_X1 U7089 ( .A(n6044), .ZN(n6049) );
  OAI21_X1 U7090 ( .B1(n6046), .B2(n6045), .A(n6537), .ZN(n6048) );
  AOI22_X1 U7091 ( .A1(n6049), .A2(n6048), .B1(EBX_REG_5__SCAN_IN), .B2(n6047), 
        .ZN(n6061) );
  AOI22_X1 U7092 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6051), .B1(n6050), 
        .B2(n6215), .ZN(n6060) );
  INV_X1 U7093 ( .A(n6052), .ZN(n6056) );
  INV_X1 U7094 ( .A(n6053), .ZN(n6055) );
  AOI22_X1 U7095 ( .A1(n6057), .A2(n6056), .B1(n6055), .B2(n6054), .ZN(n6059)
         );
  NAND4_X1 U7096 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(U2822)
         );
  AOI22_X1 U7097 ( .A1(n6131), .A2(n6063), .B1(n6062), .B2(n6163), .ZN(n6064)
         );
  OAI21_X1 U7098 ( .B1(n6066), .B2(n6065), .A(n6064), .ZN(U2848) );
  AOI22_X1 U7099 ( .A1(n6067), .A2(n6071), .B1(n6070), .B2(DATAI_18_), .ZN(
        n6069) );
  AOI22_X1 U7100 ( .A1(n6074), .A2(DATAI_2_), .B1(n6073), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7101 ( .A1(n6069), .A2(n6068), .ZN(U2873) );
  AOI22_X1 U7102 ( .A1(n6072), .A2(n6071), .B1(n6070), .B2(DATAI_16_), .ZN(
        n6076) );
  AOI22_X1 U7103 ( .A1(n6074), .A2(DATAI_0_), .B1(n6073), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7104 ( .A1(n6076), .A2(n6075), .ZN(U2875) );
  AOI22_X1 U7105 ( .A1(n6603), .A2(LWORD_REG_15__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U7106 ( .B1(n6078), .B2(n6108), .A(n6077), .ZN(U2908) );
  INV_X1 U7107 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6080) );
  AOI22_X1 U7108 ( .A1(n6603), .A2(LWORD_REG_14__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U7109 ( .B1(n6080), .B2(n6108), .A(n6079), .ZN(U2909) );
  INV_X1 U7110 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6082) );
  AOI22_X1 U7111 ( .A1(n6603), .A2(LWORD_REG_13__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U7112 ( .B1(n6082), .B2(n6108), .A(n6081), .ZN(U2910) );
  INV_X1 U7113 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6084) );
  AOI22_X1 U7114 ( .A1(n6603), .A2(LWORD_REG_12__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6083) );
  OAI21_X1 U7115 ( .B1(n6084), .B2(n6108), .A(n6083), .ZN(U2911) );
  INV_X1 U7116 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6086) );
  AOI22_X1 U7117 ( .A1(n6603), .A2(LWORD_REG_11__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6085) );
  OAI21_X1 U7118 ( .B1(n6086), .B2(n6108), .A(n6085), .ZN(U2912) );
  INV_X1 U7119 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6088) );
  AOI22_X1 U7120 ( .A1(n6603), .A2(LWORD_REG_10__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7121 ( .B1(n6088), .B2(n6108), .A(n6087), .ZN(U2913) );
  INV_X1 U7122 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6090) );
  AOI22_X1 U7123 ( .A1(n6603), .A2(LWORD_REG_9__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7124 ( .B1(n6090), .B2(n6108), .A(n6089), .ZN(U2914) );
  INV_X1 U7125 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6092) );
  AOI22_X1 U7126 ( .A1(n6603), .A2(LWORD_REG_8__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7127 ( .B1(n6092), .B2(n6108), .A(n6091), .ZN(U2915) );
  AOI22_X1 U7128 ( .A1(n6106), .A2(LWORD_REG_7__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7129 ( .B1(n4954), .B2(n6108), .A(n6093), .ZN(U2916) );
  INV_X1 U7130 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6095) );
  AOI22_X1 U7131 ( .A1(n6106), .A2(LWORD_REG_6__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6094) );
  OAI21_X1 U7132 ( .B1(n6095), .B2(n6108), .A(n6094), .ZN(U2917) );
  AOI22_X1 U7133 ( .A1(n6106), .A2(LWORD_REG_5__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7134 ( .B1(n3466), .B2(n6108), .A(n6096), .ZN(U2918) );
  AOI22_X1 U7135 ( .A1(n6106), .A2(LWORD_REG_4__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7136 ( .B1(n6098), .B2(n6108), .A(n6097), .ZN(U2919) );
  AOI22_X1 U7137 ( .A1(n6106), .A2(LWORD_REG_3__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6099) );
  OAI21_X1 U7138 ( .B1(n6100), .B2(n6108), .A(n6099), .ZN(U2920) );
  AOI22_X1 U7139 ( .A1(n6106), .A2(LWORD_REG_2__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7140 ( .B1(n6102), .B2(n6108), .A(n6101), .ZN(U2921) );
  AOI22_X1 U7141 ( .A1(n6106), .A2(LWORD_REG_1__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7142 ( .B1(n6104), .B2(n6108), .A(n6103), .ZN(U2922) );
  AOI22_X1 U7143 ( .A1(n6106), .A2(LWORD_REG_0__SCAN_IN), .B1(n6105), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7144 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(U2923) );
  AOI22_X1 U7145 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6122), .B1(n6121), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7146 ( .B1(n6124), .B2(n6782), .A(n6111), .ZN(U2945) );
  AOI22_X1 U7147 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6122), .B1(n6121), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7148 ( .B1(n6124), .B2(n6648), .A(n6112), .ZN(U2946) );
  INV_X1 U7149 ( .A(DATAI_8_), .ZN(n6720) );
  AOI22_X1 U7150 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6118), .B1(n6121), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7151 ( .B1(n6124), .B2(n6720), .A(n6113), .ZN(U2947) );
  INV_X1 U7152 ( .A(DATAI_9_), .ZN(n6672) );
  AOI22_X1 U7153 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6118), .B1(n6121), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7154 ( .B1(n6124), .B2(n6672), .A(n6114), .ZN(U2948) );
  INV_X1 U7155 ( .A(DATAI_10_), .ZN(n6735) );
  AOI22_X1 U7156 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6118), .B1(n6121), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7157 ( .B1(n6124), .B2(n6735), .A(n6115), .ZN(U2949) );
  INV_X1 U7158 ( .A(DATAI_11_), .ZN(n6117) );
  AOI22_X1 U7159 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6118), .B1(n6121), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7160 ( .B1(n6124), .B2(n6117), .A(n6116), .ZN(U2950) );
  INV_X1 U7161 ( .A(DATAI_12_), .ZN(n6644) );
  AOI22_X1 U7162 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6118), .B1(n6121), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7163 ( .B1(n6124), .B2(n6644), .A(n6119), .ZN(U2951) );
  INV_X1 U7164 ( .A(DATAI_13_), .ZN(n6683) );
  AOI22_X1 U7165 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6122), .B1(n6121), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7166 ( .B1(n6124), .B2(n6683), .A(n6120), .ZN(U2952) );
  INV_X1 U7167 ( .A(DATAI_14_), .ZN(n6774) );
  AOI22_X1 U7168 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6122), .B1(n6121), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7169 ( .B1(n6124), .B2(n6774), .A(n6123), .ZN(U2953) );
  NAND2_X1 U7170 ( .A1(n6125), .A2(n6126), .ZN(n6128) );
  XNOR2_X1 U7171 ( .A(n2985), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6127)
         );
  XNOR2_X1 U7172 ( .A(n6128), .B(n6127), .ZN(n6170) );
  AOI22_X1 U7173 ( .A1(n6221), .A2(REIP_REG_11__SCAN_IN), .B1(n6153), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6133) );
  AOI22_X1 U7174 ( .A1(n6131), .A2(n6149), .B1(n6130), .B2(n6129), .ZN(n6132)
         );
  OAI211_X1 U7175 ( .C1(n6170), .C2(n6134), .A(n6133), .B(n6132), .ZN(U2975)
         );
  AOI22_X1 U7176 ( .A1(n6221), .A2(REIP_REG_6__SCAN_IN), .B1(n6153), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6141) );
  OAI21_X1 U7177 ( .B1(n6135), .B2(n6137), .A(n6136), .ZN(n6138) );
  INV_X1 U7178 ( .A(n6138), .ZN(n6206) );
  AOI22_X1 U7179 ( .A1(n6206), .A2(n6158), .B1(n6149), .B2(n6139), .ZN(n6140)
         );
  OAI211_X1 U7180 ( .C1(n6162), .C2(n6142), .A(n6141), .B(n6140), .ZN(U2980)
         );
  AOI22_X1 U7181 ( .A1(n6221), .A2(REIP_REG_3__SCAN_IN), .B1(n6153), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6151) );
  OAI21_X1 U7182 ( .B1(n6143), .B2(n6145), .A(n6144), .ZN(n6146) );
  INV_X1 U7183 ( .A(n6146), .ZN(n6226) );
  INV_X1 U7184 ( .A(n6147), .ZN(n6148) );
  AOI22_X1 U7185 ( .A1(n6226), .A2(n6158), .B1(n6149), .B2(n6148), .ZN(n6150)
         );
  OAI211_X1 U7186 ( .C1(n6162), .C2(n6152), .A(n6151), .B(n6150), .ZN(U2983)
         );
  AOI22_X1 U7187 ( .A1(n6221), .A2(REIP_REG_2__SCAN_IN), .B1(n6153), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6160) );
  XOR2_X1 U7188 ( .A(n6154), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6156) );
  XNOR2_X1 U7189 ( .A(n6156), .B(n6155), .ZN(n6240) );
  AOI22_X1 U7190 ( .A1(n6240), .A2(n6158), .B1(n6157), .B2(n6149), .ZN(n6159)
         );
  OAI211_X1 U7191 ( .C1(n6162), .C2(n6161), .A(n6160), .B(n6159), .ZN(U2984)
         );
  AOI22_X1 U7192 ( .A1(n6238), .A2(n6163), .B1(n6221), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6168) );
  AOI22_X1 U7193 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6166), .B1(n6165), .B2(n6164), .ZN(n6167) );
  OAI211_X1 U7194 ( .C1(n6170), .C2(n6169), .A(n6168), .B(n6167), .ZN(U3007)
         );
  AOI21_X1 U7195 ( .B1(n6238), .B2(n6172), .A(n6171), .ZN(n6179) );
  AOI22_X1 U7196 ( .A1(n6174), .A2(n6241), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6173), .ZN(n6178) );
  OAI211_X1 U7197 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6176), .B(n6175), .ZN(n6177) );
  NAND3_X1 U7198 ( .A1(n6179), .A2(n6178), .A3(n6177), .ZN(U3008) );
  INV_X1 U7199 ( .A(n6180), .ZN(n6188) );
  AOI211_X1 U7200 ( .C1(n6182), .C2(n6190), .A(n6181), .B(n6200), .ZN(n6187)
         );
  INV_X1 U7201 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6543) );
  OAI22_X1 U7202 ( .A1(n6185), .A2(n6184), .B1(n6543), .B2(n6183), .ZN(n6186)
         );
  AOI211_X1 U7203 ( .C1(n6188), .C2(n6241), .A(n6187), .B(n6186), .ZN(n6189)
         );
  OAI21_X1 U7204 ( .B1(n6191), .B2(n6190), .A(n6189), .ZN(U3010) );
  INV_X1 U7205 ( .A(n6192), .ZN(n6193) );
  AOI21_X1 U7206 ( .B1(n6238), .B2(n6194), .A(n6193), .ZN(n6199) );
  INV_X1 U7207 ( .A(n6195), .ZN(n6197) );
  AOI22_X1 U7208 ( .A1(n6197), .A2(n6241), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6196), .ZN(n6198) );
  OAI211_X1 U7209 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6200), .A(n6199), 
        .B(n6198), .ZN(U3011) );
  OR2_X1 U7210 ( .A1(n6204), .A2(n6210), .ZN(n6201) );
  AOI21_X1 U7211 ( .B1(n6202), .B2(n6201), .A(n6239), .ZN(n6220) );
  AOI22_X1 U7212 ( .A1(n6238), .A2(n6203), .B1(n6221), .B2(REIP_REG_6__SCAN_IN), .ZN(n6208) );
  NOR3_X1 U7213 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6204), .A3(n6210), 
        .ZN(n6205) );
  AOI22_X1 U7214 ( .A1(n6206), .A2(n6241), .B1(n6205), .B2(n6223), .ZN(n6207)
         );
  OAI211_X1 U7215 ( .C1(n6220), .C2(n6209), .A(n6208), .B(n6207), .ZN(U3012)
         );
  OAI22_X1 U7216 ( .A1(n6242), .A2(n6212), .B1(n6211), .B2(n6210), .ZN(n6213)
         );
  NOR2_X1 U7217 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6213), .ZN(n6219)
         );
  INV_X1 U7218 ( .A(n6214), .ZN(n6216) );
  AOI22_X1 U7219 ( .A1(n6216), .A2(n6241), .B1(n6238), .B2(n6215), .ZN(n6218)
         );
  NAND2_X1 U7220 ( .A1(n6221), .A2(REIP_REG_5__SCAN_IN), .ZN(n6217) );
  OAI211_X1 U7221 ( .C1(n6220), .C2(n6219), .A(n6218), .B(n6217), .ZN(U3013)
         );
  AOI22_X1 U7222 ( .A1(n6238), .A2(n6222), .B1(n6221), .B2(REIP_REG_3__SCAN_IN), .ZN(n6229) );
  INV_X1 U7223 ( .A(n6223), .ZN(n6224) );
  NOR2_X1 U7224 ( .A1(n6225), .A2(n6224), .ZN(n6227) );
  AOI22_X1 U7225 ( .A1(n6227), .A2(n6230), .B1(n6226), .B2(n6241), .ZN(n6228)
         );
  OAI211_X1 U7226 ( .C1(n6231), .C2(n6230), .A(n6229), .B(n6228), .ZN(U3015)
         );
  INV_X1 U7227 ( .A(n6232), .ZN(n6237) );
  OAI21_X1 U7228 ( .B1(n6234), .B2(n6243), .A(n6233), .ZN(n6235) );
  AOI22_X1 U7229 ( .A1(n6238), .A2(n6237), .B1(n6236), .B2(n6235), .ZN(n6248)
         );
  AOI22_X1 U7230 ( .A1(n6241), .A2(n6240), .B1(n6239), .B2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7231 ( .A1(n6221), .A2(REIP_REG_2__SCAN_IN), .ZN(n6246) );
  INV_X1 U7232 ( .A(n6242), .ZN(n6244) );
  NAND3_X1 U7233 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6244), .A3(n6243), 
        .ZN(n6245) );
  NAND4_X1 U7234 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(U3016)
         );
  INV_X1 U7235 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6250) );
  NOR2_X1 U7236 ( .A1(n6250), .A2(n6249), .ZN(U3019) );
  INV_X1 U7237 ( .A(n6251), .ZN(n6380) );
  NAND2_X1 U7238 ( .A1(n6380), .A2(n6252), .ZN(n6285) );
  OAI22_X1 U7239 ( .A1(n6286), .A2(n6399), .B1(n6381), .B2(n6285), .ZN(n6253)
         );
  INV_X1 U7240 ( .A(n6253), .ZN(n6266) );
  NAND2_X1 U7241 ( .A1(n6254), .A2(n4585), .ZN(n6255) );
  OAI21_X1 U7242 ( .B1(n6256), .B2(n6255), .A(n6384), .ZN(n6264) );
  OR2_X1 U7243 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  AND2_X1 U7244 ( .A1(n6259), .A2(n6285), .ZN(n6263) );
  INV_X1 U7245 ( .A(n6263), .ZN(n6261) );
  AOI21_X1 U7246 ( .B1(n6262), .B2(n6390), .A(n6389), .ZN(n6260) );
  OAI22_X1 U7247 ( .A1(n6264), .A2(n6263), .B1(n6262), .B2(n6503), .ZN(n6288)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6289), .B1(n6396), 
        .B2(n6288), .ZN(n6265) );
  OAI211_X1 U7249 ( .C1(n6382), .C2(n6305), .A(n6266), .B(n6265), .ZN(U3044)
         );
  OAI22_X1 U7250 ( .A1(n6305), .A2(n6406), .B1(n6400), .B2(n6285), .ZN(n6267)
         );
  INV_X1 U7251 ( .A(n6267), .ZN(n6269) );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6289), .B1(n6403), 
        .B2(n6288), .ZN(n6268) );
  OAI211_X1 U7253 ( .C1(n6286), .C2(n6401), .A(n6269), .B(n6268), .ZN(U3045)
         );
  OAI22_X1 U7254 ( .A1(n6286), .A2(n6408), .B1(n6407), .B2(n6285), .ZN(n6270)
         );
  INV_X1 U7255 ( .A(n6270), .ZN(n6272) );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6289), .B1(n6410), 
        .B2(n6288), .ZN(n6271) );
  OAI211_X1 U7257 ( .C1(n6413), .C2(n6305), .A(n6272), .B(n6271), .ZN(U3046)
         );
  OAI22_X1 U7258 ( .A1(n6305), .A2(n6415), .B1(n6414), .B2(n6285), .ZN(n6273)
         );
  INV_X1 U7259 ( .A(n6273), .ZN(n6275) );
  AOI22_X1 U7260 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6289), .B1(n6417), 
        .B2(n6288), .ZN(n6274) );
  OAI211_X1 U7261 ( .C1(n6286), .C2(n6420), .A(n6275), .B(n6274), .ZN(U3047)
         );
  OAI22_X1 U7262 ( .A1(n6305), .A2(n6427), .B1(n6421), .B2(n6285), .ZN(n6276)
         );
  INV_X1 U7263 ( .A(n6276), .ZN(n6278) );
  AOI22_X1 U7264 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6289), .B1(n6424), 
        .B2(n6288), .ZN(n6277) );
  OAI211_X1 U7265 ( .C1(n6286), .C2(n6422), .A(n6278), .B(n6277), .ZN(U3048)
         );
  OAI22_X1 U7266 ( .A1(n6305), .A2(n6429), .B1(n6428), .B2(n6285), .ZN(n6279)
         );
  INV_X1 U7267 ( .A(n6279), .ZN(n6281) );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6289), .B1(n6431), 
        .B2(n6288), .ZN(n6280) );
  OAI211_X1 U7269 ( .C1(n6286), .C2(n6434), .A(n6281), .B(n6280), .ZN(U3049)
         );
  OAI22_X1 U7270 ( .A1(n6286), .A2(n6441), .B1(n6435), .B2(n6285), .ZN(n6282)
         );
  INV_X1 U7271 ( .A(n6282), .ZN(n6284) );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6289), .B1(n6438), 
        .B2(n6288), .ZN(n6283) );
  OAI211_X1 U7273 ( .C1(n6436), .C2(n6305), .A(n6284), .B(n6283), .ZN(U3050)
         );
  OAI22_X1 U7274 ( .A1(n6286), .A2(n6453), .B1(n6443), .B2(n6285), .ZN(n6287)
         );
  INV_X1 U7275 ( .A(n6287), .ZN(n6291) );
  AOI22_X1 U7276 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6289), .B1(n6448), 
        .B2(n6288), .ZN(n6290) );
  OAI211_X1 U7277 ( .C1(n6444), .C2(n6305), .A(n6291), .B(n6290), .ZN(U3051)
         );
  OAI22_X1 U7278 ( .A1(n6400), .A2(n6299), .B1(n6298), .B2(n6360), .ZN(n6292)
         );
  INV_X1 U7279 ( .A(n6292), .ZN(n6294) );
  AOI22_X1 U7280 ( .A1(n6302), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6362), 
        .B2(n6301), .ZN(n6293) );
  OAI211_X1 U7281 ( .C1(n6401), .C2(n6305), .A(n6294), .B(n6293), .ZN(U3053)
         );
  OAI22_X1 U7282 ( .A1(n6414), .A2(n6299), .B1(n6298), .B2(n6365), .ZN(n6295)
         );
  INV_X1 U7283 ( .A(n6295), .ZN(n6297) );
  AOI22_X1 U7284 ( .A1(n6302), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6367), 
        .B2(n6301), .ZN(n6296) );
  OAI211_X1 U7285 ( .C1(n6420), .C2(n6305), .A(n6297), .B(n6296), .ZN(U3055)
         );
  OAI22_X1 U7286 ( .A1(n6421), .A2(n6299), .B1(n6298), .B2(n6370), .ZN(n6300)
         );
  INV_X1 U7287 ( .A(n6300), .ZN(n6304) );
  AOI22_X1 U7288 ( .A1(n6302), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6375), 
        .B2(n6301), .ZN(n6303) );
  OAI211_X1 U7289 ( .C1(n6422), .C2(n6305), .A(n6304), .B(n6303), .ZN(U3056)
         );
  NOR2_X1 U7290 ( .A1(n6306), .A2(n6390), .ZN(n6311) );
  NAND3_X1 U7291 ( .A1(n6308), .A2(n6307), .A3(n3383), .ZN(n6309) );
  NAND2_X1 U7292 ( .A1(n6309), .A2(n6343), .ZN(n6314) );
  OAI22_X1 U7293 ( .A1(n6379), .A2(n6382), .B1(n6381), .B2(n6343), .ZN(n6310)
         );
  INV_X1 U7294 ( .A(n6310), .ZN(n6318) );
  INV_X1 U7295 ( .A(n6311), .ZN(n6315) );
  AOI21_X1 U7296 ( .B1(n6312), .B2(n6390), .A(n6389), .ZN(n6313) );
  AOI22_X1 U7297 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6355), .B1(n6316), 
        .B2(n6352), .ZN(n6317) );
  OAI211_X1 U7298 ( .C1(n6359), .C2(n6319), .A(n6318), .B(n6317), .ZN(U3076)
         );
  OAI22_X1 U7299 ( .A1(n6379), .A2(n6406), .B1(n6400), .B2(n6343), .ZN(n6320)
         );
  INV_X1 U7300 ( .A(n6320), .ZN(n6323) );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6355), .B1(n6321), 
        .B2(n6352), .ZN(n6322) );
  OAI211_X1 U7302 ( .C1(n6359), .C2(n6360), .A(n6323), .B(n6322), .ZN(U3077)
         );
  OAI22_X1 U7303 ( .A1(n6379), .A2(n6413), .B1(n6407), .B2(n6343), .ZN(n6324)
         );
  INV_X1 U7304 ( .A(n6324), .ZN(n6327) );
  AOI22_X1 U7305 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6355), .B1(n6325), 
        .B2(n6352), .ZN(n6326) );
  OAI211_X1 U7306 ( .C1(n6359), .C2(n6328), .A(n6327), .B(n6326), .ZN(U3078)
         );
  INV_X1 U7307 ( .A(n6343), .ZN(n6349) );
  AOI22_X1 U7308 ( .A1(n6352), .A2(n6330), .B1(n6329), .B2(n6349), .ZN(n6332)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6355), .B1(n6367), 
        .B2(n6353), .ZN(n6331) );
  OAI211_X1 U7310 ( .C1(n6359), .C2(n6365), .A(n6332), .B(n6331), .ZN(U3079)
         );
  AOI22_X1 U7311 ( .A1(n6352), .A2(n6334), .B1(n6333), .B2(n6349), .ZN(n6336)
         );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6355), .B1(n6375), 
        .B2(n6353), .ZN(n6335) );
  OAI211_X1 U7313 ( .C1(n6359), .C2(n6370), .A(n6336), .B(n6335), .ZN(U3080)
         );
  AOI22_X1 U7314 ( .A1(n6352), .A2(n6338), .B1(n6337), .B2(n6349), .ZN(n6341)
         );
  AOI22_X1 U7315 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6355), .B1(n6339), 
        .B2(n6353), .ZN(n6340) );
  OAI211_X1 U7316 ( .C1(n6359), .C2(n6342), .A(n6341), .B(n6340), .ZN(U3081)
         );
  OAI22_X1 U7317 ( .A1(n6379), .A2(n6436), .B1(n6435), .B2(n6343), .ZN(n6344)
         );
  INV_X1 U7318 ( .A(n6344), .ZN(n6347) );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6355), .B1(n6345), 
        .B2(n6352), .ZN(n6346) );
  OAI211_X1 U7320 ( .C1(n6359), .C2(n6348), .A(n6347), .B(n6346), .ZN(U3082)
         );
  AOI22_X1 U7321 ( .A1(n6352), .A2(n6351), .B1(n6350), .B2(n6349), .ZN(n6357)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6355), .B1(n6354), 
        .B2(n6353), .ZN(n6356) );
  OAI211_X1 U7323 ( .C1(n6359), .C2(n6358), .A(n6357), .B(n6356), .ZN(U3083)
         );
  OAI22_X1 U7324 ( .A1(n6400), .A2(n6372), .B1(n6371), .B2(n6360), .ZN(n6361)
         );
  INV_X1 U7325 ( .A(n6361), .ZN(n6364) );
  AOI22_X1 U7326 ( .A1(n6376), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6362), 
        .B2(n6374), .ZN(n6363) );
  OAI211_X1 U7327 ( .C1(n6401), .C2(n6379), .A(n6364), .B(n6363), .ZN(U3085)
         );
  OAI22_X1 U7328 ( .A1(n6414), .A2(n6372), .B1(n6371), .B2(n6365), .ZN(n6366)
         );
  INV_X1 U7329 ( .A(n6366), .ZN(n6369) );
  AOI22_X1 U7330 ( .A1(n6376), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6367), 
        .B2(n6374), .ZN(n6368) );
  OAI211_X1 U7331 ( .C1(n6420), .C2(n6379), .A(n6369), .B(n6368), .ZN(U3087)
         );
  OAI22_X1 U7332 ( .A1(n6421), .A2(n6372), .B1(n6371), .B2(n6370), .ZN(n6373)
         );
  INV_X1 U7333 ( .A(n6373), .ZN(n6378) );
  AOI22_X1 U7334 ( .A1(n6376), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6375), 
        .B2(n6374), .ZN(n6377) );
  OAI211_X1 U7335 ( .C1(n6422), .C2(n6379), .A(n6378), .B(n6377), .ZN(U3088)
         );
  NAND2_X1 U7336 ( .A1(n6380), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6442) );
  OAI22_X1 U7337 ( .A1(n6445), .A2(n6382), .B1(n6381), .B2(n6442), .ZN(n6383)
         );
  INV_X1 U7338 ( .A(n6383), .ZN(n6398) );
  OAI21_X1 U7339 ( .B1(n6386), .B2(n6385), .A(n6384), .ZN(n6395) );
  NAND2_X1 U7340 ( .A1(n6387), .A2(n3383), .ZN(n6388) );
  NAND2_X1 U7341 ( .A1(n6388), .A2(n6442), .ZN(n6392) );
  AOI21_X1 U7342 ( .B1(n6393), .B2(n6390), .A(n6389), .ZN(n6391) );
  OAI21_X1 U7343 ( .B1(n6395), .B2(n6392), .A(n6391), .ZN(n6449) );
  INV_X1 U7344 ( .A(n6392), .ZN(n6394) );
  OAI22_X1 U7345 ( .A1(n6395), .A2(n6394), .B1(n6393), .B2(n6503), .ZN(n6447)
         );
  AOI22_X1 U7346 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6449), .B1(n6396), 
        .B2(n6447), .ZN(n6397) );
  OAI211_X1 U7347 ( .C1(n6399), .C2(n6452), .A(n6398), .B(n6397), .ZN(U3108)
         );
  OAI22_X1 U7348 ( .A1(n6452), .A2(n6401), .B1(n6400), .B2(n6442), .ZN(n6402)
         );
  INV_X1 U7349 ( .A(n6402), .ZN(n6405) );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6449), .B1(n6403), 
        .B2(n6447), .ZN(n6404) );
  OAI211_X1 U7351 ( .C1(n6406), .C2(n6445), .A(n6405), .B(n6404), .ZN(U3109)
         );
  OAI22_X1 U7352 ( .A1(n6452), .A2(n6408), .B1(n6407), .B2(n6442), .ZN(n6409)
         );
  INV_X1 U7353 ( .A(n6409), .ZN(n6412) );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6449), .B1(n6410), 
        .B2(n6447), .ZN(n6411) );
  OAI211_X1 U7355 ( .C1(n6413), .C2(n6445), .A(n6412), .B(n6411), .ZN(U3110)
         );
  OAI22_X1 U7356 ( .A1(n6445), .A2(n6415), .B1(n6414), .B2(n6442), .ZN(n6416)
         );
  INV_X1 U7357 ( .A(n6416), .ZN(n6419) );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6449), .B1(n6417), 
        .B2(n6447), .ZN(n6418) );
  OAI211_X1 U7359 ( .C1(n6420), .C2(n6452), .A(n6419), .B(n6418), .ZN(U3111)
         );
  OAI22_X1 U7360 ( .A1(n6452), .A2(n6422), .B1(n6421), .B2(n6442), .ZN(n6423)
         );
  INV_X1 U7361 ( .A(n6423), .ZN(n6426) );
  AOI22_X1 U7362 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6449), .B1(n6424), 
        .B2(n6447), .ZN(n6425) );
  OAI211_X1 U7363 ( .C1(n6427), .C2(n6445), .A(n6426), .B(n6425), .ZN(U3112)
         );
  OAI22_X1 U7364 ( .A1(n6445), .A2(n6429), .B1(n6428), .B2(n6442), .ZN(n6430)
         );
  INV_X1 U7365 ( .A(n6430), .ZN(n6433) );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6449), .B1(n6431), 
        .B2(n6447), .ZN(n6432) );
  OAI211_X1 U7367 ( .C1(n6434), .C2(n6452), .A(n6433), .B(n6432), .ZN(U3113)
         );
  OAI22_X1 U7368 ( .A1(n6445), .A2(n6436), .B1(n6435), .B2(n6442), .ZN(n6437)
         );
  INV_X1 U7369 ( .A(n6437), .ZN(n6440) );
  AOI22_X1 U7370 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6449), .B1(n6438), 
        .B2(n6447), .ZN(n6439) );
  OAI211_X1 U7371 ( .C1(n6441), .C2(n6452), .A(n6440), .B(n6439), .ZN(U3114)
         );
  OAI22_X1 U7372 ( .A1(n6445), .A2(n6444), .B1(n6443), .B2(n6442), .ZN(n6446)
         );
  INV_X1 U7373 ( .A(n6446), .ZN(n6451) );
  AOI22_X1 U7374 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6449), .B1(n6448), 
        .B2(n6447), .ZN(n6450) );
  OAI211_X1 U7375 ( .C1(n6453), .C2(n6452), .A(n6451), .B(n6450), .ZN(U3115)
         );
  AOI21_X1 U7376 ( .B1(n6469), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6486) );
  INV_X1 U7377 ( .A(n6454), .ZN(n6456) );
  NOR3_X1 U7378 ( .A1(n6457), .A2(n6456), .A3(n6455), .ZN(n6463) );
  INV_X1 U7379 ( .A(n6463), .ZN(n6460) );
  OAI211_X1 U7380 ( .C1(n6461), .C2(n6460), .A(n6459), .B(n6458), .ZN(n6462)
         );
  OAI21_X1 U7381 ( .B1(n6463), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6462), 
        .ZN(n6465) );
  AOI21_X1 U7382 ( .B1(n6465), .B2(n6466), .A(n6464), .ZN(n6468) );
  NOR2_X1 U7383 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  OAI22_X1 U7384 ( .A1(n6469), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6468), .B2(n6467), .ZN(n6485) );
  INV_X1 U7385 ( .A(n6470), .ZN(n6482) );
  OAI21_X1 U7386 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6471), 
        .ZN(n6481) );
  INV_X1 U7387 ( .A(n3999), .ZN(n6472) );
  NOR3_X1 U7388 ( .A1(n6474), .A2(n6473), .A3(n6472), .ZN(n6477) );
  OAI22_X1 U7389 ( .A1(n6480), .A2(n6477), .B1(n6476), .B2(n6475), .ZN(n6478)
         );
  AOI21_X1 U7390 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n6599) );
  NAND4_X1 U7391 ( .A1(n6482), .A2(n6481), .A3(n4293), .A4(n6599), .ZN(n6484)
         );
  AOI211_X1 U7392 ( .C1(n6486), .C2(n6485), .A(n6484), .B(n6483), .ZN(n6500)
         );
  NOR3_X1 U7394 ( .A1(n6488), .A2(n6605), .A3(n6487), .ZN(n6490) );
  AOI21_X1 U7395 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6489) );
  NOR3_X1 U7396 ( .A1(n6490), .A2(n6489), .A3(n6503), .ZN(n6492) );
  AOI21_X1 U7397 ( .B1(n6491), .B2(n6606), .A(n6492), .ZN(n6495) );
  OAI221_X1 U7398 ( .B1(n6504), .B2(n6500), .C1(n6504), .C2(n6493), .A(n6492), 
        .ZN(n6588) );
  OAI21_X1 U7399 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6708), .A(n6588), .ZN(
        n6505) );
  OAI33_X1 U7400 ( .A1(1'b0), .A2(n6495), .A3(STATE2_REG_0__SCAN_IN), .B1(
        n6504), .B2(n6494), .B3(n6505), .ZN(n6498) );
  OAI211_X1 U7401 ( .C1(n6500), .C2(n6499), .A(n6498), .B(n6497), .ZN(U3148)
         );
  INV_X1 U7402 ( .A(n6588), .ZN(n6509) );
  AOI21_X1 U7403 ( .B1(n6502), .B2(n6708), .A(n6501), .ZN(n6508) );
  NAND2_X1 U7404 ( .A1(n6504), .A2(n6503), .ZN(n6510) );
  NAND3_X1 U7405 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6510), .A3(n6505), .ZN(
        n6506) );
  OAI211_X1 U7406 ( .C1(n6509), .C2(n6508), .A(n6507), .B(n6506), .ZN(U3149)
         );
  OAI211_X1 U7407 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6708), .A(n6586), .B(
        n6510), .ZN(n6512) );
  OAI21_X1 U7408 ( .B1(n6606), .B2(n6512), .A(n6511), .ZN(U3150) );
  INV_X1 U7409 ( .A(n6585), .ZN(n6581) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6581), .ZN(U3151) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6581), .ZN(U3152) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6581), .ZN(U3153) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6581), .ZN(U3154) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6581), .ZN(U3155) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6581), .ZN(U3156) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6581), .ZN(U3157) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6581), .ZN(U3158) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6581), .ZN(U3159) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6581), .ZN(U3160) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6581), .ZN(U3161) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6581), .ZN(U3162) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6581), .ZN(U3163) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6581), .ZN(U3164) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6581), .ZN(U3165) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6581), .ZN(U3166) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6581), .ZN(U3167) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6581), .ZN(U3168) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6581), .ZN(U3169) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6581), .ZN(U3170) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6581), .ZN(U3171) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6581), .ZN(U3172) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6581), .ZN(U3173) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6581), .ZN(U3174) );
  AND2_X1 U7434 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6581), .ZN(U3175) );
  AND2_X1 U7435 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6581), .ZN(U3176) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6581), .ZN(U3177) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6581), .ZN(U3178) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6581), .ZN(U3179) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6581), .ZN(U3180) );
  NOR2_X1 U7440 ( .A1(n6519), .A2(n6513), .ZN(n6520) );
  AOI22_X1 U7441 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6528) );
  INV_X1 U7442 ( .A(HOLD), .ZN(n6740) );
  NOR2_X1 U7443 ( .A1(n6519), .A2(n6740), .ZN(n6516) );
  INV_X2 U7444 ( .A(n6812), .ZN(n6811) );
  INV_X1 U7445 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6716) );
  INV_X1 U7446 ( .A(NA_N), .ZN(n6521) );
  AOI221_X1 U7447 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6521), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6525) );
  AOI221_X1 U7448 ( .B1(n6516), .B2(n6811), .C1(n6716), .C2(n6811), .A(n6525), 
        .ZN(n6514) );
  OAI21_X1 U7449 ( .B1(n6520), .B2(n6528), .A(n6514), .ZN(U3181) );
  NOR2_X1 U7450 ( .A1(n6523), .A2(n6716), .ZN(n6522) );
  NAND2_X1 U7451 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6515) );
  OAI21_X1 U7452 ( .B1(n6522), .B2(n6516), .A(n6515), .ZN(n6517) );
  OAI211_X1 U7453 ( .C1(n6519), .C2(n6708), .A(n6518), .B(n6517), .ZN(U3182)
         );
  AOI21_X1 U7454 ( .B1(n6522), .B2(n6521), .A(n6520), .ZN(n6527) );
  AOI221_X1 U7455 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6708), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6524) );
  AOI221_X1 U7456 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6524), .C2(HOLD), .A(n6523), .ZN(n6526) );
  OAI22_X1 U7457 ( .A1(n6528), .A2(n6527), .B1(n6526), .B2(n6525), .ZN(U3183)
         );
  NAND2_X2 U7458 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6812), .ZN(n6575) );
  AOI22_X1 U7459 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6811), .ZN(n6529) );
  OAI21_X1 U7460 ( .B1(n6590), .B2(n6575), .A(n6529), .ZN(U3184) );
  AOI22_X1 U7461 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6811), .ZN(n6530) );
  OAI21_X1 U7462 ( .B1(n6531), .B2(n6575), .A(n6530), .ZN(U3185) );
  AOI22_X1 U7463 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6811), .ZN(n6532) );
  OAI21_X1 U7464 ( .B1(n6533), .B2(n6575), .A(n6532), .ZN(U3186) );
  AOI22_X1 U7465 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6811), .ZN(n6534) );
  OAI21_X1 U7466 ( .B1(n6535), .B2(n6575), .A(n6534), .ZN(U3187) );
  AOI22_X1 U7467 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6811), .ZN(n6536) );
  OAI21_X1 U7468 ( .B1(n6537), .B2(n6575), .A(n6536), .ZN(U3188) );
  AOI22_X1 U7469 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6811), .ZN(n6538) );
  OAI21_X1 U7470 ( .B1(n6539), .B2(n6575), .A(n6538), .ZN(U3189) );
  AOI22_X1 U7471 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6811), .ZN(n6540) );
  OAI21_X1 U7472 ( .B1(n6541), .B2(n6575), .A(n6540), .ZN(U3190) );
  AOI22_X1 U7473 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6811), .ZN(n6542) );
  OAI21_X1 U7474 ( .B1(n6543), .B2(n6575), .A(n6542), .ZN(U3191) );
  AOI22_X1 U7475 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6811), .ZN(n6544) );
  OAI21_X1 U7476 ( .B1(n6545), .B2(n6575), .A(n6544), .ZN(U3192) );
  AOI22_X1 U7477 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6811), .ZN(n6546) );
  OAI21_X1 U7478 ( .B1(n6547), .B2(n6575), .A(n6546), .ZN(U3193) );
  AOI22_X1 U7479 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6811), .ZN(n6548) );
  OAI21_X1 U7480 ( .B1(n6549), .B2(n6575), .A(n6548), .ZN(U3194) );
  AOI22_X1 U7481 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6811), .ZN(n6550) );
  OAI21_X1 U7482 ( .B1(n6551), .B2(n6575), .A(n6550), .ZN(U3195) );
  INV_X2 U7483 ( .A(n6579), .ZN(n6573) );
  AOI22_X1 U7484 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6811), .ZN(n6552) );
  OAI21_X1 U7485 ( .B1(n6553), .B2(n6575), .A(n6552), .ZN(U3196) );
  AOI22_X1 U7486 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6811), .ZN(n6554) );
  OAI21_X1 U7487 ( .B1(n6555), .B2(n6575), .A(n6554), .ZN(U3197) );
  AOI22_X1 U7488 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6811), .ZN(n6556) );
  OAI21_X1 U7489 ( .B1(n6557), .B2(n6575), .A(n6556), .ZN(U3198) );
  AOI22_X1 U7490 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6811), .ZN(n6558) );
  OAI21_X1 U7491 ( .B1(n6559), .B2(n6575), .A(n6558), .ZN(U3199) );
  AOI22_X1 U7492 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6811), .ZN(n6560) );
  OAI21_X1 U7493 ( .B1(n6561), .B2(n6575), .A(n6560), .ZN(U3200) );
  AOI22_X1 U7494 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6811), .ZN(n6562) );
  OAI21_X1 U7495 ( .B1(n6563), .B2(n6575), .A(n6562), .ZN(U3201) );
  INV_X1 U7496 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U7497 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6811), .ZN(n6564) );
  OAI21_X1 U7498 ( .B1(n6810), .B2(n6575), .A(n6564), .ZN(U3202) );
  AOI22_X1 U7499 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6811), .ZN(n6565) );
  OAI21_X1 U7500 ( .B1(n6705), .B2(n6575), .A(n6565), .ZN(U3203) );
  AOI22_X1 U7501 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6811), .ZN(n6566) );
  OAI21_X1 U7502 ( .B1(n6751), .B2(n6575), .A(n6566), .ZN(U3204) );
  AOI22_X1 U7503 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6811), .ZN(n6567) );
  OAI21_X1 U7504 ( .B1(n6750), .B2(n6575), .A(n6567), .ZN(U3205) );
  AOI22_X1 U7505 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6811), .ZN(n6568) );
  OAI21_X1 U7506 ( .B1(n6723), .B2(n6575), .A(n6568), .ZN(U3206) );
  AOI22_X1 U7507 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6811), .ZN(n6569) );
  OAI21_X1 U7508 ( .B1(n6628), .B2(n6575), .A(n6569), .ZN(U3207) );
  AOI22_X1 U7509 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6811), .ZN(n6570) );
  OAI21_X1 U7510 ( .B1(n6785), .B2(n6575), .A(n6570), .ZN(U3208) );
  AOI22_X1 U7511 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6811), .ZN(n6571) );
  OAI21_X1 U7512 ( .B1(n6726), .B2(n6579), .A(n6571), .ZN(U3209) );
  AOI22_X1 U7513 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6811), .ZN(n6572) );
  OAI21_X1 U7514 ( .B1(n6726), .B2(n6575), .A(n6572), .ZN(U3210) );
  AOI22_X1 U7515 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6573), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6811), .ZN(n6574) );
  OAI21_X1 U7516 ( .B1(n6733), .B2(n6575), .A(n6574), .ZN(U3211) );
  AOI22_X1 U7517 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6811), .ZN(n6576) );
  OAI21_X1 U7518 ( .B1(n6748), .B2(n6579), .A(n6576), .ZN(U3212) );
  AOI22_X1 U7519 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6811), .ZN(n6578) );
  OAI21_X1 U7520 ( .B1(n6688), .B2(n6579), .A(n6578), .ZN(U3213) );
  MUX2_X1 U7521 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6812), .Z(U3446) );
  MUX2_X1 U7522 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6812), .Z(U3447) );
  MUX2_X1 U7523 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6812), .Z(U3448) );
  INV_X1 U7524 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6582) );
  INV_X1 U7525 ( .A(n6583), .ZN(n6580) );
  AOI21_X1 U7526 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(U3451) );
  OAI21_X1 U7527 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(U3452) );
  OAI211_X1 U7528 ( .C1(n6589), .C2(n6588), .A(n6587), .B(n6586), .ZN(U3453)
         );
  AOI21_X1 U7529 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6591) );
  AOI22_X1 U7530 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6591), .B2(n6590), .ZN(n6594) );
  INV_X1 U7531 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U7532 ( .A1(n6597), .A2(n6594), .B1(n6593), .B2(n6592), .ZN(U3468)
         );
  INV_X1 U7533 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6596) );
  OAI21_X1 U7534 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6597), .ZN(n6595) );
  OAI21_X1 U7535 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(U3469) );
  INV_X1 U7536 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6673) );
  AOI22_X1 U7537 ( .A1(n6812), .A2(READREQUEST_REG_SCAN_IN), .B1(n6673), .B2(
        n6811), .ZN(U3470) );
  INV_X1 U7538 ( .A(MORE_REG_SCAN_IN), .ZN(n6756) );
  INV_X1 U7539 ( .A(n6600), .ZN(n6598) );
  AOI22_X1 U7540 ( .A1(n6600), .A2(n6599), .B1(n6756), .B2(n6598), .ZN(U3471)
         );
  AOI211_X1 U7541 ( .C1(n6603), .C2(n6708), .A(n6602), .B(n6601), .ZN(n6610)
         );
  OAI211_X1 U7542 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6605), .A(n6604), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6607) );
  AOI21_X1 U7543 ( .B1(n6607), .B2(STATE2_REG_0__SCAN_IN), .A(n6606), .ZN(
        n6609) );
  NAND2_X1 U7544 ( .A1(n6610), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6608) );
  OAI21_X1 U7545 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(U3472) );
  INV_X1 U7546 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6643) );
  AOI22_X1 U7547 ( .A1(n6812), .A2(n6707), .B1(n6643), .B2(n6811), .ZN(U3473)
         );
  AOI22_X1 U7548 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(REIP_REG_23__SCAN_IN), 
        .B2(keyinput_f59), .ZN(n6611) );
  OAI221_X1 U7549 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(REIP_REG_23__SCAN_IN), .C2(keyinput_f59), .A(n6611), .ZN(n6670) );
  AOI22_X1 U7550 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_f37), .B1(
        DATAI_16_), .B2(keyinput_f15), .ZN(n6612) );
  OAI221_X1 U7551 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_f37), .C1(
        DATAI_16_), .C2(keyinput_f15), .A(n6612), .ZN(n6669) );
  INV_X1 U7552 ( .A(DATAI_31_), .ZN(n6738) );
  AOI22_X1 U7553 ( .A1(keyinput_f49), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        n6738), .B2(keyinput_f0), .ZN(n6613) );
  OAI221_X1 U7554 ( .B1(keyinput_f49), .B2(BYTEENABLE_REG_2__SCAN_IN), .C1(
        n6738), .C2(keyinput_f0), .A(n6613), .ZN(n6623) );
  OAI22_X1 U7555 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(
        keyinput_f9), .B2(DATAI_22_), .ZN(n6614) );
  AOI221_X1 U7556 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        DATAI_22_), .C2(keyinput_f9), .A(n6614), .ZN(n6621) );
  OAI22_X1 U7557 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_f55), .B1(
        keyinput_f57), .B2(REIP_REG_25__SCAN_IN), .ZN(n6615) );
  AOI221_X1 U7558 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_f55), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_f57), .A(n6615), .ZN(n6620) );
  OAI22_X1 U7559 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n6616) );
  AOI221_X1 U7560 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(keyinput_f42), .C2(
        REQUESTPENDING_REG_SCAN_IN), .A(n6616), .ZN(n6619) );
  OAI22_X1 U7561 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(keyinput_f30), .B2(
        DATAI_1_), .ZN(n6617) );
  AOI221_X1 U7562 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(DATAI_1_), .C2(
        keyinput_f30), .A(n6617), .ZN(n6618) );
  NAND4_X1 U7563 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6622)
         );
  AOI211_X1 U7564 ( .C1(keyinput_f56), .C2(REIP_REG_26__SCAN_IN), .A(n6623), 
        .B(n6622), .ZN(n6624) );
  OAI21_X1 U7565 ( .B1(keyinput_f56), .B2(REIP_REG_26__SCAN_IN), .A(n6624), 
        .ZN(n6668) );
  AOI22_X1 U7566 ( .A1(keyinput_f36), .A2(HOLD), .B1(DATAI_5_), .B2(
        keyinput_f26), .ZN(n6625) );
  OAI221_X1 U7567 ( .B1(keyinput_f36), .B2(HOLD), .C1(DATAI_5_), .C2(
        keyinput_f26), .A(n6625), .ZN(n6633) );
  AOI22_X1 U7568 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        DATAI_11_), .B2(keyinput_f20), .ZN(n6626) );
  OAI221_X1 U7569 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        DATAI_11_), .C2(keyinput_f20), .A(n6626), .ZN(n6632) );
  AOI22_X1 U7570 ( .A1(n6628), .A2(keyinput_f58), .B1(keyinput_f17), .B2(n6774), .ZN(n6627) );
  OAI221_X1 U7571 ( .B1(n6628), .B2(keyinput_f58), .C1(n6774), .C2(
        keyinput_f17), .A(n6627), .ZN(n6631) );
  AOI22_X1 U7572 ( .A1(keyinput_f33), .A2(NA_N), .B1(REIP_REG_20__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n6629) );
  OAI221_X1 U7573 ( .B1(keyinput_f33), .B2(NA_N), .C1(REIP_REG_20__SCAN_IN), 
        .C2(keyinput_f62), .A(n6629), .ZN(n6630) );
  NOR4_X1 U7574 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6666)
         );
  AOI22_X1 U7575 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_f44), .B1(DATAI_8_), 
        .B2(keyinput_f23), .ZN(n6634) );
  OAI221_X1 U7576 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_f44), .C1(DATAI_8_), 
        .C2(keyinput_f23), .A(n6634), .ZN(n6641) );
  AOI22_X1 U7577 ( .A1(keyinput_f38), .A2(ADS_N_REG_SCAN_IN), .B1(DATAI_4_), 
        .B2(keyinput_f27), .ZN(n6635) );
  OAI221_X1 U7578 ( .B1(keyinput_f38), .B2(ADS_N_REG_SCAN_IN), .C1(DATAI_4_), 
        .C2(keyinput_f27), .A(n6635), .ZN(n6640) );
  AOI22_X1 U7579 ( .A1(keyinput_f34), .A2(BS16_N), .B1(DATAI_26_), .B2(
        keyinput_f5), .ZN(n6636) );
  OAI221_X1 U7580 ( .B1(keyinput_f34), .B2(BS16_N), .C1(DATAI_26_), .C2(
        keyinput_f5), .A(n6636), .ZN(n6639) );
  AOI22_X1 U7581 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n6637) );
  OAI221_X1 U7582 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n6637), .ZN(n6638) );
  NOR4_X1 U7583 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n6665)
         );
  AOI22_X1 U7584 ( .A1(n6644), .A2(keyinput_f19), .B1(keyinput_f40), .B2(n6643), .ZN(n6642) );
  OAI221_X1 U7585 ( .B1(n6644), .B2(keyinput_f19), .C1(n6643), .C2(
        keyinput_f40), .A(n6642), .ZN(n6652) );
  AOI22_X1 U7586 ( .A1(n6750), .A2(keyinput_f60), .B1(keyinput_f45), .B2(n6741), .ZN(n6645) );
  OAI221_X1 U7587 ( .B1(n6750), .B2(keyinput_f60), .C1(n6741), .C2(
        keyinput_f45), .A(n6645), .ZN(n6651) );
  AOI22_X1 U7588 ( .A1(n6733), .A2(keyinput_f54), .B1(keyinput_f31), .B2(n6747), .ZN(n6646) );
  OAI221_X1 U7589 ( .B1(n6733), .B2(keyinput_f54), .C1(n6747), .C2(
        keyinput_f31), .A(n6646), .ZN(n6650) );
  AOI22_X1 U7590 ( .A1(n6648), .A2(keyinput_f24), .B1(keyinput_f32), .B2(n6707), .ZN(n6647) );
  OAI221_X1 U7591 ( .B1(n6648), .B2(keyinput_f24), .C1(n6707), .C2(
        keyinput_f32), .A(n6647), .ZN(n6649) );
  NOR4_X1 U7592 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6664)
         );
  AOI22_X1 U7593 ( .A1(n6717), .A2(keyinput_f8), .B1(n6748), .B2(keyinput_f52), 
        .ZN(n6653) );
  OAI221_X1 U7594 ( .B1(n6717), .B2(keyinput_f8), .C1(n6748), .C2(keyinput_f52), .A(n6653), .ZN(n6662) );
  INV_X1 U7595 ( .A(DATAI_28_), .ZN(n6655) );
  AOI22_X1 U7596 ( .A1(n6655), .A2(keyinput_f3), .B1(n6751), .B2(keyinput_f61), 
        .ZN(n6654) );
  OAI221_X1 U7597 ( .B1(n6655), .B2(keyinput_f3), .C1(n6751), .C2(keyinput_f61), .A(n6654), .ZN(n6661) );
  AOI22_X1 U7598 ( .A1(n6788), .A2(keyinput_f10), .B1(n6782), .B2(keyinput_f25), .ZN(n6656) );
  OAI221_X1 U7599 ( .B1(n6788), .B2(keyinput_f10), .C1(n6782), .C2(
        keyinput_f25), .A(n6656), .ZN(n6660) );
  INV_X1 U7600 ( .A(DATAI_17_), .ZN(n6658) );
  AOI22_X1 U7601 ( .A1(n6786), .A2(keyinput_f28), .B1(keyinput_f14), .B2(n6658), .ZN(n6657) );
  OAI221_X1 U7602 ( .B1(n6786), .B2(keyinput_f28), .C1(n6658), .C2(
        keyinput_f14), .A(n6657), .ZN(n6659) );
  NOR4_X1 U7603 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6663)
         );
  NAND4_X1 U7604 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6667)
         );
  NOR4_X1 U7605 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6699)
         );
  XOR2_X1 U7606 ( .A(keyinput_f47), .B(BYTEENABLE_REG_0__SCAN_IN), .Z(n6675)
         );
  AOI22_X1 U7607 ( .A1(n6673), .A2(keyinput_f46), .B1(n6672), .B2(keyinput_f22), .ZN(n6671) );
  OAI221_X1 U7608 ( .B1(n6673), .B2(keyinput_f46), .C1(n6672), .C2(
        keyinput_f22), .A(n6671), .ZN(n6674) );
  AOI211_X1 U7609 ( .C1(n6710), .C2(keyinput_f48), .A(n6675), .B(n6674), .ZN(
        n6676) );
  OAI21_X1 U7610 ( .B1(n6710), .B2(keyinput_f48), .A(n6676), .ZN(n6696) );
  AOI22_X1 U7611 ( .A1(n6679), .A2(keyinput_f12), .B1(keyinput_f41), .B2(n6678), .ZN(n6677) );
  OAI221_X1 U7612 ( .B1(n6679), .B2(keyinput_f12), .C1(n6678), .C2(
        keyinput_f41), .A(n6677), .ZN(n6695) );
  AOI22_X1 U7613 ( .A1(n6719), .A2(keyinput_f29), .B1(n4617), .B2(keyinput_f7), 
        .ZN(n6680) );
  OAI221_X1 U7614 ( .B1(n6719), .B2(keyinput_f29), .C1(n4617), .C2(keyinput_f7), .A(n6680), .ZN(n6694) );
  OAI22_X1 U7615 ( .A1(n6683), .A2(keyinput_f18), .B1(n6682), .B2(keyinput_f11), .ZN(n6681) );
  AOI221_X1 U7616 ( .B1(n6683), .B2(keyinput_f18), .C1(keyinput_f11), .C2(
        n6682), .A(n6681), .ZN(n6692) );
  OAI22_X1 U7617 ( .A1(n6685), .A2(keyinput_f53), .B1(n6735), .B2(keyinput_f21), .ZN(n6684) );
  AOI221_X1 U7618 ( .B1(n6685), .B2(keyinput_f53), .C1(keyinput_f21), .C2(
        n6735), .A(n6684), .ZN(n6691) );
  OAI22_X1 U7619 ( .A1(n6708), .A2(keyinput_f35), .B1(n6755), .B2(keyinput_f50), .ZN(n6686) );
  AOI221_X1 U7620 ( .B1(n6708), .B2(keyinput_f35), .C1(keyinput_f50), .C2(
        n6755), .A(n6686), .ZN(n6690) );
  INV_X1 U7621 ( .A(DATAI_15_), .ZN(n6789) );
  OAI22_X1 U7622 ( .A1(n6688), .A2(keyinput_f51), .B1(n6789), .B2(keyinput_f16), .ZN(n6687) );
  AOI221_X1 U7623 ( .B1(n6688), .B2(keyinput_f51), .C1(keyinput_f16), .C2(
        n6789), .A(n6687), .ZN(n6689) );
  NAND4_X1 U7624 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6693)
         );
  NOR4_X1 U7625 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n6698)
         );
  NOR2_X1 U7626 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_f63), .ZN(n6697) );
  AOI221_X1 U7627 ( .B1(n6699), .B2(n6698), .C1(keyinput_f63), .C2(
        REIP_REG_19__SCAN_IN), .A(n6697), .ZN(n6809) );
  INV_X1 U7628 ( .A(DATAI_27_), .ZN(n6702) );
  INV_X1 U7629 ( .A(DATAI_18_), .ZN(n6701) );
  AOI22_X1 U7630 ( .A1(n6702), .A2(keyinput_g4), .B1(keyinput_g13), .B2(n6701), 
        .ZN(n6700) );
  OAI221_X1 U7631 ( .B1(n6702), .B2(keyinput_g4), .C1(n6701), .C2(keyinput_g13), .A(n6700), .ZN(n6714) );
  INV_X1 U7632 ( .A(BS16_N), .ZN(n6704) );
  AOI22_X1 U7633 ( .A1(n6705), .A2(keyinput_g62), .B1(keyinput_g34), .B2(n6704), .ZN(n6703) );
  OAI221_X1 U7634 ( .B1(n6705), .B2(keyinput_g62), .C1(n6704), .C2(
        keyinput_g34), .A(n6703), .ZN(n6713) );
  AOI22_X1 U7635 ( .A1(n6708), .A2(keyinput_g35), .B1(keyinput_g32), .B2(n6707), .ZN(n6706) );
  OAI221_X1 U7636 ( .B1(n6708), .B2(keyinput_g35), .C1(n6707), .C2(
        keyinput_g32), .A(n6706), .ZN(n6712) );
  AOI22_X1 U7637 ( .A1(n6710), .A2(keyinput_g48), .B1(n4620), .B2(keyinput_g1), 
        .ZN(n6709) );
  OAI221_X1 U7638 ( .B1(n6710), .B2(keyinput_g48), .C1(n4620), .C2(keyinput_g1), .A(n6709), .ZN(n6711) );
  NOR4_X1 U7639 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6764)
         );
  AOI22_X1 U7640 ( .A1(n6717), .A2(keyinput_g8), .B1(keyinput_g42), .B2(n6716), 
        .ZN(n6715) );
  OAI221_X1 U7641 ( .B1(n6717), .B2(keyinput_g8), .C1(n6716), .C2(keyinput_g42), .A(n6715), .ZN(n6730) );
  AOI22_X1 U7642 ( .A1(n6720), .A2(keyinput_g23), .B1(keyinput_g29), .B2(n6719), .ZN(n6718) );
  OAI221_X1 U7643 ( .B1(n6720), .B2(keyinput_g23), .C1(n6719), .C2(
        keyinput_g29), .A(n6718), .ZN(n6729) );
  INV_X1 U7644 ( .A(DATAI_22_), .ZN(n6722) );
  AOI22_X1 U7645 ( .A1(n6723), .A2(keyinput_g59), .B1(keyinput_g9), .B2(n6722), 
        .ZN(n6721) );
  OAI221_X1 U7646 ( .B1(n6723), .B2(keyinput_g59), .C1(n6722), .C2(keyinput_g9), .A(n6721), .ZN(n6728) );
  AOI22_X1 U7647 ( .A1(n6726), .A2(keyinput_g55), .B1(keyinput_g26), .B2(n6725), .ZN(n6724) );
  OAI221_X1 U7648 ( .B1(n6726), .B2(keyinput_g55), .C1(n6725), .C2(
        keyinput_g26), .A(n6724), .ZN(n6727) );
  NOR4_X1 U7649 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6763)
         );
  INV_X1 U7650 ( .A(DATAI_16_), .ZN(n6732) );
  AOI22_X1 U7651 ( .A1(n6733), .A2(keyinput_g54), .B1(keyinput_g15), .B2(n6732), .ZN(n6731) );
  OAI221_X1 U7652 ( .B1(n6733), .B2(keyinput_g54), .C1(n6732), .C2(
        keyinput_g15), .A(n6731), .ZN(n6745) );
  AOI22_X1 U7653 ( .A1(n6735), .A2(keyinput_g21), .B1(keyinput_g6), .B2(n4606), 
        .ZN(n6734) );
  OAI221_X1 U7654 ( .B1(n6735), .B2(keyinput_g21), .C1(n4606), .C2(keyinput_g6), .A(n6734), .ZN(n6744) );
  AOI22_X1 U7655 ( .A1(n6738), .A2(keyinput_g0), .B1(keyinput_g30), .B2(n6737), 
        .ZN(n6736) );
  OAI221_X1 U7656 ( .B1(n6738), .B2(keyinput_g0), .C1(n6737), .C2(keyinput_g30), .A(n6736), .ZN(n6743) );
  AOI22_X1 U7657 ( .A1(n6741), .A2(keyinput_g45), .B1(keyinput_g36), .B2(n6740), .ZN(n6739) );
  OAI221_X1 U7658 ( .B1(n6741), .B2(keyinput_g45), .C1(n6740), .C2(
        keyinput_g36), .A(n6739), .ZN(n6742) );
  NOR4_X1 U7659 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n6762)
         );
  AOI22_X1 U7660 ( .A1(n6748), .A2(keyinput_g52), .B1(keyinput_g31), .B2(n6747), .ZN(n6746) );
  OAI221_X1 U7661 ( .B1(n6748), .B2(keyinput_g52), .C1(n6747), .C2(
        keyinput_g31), .A(n6746), .ZN(n6760) );
  AOI22_X1 U7662 ( .A1(n6751), .A2(keyinput_g61), .B1(n6750), .B2(keyinput_g60), .ZN(n6749) );
  OAI221_X1 U7663 ( .B1(n6751), .B2(keyinput_g61), .C1(n6750), .C2(
        keyinput_g60), .A(n6749), .ZN(n6759) );
  INV_X1 U7664 ( .A(DATAI_29_), .ZN(n6753) );
  AOI22_X1 U7665 ( .A1(n6753), .A2(keyinput_g2), .B1(keyinput_g5), .B2(n4612), 
        .ZN(n6752) );
  OAI221_X1 U7666 ( .B1(n6753), .B2(keyinput_g2), .C1(n4612), .C2(keyinput_g5), 
        .A(n6752), .ZN(n6758) );
  AOI22_X1 U7667 ( .A1(n6756), .A2(keyinput_g44), .B1(keyinput_g50), .B2(n6755), .ZN(n6754) );
  OAI221_X1 U7668 ( .B1(n6756), .B2(keyinput_g44), .C1(n6755), .C2(
        keyinput_g50), .A(n6754), .ZN(n6757) );
  NOR4_X1 U7669 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6761)
         );
  NAND4_X1 U7670 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6807)
         );
  AOI22_X1 U7671 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        DATAI_17_), .B2(keyinput_g14), .ZN(n6765) );
  OAI221_X1 U7672 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        DATAI_17_), .C2(keyinput_g14), .A(n6765), .ZN(n6772) );
  AOI22_X1 U7673 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6766) );
  OAI221_X1 U7674 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6766), .ZN(n6771) );
  AOI22_X1 U7675 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(NA_N), .B2(
        keyinput_g33), .ZN(n6767) );
  OAI221_X1 U7676 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(NA_N), .C2(
        keyinput_g33), .A(n6767), .ZN(n6770) );
  AOI22_X1 U7677 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(REIP_REG_24__SCAN_IN), 
        .B2(keyinput_g58), .ZN(n6768) );
  OAI221_X1 U7678 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6768), .ZN(n6769) );
  NOR4_X1 U7679 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6805)
         );
  XNOR2_X1 U7680 ( .A(DATAI_20_), .B(keyinput_g11), .ZN(n6780) );
  AOI22_X1 U7681 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g49), .B1(
        n6774), .B2(keyinput_g17), .ZN(n6773) );
  OAI221_X1 U7682 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g49), .C1(
        n6774), .C2(keyinput_g17), .A(n6773), .ZN(n6779) );
  AOI22_X1 U7683 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(REIP_REG_31__SCAN_IN), 
        .B2(keyinput_g51), .ZN(n6775) );
  OAI221_X1 U7684 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_g51), .A(n6775), .ZN(n6778) );
  AOI22_X1 U7685 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(DATAI_28_), 
        .B2(keyinput_g3), .ZN(n6776) );
  OAI221_X1 U7686 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(DATAI_28_), 
        .C2(keyinput_g3), .A(n6776), .ZN(n6777) );
  NOR4_X1 U7687 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6804)
         );
  AOI22_X1 U7688 ( .A1(n4617), .A2(keyinput_g7), .B1(keyinput_g25), .B2(n6782), 
        .ZN(n6781) );
  OAI221_X1 U7689 ( .B1(n4617), .B2(keyinput_g7), .C1(n6782), .C2(keyinput_g25), .A(n6781), .ZN(n6793) );
  AOI22_X1 U7690 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_g39), .B1(DATAI_7_), .B2(keyinput_g24), .ZN(n6783) );
  OAI221_X1 U7691 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_7_), .C2(keyinput_g24), .A(n6783), .ZN(n6792) );
  AOI22_X1 U7692 ( .A1(n6786), .A2(keyinput_g28), .B1(n6785), .B2(keyinput_g57), .ZN(n6784) );
  OAI221_X1 U7693 ( .B1(n6786), .B2(keyinput_g28), .C1(n6785), .C2(
        keyinput_g57), .A(n6784), .ZN(n6791) );
  AOI22_X1 U7694 ( .A1(n6789), .A2(keyinput_g16), .B1(n6788), .B2(keyinput_g10), .ZN(n6787) );
  OAI221_X1 U7695 ( .B1(n6789), .B2(keyinput_g16), .C1(n6788), .C2(
        keyinput_g10), .A(n6787), .ZN(n6790) );
  NOR4_X1 U7696 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6803)
         );
  AOI22_X1 U7697 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6794) );
  OAI221_X1 U7698 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6794), .ZN(n6801) );
  AOI22_X1 U7699 ( .A1(DATAI_12_), .A2(keyinput_g19), .B1(DATAI_13_), .B2(
        keyinput_g18), .ZN(n6795) );
  OAI221_X1 U7700 ( .B1(DATAI_12_), .B2(keyinput_g19), .C1(DATAI_13_), .C2(
        keyinput_g18), .A(n6795), .ZN(n6800) );
  AOI22_X1 U7701 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_g40), .B1(DATAI_11_), 
        .B2(keyinput_g20), .ZN(n6796) );
  OAI221_X1 U7702 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .C1(DATAI_11_), 
        .C2(keyinput_g20), .A(n6796), .ZN(n6799) );
  AOI22_X1 U7703 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_g53), .ZN(n6797) );
  OAI221_X1 U7704 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_g53), .A(n6797), .ZN(n6798) );
  NOR4_X1 U7705 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6802)
         );
  NAND4_X1 U7706 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6806)
         );
  OAI22_X1 U7707 ( .A1(keyinput_g63), .A2(n6810), .B1(n6807), .B2(n6806), .ZN(
        n6808) );
  AOI211_X1 U7708 ( .C1(keyinput_g63), .C2(n6810), .A(n6809), .B(n6808), .ZN(
        n6814) );
  AOI22_X1 U7709 ( .A1(n6812), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6811), .ZN(n6813) );
  XNOR2_X1 U7710 ( .A(n6814), .B(n6813), .ZN(U3445) );
  AND2_X1 U3927 ( .A1(n4180), .A2(n4201), .ZN(n3035) );
  CLKBUF_X1 U34460 ( .A(n3150), .Z(n3875) );
  CLKBUF_X1 U34470 ( .A(n3298), .Z(n3016) );
  CLKBUF_X1 U3576 ( .A(n3269), .Z(n4190) );
  AND2_X1 U3584 ( .A1(n4391), .A2(n4009), .ZN(n3247) );
  CLKBUF_X1 U3925 ( .A(n5612), .Z(n3000) );
  CLKBUF_X1 U4191 ( .A(n5342), .Z(n2997) );
endmodule

