

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806;

  AOI21_X1 U11138 ( .B1(n10692), .B2(n16500), .A(n16499), .ZN(n16714) );
  XNOR2_X1 U11139 ( .A(n14904), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14974) );
  NOR2_X1 U11140 ( .A1(n16632), .A2(n16595), .ZN(n16610) );
  NOR2_X1 U11141 ( .A1(n9836), .A2(n21707), .ZN(n16557) );
  NAND2_X1 U11142 ( .A1(n16643), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16642) );
  OR3_X1 U11143 ( .A1(n16718), .A2(n10692), .A3(n16705), .ZN(n16693) );
  INV_X1 U11144 ( .A(n20625), .ZN(n20588) );
  INV_X1 U11145 ( .A(n17846), .ZN(n17857) );
  NOR2_X1 U11146 ( .A1(n12923), .A2(n12922), .ZN(n16298) );
  INV_X1 U11147 ( .A(n20124), .ZN(n20486) );
  AND2_X1 U11148 ( .A1(n10807), .A2(n10808), .ZN(n19892) );
  AND2_X1 U11149 ( .A1(n10807), .A2(n10806), .ZN(n19926) );
  CLKBUF_X2 U11150 ( .A(n13368), .Z(n13375) );
  NOR2_X1 U11151 ( .A1(n10803), .A2(n19802), .ZN(n10878) );
  INV_X2 U11152 ( .A(n10961), .ZN(n11177) );
  CLKBUF_X1 U11153 ( .A(n10810), .Z(n19802) );
  INV_X1 U11154 ( .A(n14388), .ZN(n18220) );
  INV_X2 U11155 ( .A(n13142), .ZN(n14395) );
  INV_X1 U11157 ( .A(n13087), .ZN(n11711) );
  AND2_X2 U11158 ( .A1(n12996), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11209) );
  INV_X2 U11159 ( .A(n18198), .ZN(n18174) );
  INV_X2 U11160 ( .A(n18186), .ZN(n18221) );
  INV_X1 U11161 ( .A(n13047), .ZN(n18198) );
  INV_X2 U11162 ( .A(n10848), .ZN(n12840) );
  INV_X1 U11163 ( .A(n12035), .ZN(n11812) );
  CLKBUF_X1 U11164 ( .A(n11698), .Z(n18153) );
  CLKBUF_X2 U11165 ( .A(n11913), .Z(n12596) );
  INV_X2 U11166 ( .A(n18200), .ZN(n18175) );
  BUF_X1 U11167 ( .A(n11937), .Z(n20800) );
  INV_X1 U11168 ( .A(n20776), .ZN(n14727) );
  AND2_X2 U11169 ( .A1(n11922), .A2(n13823), .ZN(n11926) );
  NOR2_X2 U11170 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U11171 ( .A1(n11609), .A2(n13884), .ZN(n18203) );
  OR2_X1 U11172 ( .A1(n11869), .A2(n11868), .ZN(n11931) );
  NAND4_X1 U11173 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11949) );
  AND4_X1 U11174 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11893) );
  NAND2_X1 U11175 ( .A1(n9748), .A2(n11858), .ZN(n11925) );
  CLKBUF_X1 U11176 ( .A(n21470), .Z(n9694) );
  NOR2_X1 U11177 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21470) );
  AND2_X2 U11178 ( .A1(n10228), .A2(n14181), .ZN(n12549) );
  AOI21_X1 U11179 ( .B1(n11912), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11882), .ZN(n11884) );
  NOR2_X1 U11180 ( .A1(n12222), .A2(n13344), .ZN(n12240) );
  NOR2_X1 U11181 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U11182 ( .A1(n10083), .A2(n10082), .ZN(n10003) );
  INV_X1 U11183 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10317) );
  AND2_X1 U11184 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  NOR3_X1 U11185 ( .A1(n16297), .A2(n16299), .A3(n16308), .ZN(n12926) );
  INV_X1 U11186 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14462) );
  INV_X1 U11187 ( .A(n18224), .ZN(n18180) );
  INV_X1 U11188 ( .A(n13676), .ZN(n14723) );
  INV_X2 U11190 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10715) );
  OR2_X1 U11191 ( .A1(n16902), .A2(n11474), .ZN(n16872) );
  AND2_X1 U11192 ( .A1(n10807), .A2(n10799), .ZN(n10865) );
  BUF_X1 U11193 ( .A(n10878), .Z(n20225) );
  INV_X1 U11194 ( .A(n11451), .ZN(n10101) );
  INV_X1 U11195 ( .A(n13086), .ZN(n13142) );
  INV_X1 U11196 ( .A(n18200), .ZN(n9697) );
  INV_X2 U11197 ( .A(n14359), .ZN(n18158) );
  BUF_X1 U11198 ( .A(n11949), .Z(n20792) );
  NOR2_X1 U11199 ( .A1(n17356), .A2(n15401), .ZN(n17340) );
  NOR2_X1 U11200 ( .A1(n13317), .A2(n12664), .ZN(n16565) );
  INV_X2 U11201 ( .A(n11124), .ZN(n11131) );
  AND2_X1 U11202 ( .A1(n10807), .A2(n10796), .ZN(n17033) );
  AND2_X1 U11203 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13906) );
  INV_X1 U11204 ( .A(n20818), .ZN(n14956) );
  NAND2_X2 U11205 ( .A1(n9881), .A2(n9879), .ZN(n14524) );
  INV_X1 U11206 ( .A(n15037), .ZN(n15049) );
  NOR2_X1 U11207 ( .A1(n9836), .A2(n16730), .ZN(n16526) );
  NAND2_X1 U11208 ( .A1(n14760), .A2(n14851), .ZN(n16596) );
  NOR2_X1 U11209 ( .A1(n16642), .A2(n11525), .ZN(n16633) );
  OAI21_X1 U11210 ( .B1(n20096), .B2(n20116), .A(n20298), .ZN(n20118) );
  INV_X1 U11212 ( .A(n18364), .ZN(n19065) );
  NAND2_X1 U11213 ( .A1(n10283), .A2(n13283), .ZN(n18489) );
  OR2_X1 U11214 ( .A1(n14712), .A2(n14711), .ZN(n14753) );
  NAND2_X1 U11215 ( .A1(n14038), .A2(n17277), .ZN(n20537) );
  AOI211_X1 U11216 ( .C1(n16415), .C2(BUF2_REG_28__SCAN_IN), .A(n16375), .B(
        n16374), .ZN(n16376) );
  NAND2_X1 U11217 ( .A1(n20251), .A2(n20123), .ZN(n20182) );
  INV_X2 U11218 ( .A(n14388), .ZN(n9707) );
  MUX2_X1 U11219 ( .A(n11032), .B(n10491), .S(n19834), .Z(n10911) );
  NOR2_X2 U11220 ( .A1(n18592), .A2(n18594), .ZN(n18566) );
  AND2_X2 U11221 ( .A1(n10444), .A2(n14462), .ZN(n9704) );
  BUF_X1 U11222 ( .A(n14070), .Z(n10100) );
  NAND2_X2 U11223 ( .A1(n11849), .A2(n11848), .ZN(n12266) );
  NAND2_X2 U11224 ( .A1(n11893), .A2(n11892), .ZN(n11940) );
  INV_X2 U11225 ( .A(n9942), .ZN(n9869) );
  AOI211_X2 U11226 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17553), .A(n17532), 
        .B(n17531), .ZN(n17533) );
  NOR2_X2 U11227 ( .A1(n13560), .A2(n13561), .ZN(n13559) );
  NAND2_X2 U11228 ( .A1(n18671), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17226) );
  NOR2_X2 U11229 ( .A1(n13537), .A2(n10162), .ZN(n18671) );
  AND2_X4 U11230 ( .A1(n11775), .A2(n13841), .ZN(n11887) );
  NOR2_X2 U11231 ( .A1(n16119), .A2(n16117), .ZN(n16108) );
  AND2_X4 U11232 ( .A1(n11781), .A2(n14182), .ZN(n12009) );
  NAND3_X2 U11233 ( .A1(n10834), .A2(n10425), .A3(n10833), .ZN(n10863) );
  AND4_X2 U11234 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10834) );
  INV_X2 U11235 ( .A(n10755), .ZN(n10132) );
  NOR2_X4 U11236 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14181) );
  NAND2_X2 U11237 ( .A1(n13203), .A2(n18734), .ZN(n18568) );
  XOR2_X2 U11238 ( .A(n14759), .B(n14758), .Z(n14857) );
  NAND2_X2 U11239 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  AOI211_X2 U11240 ( .C1(n17052), .C2(n19465), .A(n13532), .B(n13531), .ZN(
        n13533) );
  AND2_X4 U11241 ( .A1(n11047), .A2(n10344), .ZN(n12911) );
  INV_X2 U11242 ( .A(n11022), .ZN(n10734) );
  NAND2_X2 U11243 ( .A1(n10194), .A2(n10193), .ZN(n11022) );
  NOR2_X2 U11244 ( .A1(n15267), .A2(n15256), .ZN(n15255) );
  NOR2_X2 U11245 ( .A1(n17140), .A2(n13281), .ZN(n13537) );
  NOR2_X2 U11246 ( .A1(n17141), .A2(n18993), .ZN(n17140) );
  CLKBUF_X2 U11247 ( .A(n13336), .Z(n15514) );
  NOR2_X1 U11248 ( .A1(n16565), .A2(n9884), .ZN(n9883) );
  NOR2_X1 U11249 ( .A1(n16561), .A2(n16562), .ZN(n16560) );
  NAND2_X1 U11250 ( .A1(n10006), .A2(n12187), .ZN(n15583) );
  INV_X2 U11251 ( .A(n20582), .ZN(n15350) );
  NAND2_X1 U11252 ( .A1(n17318), .A2(n17317), .ZN(n17320) );
  NAND2_X1 U11253 ( .A1(n20251), .A2(n20250), .ZN(n20326) );
  NAND2_X1 U11254 ( .A1(n14630), .A2(n14629), .ZN(n14631) );
  NAND2_X1 U11255 ( .A1(n14069), .A2(n14068), .ZN(n14067) );
  NOR2_X1 U11256 ( .A1(n18286), .A2(n18415), .ZN(n18351) );
  BUF_X1 U11257 ( .A(n10867), .Z(n20186) );
  INV_X4 U11258 ( .A(n20714), .ZN(n15586) );
  NAND2_X1 U11259 ( .A1(n12276), .A2(n12275), .ZN(n20971) );
  CLKBUF_X1 U11260 ( .A(n10643), .Z(n10645) );
  NAND2_X1 U11261 ( .A1(n10655), .A2(n10959), .ZN(n10671) );
  AND2_X1 U11262 ( .A1(n9959), .A2(n18783), .ZN(n9958) );
  XNOR2_X1 U11263 ( .A(n13262), .B(n13261), .ZN(n18789) );
  INV_X2 U11264 ( .A(n11593), .ZN(n17820) );
  NAND2_X2 U11265 ( .A1(n10129), .A2(n10068), .ZN(n10757) );
  NAND2_X1 U11266 ( .A1(n11945), .A2(n20800), .ZN(n11948) );
  INV_X1 U11267 ( .A(n11926), .ZN(n15351) );
  NOR2_X1 U11268 ( .A1(n13742), .A2(n14956), .ZN(n13730) );
  NAND4_X1 U11269 ( .A1(n11958), .A2(n14146), .A3(n14143), .A4(n11926), .ZN(
        n13363) );
  CLKBUF_X3 U11270 ( .A(n13369), .Z(n14064) );
  CLKBUF_X2 U11271 ( .A(n11131), .Z(n11051) );
  INV_X1 U11272 ( .A(n14983), .ZN(n14979) );
  AND2_X1 U11273 ( .A1(n11923), .A2(n11931), .ZN(n11959) );
  CLKBUF_X1 U11274 ( .A(n11895), .Z(n20804) );
  BUF_X2 U11275 ( .A(n11936), .Z(n20776) );
  NAND2_X1 U11276 ( .A1(n13874), .A2(n11925), .ZN(n11942) );
  AND2_X1 U11277 ( .A1(n11895), .A2(n11931), .ZN(n11894) );
  INV_X2 U11278 ( .A(n11895), .ZN(n13874) );
  BUF_X1 U11279 ( .A(n11925), .Z(n20808) );
  INV_X2 U11280 ( .A(n11925), .ZN(n14143) );
  NAND4_X1 U11281 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11895) );
  NOR2_X1 U11282 ( .A1(n11780), .A2(n11779), .ZN(n11788) );
  AND4_X1 U11283 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n11849) );
  INV_X4 U11284 ( .A(n11711), .ZN(n18229) );
  CLKBUF_X2 U11285 ( .A(n11974), .Z(n13633) );
  CLKBUF_X2 U11286 ( .A(n12549), .Z(n11824) );
  INV_X2 U11287 ( .A(n18085), .ZN(n17897) );
  CLKBUF_X2 U11288 ( .A(n14776), .Z(n13615) );
  CLKBUF_X2 U11290 ( .A(n11906), .Z(n14774) );
  BUF_X2 U11291 ( .A(n12636), .Z(n14782) );
  BUF_X2 U11292 ( .A(n12010), .Z(n13632) );
  INV_X1 U11293 ( .A(n18186), .ZN(n13105) );
  AND2_X2 U11294 ( .A1(n11775), .A2(n13859), .ZN(n12636) );
  AND2_X2 U11295 ( .A1(n11782), .A2(n13859), .ZN(n11974) );
  INV_X4 U11296 ( .A(n13929), .ZN(n14359) );
  INV_X1 U11297 ( .A(n13041), .ZN(n9695) );
  BUF_X2 U11298 ( .A(n11896), .Z(n14775) );
  INV_X1 U11299 ( .A(n10391), .ZN(n9701) );
  CLKBUF_X2 U11300 ( .A(n11698), .Z(n18216) );
  AND2_X2 U11301 ( .A1(n13859), .A2(n14182), .ZN(n11907) );
  AND2_X2 U11302 ( .A1(n13859), .A2(n14181), .ZN(n11896) );
  NOR2_X4 U11303 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13859) );
  NOR2_X4 U11304 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10353) );
  NOR2_X4 U11305 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13884) );
  XNOR2_X1 U11306 ( .A(n13582), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14713) );
  NOR2_X1 U11307 ( .A1(n10388), .A2(n12671), .ZN(n12672) );
  AND2_X1 U11308 ( .A1(n10054), .A2(n16566), .ZN(n16767) );
  AOI21_X1 U11309 ( .B1(n14770), .B2(n9715), .A(n14769), .ZN(n14771) );
  AOI21_X1 U11310 ( .B1(n9883), .B2(n19781), .A(n14938), .ZN(n14939) );
  NOR2_X1 U11311 ( .A1(n16633), .A2(n9744), .ZN(n11515) );
  NAND2_X1 U11312 ( .A1(n9876), .A2(n9877), .ZN(n16566) );
  NAND2_X1 U11313 ( .A1(n15546), .A2(n9860), .ZN(n13336) );
  OAI21_X1 U11314 ( .B1(n14888), .B2(n14887), .A(n9773), .ZN(n14894) );
  AND2_X1 U11315 ( .A1(n15625), .A2(n15596), .ZN(n15615) );
  NOR2_X1 U11316 ( .A1(n15566), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15556) );
  NAND2_X1 U11317 ( .A1(n15158), .A2(n15157), .ZN(n15561) );
  AND2_X1 U11318 ( .A1(n15926), .A2(n15925), .ZN(n16699) );
  OR2_X1 U11319 ( .A1(n16647), .A2(n11501), .ZN(n16644) );
  NAND2_X1 U11320 ( .A1(n11553), .A2(n11554), .ZN(n16617) );
  AOI21_X1 U11321 ( .B1(n11365), .B2(n15926), .A(n14964), .ZN(n15908) );
  AND2_X1 U11322 ( .A1(n9848), .A2(n9847), .ZN(n10030) );
  AND2_X1 U11323 ( .A1(n16298), .A2(n16301), .ZN(n12925) );
  NOR2_X1 U11324 ( .A1(n9850), .A2(n16908), .ZN(n9849) );
  XNOR2_X1 U11325 ( .A(n12921), .B(n12903), .ZN(n16297) );
  NAND2_X1 U11326 ( .A1(n10332), .A2(n12884), .ZN(n12921) );
  AND2_X1 U11327 ( .A1(n15279), .A2(n12429), .ZN(n15264) );
  XNOR2_X1 U11328 ( .A(n14900), .B(n14899), .ZN(n15053) );
  NOR2_X1 U11329 ( .A1(n15485), .A2(n15486), .ZN(n15279) );
  NAND2_X1 U11330 ( .A1(n10940), .A2(n10406), .ZN(n16921) );
  XNOR2_X1 U11331 ( .A(n11101), .B(n10961), .ZN(n16657) );
  AOI21_X1 U11332 ( .B1(n18552), .B2(n18734), .A(n9796), .ZN(n9961) );
  NOR2_X2 U11333 ( .A1(n16040), .A2(n12659), .ZN(n16431) );
  CLKBUF_X1 U11334 ( .A(n14619), .Z(n14639) );
  AND2_X1 U11335 ( .A1(n17211), .A2(n13304), .ZN(n17087) );
  OR2_X1 U11336 ( .A1(n15657), .A2(n15592), .ZN(n15679) );
  AND2_X1 U11337 ( .A1(n18745), .A2(n18888), .ZN(n18601) );
  NAND2_X1 U11338 ( .A1(n20251), .A2(n20477), .ZN(n20249) );
  NAND2_X1 U11339 ( .A1(n11343), .A2(n10412), .ZN(n16040) );
  AND2_X1 U11340 ( .A1(n10239), .A2(n18830), .ZN(n9964) );
  NOR2_X2 U11341 ( .A1(n20292), .A2(n20125), .ZN(n20145) );
  INV_X1 U11342 ( .A(n20122), .ZN(n20251) );
  NOR2_X2 U11343 ( .A1(n20125), .A2(n20032), .ZN(n19880) );
  NOR2_X2 U11344 ( .A1(n20122), .A2(n20333), .ZN(n20389) );
  NAND2_X1 U11345 ( .A1(n20486), .A2(n20090), .ZN(n20292) );
  NAND2_X1 U11346 ( .A1(n9981), .A2(n12318), .ZN(n15490) );
  OR2_X1 U11347 ( .A1(n10900), .A2(n10899), .ZN(n10903) );
  AND2_X1 U11348 ( .A1(n13204), .A2(n13202), .ZN(n17129) );
  NAND2_X1 U11349 ( .A1(n12064), .A2(n10382), .ZN(n12302) );
  NAND4_X1 U11350 ( .A1(n10816), .A2(n10426), .A3(n10427), .A4(n10424), .ZN(
        n10053) );
  NAND2_X1 U11351 ( .A1(n13200), .A2(n18734), .ZN(n13204) );
  OAI21_X1 U11352 ( .B1(n14057), .B2(n14055), .A(n12695), .ZN(n14068) );
  OR2_X1 U11353 ( .A1(n18728), .A2(n9827), .ZN(n13200) );
  AND2_X1 U11354 ( .A1(n12680), .A2(n14157), .ZN(n14069) );
  NAND2_X1 U11355 ( .A1(n18360), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18359) );
  CLKBUF_X1 U11356 ( .A(n15905), .Z(n21065) );
  NOR3_X2 U11357 ( .A1(n14309), .A2(n11399), .A3(n10359), .ZN(n14617) );
  OAI21_X1 U11358 ( .B1(n12685), .B2(n12684), .A(n12695), .ZN(n14057) );
  INV_X1 U11359 ( .A(n14863), .ZN(n16884) );
  OR2_X1 U11360 ( .A1(n17139), .A2(n13197), .ZN(n18728) );
  AND2_X1 U11361 ( .A1(n10638), .A2(n10637), .ZN(n16073) );
  NAND2_X1 U11362 ( .A1(n10240), .A2(n13195), .ZN(n9967) );
  OR2_X1 U11363 ( .A1(n11504), .A2(n11505), .ZN(n14309) );
  AND2_X1 U11364 ( .A1(n16952), .A2(n11471), .ZN(n16936) );
  NAND2_X2 U11366 ( .A1(n16246), .A2(n10783), .ZN(n10868) );
  NAND2_X1 U11367 ( .A1(n16246), .A2(n10780), .ZN(n10867) );
  NAND2_X1 U11368 ( .A1(n14690), .A2(n14689), .ZN(n19501) );
  OAI21_X1 U11369 ( .B1(n10100), .B2(n14608), .A(n12676), .ZN(n12697) );
  AND2_X2 U11370 ( .A1(n14217), .A2(n19509), .ZN(n18282) );
  AND2_X1 U11371 ( .A1(n16966), .A2(n17401), .ZN(n10808) );
  OR2_X1 U11372 ( .A1(n16007), .A2(n16011), .ZN(n15992) );
  OAI22_X1 U11373 ( .A1(n19816), .A2(n19851), .B1(n19815), .B2(n19850), .ZN(
        n20341) );
  AND2_X1 U11374 ( .A1(n10646), .A2(n10648), .ZN(n16092) );
  AND2_X1 U11375 ( .A1(n14161), .A2(n14162), .ZN(n14160) );
  OAI22_X1 U11376 ( .A1(n19826), .A2(n19851), .B1(n16440), .B2(n19850), .ZN(
        n20360) );
  AND2_X2 U11377 ( .A1(n20537), .A2(n12252), .ZN(n20703) );
  NAND2_X2 U11378 ( .A1(n10791), .A2(n10795), .ZN(n16966) );
  AND2_X1 U11379 ( .A1(n19788), .A2(n10793), .ZN(n10799) );
  NAND2_X1 U11380 ( .A1(n12003), .A2(n12002), .ZN(n12026) );
  NOR2_X1 U11381 ( .A1(n10779), .A2(n10791), .ZN(n10806) );
  AND2_X2 U11382 ( .A1(n11070), .A2(n17047), .ZN(n11467) );
  OAI21_X1 U11383 ( .B1(n13155), .B2(n10246), .A(n13174), .ZN(n10242) );
  AND2_X1 U11384 ( .A1(n10364), .A2(n10363), .ZN(n10362) );
  OR2_X1 U11385 ( .A1(n13887), .A2(n13886), .ZN(n9990) );
  AND2_X2 U11386 ( .A1(n10781), .A2(n10792), .ZN(n19788) );
  OR2_X1 U11387 ( .A1(n17295), .A2(n20531), .ZN(n13359) );
  OR2_X2 U11388 ( .A1(n11968), .A2(n20894), .ZN(n20826) );
  NAND2_X1 U11389 ( .A1(n20894), .A2(n11968), .ZN(n12007) );
  OAI21_X1 U11390 ( .B1(n10155), .B2(n18789), .A(n10154), .ZN(n14108) );
  AND2_X1 U11391 ( .A1(n11382), .A2(n14207), .ZN(n10364) );
  NAND2_X1 U11392 ( .A1(n13285), .A2(n11728), .ZN(n13887) );
  XNOR2_X1 U11393 ( .A(n11366), .B(n9916), .ZN(n9871) );
  OR2_X1 U11394 ( .A1(n10778), .A2(n10777), .ZN(n10781) );
  NAND2_X1 U11395 ( .A1(n10021), .A2(n10016), .ZN(n20894) );
  NAND2_X2 U11396 ( .A1(n13190), .A2(n14692), .ZN(n18734) );
  OAI21_X1 U11397 ( .B1(n14134), .B2(n9960), .A(n9958), .ZN(n13135) );
  AND2_X1 U11398 ( .A1(n11972), .A2(n11970), .ZN(n11968) );
  OR2_X1 U11399 ( .A1(n17606), .A2(n17607), .ZN(n17604) );
  NOR2_X2 U11400 ( .A1(n16076), .A2(n16588), .ZN(n16075) );
  NOR2_X1 U11401 ( .A1(n10200), .A2(n10768), .ZN(n9940) );
  NOR2_X2 U11402 ( .A1(n11026), .A2(n11025), .ZN(n14605) );
  AOI21_X1 U11403 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10773), .ZN(n11366) );
  AND2_X1 U11404 ( .A1(n10764), .A2(n10763), .ZN(n10348) );
  NOR2_X1 U11405 ( .A1(n13891), .A2(n10282), .ZN(n13284) );
  AND2_X1 U11406 ( .A1(n10757), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10200) );
  OR2_X1 U11407 ( .A1(n14131), .A2(n13258), .ZN(n13262) );
  AND2_X1 U11408 ( .A1(n13228), .A2(n18489), .ZN(n13891) );
  AND2_X1 U11409 ( .A1(n9873), .A2(n9872), .ZN(n10045) );
  AND2_X1 U11410 ( .A1(n10055), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U11411 ( .A1(n10067), .A2(n14514), .ZN(n14476) );
  NAND2_X1 U11412 ( .A1(n13097), .A2(n13096), .ZN(n13112) );
  NAND2_X1 U11413 ( .A1(n9875), .A2(n9874), .ZN(n10732) );
  NAND2_X1 U11414 ( .A1(n10328), .A2(n13718), .ZN(n10069) );
  INV_X2 U11415 ( .A(n11140), .ZN(n14962) );
  INV_X1 U11416 ( .A(n11149), .ZN(n11335) );
  AND2_X1 U11417 ( .A1(n17114), .A2(n10085), .ZN(n11591) );
  NAND2_X1 U11418 ( .A1(n10327), .A2(n9770), .ZN(n13718) );
  NOR2_X1 U11419 ( .A1(n19055), .A2(n13231), .ZN(n14218) );
  NOR2_X1 U11420 ( .A1(n18539), .A2(n18542), .ZN(n17114) );
  AND3_X1 U11421 ( .A1(n10329), .A2(n10752), .A3(n20510), .ZN(n10327) );
  NAND2_X1 U11422 ( .A1(n11005), .A2(n14983), .ZN(n13726) );
  AND3_X1 U11423 ( .A1(n9996), .A2(n19846), .A3(n20511), .ZN(n9995) );
  NAND2_X1 U11424 ( .A1(n11939), .A2(n14064), .ZN(n13470) );
  NAND2_X1 U11425 ( .A1(n10393), .A2(n9750), .ZN(n14223) );
  OR2_X1 U11426 ( .A1(n13131), .A2(n13130), .ZN(n13259) );
  AND3_X1 U11427 ( .A1(n9699), .A2(n10734), .A3(n10336), .ZN(n10337) );
  AND2_X1 U11428 ( .A1(n10338), .A2(n14498), .ZN(n9854) );
  INV_X1 U11429 ( .A(n10738), .ZN(n10329) );
  NAND2_X1 U11430 ( .A1(n11131), .A2(n20510), .ZN(n11005) );
  NAND2_X1 U11431 ( .A1(n11130), .A2(n19839), .ZN(n11133) );
  NOR2_X1 U11432 ( .A1(n11131), .A2(n17044), .ZN(n10422) );
  INV_X1 U11433 ( .A(n11024), .ZN(n20511) );
  AND2_X1 U11434 ( .A1(n11615), .A2(n11614), .ZN(n19035) );
  OR2_X1 U11435 ( .A1(n11691), .A2(n11690), .ZN(n13230) );
  CLKBUF_X2 U11436 ( .A(n11340), .Z(n14961) );
  INV_X1 U11437 ( .A(n10606), .ZN(n10961) );
  INV_X2 U11438 ( .A(U212), .ZN(n17443) );
  CLKBUF_X1 U11439 ( .A(n11942), .Z(n13487) );
  AND4_X1 U11440 ( .A1(n13085), .A2(n13084), .A3(n13083), .A4(n13082), .ZN(
        n10393) );
  OR2_X1 U11441 ( .A1(n13111), .A2(n13110), .ZN(n13255) );
  OR2_X1 U11442 ( .A1(n13151), .A2(n13150), .ZN(n13250) );
  INV_X1 U11443 ( .A(n11130), .ZN(n9699) );
  AND2_X1 U11444 ( .A1(n14524), .A2(n11451), .ZN(n10338) );
  INV_X1 U11445 ( .A(n14498), .ZN(n20510) );
  NAND2_X1 U11446 ( .A1(n14498), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U11447 ( .A1(n11124), .A2(n14498), .ZN(n14983) );
  AND2_X1 U11448 ( .A1(n10741), .A2(n14524), .ZN(n11117) );
  CLKBUF_X1 U11449 ( .A(n10746), .Z(n14523) );
  INV_X2 U11450 ( .A(n11130), .ZN(n19834) );
  NAND4_X2 U11451 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n18364) );
  AND2_X1 U11452 ( .A1(n10860), .A2(n10392), .ZN(n11137) );
  CLKBUF_X2 U11453 ( .A(n11931), .Z(n20818) );
  CLKBUF_X1 U11454 ( .A(n12266), .Z(n20812) );
  AND2_X2 U11455 ( .A1(n11931), .A2(n12266), .ZN(n14146) );
  NAND2_X1 U11456 ( .A1(n9929), .A2(n9918), .ZN(n10746) );
  NAND2_X2 U11457 ( .A1(n10171), .A2(n10173), .ZN(n11130) );
  NAND2_X2 U11458 ( .A1(n10490), .A2(n10489), .ZN(n14498) );
  NAND2_X1 U11459 ( .A1(n10117), .A2(n10106), .ZN(n11451) );
  NAND4_X2 U11460 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11936) );
  OR2_X2 U11461 ( .A1(n11881), .A2(n11880), .ZN(n11937) );
  AND4_X1 U11462 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        n13073) );
  AND4_X1 U11463 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        n13074) );
  AND4_X1 U11464 ( .A1(n13063), .A2(n13062), .A3(n13061), .A4(n13060), .ZN(
        n13075) );
  NAND2_X1 U11465 ( .A1(n10174), .A2(n10715), .ZN(n10173) );
  AND4_X1 U11466 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11892) );
  AND4_X1 U11467 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11920) );
  AND4_X1 U11468 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n11848) );
  AOI21_X1 U11469 ( .B1(n11912), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11871), .ZN(n11874) );
  AND4_X1 U11470 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11810) );
  AND4_X1 U11471 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11808) );
  AND2_X1 U11472 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11882) );
  INV_X2 U11473 ( .A(n10420), .ZN(n9696) );
  INV_X2 U11474 ( .A(n13041), .ZN(n18222) );
  INV_X2 U11475 ( .A(n13068), .ZN(n14388) );
  AND2_X1 U11476 ( .A1(n12012), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11871) );
  AND2_X1 U11477 ( .A1(n11912), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11780) );
  BUF_X2 U11478 ( .A(n11912), .Z(n13610) );
  NAND2_X1 U11479 ( .A1(n11600), .A2(n11607), .ZN(n18085) );
  NAND2_X2 U11480 ( .A1(n11601), .A2(n13926), .ZN(n13041) );
  AND2_X2 U11481 ( .A1(n10228), .A2(n11775), .ZN(n11906) );
  BUF_X2 U11482 ( .A(n11698), .Z(n18058) );
  AND2_X2 U11483 ( .A1(n14181), .A2(n11781), .ZN(n14776) );
  BUF_X2 U11484 ( .A(n12012), .Z(n9698) );
  INV_X2 U11485 ( .A(n17478), .ZN(n17480) );
  OR2_X2 U11486 ( .A1(n12264), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20576) );
  AND2_X2 U11487 ( .A1(n10721), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10839) );
  AND2_X2 U11488 ( .A1(n11775), .A2(n11781), .ZN(n12010) );
  AND2_X2 U11489 ( .A1(n10072), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11775) );
  AND2_X1 U11490 ( .A1(n11598), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11608) );
  AND2_X1 U11491 ( .A1(n19488), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11606) );
  AND2_X1 U11492 ( .A1(n13888), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11600) );
  AND2_X2 U11493 ( .A1(n10353), .A2(n16991), .ZN(n10721) );
  AND2_X1 U11494 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11770), .ZN(
        n11782) );
  NOR3_X2 U11495 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17833) );
  INV_X1 U11496 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10072) );
  INV_X1 U11497 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11598) );
  AND2_X1 U11498 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11607) );
  INV_X1 U11499 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13888) );
  NAND2_X1 U11500 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13913) );
  AND2_X1 U11501 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10444) );
  AND2_X1 U11502 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11047) );
  INV_X1 U11503 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13907) );
  NOR2_X2 U11504 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11599) );
  AND2_X1 U11505 ( .A1(n13686), .A2(n15154), .ZN(n14951) );
  NOR2_X4 U11506 ( .A1(n15181), .A2(n10236), .ZN(n15154) );
  XNOR2_X2 U11507 ( .A(n13194), .B(n13192), .ZN(n14123) );
  AOI21_X1 U11508 ( .B1(n15028), .B2(n16146), .A(n15928), .ZN(n15920) );
  NOR2_X2 U11509 ( .A1(n16745), .A2(n11476), .ZN(n16719) );
  OR2_X2 U11510 ( .A1(n12327), .A2(n12329), .ZN(n12375) );
  NOR2_X2 U11511 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17611), .ZN(n17593) );
  AOI21_X2 U11512 ( .B1(n15667), .B2(n15595), .A(n15594), .ZN(n15625) );
  NAND2_X2 U11513 ( .A1(n15668), .A2(n15678), .ZN(n15667) );
  NOR2_X2 U11514 ( .A1(n14517), .A2(n14518), .ZN(n14516) );
  INV_X2 U11515 ( .A(n11130), .ZN(n9700) );
  INV_X2 U11516 ( .A(n10741), .ZN(n10739) );
  NOR2_X2 U11517 ( .A1(n13212), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17072) );
  AND2_X4 U11518 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10445) );
  OAI21_X2 U11519 ( .B1(n14069), .B2(n14068), .A(n14067), .ZN(n20124) );
  NAND2_X1 U11520 ( .A1(n11609), .A2(n13906), .ZN(n18200) );
  INV_X1 U11521 ( .A(n13080), .ZN(n9702) );
  INV_X1 U11522 ( .A(n10391), .ZN(n13080) );
  NAND2_X1 U11523 ( .A1(n13884), .A2(n11599), .ZN(n10391) );
  AND2_X1 U11524 ( .A1(n10444), .A2(n14462), .ZN(n9703) );
  AND2_X1 U11525 ( .A1(n10444), .A2(n14462), .ZN(n9705) );
  AND2_X1 U11526 ( .A1(n10444), .A2(n14462), .ZN(n9706) );
  AND2_X1 U11527 ( .A1(n11606), .A2(n13884), .ZN(n13068) );
  XNOR2_X1 U11528 ( .A(n13112), .B(n13113), .ZN(n14134) );
  NOR2_X2 U11529 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17585), .ZN(n17571) );
  AND2_X1 U11530 ( .A1(n10353), .A2(n16991), .ZN(n9710) );
  INV_X2 U11532 ( .A(n12858), .ZN(n9709) );
  AND2_X2 U11533 ( .A1(n14617), .A2(n14664), .ZN(n14663) );
  AND2_X1 U11534 ( .A1(n10353), .A2(n16991), .ZN(n9711) );
  NOR2_X2 U11535 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17563), .ZN(n17547) );
  AND2_X2 U11536 ( .A1(n13555), .A2(n15938), .ZN(n11540) );
  NOR2_X4 U11537 ( .A1(n13556), .A2(n13557), .ZN(n13555) );
  NOR2_X2 U11538 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17728), .ZN(n17727) );
  NOR2_X2 U11539 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17542), .ZN(n17525) );
  NOR2_X1 U11540 ( .A1(n11131), .A2(n11024), .ZN(n10376) );
  AND2_X1 U11541 ( .A1(n20510), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U11542 ( .A1(n10729), .A2(n10715), .ZN(n10193) );
  NAND2_X1 U11543 ( .A1(n10720), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10194) );
  NAND2_X1 U11544 ( .A1(n15583), .A2(n9719), .ZN(n10043) );
  OAI21_X1 U11545 ( .B1(n15583), .B2(n12192), .A(n9858), .ZN(n9860) );
  AND2_X1 U11546 ( .A1(n9859), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9858) );
  OR2_X1 U11547 ( .A1(n9713), .A2(n12192), .ZN(n9859) );
  AND2_X1 U11548 ( .A1(n11936), .A2(n11949), .ZN(n13369) );
  AND2_X2 U11549 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14182) );
  NAND2_X1 U11550 ( .A1(n10368), .A2(n10000), .ZN(n10002) );
  NOR2_X1 U11551 ( .A1(n9734), .A2(n10001), .ZN(n10000) );
  INV_X1 U11552 ( .A(n10366), .ZN(n10001) );
  NAND2_X1 U11553 ( .A1(n9854), .A2(n10337), .ZN(n10755) );
  NOR2_X1 U11554 ( .A1(n10284), .A2(n13231), .ZN(n11720) );
  OR2_X1 U11555 ( .A1(n13230), .A2(n13223), .ZN(n10284) );
  NOR2_X1 U11556 ( .A1(n19065), .A2(n19046), .ZN(n13283) );
  INV_X1 U11557 ( .A(n11023), .ZN(n11040) );
  AND2_X2 U11558 ( .A1(n11996), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10228) );
  NAND2_X1 U11559 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10109) );
  NAND2_X1 U11560 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10115) );
  NAND2_X1 U11561 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10126) );
  NAND2_X1 U11562 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n9927) );
  NAND2_X1 U11563 ( .A1(n12993), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n9921) );
  NAND2_X1 U11564 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n9938) );
  CLKBUF_X1 U11565 ( .A(n12011), .Z(n12548) );
  CLKBUF_X2 U11566 ( .A(n11901), .Z(n13609) );
  CLKBUF_X2 U11567 ( .A(n11907), .Z(n14783) );
  NAND2_X1 U11568 ( .A1(n12063), .A2(n12062), .ZN(n12086) );
  OR2_X1 U11569 ( .A1(n12222), .A2(n12061), .ZN(n12062) );
  XNOR2_X1 U11570 ( .A(n9974), .B(n9973), .ZN(n12025) );
  INV_X1 U11571 ( .A(n12024), .ZN(n9973) );
  NAND2_X1 U11572 ( .A1(n9975), .A2(n9757), .ZN(n9974) );
  OAI22_X1 U11573 ( .A1(n12222), .A2(n12023), .B1(n12094), .B2(n12034), .ZN(
        n12024) );
  NAND2_X1 U11574 ( .A1(n12114), .A2(n11993), .ZN(n11995) );
  NAND2_X1 U11575 ( .A1(n11935), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12000) );
  AND4_X1 U11576 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11809) );
  AND4_X1 U11577 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11807) );
  NOR2_X1 U11578 ( .A1(n12248), .A2(n12250), .ZN(n13486) );
  OR2_X1 U11579 ( .A1(n10592), .A2(n10591), .ZN(n10606) );
  AND2_X1 U11580 ( .A1(n10737), .A2(n9787), .ZN(n10044) );
  NAND2_X1 U11581 ( .A1(n10733), .A2(n11453), .ZN(n11455) );
  AND2_X1 U11582 ( .A1(n10730), .A2(n10734), .ZN(n9875) );
  OAI21_X1 U11583 ( .B1(n10753), .B2(n10329), .A(n9942), .ZN(n9874) );
  NOR2_X1 U11584 ( .A1(n10746), .A2(n10741), .ZN(n10336) );
  OAI21_X1 U11585 ( .B1(n12156), .B2(n12222), .A(n12155), .ZN(n12157) );
  NAND2_X1 U11586 ( .A1(n10011), .A2(n10008), .ZN(n10007) );
  NAND2_X1 U11587 ( .A1(n15688), .A2(n10012), .ZN(n10011) );
  NAND2_X1 U11588 ( .A1(n10014), .A2(n10013), .ZN(n10012) );
  INV_X1 U11589 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10013) );
  INV_X1 U11590 ( .A(n15689), .ZN(n10014) );
  AND2_X1 U11591 ( .A1(n9862), .A2(n12184), .ZN(n10084) );
  OAI21_X1 U11592 ( .B1(n15594), .B2(n12181), .A(n12183), .ZN(n9862) );
  AND2_X2 U11593 ( .A1(n12171), .A2(n12170), .ZN(n12190) );
  NAND2_X1 U11594 ( .A1(n17295), .A2(n9802), .ZN(n13356) );
  AND4_X1 U11595 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11790) );
  AND4_X1 U11596 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11787) );
  AND4_X1 U11597 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11789) );
  AND4_X1 U11598 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11858) );
  NAND2_X1 U11599 ( .A1(n9714), .A2(n10329), .ZN(n11035) );
  AND2_X1 U11600 ( .A1(n14991), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15015) );
  NAND2_X1 U11601 ( .A1(n10069), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10068) );
  AND2_X1 U11602 ( .A1(n13021), .A2(n10615), .ZN(n11530) );
  NOR2_X1 U11603 ( .A1(n16001), .A2(n10303), .ZN(n10302) );
  INV_X1 U11604 ( .A(n13033), .ZN(n10303) );
  INV_X1 U11605 ( .A(n12651), .ZN(n12654) );
  AND2_X1 U11606 ( .A1(n10370), .A2(n10955), .ZN(n10369) );
  AND2_X1 U11607 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  INV_X1 U11608 ( .A(n11465), .ZN(n11132) );
  INV_X1 U11609 ( .A(n14608), .ZN(n12691) );
  INV_X1 U11610 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19889) );
  NOR2_X1 U11611 ( .A1(n20509), .A2(n20513), .ZN(n14445) );
  NOR2_X1 U11612 ( .A1(n11722), .A2(n10285), .ZN(n11728) );
  NAND2_X1 U11613 ( .A1(n10287), .A2(n10286), .ZN(n10285) );
  INV_X1 U11614 ( .A(n11730), .ZN(n10287) );
  NOR2_X1 U11615 ( .A1(n11727), .A2(n13223), .ZN(n10286) );
  OR2_X1 U11616 ( .A1(n11729), .A2(n13909), .ZN(n14214) );
  AND2_X1 U11617 ( .A1(n18489), .A2(n13892), .ZN(n10282) );
  NOR2_X1 U11618 ( .A1(n13913), .A2(n19488), .ZN(n14675) );
  NAND2_X1 U11619 ( .A1(n11695), .A2(n9992), .ZN(n13231) );
  NOR2_X1 U11620 ( .A1(n9994), .A2(n9993), .ZN(n9992) );
  INV_X1 U11621 ( .A(n14064), .ZN(n13819) );
  NAND2_X1 U11622 ( .A1(n13400), .A2(n13375), .ZN(n13870) );
  NAND2_X1 U11623 ( .A1(n15130), .A2(n10223), .ZN(n15086) );
  NOR2_X1 U11624 ( .A1(n10226), .A2(n10224), .ZN(n10223) );
  INV_X1 U11625 ( .A(n13462), .ZN(n10224) );
  OR3_X1 U11626 ( .A1(n15103), .A2(n15112), .A3(n10227), .ZN(n10226) );
  AND2_X1 U11627 ( .A1(n13332), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13334) );
  CLKBUF_X1 U11628 ( .A(n12190), .Z(n12192) );
  NAND2_X1 U11629 ( .A1(n10483), .A2(n10715), .ZN(n10490) );
  NAND2_X1 U11630 ( .A1(n15042), .A2(n15041), .ZN(n19664) );
  OAI21_X1 U11631 ( .B1(n14605), .B2(n14490), .A(n13759), .ZN(n14521) );
  NOR2_X1 U11632 ( .A1(n15032), .A2(n20509), .ZN(n13935) );
  OR2_X1 U11633 ( .A1(n15023), .A2(n15956), .ZN(n15025) );
  AND2_X1 U11634 ( .A1(n13555), .A2(n10304), .ZN(n14964) );
  AND2_X1 U11635 ( .A1(n10307), .A2(n15938), .ZN(n10304) );
  NOR2_X1 U11636 ( .A1(n11365), .A2(n10308), .ZN(n10307) );
  AND2_X1 U11637 ( .A1(n10306), .A2(n15938), .ZN(n10305) );
  INV_X1 U11638 ( .A(n10308), .ZN(n10306) );
  NAND2_X1 U11639 ( .A1(n9972), .A2(n9971), .ZN(n16561) );
  AND2_X1 U11640 ( .A1(n12657), .A2(n13314), .ZN(n9971) );
  OAI21_X1 U11641 ( .B1(n16609), .B2(n11557), .A(n9772), .ZN(n9972) );
  NAND2_X1 U11642 ( .A1(n20517), .A2(n16978), .ZN(n16979) );
  OR2_X1 U11643 ( .A1(n11677), .A2(n11676), .ZN(n18286) );
  AND2_X1 U11644 ( .A1(n18601), .A2(n18798), .ZN(n17111) );
  NOR2_X1 U11645 ( .A1(n18660), .A2(n10164), .ZN(n10163) );
  NAND2_X1 U11646 ( .A1(n14493), .A2(n13721), .ZN(n15042) );
  OAI21_X1 U11647 ( .B1(n16795), .B2(n10037), .A(n10036), .ZN(n10035) );
  NAND2_X1 U11648 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10038), .ZN(
        n10037) );
  AOI21_X1 U11649 ( .B1(n16450), .B2(n19792), .A(n14847), .ZN(n10036) );
  OR2_X1 U11650 ( .A1(n18951), .A2(n9696), .ZN(n18998) );
  NAND2_X1 U11651 ( .A1(n19892), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10060) );
  AND2_X1 U11652 ( .A1(n12076), .A2(n12075), .ZN(n12078) );
  AND2_X2 U11653 ( .A1(n14181), .A2(n13841), .ZN(n11912) );
  AND2_X1 U11654 ( .A1(n9786), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U11655 ( .A1(n10018), .A2(n10230), .ZN(n10017) );
  NAND2_X1 U11656 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U11657 ( .A1(n9869), .A2(n9761), .ZN(n10761) );
  NAND2_X1 U11658 ( .A1(n12986), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n9896) );
  NAND2_X1 U11659 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9902) );
  NAND2_X1 U11660 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n9913) );
  AND2_X1 U11661 ( .A1(n11454), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10373) );
  OR2_X1 U11662 ( .A1(n12045), .A2(n12044), .ZN(n12088) );
  NAND2_X1 U11663 ( .A1(n12106), .A2(n12281), .ZN(n12114) );
  NAND2_X1 U11664 ( .A1(n10020), .A2(n9865), .ZN(n9864) );
  NOR2_X1 U11665 ( .A1(n12034), .A2(n9866), .ZN(n9865) );
  AND2_X1 U11666 ( .A1(n13366), .A2(n13363), .ZN(n11934) );
  INV_X1 U11667 ( .A(n12033), .ZN(n11992) );
  NAND3_X1 U11668 ( .A1(n20776), .A2(n20804), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12222) );
  NAND2_X1 U11669 ( .A1(n10070), .A2(n10883), .ZN(n10946) );
  OAI21_X1 U11670 ( .B1(n10755), .B2(n9853), .A(n9806), .ZN(n10343) );
  NAND2_X1 U11671 ( .A1(n10422), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U11672 ( .A1(n10532), .A2(n10531), .ZN(n10533) );
  INV_X1 U11673 ( .A(n14153), .ZN(n12943) );
  NAND2_X1 U11674 ( .A1(n10756), .A2(n9735), .ZN(n10318) );
  NAND2_X1 U11675 ( .A1(n10749), .A2(n10748), .ZN(n9833) );
  AOI21_X1 U11676 ( .B1(n11438), .B2(P2_EBX_REG_2__SCAN_IN), .A(n9808), .ZN(
        n10769) );
  NAND2_X1 U11677 ( .A1(n10774), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10198) );
  NAND2_X1 U11678 ( .A1(n12986), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10120) );
  NAND2_X1 U11679 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10121) );
  NAND2_X1 U11680 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10119) );
  NAND2_X1 U11681 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10122) );
  NAND2_X1 U11682 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10111) );
  NAND2_X1 U11683 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10108) );
  NAND2_X1 U11684 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10110) );
  NAND2_X1 U11685 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10116) );
  NAND2_X1 U11686 ( .A1(n9704), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10114) );
  NAND2_X1 U11687 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10113) );
  NAND2_X1 U11688 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10127) );
  NAND2_X1 U11689 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10125) );
  NAND2_X1 U11690 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10124) );
  NAND2_X1 U11691 ( .A1(n10787), .A2(n16246), .ZN(n10888) );
  INV_X1 U11692 ( .A(n14079), .ZN(n10246) );
  NOR2_X1 U11693 ( .A1(n10246), .A2(n14106), .ZN(n10244) );
  NAND2_X1 U11694 ( .A1(n13374), .A2(n13373), .ZN(n13378) );
  OR2_X1 U11695 ( .A1(n13470), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n13374) );
  OR3_X1 U11696 ( .A1(n13820), .A2(n21378), .A3(n13819), .ZN(n13821) );
  AND2_X1 U11697 ( .A1(n13672), .A2(n15094), .ZN(n15081) );
  AND2_X1 U11698 ( .A1(n12546), .A2(n10238), .ZN(n10237) );
  INV_X1 U11699 ( .A(n15182), .ZN(n10238) );
  INV_X1 U11700 ( .A(n15171), .ZN(n12546) );
  NAND2_X1 U11701 ( .A1(n10237), .A2(n15155), .ZN(n10236) );
  AND2_X1 U11702 ( .A1(n12479), .A2(n12461), .ZN(n10232) );
  INV_X1 U11703 ( .A(n15251), .ZN(n12461) );
  AND2_X1 U11704 ( .A1(n15479), .A2(n15330), .ZN(n9980) );
  INV_X1 U11705 ( .A(n12320), .ZN(n14797) );
  NAND2_X1 U11706 ( .A1(n21306), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12492) );
  NOR2_X1 U11707 ( .A1(n10222), .A2(n10221), .ZN(n10220) );
  INV_X1 U11708 ( .A(n15235), .ZN(n10221) );
  INV_X1 U11709 ( .A(n15215), .ZN(n10222) );
  INV_X1 U11710 ( .A(n15332), .ZN(n10217) );
  OR2_X1 U11711 ( .A1(n11823), .A2(n11822), .ZN(n12173) );
  AND2_X1 U11712 ( .A1(n10382), .A2(n12144), .ZN(n10042) );
  INV_X1 U11713 ( .A(n14171), .ZN(n10214) );
  NAND2_X1 U11714 ( .A1(n12309), .A2(n14029), .ZN(n9861) );
  NAND2_X1 U11715 ( .A1(n14064), .A2(n13375), .ZN(n13468) );
  AND2_X1 U11716 ( .A1(n13492), .A2(n13491), .ZN(n13499) );
  OR2_X1 U11717 ( .A1(n11985), .A2(n11984), .ZN(n12107) );
  NOR2_X1 U11718 ( .A1(n13343), .A2(n20776), .ZN(n13744) );
  NAND2_X1 U11719 ( .A1(n12032), .A2(n12031), .ZN(n20939) );
  OR2_X1 U11720 ( .A1(n20937), .A2(n20936), .ZN(n21039) );
  AND4_X1 U11721 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11921) );
  AND4_X1 U11722 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11919) );
  OAI21_X1 U11723 ( .B1(n21489), .B2(n17366), .A(n21454), .ZN(n20775) );
  AND2_X1 U11724 ( .A1(n10630), .A2(n9813), .ZN(n10623) );
  NOR2_X1 U11725 ( .A1(n10657), .A2(n10209), .ZN(n10208) );
  INV_X1 U11726 ( .A(n10631), .ZN(n10209) );
  OR2_X1 U11727 ( .A1(n10595), .A2(n9700), .ZN(n10959) );
  AND2_X1 U11728 ( .A1(n10904), .A2(n9782), .ZN(n10957) );
  AND2_X1 U11729 ( .A1(n10931), .A2(n10911), .ZN(n10540) );
  CLKBUF_X1 U11730 ( .A(n12911), .Z(n12989) );
  AND2_X1 U11731 ( .A1(n10334), .A2(n16336), .ZN(n10333) );
  NAND2_X1 U11732 ( .A1(n11261), .A2(n10315), .ZN(n10314) );
  INV_X1 U11733 ( .A(n14585), .ZN(n10315) );
  INV_X1 U11734 ( .A(n16006), .ZN(n10354) );
  AND2_X1 U11735 ( .A1(n10357), .A2(n10356), .ZN(n10355) );
  NOR2_X1 U11736 ( .A1(n10361), .A2(n14308), .ZN(n10360) );
  INV_X1 U11737 ( .A(n14549), .ZN(n10361) );
  INV_X1 U11738 ( .A(n14998), .ZN(n10281) );
  AND2_X1 U11739 ( .A1(n10539), .A2(n10538), .ZN(n10919) );
  AND2_X1 U11740 ( .A1(n13552), .A2(n10616), .ZN(n10979) );
  AND2_X1 U11741 ( .A1(n10414), .A2(n16430), .ZN(n10310) );
  OR2_X1 U11742 ( .A1(n16017), .A2(n10961), .ZN(n10663) );
  AND2_X1 U11743 ( .A1(n19677), .A2(n11177), .ZN(n10665) );
  NAND2_X1 U11744 ( .A1(n10057), .A2(n10056), .ZN(n11500) );
  OAI21_X1 U11745 ( .B1(n14861), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16667), .ZN(n10057) );
  AOI21_X1 U11746 ( .B1(n14861), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10058), .ZN(n10056) );
  INV_X1 U11747 ( .A(n10955), .ZN(n10058) );
  OR2_X1 U11748 ( .A1(n10573), .A2(n10572), .ZN(n11173) );
  NAND2_X1 U11749 ( .A1(n9945), .A2(n10771), .ZN(n10773) );
  NAND3_X1 U11750 ( .A1(n10417), .A2(n10474), .A3(n10409), .ZN(n11163) );
  AOI21_X1 U11751 ( .B1(n10839), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n10464), .ZN(n10474) );
  AND2_X1 U11752 ( .A1(n12943), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12684) );
  NOR2_X1 U11753 ( .A1(n11119), .A2(n11118), .ZN(n14467) );
  NAND2_X1 U11754 ( .A1(n12685), .A2(n12684), .ZN(n12695) );
  NAND2_X1 U11755 ( .A1(n10172), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10171) );
  OAI21_X1 U11756 ( .B1(n9935), .B2(n9930), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9929) );
  OAI21_X1 U11757 ( .B1(n9924), .B2(n9919), .A(n10715), .ZN(n9918) );
  NAND2_X1 U11758 ( .A1(n10813), .A2(n10802), .ZN(n10803) );
  INV_X1 U11759 ( .A(n19920), .ZN(n20184) );
  NOR2_X1 U11760 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14511) );
  INV_X1 U11761 ( .A(n10298), .ZN(n10296) );
  INV_X1 U11762 ( .A(n19466), .ZN(n10295) );
  NOR2_X1 U11763 ( .A1(n13252), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10148) );
  NAND2_X1 U11764 ( .A1(n14123), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10240) );
  AND2_X1 U11765 ( .A1(n9991), .A2(n9797), .ZN(n13285) );
  NAND2_X1 U11766 ( .A1(n11726), .A2(n11727), .ZN(n9991) );
  AND2_X1 U11767 ( .A1(n13225), .A2(n13224), .ZN(n13248) );
  INV_X1 U11768 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15204) );
  INV_X1 U11769 ( .A(n21485), .ZN(n15353) );
  NOR2_X1 U11770 ( .A1(n15353), .A2(n14727), .ZN(n14744) );
  AND2_X1 U11771 ( .A1(n15255), .A2(n9809), .ZN(n15161) );
  AND2_X1 U11772 ( .A1(n13875), .A2(n11958), .ZN(n14138) );
  NAND2_X1 U11773 ( .A1(n12262), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12564) );
  OR2_X1 U11774 ( .A1(n12564), .A2(n15549), .ZN(n12619) );
  AND2_X1 U11775 ( .A1(n13361), .A2(n11938), .ZN(n17277) );
  OR2_X1 U11776 ( .A1(n10186), .A2(n10185), .ZN(n14877) );
  NOR2_X1 U11777 ( .A1(n17334), .A2(n15706), .ZN(n10185) );
  NAND2_X1 U11778 ( .A1(n14822), .A2(n9771), .ZN(n13583) );
  INV_X1 U11779 ( .A(n13581), .ZN(n10029) );
  NAND2_X1 U11780 ( .A1(n13332), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13581) );
  OAI21_X1 U11781 ( .B1(n9863), .B2(n10009), .A(n10084), .ZN(n10006) );
  INV_X1 U11782 ( .A(n10011), .ZN(n9863) );
  NAND2_X1 U11783 ( .A1(n10026), .A2(n12154), .ZN(n10023) );
  INV_X1 U11784 ( .A(n12130), .ZN(n10027) );
  INV_X1 U11785 ( .A(n12152), .ZN(n10026) );
  XNOR2_X1 U11786 ( .A(n12129), .B(n17326), .ZN(n17317) );
  AND2_X1 U11787 ( .A1(n13499), .A2(n13498), .ZN(n13873) );
  OAI21_X1 U11788 ( .B1(n13359), .B2(n13358), .A(n10175), .ZN(n13502) );
  NAND2_X1 U11789 ( .A1(n13357), .A2(n14141), .ZN(n10175) );
  NAND2_X1 U11790 ( .A1(n12273), .A2(n12274), .ZN(n12276) );
  INV_X1 U11792 ( .A(n20531), .ZN(n14141) );
  INV_X1 U11793 ( .A(n21039), .ZN(n21034) );
  INV_X1 U11794 ( .A(n21461), .ZN(n21164) );
  INV_X1 U11795 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21677) );
  INV_X1 U11796 ( .A(n20974), .ZN(n21226) );
  NOR2_X1 U11797 ( .A1(n20946), .A2(n20945), .ZN(n21260) );
  CLKBUF_X1 U11798 ( .A(n13857), .Z(n13858) );
  INV_X1 U11799 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21302) );
  INV_X1 U11800 ( .A(n20996), .ZN(n21252) );
  AND2_X1 U11801 ( .A1(n21065), .A2(n12049), .ZN(n21311) );
  NAND2_X1 U11802 ( .A1(n21369), .A2(n20775), .ZN(n20945) );
  NAND2_X1 U11803 ( .A1(n10176), .A2(n12247), .ZN(n17295) );
  OAI21_X1 U11804 ( .B1(n12244), .B2(n12243), .A(n12245), .ZN(n10176) );
  OR2_X1 U11805 ( .A1(n13820), .A2(n11957), .ZN(n17288) );
  NAND2_X1 U11806 ( .A1(n10990), .A2(n10989), .ZN(n14889) );
  NAND2_X1 U11807 ( .A1(n14891), .A2(n10604), .ZN(n10608) );
  OAI211_X1 U11808 ( .C1(n10613), .C2(P2_EBX_REG_25__SCAN_IN), .A(n9700), .B(
        P2_EBX_REG_26__SCAN_IN), .ZN(n10604) );
  AND2_X1 U11809 ( .A1(n13321), .A2(n9826), .ZN(n14991) );
  AND2_X1 U11810 ( .A1(n10957), .A2(n16132), .ZN(n10672) );
  INV_X1 U11811 ( .A(n19671), .ZN(n16202) );
  INV_X1 U11812 ( .A(n16219), .ZN(n16273) );
  NAND2_X1 U11813 ( .A1(n14304), .A2(n10401), .ZN(n14619) );
  NAND2_X1 U11814 ( .A1(n13812), .A2(n11002), .ZN(n14153) );
  NAND2_X1 U11815 ( .A1(n14067), .A2(n10331), .ZN(n14154) );
  AND2_X1 U11816 ( .A1(n12698), .A2(n12696), .ZN(n10331) );
  NOR2_X1 U11817 ( .A1(n10323), .A2(n10321), .ZN(n10320) );
  INV_X1 U11818 ( .A(n10325), .ZN(n10323) );
  NOR2_X1 U11819 ( .A1(n10326), .A2(n16288), .ZN(n10325) );
  INV_X1 U11820 ( .A(n16281), .ZN(n10326) );
  NOR2_X1 U11821 ( .A1(n9767), .A2(n10312), .ZN(n10311) );
  NAND2_X1 U11822 ( .A1(n9880), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9879) );
  NAND2_X1 U11823 ( .A1(n9882), .A2(n10715), .ZN(n9881) );
  NOR2_X1 U11824 ( .A1(n15025), .A2(n15944), .ZN(n15024) );
  NAND2_X1 U11825 ( .A1(n15015), .A2(n9729), .ZN(n15021) );
  NAND2_X1 U11826 ( .A1(n9948), .A2(n11385), .ZN(n11386) );
  INV_X1 U11827 ( .A(n14545), .ZN(n10363) );
  INV_X1 U11828 ( .A(n10345), .ZN(n14895) );
  NAND2_X1 U11829 ( .A1(n11420), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U11830 ( .A1(n16479), .A2(n16477), .ZN(n14888) );
  OAI211_X1 U11831 ( .C1(n10002), .C2(n9999), .A(n9998), .B(n11532), .ZN(
        n11534) );
  OR2_X1 U11832 ( .A1(n10694), .A2(n9999), .ZN(n9998) );
  NAND2_X1 U11833 ( .A1(n9776), .A2(n11530), .ZN(n9999) );
  NAND2_X1 U11834 ( .A1(n10621), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13022) );
  NAND2_X1 U11835 ( .A1(n16643), .A2(n13014), .ZN(n16514) );
  INV_X1 U11836 ( .A(n10002), .ZN(n13017) );
  AND2_X1 U11837 ( .A1(n11354), .A2(n11353), .ZN(n16001) );
  NOR2_X1 U11838 ( .A1(n15999), .A2(n16001), .ZN(n16000) );
  NOR2_X1 U11839 ( .A1(n12664), .A2(n16758), .ZN(n9877) );
  OR2_X1 U11840 ( .A1(n16028), .A2(n10961), .ZN(n10666) );
  INV_X1 U11841 ( .A(n10140), .ZN(n10138) );
  OAI21_X1 U11842 ( .B1(n10144), .B2(n10141), .A(n13314), .ZN(n10140) );
  INV_X1 U11843 ( .A(n16543), .ZN(n10141) );
  NAND2_X1 U11844 ( .A1(n9807), .A2(n10146), .ZN(n10136) );
  NAND2_X1 U11845 ( .A1(n10143), .A2(n10142), .ZN(n16574) );
  OR2_X1 U11846 ( .A1(n10146), .A2(n16572), .ZN(n10142) );
  INV_X1 U11847 ( .A(n14527), .ZN(n14596) );
  AND3_X1 U11848 ( .A1(n11238), .A2(n11237), .A3(n11236), .ZN(n11519) );
  NAND2_X1 U11849 ( .A1(n10782), .A2(n10792), .ZN(n10791) );
  NOR2_X1 U11850 ( .A1(n14523), .A2(n17044), .ZN(n13812) );
  NAND2_X1 U11851 ( .A1(n12687), .A2(n12686), .ZN(n13814) );
  NAND2_X1 U11852 ( .A1(n19788), .A2(n12691), .ZN(n12687) );
  MUX2_X1 U11853 ( .A(n14986), .B(n14985), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n17002) );
  INV_X1 U11854 ( .A(n11005), .ZN(n13768) );
  NAND2_X1 U11855 ( .A1(n13764), .A2(n13763), .ZN(n14496) );
  NAND2_X1 U11856 ( .A1(n20124), .A2(n20090), .ZN(n20032) );
  AND2_X1 U11857 ( .A1(n20491), .A2(n20479), .ZN(n20065) );
  NOR2_X1 U11858 ( .A1(n21570), .A2(n20497), .ZN(n20288) );
  NAND2_X1 U11859 ( .A1(n20491), .A2(n19957), .ZN(n20257) );
  OR2_X1 U11860 ( .A1(n20124), .A2(n20090), .ZN(n20122) );
  NOR2_X1 U11861 ( .A1(n11024), .A2(n11040), .ZN(n11025) );
  AND2_X1 U11862 ( .A1(n11000), .A2(n10999), .ZN(n11042) );
  NAND2_X1 U11863 ( .A1(n17527), .A2(n11593), .ZN(n17511) );
  OAI21_X1 U11864 ( .B1(n17604), .B2(n18589), .A(n11593), .ZN(n10092) );
  NAND2_X1 U11865 ( .A1(n17604), .A2(n11593), .ZN(n17594) );
  NAND2_X1 U11866 ( .A1(n11593), .A2(n10095), .ZN(n10094) );
  NAND2_X1 U11867 ( .A1(n17667), .A2(n18590), .ZN(n10095) );
  OAI21_X1 U11868 ( .B1(n14214), .B2(n14213), .A(n14212), .ZN(n14322) );
  NAND2_X1 U11869 ( .A1(n9989), .A2(n9988), .ZN(n14216) );
  AND2_X1 U11870 ( .A1(n19469), .A2(n19627), .ZN(n9988) );
  NAND2_X1 U11871 ( .A1(n9990), .A2(n9818), .ZN(n9989) );
  INV_X1 U11872 ( .A(n19035), .ZN(n18428) );
  NAND2_X1 U11873 ( .A1(n19509), .A2(n19469), .ZN(n18488) );
  AND2_X1 U11874 ( .A1(n9726), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10085) );
  INV_X1 U11875 ( .A(n10148), .ZN(n10147) );
  NAND2_X1 U11876 ( .A1(n10152), .A2(n9762), .ZN(n14087) );
  OAI21_X1 U11877 ( .B1(n17175), .B2(n13253), .A(n14222), .ZN(n10152) );
  NAND2_X1 U11878 ( .A1(n13253), .A2(n10151), .ZN(n10150) );
  OR2_X1 U11879 ( .A1(n11628), .A2(n11627), .ZN(n18490) );
  OR2_X1 U11880 ( .A1(n18224), .A2(n18197), .ZN(n11619) );
  NAND2_X1 U11881 ( .A1(n10163), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10162) );
  NAND2_X1 U11882 ( .A1(n13198), .A2(n10248), .ZN(n10247) );
  OR2_X1 U11883 ( .A1(n13189), .A2(n13188), .ZN(n14692) );
  NAND2_X1 U11884 ( .A1(n10156), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10155) );
  INV_X1 U11885 ( .A(n14109), .ZN(n10156) );
  INV_X1 U11886 ( .A(n18490), .ZN(n19626) );
  INV_X1 U11887 ( .A(n13231), .ZN(n19058) );
  AND2_X1 U11888 ( .A1(n13702), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20771)
         );
  OR2_X1 U11889 ( .A1(n21370), .A2(n21369), .ZN(n20531) );
  NAND2_X1 U11890 ( .A1(n13480), .A2(n13479), .ZN(n13482) );
  AND2_X1 U11891 ( .A1(n20653), .A2(n14956), .ZN(n20648) );
  INV_X1 U11892 ( .A(n15631), .ZN(n15470) );
  OR2_X1 U11893 ( .A1(n14039), .A2(n20662), .ZN(n20675) );
  INV_X1 U11894 ( .A(n20683), .ZN(n14039) );
  INV_X2 U11895 ( .A(n14294), .ZN(n21497) );
  XNOR2_X1 U11896 ( .A(n14724), .B(n14812), .ZN(n15056) );
  OR2_X1 U11897 ( .A1(n14773), .A2(n15509), .ZN(n14724) );
  INV_X1 U11898 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15549) );
  INV_X1 U11899 ( .A(n20770), .ZN(n20709) );
  INV_X1 U11900 ( .A(n20757), .ZN(n17334) );
  INV_X1 U11901 ( .A(n15054), .ZN(n10180) );
  OAI21_X1 U11902 ( .B1(n15528), .B2(n10190), .A(n10188), .ZN(n15060) );
  XNOR2_X1 U11903 ( .A(n10403), .B(n13338), .ZN(n10190) );
  NAND2_X1 U11904 ( .A1(n15528), .A2(n10189), .ZN(n10188) );
  NOR2_X1 U11905 ( .A1(n14877), .A2(n10183), .ZN(n15697) );
  NAND2_X1 U11906 ( .A1(n10184), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10183) );
  NAND2_X1 U11907 ( .A1(n20757), .A2(n14881), .ZN(n10184) );
  NAND2_X1 U11908 ( .A1(n13507), .A2(n10177), .ZN(n15767) );
  NAND2_X1 U11909 ( .A1(n20757), .A2(n13506), .ZN(n10177) );
  INV_X1 U11910 ( .A(n20576), .ZN(n20718) );
  NAND2_X1 U11911 ( .A1(n12026), .A2(n12008), .ZN(n13843) );
  INV_X1 U11912 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17370) );
  INV_X1 U11913 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21369) );
  OR2_X1 U11914 ( .A1(n13719), .A2(n14514), .ZN(n15032) );
  NAND2_X1 U11915 ( .A1(n15916), .A2(n10269), .ZN(n10268) );
  INV_X1 U11916 ( .A(n10270), .ZN(n10269) );
  OAI21_X1 U11917 ( .B1(n15917), .B2(n16254), .A(n10271), .ZN(n10270) );
  OAI21_X1 U11918 ( .B1(n16697), .B2(n16254), .A(n9839), .ZN(n9838) );
  AOI21_X1 U11919 ( .B1(n15923), .B2(n19676), .A(n9840), .ZN(n9839) );
  NAND2_X1 U11920 ( .A1(n15921), .A2(n15922), .ZN(n9840) );
  XNOR2_X1 U11921 ( .A(n15920), .B(n16482), .ZN(n9842) );
  AND2_X1 U11922 ( .A1(n17002), .A2(n19681), .ZN(n19669) );
  AND2_X1 U11923 ( .A1(n15049), .A2(n15048), .ZN(n19674) );
  INV_X1 U11924 ( .A(n20090), .ZN(n19858) );
  AOI21_X1 U11925 ( .B1(n13576), .B2(n19787), .A(n13575), .ZN(n13577) );
  NAND2_X1 U11926 ( .A1(n10139), .A2(n10144), .ZN(n13316) );
  NAND2_X1 U11927 ( .A1(n10134), .A2(n10133), .ZN(n10139) );
  NAND2_X1 U11928 ( .A1(n9856), .A2(n16776), .ZN(n9855) );
  AND2_X1 U11929 ( .A1(n17388), .A2(n16984), .ZN(n19787) );
  NAND2_X1 U11930 ( .A1(n16514), .A2(n10607), .ZN(n10104) );
  NAND2_X1 U11931 ( .A1(n16717), .A2(n10607), .ZN(n10105) );
  NAND2_X1 U11932 ( .A1(n9836), .A2(n21707), .ZN(n16753) );
  INV_X1 U11933 ( .A(n16785), .ZN(n9852) );
  NAND2_X1 U11934 ( .A1(n10039), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16795) );
  OAI21_X1 U11935 ( .B1(n16596), .B2(n16942), .A(n14846), .ZN(n10039) );
  OAI21_X1 U11936 ( .B1(n10052), .B2(n10049), .A(n10046), .ZN(n16792) );
  INV_X1 U11937 ( .A(n14849), .ZN(n10049) );
  AND2_X1 U11938 ( .A1(n14853), .A2(n10047), .ZN(n10046) );
  NAND2_X1 U11939 ( .A1(n14849), .A2(n10048), .ZN(n10047) );
  AOI21_X1 U11940 ( .B1(n16643), .B2(n10201), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16611) );
  NOR2_X1 U11941 ( .A1(n10204), .A2(n10203), .ZN(n10201) );
  OR2_X1 U11942 ( .A1(n11516), .A2(n17400), .ZN(n11529) );
  INV_X1 U11943 ( .A(n19792), .ZN(n16958) );
  INV_X1 U11944 ( .A(n19803), .ZN(n16967) );
  NOR2_X2 U11945 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20484) );
  OR2_X1 U11946 ( .A1(n20298), .A2(n16982), .ZN(n20495) );
  NAND2_X1 U11947 ( .A1(n15031), .A2(n15030), .ZN(n17049) );
  NOR2_X1 U11948 ( .A1(n19468), .A2(n18488), .ZN(n19642) );
  NAND2_X1 U11949 ( .A1(n19642), .A2(n18428), .ZN(n19640) );
  INV_X1 U11950 ( .A(n19642), .ZN(n19638) );
  NAND2_X1 U11951 ( .A1(n19501), .A2(n19509), .ZN(n17488) );
  AND2_X1 U11952 ( .A1(n17512), .A2(n11593), .ZN(n17503) );
  XNOR2_X1 U11953 ( .A(n17503), .B(n10091), .ZN(n10090) );
  INV_X1 U11954 ( .A(n17504), .ZN(n10091) );
  INV_X1 U11955 ( .A(n17829), .ZN(n17864) );
  NAND2_X1 U11956 ( .A1(n18300), .A2(n9982), .ZN(n9987) );
  NOR2_X1 U11957 ( .A1(n18431), .A2(n9985), .ZN(n9982) );
  NAND2_X1 U11958 ( .A1(n18300), .A2(n9983), .ZN(n18287) );
  AND2_X1 U11959 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n9984), .ZN(n9983) );
  NOR2_X1 U11960 ( .A1(n21561), .A2(n9985), .ZN(n9984) );
  AND4_X1 U11961 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11648) );
  AND4_X1 U11962 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11646) );
  AND4_X1 U11963 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n11649) );
  NAND2_X2 U11964 ( .A1(n18282), .A2(n18364), .ZN(n18415) );
  NAND2_X1 U11965 ( .A1(n14218), .A2(n18282), .ZN(n18421) );
  AND2_X1 U11966 ( .A1(n17111), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14697) );
  NAND2_X1 U11967 ( .A1(n10293), .A2(n10291), .ZN(n10290) );
  INV_X1 U11968 ( .A(n10292), .ZN(n10291) );
  NAND2_X1 U11969 ( .A1(n17107), .A2(n17106), .ZN(n10293) );
  OAI21_X1 U11970 ( .B1(n18696), .B2(n17109), .A(n17108), .ZN(n10292) );
  OR2_X1 U11971 ( .A1(n18786), .A2(n14692), .ZN(n18700) );
  NOR2_X2 U11972 ( .A1(n18786), .A2(n18405), .ZN(n18760) );
  INV_X1 U11973 ( .A(n18760), .ZN(n18748) );
  OR2_X1 U11974 ( .A1(n17488), .A2(n18490), .ZN(n18701) );
  INV_X1 U11975 ( .A(n17051), .ZN(n10159) );
  AOI21_X1 U11976 ( .B1(n17087), .B2(n19015), .A(n13297), .ZN(n17204) );
  AND2_X1 U11977 ( .A1(n17219), .A2(n17218), .ZN(n18804) );
  AND2_X1 U11978 ( .A1(n10297), .A2(n10298), .ZN(n19465) );
  AND2_X1 U11979 ( .A1(n17252), .A2(n14692), .ZN(n19002) );
  INV_X1 U11980 ( .A(n18998), .ZN(n19008) );
  AND2_X1 U11981 ( .A1(n13245), .A2(n19509), .ZN(n18951) );
  INV_X1 U11982 ( .A(n20771), .ZN(n20769) );
  INV_X1 U11983 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21567) );
  INV_X1 U11984 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21549) );
  INV_X1 U11985 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21789) );
  INV_X1 U11986 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21445) );
  NAND2_X1 U11987 ( .A1(n11894), .A2(n12282), .ZN(n10082) );
  NAND2_X1 U11988 ( .A1(n12102), .A2(n14146), .ZN(n10083) );
  NAND2_X1 U11989 ( .A1(n20933), .A2(n12025), .ZN(n12082) );
  AND2_X1 U11990 ( .A1(n12205), .A2(n12204), .ZN(n12214) );
  NAND2_X1 U11991 ( .A1(n11938), .A2(n12282), .ZN(n11943) );
  NAND2_X1 U11992 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  NAND2_X1 U11993 ( .A1(n17033), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10061) );
  INV_X1 U11994 ( .A(n11086), .ZN(n10885) );
  NAND2_X1 U11995 ( .A1(n9700), .A2(n19839), .ZN(n10750) );
  AOI22_X1 U11996 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10719) );
  AND2_X1 U11997 ( .A1(n12231), .A2(n12230), .ZN(n12233) );
  AND2_X1 U11998 ( .A1(n12195), .A2(n12194), .ZN(n12218) );
  AND2_X1 U11999 ( .A1(n12142), .A2(n12141), .ZN(n12143) );
  INV_X1 U12000 ( .A(n12087), .ZN(n12064) );
  AND2_X1 U12001 ( .A1(n12077), .A2(n12086), .ZN(n10382) );
  INV_X1 U12002 ( .A(n12078), .ZN(n12077) );
  OR2_X1 U12003 ( .A1(n12074), .A2(n12073), .ZN(n12159) );
  INV_X1 U12004 ( .A(n12086), .ZN(n10005) );
  OR2_X1 U12005 ( .A1(n12060), .A2(n12059), .ZN(n12090) );
  CLKBUF_X1 U12006 ( .A(n12011), .Z(n11817) );
  INV_X1 U12007 ( .A(n12107), .ZN(n12101) );
  OAI21_X1 U12008 ( .B1(n13857), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11969), 
        .ZN(n12099) );
  INV_X1 U12009 ( .A(n10017), .ZN(n9976) );
  AND2_X1 U12010 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11838) );
  AOI22_X1 U12011 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10166) );
  AND2_X1 U12012 ( .A1(n12012), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11861) );
  AOI22_X1 U12013 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11896), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11866) );
  AOI21_X1 U12014 ( .B1(n14175), .B2(n21369), .A(n12048), .ZN(n20773) );
  INV_X1 U12015 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U12016 ( .A1(n10381), .A2(n10022), .ZN(n10021) );
  OR2_X1 U12017 ( .A1(n20804), .A2(n21369), .ZN(n12033) );
  AOI21_X1 U12018 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21474), .A(
        n12233), .ZN(n12228) );
  INV_X1 U12019 ( .A(n12222), .ZN(n12234) );
  INV_X1 U12020 ( .A(n13350), .ZN(n12226) );
  XNOR2_X1 U12021 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U12022 ( .A1(n9704), .A2(n10715), .ZN(n10848) );
  NOR2_X1 U12023 ( .A1(n12885), .A2(n10335), .ZN(n10334) );
  INV_X1 U12024 ( .A(n12826), .ZN(n10335) );
  NAND2_X1 U12025 ( .A1(n19834), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10517) );
  NOR2_X1 U12026 ( .A1(n10753), .A2(n17044), .ZN(n9885) );
  NAND2_X1 U12027 ( .A1(n10132), .A2(n9760), .ZN(n10131) );
  AND2_X1 U12028 ( .A1(n10371), .A2(n16635), .ZN(n10370) );
  AND2_X1 U12029 ( .A1(n16655), .A2(n11103), .ZN(n9969) );
  AND2_X1 U12030 ( .A1(n9868), .A2(n9867), .ZN(n10814) );
  AND2_X1 U12031 ( .A1(n10495), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10464) );
  OR2_X1 U12032 ( .A1(n10856), .A2(n10855), .ZN(n10857) );
  OAI22_X1 U12033 ( .A1(n9736), .A2(n10854), .B1(n19971), .B2(n10853), .ZN(
        n10855) );
  NAND2_X1 U12034 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n9908) );
  NAND2_X1 U12035 ( .A1(n12986), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n9907) );
  NAND2_X1 U12036 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n9906) );
  NAND2_X1 U12037 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9898) );
  NAND2_X1 U12038 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9895) );
  NAND2_X1 U12039 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9897) );
  NAND2_X1 U12040 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9900) );
  NAND2_X1 U12041 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9903) );
  NAND2_X1 U12042 ( .A1(n9703), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n9901) );
  NAND2_X1 U12043 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n9911) );
  NAND2_X1 U12044 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n9914) );
  NAND2_X1 U12045 ( .A1(n10774), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10749) );
  NAND2_X1 U12046 ( .A1(n10757), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10756) );
  AND2_X1 U12047 ( .A1(n10372), .A2(n9817), .ZN(n10375) );
  AND2_X1 U12048 ( .A1(n10422), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U12049 ( .A1(n12986), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n9932) );
  NAND2_X1 U12050 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n9933) );
  NAND2_X1 U12051 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n9931) );
  NAND2_X1 U12052 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n9934) );
  NAND2_X1 U12053 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n9928) );
  NAND2_X1 U12054 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12055 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n9925) );
  NAND2_X1 U12056 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n9923) );
  NAND2_X1 U12057 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n9920) );
  NAND2_X1 U12058 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n9922) );
  NAND2_X1 U12059 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n9939) );
  NAND2_X1 U12060 ( .A1(n9703), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n9937) );
  NAND2_X1 U12061 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n9936) );
  AOI22_X1 U12062 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10698) );
  AND2_X1 U12063 ( .A1(n11599), .A2(n13906), .ZN(n11698) );
  NAND2_X1 U12064 ( .A1(n18286), .A2(n13231), .ZN(n11722) );
  AND2_X1 U12065 ( .A1(n15081), .A2(n15083), .ZN(n13684) );
  AND2_X1 U12066 ( .A1(n13671), .A2(n13670), .ZN(n15094) );
  NAND2_X1 U12067 ( .A1(n13860), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13666) );
  NOR2_X1 U12068 ( .A1(n12022), .A2(n12021), .ZN(n12094) );
  AND2_X1 U12069 ( .A1(n14146), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12297) );
  INV_X1 U12070 ( .A(n15084), .ZN(n10227) );
  NOR2_X1 U12071 ( .A1(n10219), .A2(n13443), .ZN(n10218) );
  INV_X1 U12072 ( .A(n10220), .ZN(n10219) );
  NAND2_X1 U12073 ( .A1(n15689), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10010) );
  INV_X1 U12074 ( .A(n15644), .ZN(n10040) );
  OAI21_X1 U12075 ( .B1(n12126), .B2(n12123), .A(n10076), .ZN(n10079) );
  INV_X1 U12076 ( .A(n10077), .ZN(n10076) );
  OAI21_X1 U12077 ( .B1(n12124), .B2(n12123), .A(n20716), .ZN(n10077) );
  NAND2_X1 U12078 ( .A1(n9861), .A2(n10074), .ZN(n10073) );
  AND2_X1 U12079 ( .A1(n12093), .A2(n20716), .ZN(n10074) );
  OR2_X1 U12080 ( .A1(n14030), .A2(n20767), .ZN(n12117) );
  NAND2_X1 U12081 ( .A1(n12126), .A2(n12124), .ZN(n14574) );
  NAND2_X1 U12082 ( .A1(n20792), .A2(n20808), .ZN(n13344) );
  NAND2_X1 U12083 ( .A1(n11935), .A2(n9804), .ZN(n10229) );
  OAI211_X1 U12084 ( .C1(n12222), .C2(n11991), .A(n11990), .B(n11989), .ZN(
        n12281) );
  INV_X1 U12085 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11991) );
  INV_X1 U12086 ( .A(n12025), .ZN(n20935) );
  XNOR2_X1 U12087 ( .A(n12026), .B(n20939), .ZN(n14175) );
  AND2_X1 U12088 ( .A1(n13347), .A2(n13494), .ZN(n13828) );
  NAND2_X1 U12089 ( .A1(n20826), .A2(n12007), .ZN(n13857) );
  NAND2_X1 U12090 ( .A1(n12034), .A2(n12033), .ZN(n12246) );
  XNOR2_X1 U12091 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11001) );
  AND2_X1 U12092 ( .A1(n11019), .A2(n11018), .ZN(n11023) );
  OR2_X1 U12093 ( .A1(n11017), .A2(n11016), .ZN(n11019) );
  NAND2_X1 U12094 ( .A1(n10690), .A2(n10959), .ZN(n10687) );
  NOR2_X1 U12095 ( .A1(n15981), .A2(n16519), .ZN(n15968) );
  NOR2_X1 U12096 ( .A1(n16096), .A2(n16098), .ZN(n16085) );
  NAND2_X1 U12097 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10266) );
  INV_X1 U12098 ( .A(n10951), .ZN(n10594) );
  MUX2_X1 U12099 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n10882), .S(n10980), .Z(
        n10941) );
  INV_X1 U12100 ( .A(n12832), .ZN(n11284) );
  INV_X1 U12101 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10443) );
  INV_X1 U12102 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10442) );
  AND2_X1 U12103 ( .A1(n12866), .A2(n12865), .ZN(n16312) );
  NAND2_X1 U12104 ( .A1(n10313), .A2(n11315), .ZN(n10312) );
  INV_X1 U12105 ( .A(n10314), .ZN(n10313) );
  NAND2_X1 U12106 ( .A1(n9869), .A2(n19846), .ZN(n11453) );
  NOR2_X1 U12107 ( .A1(n16530), .A2(n10277), .ZN(n10276) );
  NAND2_X1 U12108 ( .A1(n15015), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15018) );
  AND2_X1 U12109 ( .A1(n11412), .A2(n14762), .ZN(n10357) );
  AND2_X1 U12110 ( .A1(n14663), .A2(n14762), .ZN(n12666) );
  NAND2_X1 U12111 ( .A1(n15011), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15010) );
  NAND2_X1 U12112 ( .A1(n10265), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10264) );
  INV_X1 U12113 ( .A(n10266), .ZN(n10265) );
  NAND2_X1 U12114 ( .A1(n16926), .A2(n16937), .ZN(n9832) );
  NAND2_X1 U12115 ( .A1(n10309), .A2(n11541), .ZN(n10308) );
  INV_X1 U12116 ( .A(n15924), .ZN(n10309) );
  AOI22_X1 U12117 ( .A1(n10694), .A2(n9734), .B1(n10693), .B2(n10692), .ZN(
        n10978) );
  OR2_X1 U12118 ( .A1(n16014), .A2(n10961), .ZN(n10686) );
  NAND2_X1 U12119 ( .A1(n10685), .A2(n10684), .ZN(n16540) );
  INV_X1 U12120 ( .A(n11561), .ZN(n10685) );
  NOR2_X1 U12121 ( .A1(n16562), .A2(n10683), .ZN(n10684) );
  AND2_X1 U12122 ( .A1(n11345), .A2(n11344), .ZN(n12659) );
  AND2_X1 U12123 ( .A1(n16773), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12662) );
  NAND2_X1 U12124 ( .A1(n10360), .A2(n14648), .ZN(n10359) );
  AND2_X1 U12125 ( .A1(n16103), .A2(n11177), .ZN(n10668) );
  AND2_X1 U12126 ( .A1(n10668), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16542) );
  NAND2_X1 U12127 ( .A1(n10370), .A2(n10367), .ZN(n10366) );
  INV_X1 U12128 ( .A(n10974), .ZN(n10367) );
  AND2_X1 U12129 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16813) );
  OR2_X1 U12130 ( .A1(n16133), .A2(n10972), .ZN(n11497) );
  AND2_X1 U12131 ( .A1(n14160), .A2(n14207), .ZN(n14316) );
  OR2_X1 U12132 ( .A1(n10557), .A2(n10556), .ZN(n11169) );
  OR2_X1 U12133 ( .A1(n10451), .A2(n10450), .ZN(n11159) );
  INV_X1 U12134 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16928) );
  NAND2_X1 U12135 ( .A1(n11438), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10349) );
  NAND3_X1 U12136 ( .A1(n10342), .A2(n10340), .A3(n10766), .ZN(n10778) );
  NAND2_X1 U12137 ( .A1(n10346), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10340) );
  NOR2_X1 U12138 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  AND2_X1 U12139 ( .A1(n14467), .A2(n11466), .ZN(n13756) );
  AND2_X1 U12140 ( .A1(n11051), .A2(n10861), .ZN(n17396) );
  OR2_X1 U12141 ( .A1(n14153), .A2(n19824), .ZN(n12692) );
  AND2_X1 U12142 ( .A1(n11053), .A2(n14524), .ZN(n10742) );
  NAND2_X1 U12143 ( .A1(n10195), .A2(n10199), .ZN(n10032) );
  NAND2_X1 U12144 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  NAND2_X1 U12145 ( .A1(n9944), .A2(n10732), .ZN(n11457) );
  AND2_X1 U12146 ( .A1(n10731), .A2(n20510), .ZN(n9944) );
  OR2_X1 U12147 ( .A1(n14153), .A2(n19829), .ZN(n12678) );
  CLKBUF_X1 U12148 ( .A(n11047), .Z(n14475) );
  AND3_X1 U12149 ( .A1(n11063), .A2(n11062), .A3(n11061), .ZN(n13760) );
  OAI21_X1 U12150 ( .B1(n10123), .B2(n10118), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10117) );
  OAI21_X1 U12151 ( .B1(n10112), .B2(n10107), .A(n10715), .ZN(n10106) );
  NAND2_X1 U12152 ( .A1(n20476), .A2(n20298), .ZN(n17028) );
  AND2_X1 U12153 ( .A1(n11576), .A2(n10097), .ZN(n10096) );
  INV_X1 U12154 ( .A(n18652), .ZN(n10097) );
  INV_X1 U12155 ( .A(n18651), .ZN(n11576) );
  AND2_X1 U12156 ( .A1(n18754), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18720) );
  NAND2_X1 U12157 ( .A1(n14223), .A2(n13249), .ZN(n13254) );
  NAND2_X1 U12158 ( .A1(n13310), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10257) );
  NAND2_X1 U12159 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10256) );
  NOR2_X1 U12160 ( .A1(n21581), .A2(n17192), .ZN(n10255) );
  INV_X1 U12161 ( .A(n10242), .ZN(n10241) );
  NAND2_X1 U12162 ( .A1(n11728), .A2(n13230), .ZN(n13228) );
  NOR3_X1 U12163 ( .A1(n13291), .A2(n13290), .A3(n13910), .ZN(n13890) );
  OR2_X1 U12164 ( .A1(n18224), .A2(n11594), .ZN(n11595) );
  OR2_X1 U12165 ( .A1(n11662), .A2(n11661), .ZN(n11727) );
  OR2_X1 U12166 ( .A1(n11717), .A2(n11716), .ZN(n13223) );
  AOI21_X1 U12167 ( .B1(n19020), .B2(n14680), .A(n19506), .ZN(n19032) );
  NAND2_X1 U12168 ( .A1(n14944), .A2(n21369), .ZN(n12264) );
  AND2_X1 U12169 ( .A1(n14744), .A2(n14742), .ZN(n20612) );
  INV_X1 U12170 ( .A(n14168), .ZN(n12290) );
  INV_X1 U12171 ( .A(n20612), .ZN(n20595) );
  OR2_X1 U12172 ( .A1(n15062), .A2(n11939), .ZN(n13480) );
  AND2_X1 U12173 ( .A1(n13826), .A2(n13825), .ZN(n14140) );
  AND2_X1 U12174 ( .A1(n13844), .A2(n13821), .ZN(n13822) );
  INV_X1 U12175 ( .A(n12492), .ZN(n14803) );
  NAND2_X1 U12176 ( .A1(n14723), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14773) );
  NAND2_X1 U12177 ( .A1(n12263), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12580) );
  INV_X1 U12178 ( .A(n12619), .ZN(n12263) );
  AND2_X1 U12179 ( .A1(n12629), .A2(n12647), .ZN(n14711) );
  NAND2_X1 U12180 ( .A1(n15144), .A2(n10234), .ZN(n10233) );
  INV_X1 U12181 ( .A(n10236), .ZN(n10234) );
  INV_X1 U12182 ( .A(n10237), .ZN(n10235) );
  NAND2_X1 U12183 ( .A1(n12261), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12530) );
  INV_X1 U12184 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12529) );
  OR2_X1 U12185 ( .A1(n12497), .A2(n15204), .ZN(n12513) );
  NAND2_X1 U12186 ( .A1(n12260), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12497) );
  INV_X1 U12187 ( .A(n12480), .ZN(n12260) );
  INV_X1 U12188 ( .A(n15214), .ZN(n10231) );
  NAND2_X1 U12189 ( .A1(n12462), .A2(n10232), .ZN(n15228) );
  NAND2_X1 U12190 ( .A1(n12259), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12463) );
  NAND2_X1 U12191 ( .A1(n12258), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12446) );
  INV_X1 U12192 ( .A(n12430), .ZN(n12258) );
  OR2_X1 U12193 ( .A1(n15282), .A2(n9980), .ZN(n9977) );
  OR2_X1 U12194 ( .A1(n15480), .A2(n15282), .ZN(n9979) );
  NAND2_X1 U12195 ( .A1(n15480), .A2(n9803), .ZN(n9978) );
  INV_X1 U12196 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12390) );
  NAND2_X1 U12197 ( .A1(n15480), .A2(n9980), .ZN(n15329) );
  AND2_X1 U12198 ( .A1(n15480), .A2(n15479), .ZN(n15482) );
  AND2_X1 U12199 ( .A1(n15280), .A2(n15343), .ZN(n15480) );
  AOI21_X1 U12200 ( .B1(n12326), .B2(n12455), .A(n12332), .ZN(n15486) );
  CLKBUF_X1 U12201 ( .A(n15279), .Z(n15280) );
  NAND2_X1 U12202 ( .A1(n15491), .A2(n10386), .ZN(n15496) );
  NAND2_X1 U12203 ( .A1(n12309), .A2(n12455), .ZN(n9981) );
  NAND2_X1 U12204 ( .A1(n14166), .A2(n12292), .ZN(n14440) );
  AND2_X2 U12205 ( .A1(n14440), .A2(n14439), .ZN(n15491) );
  XNOR2_X1 U12206 ( .A(n13337), .B(n13338), .ZN(n10189) );
  NOR2_X1 U12207 ( .A1(n15086), .A2(n14876), .ZN(n15062) );
  AND2_X1 U12208 ( .A1(n15723), .A2(n13521), .ZN(n15714) );
  NAND2_X1 U12209 ( .A1(n14824), .A2(n13508), .ZN(n10169) );
  AND2_X1 U12210 ( .A1(n15161), .A2(n13451), .ZN(n15130) );
  OR2_X1 U12211 ( .A1(n15770), .A2(n13518), .ZN(n14820) );
  NOR2_X1 U12212 ( .A1(n15767), .A2(n9766), .ZN(n14822) );
  NAND2_X1 U12213 ( .A1(n12188), .A2(n9752), .ZN(n15566) );
  NAND2_X1 U12214 ( .A1(n10007), .A2(n10084), .ZN(n12188) );
  NAND2_X1 U12215 ( .A1(n15255), .A2(n10218), .ZN(n15188) );
  AND2_X1 U12216 ( .A1(n13433), .A2(n13432), .ZN(n15215) );
  AND2_X1 U12217 ( .A1(n15255), .A2(n15235), .ZN(n15237) );
  OR2_X1 U12218 ( .A1(n15657), .A2(n15806), .ZN(n15617) );
  OR2_X1 U12219 ( .A1(n15657), .A2(n12185), .ZN(n15613) );
  OR2_X1 U12220 ( .A1(n15289), .A2(n15269), .ZN(n15267) );
  OR2_X1 U12221 ( .A1(n15306), .A2(n15287), .ZN(n15289) );
  AND2_X1 U12222 ( .A1(n13515), .A2(n13514), .ZN(n15785) );
  AND2_X1 U12223 ( .A1(n17340), .A2(n9783), .ZN(n10397) );
  AND2_X1 U12224 ( .A1(n13399), .A2(n13398), .ZN(n17339) );
  AND3_X1 U12225 ( .A1(n13394), .A2(n13402), .A3(n13393), .ZN(n15401) );
  AND2_X1 U12226 ( .A1(n13392), .A2(n10214), .ZN(n10215) );
  AND2_X1 U12227 ( .A1(n13388), .A2(n13387), .ZN(n17354) );
  OR3_X1 U12228 ( .A1(n14172), .A2(n14442), .A3(n14171), .ZN(n17355) );
  INV_X1 U12229 ( .A(n13344), .ZN(n14029) );
  NAND2_X1 U12230 ( .A1(n13502), .A2(n14186), .ZN(n15779) );
  XNOR2_X1 U12231 ( .A(n12106), .B(n12281), .ZN(n20855) );
  OR2_X1 U12232 ( .A1(n21463), .A2(n21065), .ZN(n21461) );
  INV_X1 U12233 ( .A(n11965), .ZN(n11870) );
  INV_X1 U12234 ( .A(n11945), .ZN(n13860) );
  INV_X1 U12235 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11996) );
  CLKBUF_X1 U12236 ( .A(n14175), .Z(n21464) );
  OR2_X1 U12237 ( .A1(n20971), .A2(n20774), .ZN(n20938) );
  NAND2_X1 U12238 ( .A1(n21463), .A2(n20772), .ZN(n20897) );
  AND3_X1 U12239 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21369), .A3(n20775), 
        .ZN(n20819) );
  NAND2_X1 U12240 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21166) );
  AND2_X1 U12241 ( .A1(n20971), .A2(n20774), .ZN(n21163) );
  OR3_X1 U12242 ( .A1(n11017), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n11012), .ZN(n11031) );
  INV_X1 U12243 ( .A(n11035), .ZN(n14499) );
  NOR2_X1 U12244 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  NOR2_X1 U12245 ( .A1(n19667), .A2(n15914), .ZN(n10272) );
  INV_X1 U12246 ( .A(n15913), .ZN(n10273) );
  NOR2_X1 U12247 ( .A1(n10981), .A2(n10982), .ZN(n10990) );
  NOR2_X1 U12248 ( .A1(n15955), .A2(n10421), .ZN(n15946) );
  NAND2_X1 U12249 ( .A1(n10687), .A2(n10688), .ZN(n10981) );
  AOI21_X1 U12250 ( .B1(n15968), .B2(n16511), .A(n17002), .ZN(n15955) );
  NOR2_X1 U12251 ( .A1(n10212), .A2(n10211), .ZN(n10210) );
  INV_X1 U12252 ( .A(n10416), .ZN(n10212) );
  NAND2_X1 U12253 ( .A1(n19684), .A2(n15014), .ZN(n16007) );
  AND2_X1 U12254 ( .A1(n10629), .A2(n10628), .ZN(n19677) );
  AND2_X1 U12255 ( .A1(n16051), .A2(n16045), .ZN(n16029) );
  NAND2_X1 U12256 ( .A1(n10630), .A2(n9791), .ZN(n10626) );
  AND2_X1 U12257 ( .A1(n13321), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14763) );
  NAND2_X1 U12258 ( .A1(n16075), .A2(n16070), .ZN(n16052) );
  NOR2_X1 U12259 ( .A1(n16054), .A2(n16052), .ZN(n16051) );
  NOR2_X1 U12260 ( .A1(n15010), .A2(n16590), .ZN(n15013) );
  NAND2_X1 U12261 ( .A1(n16085), .A2(n16601), .ZN(n16076) );
  NOR2_X1 U12262 ( .A1(n9733), .A2(n10266), .ZN(n15006) );
  NOR2_X1 U12263 ( .A1(n9733), .A2(n11508), .ZN(n14994) );
  NOR2_X1 U12264 ( .A1(n16145), .A2(n16147), .ZN(n16129) );
  OR2_X1 U12265 ( .A1(n16159), .A2(n16164), .ZN(n16145) );
  INV_X1 U12266 ( .A(n17002), .ZN(n16146) );
  NAND2_X1 U12267 ( .A1(n10904), .A2(n9746), .ZN(n10950) );
  OR2_X1 U12268 ( .A1(n16172), .A2(n16686), .ZN(n16159) );
  INV_X1 U12269 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n16157) );
  NAND2_X1 U12270 ( .A1(n16182), .A2(n16184), .ZN(n16172) );
  MUX2_X1 U12271 ( .A(n10574), .B(n11173), .S(n10980), .Z(n10906) );
  NAND2_X1 U12272 ( .A1(n16218), .A2(n19757), .ZN(n16204) );
  INV_X1 U12273 ( .A(n16259), .ZN(n9843) );
  NOR2_X1 U12274 ( .A1(n16995), .A2(n9845), .ZN(n9844) );
  INV_X1 U12275 ( .A(n19664), .ZN(n16249) );
  NAND2_X1 U12276 ( .A1(n11410), .A2(n9952), .ZN(n11411) );
  AND2_X1 U12277 ( .A1(n16337), .A2(n16336), .ZN(n16338) );
  NOR2_X1 U12278 ( .A1(n14589), .A2(n10314), .ZN(n14583) );
  OAI21_X1 U12279 ( .B1(n13713), .B2(n13712), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14016) );
  NOR2_X1 U12280 ( .A1(n11005), .A2(n10752), .ZN(n9887) );
  OR2_X1 U12281 ( .A1(n16451), .A2(n14525), .ZN(n14924) );
  OR2_X1 U12282 ( .A1(n16451), .A2(n14522), .ZN(n14925) );
  INV_X1 U12283 ( .A(n13718), .ZN(n13774) );
  INV_X1 U12284 ( .A(n14016), .ZN(n17029) );
  AND2_X1 U12285 ( .A1(n15024), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14989) );
  INV_X1 U12286 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15944) );
  AND2_X1 U12287 ( .A1(n9729), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10275) );
  NAND2_X1 U12288 ( .A1(n9949), .A2(n11415), .ZN(n11416) );
  INV_X1 U12289 ( .A(n10145), .ZN(n10144) );
  OAI21_X1 U12290 ( .B1(n16544), .B2(n12656), .A(n14755), .ZN(n10145) );
  NOR2_X1 U12291 ( .A1(n12653), .A2(n16544), .ZN(n10133) );
  NOR2_X1 U12292 ( .A1(n16799), .A2(n10051), .ZN(n10050) );
  INV_X1 U12293 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15008) );
  NOR3_X1 U12294 ( .A1(n9733), .A2(n15008), .A3(n10264), .ZN(n15011) );
  INV_X1 U12295 ( .A(n10360), .ZN(n10358) );
  NOR2_X1 U12296 ( .A1(n14309), .A2(n14308), .ZN(n14550) );
  INV_X1 U12297 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15003) );
  NOR2_X1 U12298 ( .A1(n16201), .A2(n10280), .ZN(n10279) );
  NOR2_X1 U12299 ( .A1(n14996), .A2(n16684), .ZN(n15001) );
  INV_X1 U12300 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16684) );
  NAND2_X1 U12301 ( .A1(n9946), .A2(n11378), .ZN(n11379) );
  AND2_X1 U12302 ( .A1(n11091), .A2(n16914), .ZN(n16908) );
  NOR2_X1 U12303 ( .A1(n14998), .A2(n17389), .ZN(n15000) );
  NAND2_X1 U12304 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14998) );
  INV_X1 U12305 ( .A(n10775), .ZN(n9916) );
  INV_X1 U12306 ( .A(n10785), .ZN(n10810) );
  NAND2_X1 U12307 ( .A1(n9950), .A2(n11429), .ZN(n11430) );
  AND2_X1 U12308 ( .A1(n10984), .A2(n10609), .ZN(n13552) );
  AND2_X1 U12309 ( .A1(n11360), .A2(n11359), .ZN(n13557) );
  INV_X1 U12310 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16717) );
  NAND2_X1 U12311 ( .A1(n11358), .A2(n10302), .ZN(n10300) );
  NAND2_X1 U12312 ( .A1(n13025), .A2(n15964), .ZN(n13560) );
  NAND2_X1 U12313 ( .A1(n10002), .A2(n10694), .ZN(n9997) );
  NOR2_X1 U12314 ( .A1(n10686), .A2(n21707), .ZN(n16538) );
  AND2_X1 U12315 ( .A1(n10686), .A2(n21707), .ZN(n16537) );
  INV_X1 U12316 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21707) );
  INV_X1 U12317 ( .A(n10050), .ZN(n10048) );
  NAND2_X1 U12318 ( .A1(n11397), .A2(n9953), .ZN(n11398) );
  INV_X1 U12319 ( .A(n16542), .ZN(n16607) );
  NAND2_X1 U12320 ( .A1(n10368), .A2(n10366), .ZN(n16539) );
  OR3_X1 U12321 ( .A1(n16106), .A2(n10961), .A3(n10204), .ZN(n16620) );
  AND3_X1 U12322 ( .A1(n11279), .A2(n11278), .A3(n11277), .ZN(n14585) );
  AND3_X1 U12323 ( .A1(n11260), .A2(n11259), .A3(n11258), .ZN(n14590) );
  CLKBUF_X1 U12324 ( .A(n11518), .Z(n14589) );
  NAND2_X1 U12325 ( .A1(n11262), .A2(n11261), .ZN(n14587) );
  AND2_X1 U12326 ( .A1(n16772), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16855) );
  INV_X1 U12327 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16886) );
  INV_X1 U12328 ( .A(n16200), .ZN(n11174) );
  NAND2_X1 U12329 ( .A1(n16927), .A2(n10934), .ZN(n10940) );
  INV_X1 U12330 ( .A(n11366), .ZN(n9917) );
  AND3_X1 U12331 ( .A1(n11168), .A2(n11167), .A3(n11166), .ZN(n16230) );
  NAND2_X1 U12332 ( .A1(n14561), .A2(n11158), .ZN(n16231) );
  NAND2_X1 U12333 ( .A1(n10778), .A2(n10777), .ZN(n10792) );
  INV_X1 U12334 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16963) );
  OAI211_X1 U12335 ( .C1(n11137), .C2(n11149), .A(n11150), .B(n11136), .ZN(
        n14535) );
  XNOR2_X1 U12336 ( .A(n13814), .B(n12692), .ZN(n13791) );
  AOI21_X1 U12337 ( .B1(n16966), .B2(n12691), .A(n12690), .ZN(n13790) );
  AND2_X1 U12338 ( .A1(n10316), .A2(n10344), .ZN(n14461) );
  INV_X1 U12339 ( .A(n10069), .ZN(n10067) );
  OR2_X1 U12340 ( .A1(n10865), .A2(n19860), .ZN(n19865) );
  NAND2_X1 U12341 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19920) );
  INV_X1 U12342 ( .A(n10746), .ZN(n19839) );
  INV_X1 U12343 ( .A(n14524), .ZN(n19846) );
  AND2_X1 U12344 ( .A1(n20124), .A2(n19858), .ZN(n20059) );
  INV_X1 U12345 ( .A(n20125), .ZN(n20123) );
  INV_X1 U12346 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20252) );
  INV_X1 U12347 ( .A(n20190), .ZN(n20477) );
  NOR2_X2 U12348 ( .A1(n17029), .A2(n17028), .ZN(n19844) );
  NOR2_X2 U12349 ( .A1(n17027), .A2(n17028), .ZN(n19845) );
  INV_X1 U12350 ( .A(n20257), .ZN(n20250) );
  INV_X1 U12351 ( .A(n19844), .ZN(n19850) );
  INV_X1 U12352 ( .A(n19845), .ZN(n19851) );
  NAND2_X1 U12353 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n16978) );
  NOR2_X1 U12354 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14446), .ZN(n15048) );
  NOR2_X1 U12355 ( .A1(n13284), .A2(n14676), .ZN(n19468) );
  NAND2_X1 U12356 ( .A1(n10297), .A2(n10294), .ZN(n14690) );
  NOR2_X1 U12357 ( .A1(n10296), .A2(n10295), .ZN(n10294) );
  NOR2_X1 U12358 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17676), .ZN(n17661) );
  NOR2_X1 U12359 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17705), .ZN(n17683) );
  OR2_X1 U12360 ( .A1(n18080), .A2(n18081), .ZN(n11633) );
  AND4_X1 U12361 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n11647) );
  OR2_X1 U12362 ( .A1(n13171), .A2(n13170), .ZN(n13269) );
  AOI21_X1 U12363 ( .B1(n13892), .B2(n19503), .A(n19624), .ZN(n18426) );
  AND2_X1 U12364 ( .A1(n11720), .A2(n9779), .ZN(n10283) );
  NOR2_X1 U12365 ( .A1(n14700), .A2(n10087), .ZN(n10086) );
  INV_X1 U12366 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U12367 ( .A1(n17123), .A2(n18629), .ZN(n18616) );
  INV_X1 U12368 ( .A(n18650), .ZN(n18593) );
  NOR2_X1 U12369 ( .A1(n17132), .A2(n17650), .ZN(n17131) );
  AND3_X1 U12370 ( .A1(n10098), .A2(n10096), .A3(n10099), .ZN(n17133) );
  NAND2_X1 U12371 ( .A1(n18689), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18651) );
  NOR2_X1 U12372 ( .A1(n17143), .A2(n17689), .ZN(n18679) );
  AND2_X1 U12373 ( .A1(n18773), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17151) );
  NAND2_X1 U12374 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17161) );
  INV_X1 U12375 ( .A(n10149), .ZN(n14133) );
  INV_X1 U12376 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17169) );
  NOR2_X1 U12377 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19512), .ZN(n18694) );
  INV_X1 U12378 ( .A(n10258), .ZN(n17073) );
  NOR2_X1 U12379 ( .A1(n10256), .A2(n10254), .ZN(n10253) );
  INV_X1 U12380 ( .A(n10255), .ZN(n10254) );
  NAND2_X1 U12381 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  INV_X1 U12382 ( .A(n10256), .ZN(n10252) );
  INV_X1 U12383 ( .A(n10257), .ZN(n10251) );
  OR3_X1 U12384 ( .A1(n17226), .A2(n9728), .A3(n10165), .ZN(n17187) );
  NAND2_X1 U12385 ( .A1(n9963), .A2(n9961), .ZN(n17110) );
  NAND2_X1 U12386 ( .A1(n18547), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9963) );
  NAND2_X1 U12387 ( .A1(n13208), .A2(n13207), .ZN(n10239) );
  AND2_X1 U12388 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17229) );
  NOR2_X1 U12389 ( .A1(n18913), .A2(n18917), .ZN(n18901) );
  NOR2_X1 U12390 ( .A1(n13287), .A2(n13286), .ZN(n13908) );
  NOR2_X1 U12391 ( .A1(n13537), .A2(n18660), .ZN(n18934) );
  NOR2_X1 U12392 ( .A1(n18728), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18727) );
  NOR2_X1 U12393 ( .A1(n18978), .A2(n18490), .ZN(n10297) );
  INV_X1 U12394 ( .A(n13263), .ZN(n13261) );
  NOR2_X1 U12395 ( .A1(n18789), .A2(n19018), .ZN(n18788) );
  AND2_X1 U12396 ( .A1(n19042), .A2(n18286), .ZN(n13289) );
  AND2_X1 U12397 ( .A1(n13240), .A2(n11749), .ZN(n19469) );
  INV_X1 U12398 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19478) );
  INV_X1 U12399 ( .A(n13913), .ZN(n13926) );
  INV_X1 U12400 ( .A(n9990), .ZN(n14676) );
  INV_X1 U12401 ( .A(n13230), .ZN(n19042) );
  INV_X1 U12402 ( .A(n11727), .ZN(n19046) );
  INV_X1 U12403 ( .A(n13223), .ZN(n19051) );
  INV_X1 U12404 ( .A(n18286), .ZN(n19055) );
  INV_X1 U12405 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19512) );
  OR2_X1 U12406 ( .A1(n18490), .A2(n18489), .ZN(n19503) );
  INV_X1 U12407 ( .A(n17029), .ZN(n17027) );
  NAND2_X1 U12408 ( .A1(n14231), .A2(n13753), .ZN(n21485) );
  AND2_X1 U12409 ( .A1(n20561), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20625) );
  AND2_X1 U12410 ( .A1(n14744), .A2(n14728), .ZN(n20608) );
  INV_X1 U12411 ( .A(n20608), .ZN(n20638) );
  AND2_X1 U12412 ( .A1(n13878), .A2(n14141), .ZN(n20653) );
  NAND2_X1 U12413 ( .A1(n15497), .A2(n14145), .ZN(n15460) );
  INV_X1 U12414 ( .A(n14960), .ZN(n15462) );
  AND2_X1 U12415 ( .A1(n14720), .A2(n20769), .ZN(n15463) );
  NOR2_X2 U12416 ( .A1(n14147), .A2(n14720), .ZN(n15499) );
  INV_X1 U12417 ( .A(n15460), .ZN(n14147) );
  NOR2_X1 U12418 ( .A1(n14145), .A2(n14146), .ZN(n14144) );
  INV_X1 U12419 ( .A(n20654), .ZN(n20658) );
  AOI21_X1 U12420 ( .B1(n14941), .B2(n17288), .A(n17306), .ZN(n14037) );
  INV_X2 U12421 ( .A(n20675), .ZN(n20681) );
  AND2_X1 U12422 ( .A1(n11957), .A2(n21378), .ZN(n14229) );
  OR2_X1 U12423 ( .A1(n14231), .A2(n14230), .ZN(n14296) );
  INV_X1 U12424 ( .A(n20700), .ZN(n21499) );
  OAI21_X1 U12425 ( .B1(n15095), .B2(n15083), .A(n15082), .ZN(n15524) );
  AND2_X1 U12426 ( .A1(n12619), .A2(n12565), .ZN(n15551) );
  AND2_X1 U12427 ( .A1(n15250), .A2(n15266), .ZN(n15631) );
  INV_X1 U12428 ( .A(n15684), .ZN(n20640) );
  OR2_X1 U12429 ( .A1(n17364), .A2(n21304), .ZN(n20770) );
  XNOR2_X1 U12430 ( .A(n10378), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15704) );
  NAND2_X1 U12431 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  NAND2_X1 U12432 ( .A1(n15528), .A2(n15504), .ZN(n10379) );
  NOR2_X1 U12433 ( .A1(n9759), .A2(n10182), .ZN(n10181) );
  INV_X1 U12434 ( .A(n13509), .ZN(n10182) );
  NAND2_X1 U12435 ( .A1(n13510), .A2(n13509), .ZN(n15731) );
  XNOR2_X1 U12436 ( .A(n10167), .B(n13335), .ZN(n15738) );
  NAND2_X1 U12437 ( .A1(n10170), .A2(n10168), .ZN(n10167) );
  OAI21_X1 U12438 ( .B1(n13581), .B2(n13508), .A(n15657), .ZN(n10170) );
  OAI21_X1 U12439 ( .B1(n15514), .B2(n10169), .A(n12192), .ZN(n10168) );
  NAND2_X1 U12440 ( .A1(n10028), .A2(n10041), .ZN(n13582) );
  NAND2_X1 U12441 ( .A1(n13581), .A2(n15657), .ZN(n10041) );
  OAI21_X1 U12442 ( .B1(n15514), .B2(n10029), .A(n12192), .ZN(n10028) );
  NAND2_X1 U12443 ( .A1(n15583), .A2(n9713), .ZN(n9857) );
  OR2_X1 U12444 ( .A1(n15815), .A2(n13517), .ZN(n15770) );
  NAND2_X1 U12445 ( .A1(n10027), .A2(n12152), .ZN(n10025) );
  INV_X1 U12446 ( .A(n10081), .ZN(n20705) );
  AND2_X1 U12447 ( .A1(n15895), .A2(n13503), .ZN(n20750) );
  NAND2_X1 U12448 ( .A1(n15781), .A2(n15779), .ZN(n20735) );
  AND2_X1 U12449 ( .A1(n13502), .A2(n13873), .ZN(n20736) );
  INV_X1 U12450 ( .A(n20753), .ZN(n20738) );
  AND2_X1 U12451 ( .A1(n13502), .A2(n13483), .ZN(n20742) );
  CLKBUF_X1 U12452 ( .A(n12284), .Z(n20893) );
  INV_X1 U12453 ( .A(n20855), .ZN(n20774) );
  OAI21_X1 U12454 ( .B1(n14203), .B2(n17372), .A(n20945), .ZN(n21475) );
  NOR2_X1 U12455 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14944) );
  CLKBUF_X1 U12456 ( .A(n11996), .Z(n11997) );
  INV_X1 U12457 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13852) );
  OR2_X1 U12458 ( .A1(n17295), .A2(n21660), .ZN(n21454) );
  OAI211_X1 U12459 ( .C1(n20787), .C2(n21306), .A(n21123), .B(n20782), .ZN(
        n20823) );
  OAI22_X1 U12460 ( .A1(n20861), .A2(n20860), .B1(n21126), .B2(n21004), .ZN(
        n20885) );
  OR2_X1 U12461 ( .A1(n20897), .A2(n20996), .ZN(n20932) );
  OAI221_X1 U12462 ( .B1(n9828), .B2(n21660), .C1(n9828), .C2(n20947), .A(
        n21260), .ZN(n20964) );
  OAI21_X1 U12463 ( .B1(n20973), .B2(n20972), .A(n21314), .ZN(n20992) );
  NAND2_X1 U12464 ( .A1(n21034), .A2(n21226), .ZN(n21028) );
  OAI211_X1 U12465 ( .C1(n10408), .C2(n21660), .A(n21123), .B(n21071), .ZN(
        n21088) );
  INV_X1 U12466 ( .A(n21157), .ZN(n21118) );
  OAI211_X1 U12467 ( .C1(n21128), .C2(n21125), .A(n21124), .B(n21123), .ZN(
        n21160) );
  INV_X1 U12468 ( .A(n21188), .ZN(n21193) );
  OAI211_X1 U12469 ( .C1(n9829), .C2(n21660), .A(n21260), .B(n21202), .ZN(
        n21222) );
  AND2_X1 U12470 ( .A1(n21311), .A2(n21197), .ZN(n21248) );
  OAI21_X1 U12471 ( .B1(n21467), .B2(n21231), .A(n21314), .ZN(n21249) );
  OAI211_X1 U12472 ( .C1(n21292), .C2(n21261), .A(n21260), .B(n21259), .ZN(
        n21295) );
  INV_X1 U12473 ( .A(n21116), .ZN(n21310) );
  INV_X1 U12474 ( .A(n21131), .ZN(n21322) );
  INV_X1 U12475 ( .A(n21135), .ZN(n21328) );
  INV_X1 U12476 ( .A(n21139), .ZN(n21334) );
  INV_X1 U12477 ( .A(n21143), .ZN(n21340) );
  INV_X1 U12478 ( .A(n21147), .ZN(n21346) );
  INV_X1 U12479 ( .A(n21151), .ZN(n21352) );
  AND2_X1 U12480 ( .A1(n21311), .A2(n21163), .ZN(n21362) );
  OAI21_X1 U12481 ( .B1(n21316), .B2(n21315), .A(n21314), .ZN(n21363) );
  INV_X1 U12482 ( .A(n21156), .ZN(n21360) );
  NOR2_X1 U12483 ( .A1(n17370), .A2(n21306), .ZN(n17366) );
  NAND2_X1 U12484 ( .A1(n17370), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21370) );
  AOI221_X1 U12485 ( .B1(n21369), .B2(n17370), .C1(n17294), .C2(n17370), .A(
        n17365), .ZN(n17371) );
  OR2_X1 U12486 ( .A1(n13340), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n17306) );
  NAND2_X1 U12487 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21380), .ZN(n21494) );
  NAND2_X1 U12488 ( .A1(n11495), .A2(n11494), .ZN(n13728) );
  INV_X1 U12489 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20499) );
  OR2_X1 U12490 ( .A1(n15986), .A2(n15987), .ZN(n10205) );
  AND2_X1 U12491 ( .A1(n16029), .A2(n16034), .ZN(n19684) );
  AND2_X1 U12492 ( .A1(n9741), .A2(n10659), .ZN(n16048) );
  NAND2_X1 U12493 ( .A1(n10630), .A2(n10631), .ZN(n10658) );
  AND2_X1 U12494 ( .A1(n10675), .A2(n10674), .ZN(n16125) );
  INV_X1 U12495 ( .A(n19669), .ZN(n16216) );
  NAND2_X1 U12496 ( .A1(n16146), .A2(n19681), .ZN(n16219) );
  INV_X1 U12497 ( .A(n19667), .ZN(n16272) );
  INV_X1 U12498 ( .A(n19674), .ZN(n16267) );
  INV_X1 U12499 ( .A(n16254), .ZN(n19678) );
  OR2_X1 U12500 ( .A1(n11235), .A2(n11234), .ZN(n14303) );
  INV_X1 U12501 ( .A(n16353), .ZN(n16357) );
  AOI21_X2 U12502 ( .B1(n13761), .B2(n14448), .A(n13010), .ZN(n16350) );
  INV_X2 U12503 ( .A(n16350), .ZN(n16360) );
  NAND2_X1 U12504 ( .A1(n16350), .A2(n14524), .ZN(n16353) );
  XNOR2_X1 U12505 ( .A(n13007), .B(n13006), .ZN(n14932) );
  OAI211_X1 U12506 ( .C1(n10323), .C2(n12963), .A(n12985), .B(n10319), .ZN(
        n13007) );
  OAI21_X1 U12507 ( .B1(n12963), .B2(n16288), .A(n10324), .ZN(n16282) );
  INV_X1 U12508 ( .A(n14925), .ZN(n16459) );
  AND2_X1 U12509 ( .A1(n14840), .A2(n14843), .ZN(n16450) );
  OR2_X1 U12510 ( .A1(n16065), .A2(n16064), .ZN(n16786) );
  AND2_X1 U12511 ( .A1(n14067), .A2(n12696), .ZN(n14158) );
  INV_X1 U12512 ( .A(n16468), .ZN(n19705) );
  NOR2_X1 U12513 ( .A1(n15049), .A2(n13935), .ZN(n13968) );
  INV_X1 U12514 ( .A(n13968), .ZN(n13971) );
  NOR2_X2 U12515 ( .A1(n13936), .A2(n11051), .ZN(n14019) );
  NAND2_X1 U12516 ( .A1(n10263), .A2(n14901), .ZN(n10259) );
  NAND2_X1 U12517 ( .A1(n15024), .A2(n9730), .ZN(n10260) );
  OR2_X1 U12518 ( .A1(n15024), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U12519 ( .A1(n10052), .A2(n10050), .ZN(n14850) );
  INV_X1 U12520 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16590) );
  AND2_X1 U12521 ( .A1(n14309), .A2(n11506), .ZN(n16142) );
  OR2_X1 U12522 ( .A1(n11516), .A2(n19785), .ZN(n11513) );
  INV_X1 U12523 ( .A(n19787), .ZN(n19774) );
  INV_X1 U12524 ( .A(n19785), .ZN(n19763) );
  INV_X1 U12525 ( .A(n19771), .ZN(n19758) );
  OR2_X1 U12526 ( .A1(n13728), .A2(n11051), .ZN(n19785) );
  INV_X1 U12527 ( .A(n17388), .ZN(n19779) );
  NAND2_X1 U12528 ( .A1(n14896), .A2(n9956), .ZN(n14897) );
  XNOR2_X1 U12529 ( .A(n10995), .B(n10994), .ZN(n14915) );
  NOR2_X1 U12530 ( .A1(n14887), .A2(n10993), .ZN(n10994) );
  AOI21_X1 U12532 ( .B1(n16499), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16487) );
  XNOR2_X1 U12533 ( .A(n16499), .B(n10350), .ZN(n16495) );
  XNOR2_X1 U12534 ( .A(n13024), .B(n13023), .ZN(n16523) );
  NOR2_X1 U12535 ( .A1(n16560), .A2(n11560), .ZN(n11562) );
  NAND2_X1 U12536 ( .A1(n16567), .A2(n16758), .ZN(n10054) );
  AND2_X1 U12537 ( .A1(n13317), .A2(n12664), .ZN(n9884) );
  NAND2_X1 U12538 ( .A1(n10137), .A2(n10135), .ZN(n12658) );
  NAND2_X1 U12539 ( .A1(n10138), .A2(n10136), .ZN(n10135) );
  AND2_X1 U12540 ( .A1(n10134), .A2(n10071), .ZN(n16573) );
  AND2_X1 U12541 ( .A1(n10146), .A2(n16572), .ZN(n10071) );
  CLKBUF_X1 U12542 ( .A(n16949), .Z(n17381) );
  OR2_X1 U12543 ( .A1(n13814), .A2(n13813), .ZN(n20090) );
  INV_X1 U12544 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20497) );
  INV_X1 U12545 ( .A(n14055), .ZN(n14056) );
  INV_X1 U12546 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21570) );
  INV_X1 U12547 ( .A(n20479), .ZN(n19957) );
  INV_X1 U12548 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13772) );
  INV_X1 U12549 ( .A(n10731), .ZN(n13769) );
  AOI21_X1 U12550 ( .B1(n14496), .B2(n17047), .A(n13767), .ZN(n17020) );
  INV_X1 U12551 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19824) );
  INV_X1 U12552 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19829) );
  AND2_X1 U12553 ( .A1(n20154), .A2(n19922), .ZN(n19913) );
  OAI211_X1 U12554 ( .C1(n19913), .C2(n19898), .A(n19897), .B(n20298), .ZN(
        n19915) );
  AND2_X1 U12555 ( .A1(n20059), .A2(n20477), .ZN(n19968) );
  INV_X1 U12556 ( .A(n19972), .ZN(n19987) );
  OAI21_X1 U12557 ( .B1(n20478), .B2(n19967), .A(n19966), .ZN(n19986) );
  OAI21_X1 U12558 ( .B1(n19999), .B2(n19998), .A(n19997), .ZN(n20026) );
  INV_X1 U12559 ( .A(n20095), .ZN(n20098) );
  NOR2_X1 U12560 ( .A1(n20064), .A2(n20063), .ZN(n20085) );
  AND2_X1 U12561 ( .A1(n20253), .A2(n20183), .ZN(n20158) );
  OAI21_X1 U12562 ( .B1(n20224), .B2(n20221), .A(n20220), .ZN(n20245) );
  INV_X1 U12563 ( .A(n20341), .ZN(n20265) );
  INV_X1 U12564 ( .A(n20347), .ZN(n20268) );
  INV_X1 U12565 ( .A(n20360), .ZN(n20274) );
  AND2_X1 U12566 ( .A1(n20298), .A2(n19814), .ZN(n20339) );
  INV_X1 U12567 ( .A(n20002), .ZN(n20344) );
  AND2_X1 U12568 ( .A1(n20298), .A2(n19820), .ZN(n20345) );
  INV_X1 U12569 ( .A(n19871), .ZN(n20351) );
  AND2_X1 U12570 ( .A1(n20298), .A2(n17037), .ZN(n20352) );
  AND2_X1 U12571 ( .A1(n20298), .A2(n19825), .ZN(n20358) );
  AND2_X1 U12572 ( .A1(n20298), .A2(n19830), .ZN(n20365) );
  INV_X1 U12573 ( .A(n19942), .ZN(n20370) );
  AND2_X1 U12574 ( .A1(n20298), .A2(n19835), .ZN(n20371) );
  INV_X1 U12575 ( .A(n20210), .ZN(n20379) );
  AND2_X1 U12576 ( .A1(n20298), .A2(n19840), .ZN(n20377) );
  INV_X1 U12577 ( .A(n20022), .ZN(n20382) );
  NOR2_X1 U12578 ( .A1(n20337), .A2(n20336), .ZN(n20385) );
  AND2_X1 U12579 ( .A1(n20298), .A2(n19849), .ZN(n20384) );
  NAND2_X1 U12580 ( .A1(n14606), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17019) );
  INV_X1 U12581 ( .A(n14605), .ZN(n14606) );
  AOI21_X1 U12582 ( .B1(n13758), .B2(n11050), .A(n16975), .ZN(n20501) );
  INV_X1 U12583 ( .A(n20520), .ZN(n20509) );
  AND3_X1 U12584 ( .A1(n16993), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17047) );
  NAND3_X1 U12585 ( .A1(n20395), .A2(n20458), .A3(n20407), .ZN(n20513) );
  INV_X1 U12586 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20414) );
  INV_X1 U12587 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n21773) );
  NOR2_X1 U12588 ( .A1(n17869), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19639) );
  NOR2_X1 U12589 ( .A1(n13891), .A2(n14688), .ZN(n19473) );
  NAND2_X1 U12590 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19627) );
  INV_X1 U12591 ( .A(n10092), .ZN(n17581) );
  NOR2_X1 U12592 ( .A1(n17615), .A2(n17820), .ZN(n17606) );
  NOR2_X1 U12593 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17631), .ZN(n17617) );
  AND2_X1 U12594 ( .A1(n10094), .A2(n10093), .ZN(n17615) );
  INV_X1 U12595 ( .A(n18621), .ZN(n10093) );
  INV_X1 U12596 ( .A(n10094), .ZN(n17616) );
  NOR2_X1 U12597 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17654), .ZN(n17639) );
  NAND2_X1 U12598 ( .A1(n11591), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11583) );
  INV_X1 U12599 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n21783) );
  NAND2_X1 U12600 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17868), .ZN(n17852) );
  NOR2_X2 U12601 ( .A1(n19640), .A2(n19502), .ZN(n17846) );
  AND2_X1 U12602 ( .A1(n19638), .A2(n11752), .ZN(n17851) );
  INV_X1 U12603 ( .A(n17851), .ZN(n17868) );
  INV_X1 U12604 ( .A(n17804), .ZN(n17865) );
  AND2_X1 U12605 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17940), .ZN(n17945) );
  NOR2_X1 U12606 ( .A1(n17997), .A2(n17996), .ZN(n17980) );
  INV_X1 U12607 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18129) );
  NOR2_X1 U12608 ( .A1(n21756), .A2(n18169), .ZN(n18131) );
  NAND3_X1 U12609 ( .A1(n18428), .A2(n14322), .A3(n14321), .ZN(n18264) );
  INV_X1 U12610 ( .A(n18264), .ZN(n18279) );
  INV_X1 U12611 ( .A(n9987), .ZN(n18291) );
  NAND2_X1 U12612 ( .A1(n18300), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n18297) );
  NAND2_X1 U12613 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18309), .ZN(n18306) );
  NOR2_X1 U12614 ( .A1(n18438), .A2(n18315), .ZN(n18309) );
  NOR2_X1 U12615 ( .A1(n18364), .A2(n18319), .ZN(n18316) );
  NAND2_X1 U12616 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18316), .ZN(n18315) );
  NOR2_X1 U12617 ( .A1(n18359), .A2(n9825), .ZN(n18320) );
  NAND2_X1 U12618 ( .A1(n18320), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18319) );
  NOR2_X1 U12619 ( .A1(n18364), .A2(n18359), .ZN(n18353) );
  NOR2_X1 U12620 ( .A1(n18373), .A2(n18372), .ZN(n18407) );
  INV_X1 U12621 ( .A(n13269), .ZN(n18409) );
  INV_X1 U12622 ( .A(n13259), .ZN(n18416) );
  INV_X1 U12623 ( .A(n18390), .ZN(n18424) );
  INV_X1 U12624 ( .A(n18421), .ZN(n18399) );
  NAND2_X1 U12625 ( .A1(n18475), .A2(n18428), .ZN(n18457) );
  INV_X1 U12626 ( .A(n18486), .ZN(n18475) );
  NAND3_X1 U12627 ( .A1(n19509), .A2(n19473), .A3(n18426), .ZN(n18486) );
  INV_X1 U12628 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18536) );
  NOR2_X1 U12629 ( .A1(n18488), .A2(n9818), .ZN(n18533) );
  INV_X1 U12630 ( .A(n18714), .ZN(n18696) );
  NOR2_X1 U12631 ( .A1(n18710), .A2(n18697), .ZN(n18689) );
  INV_X1 U12632 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18697) );
  INV_X1 U12633 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18710) );
  NOR2_X1 U12634 ( .A1(n18764), .A2(n18425), .ZN(n18714) );
  NAND2_X1 U12635 ( .A1(n14696), .A2(n10405), .ZN(n18745) );
  INV_X1 U12636 ( .A(n18745), .ZN(n18763) );
  INV_X1 U12637 ( .A(n18700), .ZN(n18725) );
  NAND2_X1 U12638 ( .A1(n10245), .A2(n13155), .ZN(n14078) );
  NAND2_X1 U12639 ( .A1(n14104), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10245) );
  NOR2_X1 U12640 ( .A1(n17161), .A2(n21640), .ZN(n18773) );
  INV_X1 U12641 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21640) );
  OR2_X1 U12642 ( .A1(n18714), .A2(n18620), .ZN(n18790) );
  OR2_X1 U12643 ( .A1(n17488), .A2(n19626), .ZN(n18786) );
  INV_X1 U12644 ( .A(n18701), .ZN(n18792) );
  NAND2_X1 U12645 ( .A1(n10147), .A2(n10153), .ZN(n14088) );
  INV_X1 U12646 ( .A(n19409), .ZN(n19313) );
  NAND2_X1 U12647 ( .A1(n18772), .A2(n18691), .ZN(n18764) );
  XNOR2_X1 U12648 ( .A(n9965), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17197) );
  NAND2_X1 U12649 ( .A1(n17086), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17085) );
  INV_X1 U12650 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21581) );
  OR3_X1 U12651 ( .A1(n17226), .A2(n17113), .A3(n18830), .ZN(n18546) );
  NOR2_X1 U12652 ( .A1(n18981), .A2(n18978), .ZN(n18822) );
  NAND2_X1 U12653 ( .A1(n10298), .A2(n18961), .ZN(n18892) );
  OR2_X1 U12654 ( .A1(n13537), .A2(n10161), .ZN(n18684) );
  INV_X1 U12655 ( .A(n10163), .ZN(n10161) );
  OR2_X1 U12656 ( .A1(n18728), .A2(n10247), .ZN(n18677) );
  INV_X1 U12657 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18947) );
  OAI21_X1 U12658 ( .B1(n18945), .B2(n18944), .A(n18951), .ZN(n18992) );
  AND2_X1 U12659 ( .A1(n19464), .A2(n18405), .ZN(n18996) );
  AND2_X1 U12660 ( .A1(n18951), .A2(n19464), .ZN(n17252) );
  INV_X1 U12661 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19477) );
  NOR3_X1 U12662 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19625), .ZN(n19090) );
  INV_X1 U12663 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19028) );
  AND2_X1 U12664 ( .A1(n13898), .A2(n13897), .ZN(n14677) );
  NOR2_X1 U12665 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19608), .ZN(
        n19506) );
  AND2_X1 U12666 ( .A1(n19621), .A2(n18425), .ZN(n19509) );
  INV_X1 U12667 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19515) );
  NAND3_X1 U12668 ( .A1(n17483), .A2(n19593), .A3(n19522), .ZN(n19624) );
  INV_X2 U12669 ( .A(n19616), .ZN(n19635) );
  NOR2_X1 U12670 ( .A1(n17027), .A2(n13714), .ZN(n17409) );
  CLKBUF_X1 U12671 ( .A(n17433), .Z(n17442) );
  NOR2_X1 U12672 ( .A1(n17445), .A2(n17409), .ZN(n17444) );
  OAI21_X1 U12673 ( .B1(n15060), .B2(n20537), .A(n15059), .ZN(P1_U2968) );
  AOI21_X1 U12674 ( .B1(n15058), .B2(n20709), .A(n15057), .ZN(n15059) );
  AOI21_X1 U12675 ( .B1(n15377), .B2(n20709), .A(n14837), .ZN(n14838) );
  OAI21_X1 U12676 ( .B1(n15060), .B2(n20753), .A(n10178), .ZN(P1_U3000) );
  NOR3_X1 U12677 ( .A1(n13523), .A2(n13522), .A3(n10179), .ZN(n10178) );
  NAND2_X1 U12678 ( .A1(n9753), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U12679 ( .A1(n10274), .A2(n10267), .ZN(P2_U2825) );
  OAI21_X1 U12680 ( .B1(n15912), .B2(n19669), .A(n15911), .ZN(n10274) );
  OR2_X1 U12681 ( .A1(n9842), .A2(n17049), .ZN(n9841) );
  INV_X1 U12682 ( .A(n9838), .ZN(n9837) );
  NOR2_X1 U12683 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  NAND2_X1 U12684 ( .A1(n16755), .A2(n9834), .ZN(P2_U3024) );
  INV_X1 U12685 ( .A(n9835), .ZN(n9834) );
  OAI21_X1 U12686 ( .B1(n16757), .B2(n17400), .A(n16756), .ZN(n9835) );
  NAND2_X1 U12687 ( .A1(n9852), .A2(n11071), .ZN(n9851) );
  INV_X1 U12688 ( .A(n10035), .ZN(n14856) );
  NAND2_X1 U12689 ( .A1(n16839), .A2(n10191), .ZN(P2_U3033) );
  INV_X1 U12690 ( .A(n10192), .ZN(n10191) );
  OAI21_X1 U12691 ( .B1(n16840), .B2(n17400), .A(n16838), .ZN(n10192) );
  OAI21_X1 U12692 ( .B1(n9870), .B2(n9744), .A(n10390), .ZN(P2_U3036) );
  OR2_X1 U12693 ( .A1(n16633), .A2(n16942), .ZN(n9870) );
  AOI21_X1 U12694 ( .B1(n10090), .B2(n17837), .A(n10089), .ZN(n17510) );
  NAND2_X1 U12695 ( .A1(n17507), .A2(n10383), .ZN(n10089) );
  NAND2_X1 U12696 ( .A1(n9987), .A2(n21561), .ZN(n9986) );
  OR2_X1 U12697 ( .A1(n17105), .A2(n10288), .ZN(P3_U2803) );
  OAI21_X1 U12698 ( .B1(n17225), .B2(n18748), .A(n10289), .ZN(n10288) );
  AOI21_X1 U12699 ( .B1(n17120), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10290), .ZN(n10289) );
  AND2_X1 U12700 ( .A1(n10160), .A2(n10157), .ZN(n13313) );
  NAND2_X1 U12701 ( .A1(n13312), .A2(n13311), .ZN(n10160) );
  AOI21_X1 U12702 ( .B1(n10159), .B2(n19015), .A(n10158), .ZN(n10157) );
  OAI21_X1 U12703 ( .B1(n13549), .B2(n18976), .A(n13548), .ZN(n13550) );
  AOI211_X1 U12704 ( .C1(n19008), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17223), .B(n17222), .ZN(n17224) );
  NOR4_X1 U12705 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(n20769), .A4(n13703), .ZN(n13704) );
  NAND2_X1 U12706 ( .A1(n17409), .A2(U214), .ZN(U212) );
  INV_X2 U12707 ( .A(n18203), .ZN(n17886) );
  INV_X1 U12708 ( .A(n11131), .ZN(n11127) );
  AND4_X1 U12709 ( .A1(n10281), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9712) );
  AND2_X2 U12710 ( .A1(n13906), .A2(n11607), .ZN(n13929) );
  INV_X1 U12711 ( .A(n13368), .ZN(n11939) );
  NAND2_X1 U12712 ( .A1(n11937), .A2(n11949), .ZN(n13368) );
  OAI21_X1 U12713 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19620), .A(n17488), 
        .ZN(n18772) );
  AND2_X1 U12714 ( .A1(n15584), .A2(n13500), .ZN(n9713) );
  AND2_X1 U12715 ( .A1(n10338), .A2(n9769), .ZN(n9714) );
  AND2_X1 U12716 ( .A1(n9856), .A2(n19781), .ZN(n9715) );
  INV_X1 U12717 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17389) );
  INV_X1 U12718 ( .A(n11130), .ZN(n10745) );
  NAND2_X1 U12719 ( .A1(n11922), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12034) );
  INV_X1 U12720 ( .A(n12034), .ZN(n10019) );
  NOR2_X1 U12721 ( .A1(n18981), .A2(n10299), .ZN(n10298) );
  NAND3_X1 U12722 ( .A1(n10745), .A2(n10739), .A3(n10746), .ZN(n9942) );
  NOR3_X1 U12723 ( .A1(n15110), .A2(n15103), .A3(n15112), .ZN(n9716) );
  NAND2_X1 U12724 ( .A1(n9857), .A2(n15641), .ZN(n15547) );
  NAND2_X1 U12725 ( .A1(n11130), .A2(n10746), .ZN(n10738) );
  AND3_X1 U12726 ( .A1(n10880), .A2(n10128), .A3(n10875), .ZN(n9717) );
  NOR2_X1 U12727 ( .A1(n16214), .A2(n16230), .ZN(n9718) );
  AND2_X1 U12728 ( .A1(n9713), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9719) );
  INV_X1 U12729 ( .A(n10752), .ZN(n11454) );
  AND2_X1 U12730 ( .A1(n9747), .A2(n10217), .ZN(n9720) );
  AND2_X1 U12731 ( .A1(n12654), .A2(n12656), .ZN(n9721) );
  AND2_X1 U12732 ( .A1(n10422), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n9722) );
  AND2_X1 U12733 ( .A1(n13195), .A2(n18993), .ZN(n9723) );
  AND2_X1 U12734 ( .A1(n10355), .A2(n10354), .ZN(n9724) );
  INV_X1 U12735 ( .A(n12653), .ZN(n10146) );
  AND2_X1 U12736 ( .A1(n15024), .A2(n9819), .ZN(n14908) );
  NAND2_X1 U12737 ( .A1(n13321), .A2(n9820), .ZN(n9725) );
  AND2_X1 U12738 ( .A1(n10622), .A2(n9811), .ZN(n15967) );
  AND2_X1 U12739 ( .A1(n10086), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9726) );
  OR2_X1 U12740 ( .A1(n17191), .A2(n13310), .ZN(n9727) );
  OR3_X1 U12741 ( .A1(n17113), .A2(n18830), .A3(n17214), .ZN(n9728) );
  AND2_X1 U12742 ( .A1(n10276), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9729) );
  AND2_X1 U12743 ( .A1(n10262), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9730) );
  AND2_X1 U12744 ( .A1(n16293), .A2(n12980), .ZN(n9731) );
  AND2_X1 U12745 ( .A1(n9820), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9732) );
  INV_X1 U12746 ( .A(n17689), .ZN(n10099) );
  OR2_X1 U12747 ( .A1(n15004), .A2(n15003), .ZN(n9733) );
  NAND2_X2 U12748 ( .A1(n13370), .A2(n20776), .ZN(n13400) );
  AND2_X4 U12749 ( .A1(n11124), .A2(n12673), .ZN(n11138) );
  AND2_X2 U12750 ( .A1(n12849), .A2(n10432), .ZN(n10496) );
  NAND2_X1 U12751 ( .A1(n10445), .A2(n12849), .ZN(n10853) );
  NAND2_X2 U12752 ( .A1(n11126), .A2(n11125), .ZN(n11140) );
  NAND2_X1 U12753 ( .A1(n11132), .A2(n12673), .ZN(n11149) );
  OR2_X1 U12754 ( .A1(n16540), .A2(n16537), .ZN(n9734) );
  OR2_X1 U12755 ( .A1(n20735), .A2(n20736), .ZN(n20757) );
  NAND2_X1 U12756 ( .A1(n15583), .A2(n15584), .ZN(n15555) );
  NAND2_X1 U12757 ( .A1(n16338), .A2(n12826), .ZN(n16311) );
  AND2_X2 U12758 ( .A1(n10722), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10519) );
  OR2_X2 U12759 ( .A1(n12858), .A2(n10715), .ZN(n10559) );
  AND2_X1 U12760 ( .A1(n10377), .A2(n10375), .ZN(n9735) );
  NAND2_X1 U12761 ( .A1(n12849), .A2(n14461), .ZN(n9736) );
  OR2_X1 U12762 ( .A1(n15181), .A2(n15182), .ZN(n9737) );
  NAND2_X1 U12763 ( .A1(n10671), .A2(n10653), .ZN(n10652) );
  OR2_X1 U12764 ( .A1(n14309), .A2(n10359), .ZN(n9738) );
  AND2_X1 U12765 ( .A1(n9997), .A2(n11530), .ZN(n9739) );
  AND2_X1 U12766 ( .A1(n10032), .A2(n10034), .ZN(n9740) );
  NOR2_X1 U12767 ( .A1(n15990), .A2(n15991), .ZN(n13026) );
  NAND2_X1 U12768 ( .A1(n16431), .A2(n16430), .ZN(n11565) );
  AND2_X1 U12769 ( .A1(n16343), .A2(n16342), .ZN(n16337) );
  AND2_X1 U12770 ( .A1(n11600), .A2(n11606), .ZN(n13087) );
  INV_X1 U12771 ( .A(n17143), .ZN(n10098) );
  NAND2_X1 U12772 ( .A1(n10630), .A2(n10208), .ZN(n9741) );
  NOR2_X1 U12773 ( .A1(n15317), .A2(n15316), .ZN(n9742) );
  OR2_X1 U12774 ( .A1(n16514), .A2(n16717), .ZN(n9743) );
  AND2_X1 U12775 ( .A1(n16642), .A2(n11525), .ZN(n9744) );
  NAND2_X1 U12776 ( .A1(n11609), .A2(n11608), .ZN(n9745) );
  AND2_X1 U12777 ( .A1(n10953), .A2(n10594), .ZN(n9746) );
  AND2_X1 U12778 ( .A1(n13409), .A2(n17339), .ZN(n9747) );
  AND2_X1 U12779 ( .A1(n10665), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11560) );
  AND4_X1 U12780 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n9748) );
  AND2_X1 U12781 ( .A1(n13026), .A2(n13027), .ZN(n13025) );
  NAND2_X1 U12782 ( .A1(n12462), .A2(n12461), .ZN(n15226) );
  NOR2_X1 U12783 ( .A1(n17226), .A2(n17113), .ZN(n9749) );
  NAND2_X1 U12784 ( .A1(n17320), .A2(n12130), .ZN(n17313) );
  AND4_X1 U12785 ( .A1(n13091), .A2(n13090), .A3(n13089), .A4(n13088), .ZN(
        n9750) );
  NAND2_X1 U12786 ( .A1(n10742), .A2(n11060), .ZN(n11449) );
  NAND2_X1 U12787 ( .A1(n10301), .A2(n10302), .ZN(n13032) );
  NAND2_X1 U12788 ( .A1(n14663), .A2(n10357), .ZN(n11568) );
  OR3_X1 U12789 ( .A1(n18623), .A2(n14693), .A3(n21581), .ZN(n9751) );
  AND2_X1 U12790 ( .A1(n12187), .A2(n12189), .ZN(n9752) );
  AND2_X1 U12791 ( .A1(n10337), .A2(n10338), .ZN(n10747) );
  OR2_X1 U12792 ( .A1(n14772), .A2(n20760), .ZN(n9753) );
  NAND2_X1 U12793 ( .A1(n14663), .A2(n10355), .ZN(n9754) );
  AND2_X1 U12794 ( .A1(n9878), .A2(n9836), .ZN(n9755) );
  AND2_X1 U12795 ( .A1(n11406), .A2(n9954), .ZN(n9756) );
  NOR2_X1 U12796 ( .A1(n14589), .A2(n10312), .ZN(n14527) );
  NAND2_X1 U12797 ( .A1(n12191), .A2(n12192), .ZN(n15546) );
  OR2_X1 U12798 ( .A1(n12094), .A2(n12033), .ZN(n9757) );
  AND2_X1 U12799 ( .A1(n9947), .A2(n11389), .ZN(n9758) );
  AND2_X1 U12800 ( .A1(n20757), .A2(n13520), .ZN(n9759) );
  AND2_X1 U12801 ( .A1(n11131), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9760) );
  AND2_X1 U12802 ( .A1(n19846), .A2(n10101), .ZN(n9761) );
  AND2_X1 U12803 ( .A1(n13254), .A2(n10150), .ZN(n9762) );
  AND2_X1 U12804 ( .A1(n16500), .A2(n10105), .ZN(n9763) );
  AND3_X1 U12805 ( .A1(n10874), .A2(n10879), .A3(n10881), .ZN(n9764) );
  AND2_X1 U12806 ( .A1(n11092), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9765) );
  AND2_X1 U12807 ( .A1(n20757), .A2(n13518), .ZN(n9766) );
  NAND2_X1 U12808 ( .A1(n14842), .A2(n14841), .ZN(n9767) );
  INV_X1 U12809 ( .A(n10186), .ZN(n15718) );
  NAND2_X1 U12810 ( .A1(n13510), .A2(n10181), .ZN(n10186) );
  AND2_X1 U12811 ( .A1(n11860), .A2(n10166), .ZN(n9768) );
  AND2_X1 U12812 ( .A1(n10739), .A2(n10734), .ZN(n9769) );
  AND3_X1 U12813 ( .A1(n10101), .A2(n10739), .A3(n14524), .ZN(n9770) );
  OR2_X1 U12814 ( .A1(n15840), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9771) );
  INV_X1 U12815 ( .A(n11438), .ZN(n10345) );
  NOR2_X1 U12816 ( .A1(n11559), .A2(n12653), .ZN(n9772) );
  INV_X1 U12817 ( .A(n10225), .ZN(n15111) );
  NOR2_X1 U12818 ( .A1(n15110), .A2(n15112), .ZN(n10225) );
  AND2_X1 U12819 ( .A1(n14886), .A2(n16478), .ZN(n9773) );
  AND2_X1 U12820 ( .A1(n9864), .A2(n11953), .ZN(n9774) );
  AND2_X1 U12821 ( .A1(n10249), .A2(n10250), .ZN(n9775) );
  AND2_X1 U12822 ( .A1(n13552), .A2(n16506), .ZN(n9776) );
  INV_X1 U12823 ( .A(n10009), .ZN(n10008) );
  NAND2_X1 U12824 ( .A1(n9777), .A2(n10010), .ZN(n10009) );
  AND2_X1 U12825 ( .A1(n12183), .A2(n15679), .ZN(n9777) );
  NAND2_X1 U12826 ( .A1(n10322), .A2(n10325), .ZN(n16283) );
  NAND2_X1 U12827 ( .A1(n11540), .A2(n11541), .ZN(n11539) );
  OR2_X1 U12828 ( .A1(n9733), .A2(n10264), .ZN(n9778) );
  AND2_X1 U12829 ( .A1(n18428), .A2(n19055), .ZN(n9779) );
  NAND2_X1 U12830 ( .A1(n16598), .A2(n16585), .ZN(n9780) );
  NAND2_X1 U12831 ( .A1(n9976), .A2(n12000), .ZN(n12027) );
  AND2_X1 U12832 ( .A1(n10410), .A2(n10653), .ZN(n9781) );
  AND2_X1 U12833 ( .A1(n9746), .A2(n10213), .ZN(n9782) );
  AND2_X1 U12834 ( .A1(n9720), .A2(n13415), .ZN(n9783) );
  AND2_X1 U12835 ( .A1(n12654), .A2(n10138), .ZN(n9784) );
  OR2_X1 U12836 ( .A1(n17582), .A2(n18589), .ZN(n9785) );
  INV_X1 U12837 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16201) );
  INV_X1 U12838 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U12839 ( .A1(n11951), .A2(n11997), .ZN(n9786) );
  NAND2_X1 U12840 ( .A1(n10376), .A2(n11454), .ZN(n9787) );
  INV_X1 U12841 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10316) );
  OR2_X1 U12842 ( .A1(n13551), .A2(n13550), .ZN(P3_U2834) );
  AND2_X2 U12843 ( .A1(n11782), .A2(n13841), .ZN(n12011) );
  INV_X1 U12844 ( .A(n18889), .ZN(n10299) );
  NAND2_X1 U12845 ( .A1(n15255), .A2(n10220), .ZN(n15184) );
  INV_X1 U12846 ( .A(n20298), .ZN(n17025) );
  OAI21_X4 U12847 ( .B1(n17019), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16979), 
        .ZN(n20298) );
  NAND2_X1 U12848 ( .A1(n17114), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11577) );
  NAND2_X1 U12849 ( .A1(n14631), .A2(n12122), .ZN(n14573) );
  NAND2_X1 U12850 ( .A1(n14160), .A2(n10364), .ZN(n14543) );
  NAND2_X1 U12851 ( .A1(n17340), .A2(n9747), .ZN(n15331) );
  INV_X1 U12852 ( .A(n11940), .ZN(n12249) );
  NAND2_X1 U12853 ( .A1(n13321), .A2(n9732), .ZN(n9789) );
  NAND2_X1 U12854 ( .A1(n10911), .A2(n10912), .ZN(n9790) );
  AND2_X1 U12855 ( .A1(n10208), .A2(n10600), .ZN(n9791) );
  AND2_X1 U12856 ( .A1(n17340), .A2(n17339), .ZN(n9792) );
  AND2_X1 U12857 ( .A1(n15015), .A2(n10276), .ZN(n9793) );
  NAND2_X1 U12858 ( .A1(n11939), .A2(n11938), .ZN(n13484) );
  INV_X1 U12859 ( .A(n20537), .ZN(n20710) );
  NAND2_X1 U12860 ( .A1(n17340), .A2(n9720), .ZN(n9794) );
  NOR2_X1 U12861 ( .A1(n14309), .A2(n10358), .ZN(n14548) );
  AND2_X1 U12862 ( .A1(n10862), .A2(n10818), .ZN(n9795) );
  INV_X1 U12863 ( .A(n11569), .ZN(n10356) );
  INV_X1 U12864 ( .A(n11453), .ZN(n11462) );
  AND2_X1 U12865 ( .A1(n18703), .A2(n9962), .ZN(n9796) );
  AND3_X1 U12866 ( .A1(n11725), .A2(n11724), .A3(n11723), .ZN(n9797) );
  AND2_X1 U12867 ( .A1(n11431), .A2(n11546), .ZN(n9798) );
  AND2_X1 U12868 ( .A1(n11400), .A2(n9955), .ZN(n9799) );
  AND2_X1 U12869 ( .A1(n9951), .A2(n11436), .ZN(n9800) );
  AND2_X1 U12870 ( .A1(n15159), .A2(n15172), .ZN(n9801) );
  INV_X1 U12871 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14130) );
  AND2_X1 U12872 ( .A1(n13860), .A2(n20792), .ZN(n9802) );
  INV_X1 U12873 ( .A(n10768), .ZN(n10197) );
  AND2_X1 U12874 ( .A1(n9980), .A2(n15282), .ZN(n9803) );
  AND2_X1 U12875 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n9804) );
  AND2_X1 U12876 ( .A1(n17594), .A2(n11586), .ZN(n9805) );
  INV_X1 U12877 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17044) );
  AND2_X1 U12878 ( .A1(n10760), .A2(n10759), .ZN(n9806) );
  AND2_X1 U12879 ( .A1(n11558), .A2(n16543), .ZN(n9807) );
  INV_X1 U12880 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9866) );
  AND2_X1 U12881 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9808) );
  INV_X1 U12882 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11508) );
  INV_X1 U12883 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n21760) );
  AND2_X1 U12884 ( .A1(n10218), .A2(n9801), .ZN(n9809) );
  AND2_X1 U12885 ( .A1(n10613), .A2(n10612), .ZN(n9810) );
  AND2_X1 U12886 ( .A1(n10210), .A2(n15979), .ZN(n9811) );
  AND2_X1 U12887 ( .A1(n10232), .A2(n10231), .ZN(n9812) );
  AND2_X1 U12888 ( .A1(n9791), .A2(n19666), .ZN(n9813) );
  INV_X1 U12889 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17860) );
  AND2_X1 U12890 ( .A1(n10239), .A2(n18568), .ZN(n9814) );
  AND2_X1 U12891 ( .A1(n9798), .A2(n15918), .ZN(n9815) );
  AND2_X1 U12892 ( .A1(n9795), .A2(n11159), .ZN(n9816) );
  NAND2_X1 U12893 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9817) );
  INV_X1 U12894 ( .A(n10973), .ZN(n10371) );
  OR3_X1 U12895 ( .A1(n19626), .A2(n19529), .A3(n18489), .ZN(n9818) );
  INV_X1 U12896 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16991) );
  NAND2_X1 U12898 ( .A1(n17114), .A2(n9726), .ZN(n17053) );
  NOR2_X1 U12899 ( .A1(n14172), .A2(n14171), .ZN(n14170) );
  AND2_X1 U12900 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9819) );
  AND2_X1 U12901 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9820) );
  INV_X1 U12902 ( .A(n10618), .ZN(n10211) );
  INV_X1 U12903 ( .A(n19781), .ZN(n16690) );
  AND2_X1 U12904 ( .A1(n11496), .A2(n11051), .ZN(n19781) );
  AND2_X1 U12905 ( .A1(n17114), .A2(n10086), .ZN(n9821) );
  NOR2_X1 U12906 ( .A1(n13265), .A2(n18788), .ZN(n9822) );
  NOR2_X1 U12907 ( .A1(n14088), .A2(n14087), .ZN(n9823) );
  NAND2_X1 U12908 ( .A1(n13199), .A2(n18913), .ZN(n9824) );
  OR2_X1 U12909 ( .A1(n18330), .A2(n18444), .ZN(n9825) );
  INV_X1 U12910 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18993) );
  AND2_X1 U12911 ( .A1(n18901), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18888) );
  INV_X1 U12912 ( .A(n10263), .ZN(n10262) );
  NAND2_X1 U12913 ( .A1(n9819), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10263) );
  AND2_X1 U12914 ( .A1(n9732), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9826) );
  OR2_X1 U12915 ( .A1(n9824), .A2(n10247), .ZN(n9827) );
  NOR2_X1 U12916 ( .A1(n21198), .A2(n20997), .ZN(n9828) );
  CLKBUF_X3 U12917 ( .A(n17890), .Z(n18152) );
  NOR2_X1 U12918 ( .A1(n21198), .A2(n21301), .ZN(n9829) );
  INV_X1 U12919 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10204) );
  INV_X1 U12920 ( .A(n9694), .ZN(n21304) );
  INV_X1 U12921 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10151) );
  INV_X1 U12922 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10278) );
  INV_X1 U12923 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10038) );
  XNOR2_X1 U12924 ( .A(n13094), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14098) );
  INV_X1 U12925 ( .A(n13305), .ZN(n10165) );
  INV_X1 U12926 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U12927 ( .A1(n10692), .A2(n10350), .ZN(n9830) );
  INV_X1 U12928 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10088) );
  INV_X1 U12929 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9962) );
  INV_X1 U12930 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10213) );
  INV_X1 U12931 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n9985) );
  INV_X1 U12932 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10164) );
  INV_X1 U12933 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10248) );
  INV_X1 U12934 ( .A(n10203), .ZN(n10202) );
  NAND2_X1 U12935 ( .A1(n16813), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10203) );
  INV_X1 U12936 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10051) );
  AND2_X1 U12937 ( .A1(n11478), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9831) );
  INV_X1 U12938 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10350) );
  AOI21_X1 U12939 ( .B1(n16767), .B2(n19796), .A(n16766), .ZN(n16768) );
  AOI21_X1 U12940 ( .B1(n16495), .B2(n19796), .A(n11551), .ZN(n11552) );
  AOI211_X1 U12941 ( .C1(n16714), .C2(n19796), .A(n16713), .B(n16712), .ZN(
        n16715) );
  AND2_X1 U12942 ( .A1(n9883), .A2(n19796), .ZN(n10388) );
  AOI22_X2 U12943 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20816), .B1(DATAI_25_), 
        .B2(n20817), .ZN(n21326) );
  AOI22_X2 U12944 ( .A1(DATAI_19_), .A2(n20817), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20816), .ZN(n21278) );
  AOI22_X2 U12945 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20816), .B1(DATAI_18_), 
        .B2(n20817), .ZN(n21274) );
  AOI22_X2 U12946 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20816), .B1(DATAI_29_), 
        .B2(n20817), .ZN(n21350) );
  NOR2_X2 U12947 ( .A1(n20770), .A2(n20769), .ZN(n20816) );
  NOR2_X2 U12948 ( .A1(n20771), .A2(n20770), .ZN(n20817) );
  NAND2_X1 U12949 ( .A1(n9832), .A2(n11090), .ZN(n16907) );
  NAND3_X1 U12950 ( .A1(n9849), .A2(n11094), .A3(n9832), .ZN(n9848) );
  NAND2_X1 U12951 ( .A1(n9833), .A2(n10318), .ZN(n9941) );
  NAND2_X2 U12952 ( .A1(n10764), .A2(n10744), .ZN(n10774) );
  NAND2_X1 U12954 ( .A1(n11455), .A2(n9943), .ZN(n9872) );
  NAND3_X1 U12955 ( .A1(n9763), .A2(n19796), .A3(n10104), .ZN(n13569) );
  NAND3_X1 U12956 ( .A1(n9841), .A2(n15927), .A3(n9837), .ZN(P2_U2826) );
  NOR2_X1 U12957 ( .A1(n16259), .A2(n16995), .ZN(n16248) );
  NAND2_X1 U12958 ( .A1(n9844), .A2(n9843), .ZN(n16237) );
  INV_X1 U12959 ( .A(n19769), .ZN(n9845) );
  NOR2_X2 U12960 ( .A1(n16237), .A2(n17380), .ZN(n16218) );
  AND2_X1 U12961 ( .A1(n9846), .A2(n9917), .ZN(n14161) );
  XNOR2_X2 U12962 ( .A(n9846), .B(n9871), .ZN(n14070) );
  NAND2_X1 U12963 ( .A1(n9889), .A2(n9890), .ZN(n9846) );
  NAND2_X1 U12964 ( .A1(n11094), .A2(n9765), .ZN(n9847) );
  INV_X1 U12965 ( .A(n11090), .ZN(n9850) );
  NAND2_X1 U12966 ( .A1(n16784), .A2(n9851), .ZN(P2_U3028) );
  NAND2_X2 U12967 ( .A1(n10132), .A2(n10422), .ZN(n11440) );
  INV_X2 U12968 ( .A(n11131), .ZN(n11002) );
  NAND2_X1 U12969 ( .A1(n9855), .A2(n13317), .ZN(n16770) );
  NAND2_X1 U12970 ( .A1(n16643), .A2(n16773), .ZN(n9856) );
  XNOR2_X1 U12971 ( .A(n20935), .B(n20933), .ZN(n15905) );
  NAND2_X2 U12972 ( .A1(n10004), .A2(n12273), .ZN(n20933) );
  NAND2_X1 U12973 ( .A1(n9861), .A2(n12093), .ZN(n10081) );
  NAND2_X2 U12974 ( .A1(n12168), .A2(n17308), .ZN(n15688) );
  NAND4_X1 U12975 ( .A1(n10003), .A2(n11947), .A3(n11948), .A4(n13823), .ZN(
        n10020) );
  NAND2_X1 U12976 ( .A1(n20156), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n9867) );
  AND2_X2 U12977 ( .A1(n10811), .A2(n10813), .ZN(n20156) );
  NAND2_X1 U12978 ( .A1(n10866), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9868) );
  AND2_X2 U12979 ( .A1(n10812), .A2(n10813), .ZN(n10866) );
  NOR2_X2 U12980 ( .A1(n14070), .A2(n19788), .ZN(n10813) );
  NAND3_X1 U12981 ( .A1(n10732), .A2(n10731), .A3(n9943), .ZN(n9873) );
  INV_X1 U12982 ( .A(n13317), .ZN(n9876) );
  NAND2_X1 U12983 ( .A1(n16566), .A2(n11564), .ZN(n9878) );
  AOI21_X1 U12984 ( .B1(n9755), .B2(n19796), .A(n11574), .ZN(n11575) );
  AND2_X2 U12985 ( .A1(n13568), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16499) );
  NAND4_X1 U12986 ( .A1(n10709), .A2(n10707), .A3(n10710), .A4(n10708), .ZN(
        n9880) );
  NAND4_X1 U12987 ( .A1(n10713), .A2(n10711), .A3(n10714), .A4(n10712), .ZN(
        n9882) );
  NAND2_X1 U12988 ( .A1(n10132), .A2(n9722), .ZN(n9945) );
  INV_X1 U12989 ( .A(n11440), .ZN(n11420) );
  NAND4_X1 U12990 ( .A1(n11454), .A2(n13726), .A3(n9885), .A4(n10754), .ZN(
        n10130) );
  NAND3_X1 U12991 ( .A1(n9886), .A2(n11084), .A3(n16948), .ZN(n16949) );
  NAND3_X1 U12992 ( .A1(n9886), .A2(n11084), .A3(n10961), .ZN(n10915) );
  NAND2_X1 U12993 ( .A1(n9886), .A2(n11084), .ZN(n10352) );
  NAND2_X1 U12994 ( .A1(n10103), .A2(n10102), .ZN(n9886) );
  NAND2_X1 U12995 ( .A1(n9887), .A2(n10396), .ZN(n10328) );
  AND2_X1 U12996 ( .A1(n11462), .A2(n9887), .ZN(n14520) );
  INV_X1 U12997 ( .A(n10032), .ZN(n9892) );
  NAND3_X1 U12998 ( .A1(n10033), .A2(n10767), .A3(n10034), .ZN(n9889) );
  NAND2_X1 U12999 ( .A1(n9941), .A2(n9888), .ZN(n10033) );
  NAND2_X1 U13000 ( .A1(n10778), .A2(n10777), .ZN(n9888) );
  NAND2_X2 U13001 ( .A1(n9891), .A2(n9940), .ZN(n10034) );
  NAND2_X1 U13002 ( .A1(n9892), .A2(n10034), .ZN(n9890) );
  AND2_X2 U13003 ( .A1(n10198), .A2(n10196), .ZN(n9891) );
  NAND2_X1 U13004 ( .A1(n9904), .A2(n9893), .ZN(n11124) );
  OAI21_X1 U13005 ( .B1(n9899), .B2(n9894), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9893) );
  NAND4_X1 U13006 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n9894)
         );
  NAND4_X1 U13007 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9899)
         );
  OAI21_X1 U13008 ( .B1(n9910), .B2(n9905), .A(n10715), .ZN(n9904) );
  NAND4_X1 U13009 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9905)
         );
  NAND2_X1 U13010 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n9909) );
  NAND4_X1 U13011 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(n9910)
         );
  NAND2_X1 U13012 ( .A1(n9704), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9912) );
  OAI211_X1 U13013 ( .C1(n14915), .C2(n17400), .A(n11493), .B(n9915), .ZN(
        P2_U3016) );
  NAND2_X1 U13014 ( .A1(n14907), .A2(n19796), .ZN(n9915) );
  XNOR2_X1 U13015 ( .A(n16485), .B(n11114), .ZN(n14907) );
  AND2_X2 U13016 ( .A1(n12681), .A2(n14070), .ZN(n10809) );
  NAND4_X1 U13017 ( .A1(n9923), .A2(n9922), .A3(n9921), .A4(n9920), .ZN(n9919)
         );
  NAND4_X1 U13018 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n9924)
         );
  NAND4_X1 U13019 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n9930)
         );
  NAND4_X1 U13020 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(n9935)
         );
  AND2_X2 U13021 ( .A1(n10045), .A2(n10737), .ZN(n10764) );
  AND2_X1 U13022 ( .A1(n9941), .A2(n10767), .ZN(n10782) );
  NAND2_X1 U13023 ( .A1(n11420), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U13024 ( .A1(n11420), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U13025 ( .A1(n11420), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U13026 ( .A1(n11420), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U13027 ( .A1(n11420), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U13028 ( .A1(n11420), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U13029 ( .A1(n11420), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U13030 ( .A1(n11420), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U13031 ( .A1(n11420), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U13032 ( .A1(n11420), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U13033 ( .A1(n9957), .A2(n13115), .ZN(n18784) );
  NAND2_X1 U13034 ( .A1(n14134), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9957) );
  NAND2_X1 U13035 ( .A1(n13115), .A2(n14130), .ZN(n9959) );
  INV_X1 U13036 ( .A(n13115), .ZN(n9960) );
  NAND3_X1 U13037 ( .A1(n18637), .A2(n13209), .A3(n18552), .ZN(n18547) );
  NAND2_X2 U13038 ( .A1(n18568), .A2(n9964), .ZN(n18552) );
  NAND2_X1 U13039 ( .A1(n9966), .A2(n10258), .ZN(n9965) );
  NAND2_X2 U13040 ( .A1(n17086), .A2(n10255), .ZN(n10258) );
  INV_X1 U13041 ( .A(n17072), .ZN(n9966) );
  NAND2_X2 U13042 ( .A1(n9967), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18956) );
  NAND2_X2 U13043 ( .A1(n9968), .A2(n11108), .ZN(n14760) );
  NAND2_X1 U13044 ( .A1(n16656), .A2(n9969), .ZN(n9968) );
  NAND2_X1 U13045 ( .A1(n10030), .A2(n11097), .ZN(n16655) );
  NAND2_X1 U13046 ( .A1(n14859), .A2(n9970), .ZN(n16656) );
  AND2_X1 U13047 ( .A1(n10030), .A2(n14858), .ZN(n9970) );
  NAND2_X1 U13048 ( .A1(n10031), .A2(n10030), .ZN(n14859) );
  NAND2_X2 U13049 ( .A1(n10705), .A2(n10706), .ZN(n10741) );
  NAND2_X2 U13050 ( .A1(n16617), .A2(n10395), .ZN(n16609) );
  NAND3_X1 U13051 ( .A1(n12026), .A2(n21369), .A3(n12008), .ZN(n9975) );
  AOI21_X2 U13052 ( .B1(n12027), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12001), .ZN(n12006) );
  NAND3_X1 U13053 ( .A1(n9979), .A2(n9978), .A3(n9977), .ZN(n15317) );
  NAND3_X1 U13054 ( .A1(n11948), .A2(n10003), .A3(n11947), .ZN(n11964) );
  NAND3_X1 U13055 ( .A1(n18287), .A2(n18415), .A3(n9986), .ZN(n18288) );
  NOR2_X2 U13056 ( .A1(n18365), .A2(n18536), .ZN(n18360) );
  NAND3_X1 U13057 ( .A1(n11702), .A2(n11700), .A3(n11701), .ZN(n9993) );
  NAND3_X1 U13058 ( .A1(n11699), .A2(n11697), .A3(n11696), .ZN(n9994) );
  XNOR2_X2 U13059 ( .A(n9740), .B(n10776), .ZN(n10785) );
  INV_X1 U13061 ( .A(n11131), .ZN(n9996) );
  AND3_X4 U13062 ( .A1(n11454), .A2(n9869), .A3(n9995), .ZN(n11438) );
  NAND3_X1 U13063 ( .A1(n10003), .A2(n11948), .A3(n11938), .ZN(n13343) );
  NAND2_X1 U13064 ( .A1(n12274), .A2(n11994), .ZN(n10004) );
  OR2_X2 U13065 ( .A1(n12099), .A2(n11995), .ZN(n12274) );
  NAND3_X1 U13066 ( .A1(n12300), .A2(n14029), .A3(n12302), .ZN(n10075) );
  OAI21_X1 U13067 ( .B1(n12087), .B2(n10005), .A(n12078), .ZN(n12300) );
  NAND2_X1 U13068 ( .A1(n15688), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15681) );
  OAI21_X1 U13069 ( .B1(n15688), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15689), .ZN(n15680) );
  NAND2_X1 U13070 ( .A1(n11935), .A2(n10015), .ZN(n10022) );
  NAND3_X1 U13071 ( .A1(n10017), .A2(n12000), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10016) );
  NAND3_X1 U13072 ( .A1(n17320), .A2(n12154), .A3(n12130), .ZN(n10024) );
  NAND3_X1 U13073 ( .A1(n10024), .A2(n17309), .A3(n10023), .ZN(n12168) );
  OAI211_X1 U13074 ( .C1(n17320), .C2(n10026), .A(n10025), .B(n12154), .ZN(
        n17307) );
  NAND2_X1 U13075 ( .A1(n16910), .A2(n11095), .ZN(n10031) );
  NAND2_X1 U13076 ( .A1(n10033), .A2(n10767), .ZN(n10776) );
  NAND3_X1 U13077 ( .A1(n10040), .A2(n12178), .A3(n15640), .ZN(n15594) );
  NAND2_X1 U13078 ( .A1(n12064), .A2(n10042), .ZN(n12171) );
  NAND2_X1 U13079 ( .A1(n10043), .A2(n15641), .ZN(n13332) );
  NAND3_X1 U13080 ( .A1(n10045), .A2(n10744), .A3(n10044), .ZN(n10346) );
  NOR2_X1 U13081 ( .A1(n16596), .A2(n16799), .ZN(n16592) );
  INV_X1 U13082 ( .A(n16596), .ZN(n10052) );
  NAND3_X1 U13083 ( .A1(n10053), .A2(n10863), .A3(n9795), .ZN(n11084) );
  NAND3_X1 U13084 ( .A1(n10053), .A2(n10863), .A3(n9816), .ZN(n11086) );
  NAND2_X1 U13085 ( .A1(n10053), .A2(n10818), .ZN(n10103) );
  NAND3_X1 U13086 ( .A1(n10742), .A2(n11451), .A3(n11060), .ZN(n10055) );
  NAND2_X1 U13087 ( .A1(n14861), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16665) );
  AOI21_X2 U13088 ( .B1(n11500), .B2(n10974), .A(n10973), .ZN(n11553) );
  OAI21_X1 U13089 ( .B1(n14861), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16667), .ZN(n10956) );
  NOR2_X1 U13090 ( .A1(n10062), .A2(n10059), .ZN(n10128) );
  NAND4_X1 U13091 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10062) );
  NAND2_X1 U13092 ( .A1(n20156), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10063) );
  NAND2_X1 U13093 ( .A1(n10866), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10064) );
  NAND2_X1 U13094 ( .A1(n20061), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10065) );
  NAND2_X1 U13096 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10066) );
  INV_X1 U13098 ( .A(n10946), .ZN(n10884) );
  NAND2_X1 U13099 ( .A1(n9764), .A2(n9717), .ZN(n10070) );
  NAND2_X1 U13100 ( .A1(n12655), .A2(n12654), .ZN(n10134) );
  INV_X1 U13101 ( .A(n16609), .ZN(n12655) );
  NAND3_X1 U13102 ( .A1(n12127), .A2(n14573), .A3(n10073), .ZN(n10080) );
  NAND2_X1 U13103 ( .A1(n10075), .A2(n12081), .ZN(n12129) );
  NAND3_X1 U13104 ( .A1(n12128), .A2(n10080), .A3(n10078), .ZN(n17318) );
  NAND2_X1 U13105 ( .A1(n10079), .A2(n10081), .ZN(n10078) );
  NAND2_X2 U13106 ( .A1(n11870), .A2(n11894), .ZN(n11945) );
  OAI22_X1 U13107 ( .A1(n17604), .A2(n9785), .B1(n11593), .B2(n17582), .ZN(
        n17580) );
  NAND4_X1 U13108 ( .A1(n10098), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        n10099), .A4(n10096), .ZN(n17123) );
  NAND3_X1 U13109 ( .A1(n10098), .A2(n10099), .A3(n11576), .ZN(n18646) );
  INV_X1 U13110 ( .A(n14070), .ZN(n16246) );
  NAND3_X1 U13111 ( .A1(n9770), .A2(n10752), .A3(n10329), .ZN(n10731) );
  NAND2_X2 U13112 ( .A1(n10101), .A2(n10734), .ZN(n10752) );
  NAND2_X1 U13113 ( .A1(n16949), .A2(n11082), .ZN(n11087) );
  NAND2_X1 U13114 ( .A1(n10863), .A2(n10862), .ZN(n10102) );
  NAND3_X1 U13116 ( .A1(n9763), .A2(n10104), .A3(n19781), .ZN(n10399) );
  NAND4_X1 U13117 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10107) );
  NAND4_X1 U13118 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10112) );
  NAND4_X1 U13119 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10118) );
  NAND4_X1 U13120 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n10123) );
  NAND4_X1 U13121 ( .A1(n11454), .A2(n13726), .A3(n11117), .A4(n10754), .ZN(
        n14447) );
  NAND2_X1 U13122 ( .A1(n12655), .A2(n9784), .ZN(n10137) );
  NAND2_X1 U13123 ( .A1(n12655), .A2(n9721), .ZN(n10143) );
  OAI21_X1 U13124 ( .B1(n14087), .B2(n10148), .A(n10153), .ZN(n10149) );
  NAND2_X1 U13125 ( .A1(n13252), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10153) );
  NAND2_X1 U13126 ( .A1(n13265), .A2(n10156), .ZN(n10154) );
  NAND3_X1 U13127 ( .A1(n13309), .A2(n17059), .A3(n9727), .ZN(n10158) );
  NOR2_X1 U13128 ( .A1(n17226), .A2(n9728), .ZN(n17211) );
  OAI211_X2 U13129 ( .C1(n13343), .C2(n15351), .A(n11934), .B(n11933), .ZN(
        n11935) );
  OR2_X2 U13130 ( .A1(n16907), .A2(n16908), .ZN(n16910) );
  NAND4_X1 U13131 ( .A1(n10454), .A2(n10452), .A3(n10455), .A4(n10453), .ZN(
        n10172) );
  NAND4_X1 U13132 ( .A1(n10456), .A2(n10457), .A3(n10459), .A4(n10458), .ZN(
        n10174) );
  NAND2_X1 U13133 ( .A1(n10374), .A2(n10132), .ZN(n10377) );
  NAND2_X2 U13134 ( .A1(n10187), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U13135 ( .A1(n11946), .A2(n11954), .ZN(n10187) );
  NAND2_X2 U13136 ( .A1(n15527), .A2(n15538), .ZN(n15528) );
  AND2_X2 U13137 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13841) );
  OR2_X1 U13138 ( .A1(n10770), .A2(n10200), .ZN(n10195) );
  INV_X1 U13139 ( .A(n10770), .ZN(n10196) );
  NAND2_X2 U13140 ( .A1(n16643), .A2(n10202), .ZN(n16632) );
  NAND3_X1 U13141 ( .A1(n10613), .A2(n10612), .A3(n11177), .ZN(n10620) );
  AOI21_X1 U13142 ( .B1(n9810), .B2(n19676), .A(n10205), .ZN(n15988) );
  NAND4_X1 U13143 ( .A1(n10207), .A2(n10206), .A3(n10365), .A4(n11532), .ZN(
        n16479) );
  NAND4_X1 U13144 ( .A1(n10978), .A2(n10977), .A3(n10979), .A4(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10206) );
  NAND4_X1 U13145 ( .A1(n10978), .A2(n10983), .A3(n10977), .A4(n10979), .ZN(
        n10207) );
  NAND2_X1 U13146 ( .A1(n10671), .A2(n9781), .ZN(n10643) );
  NAND2_X1 U13147 ( .A1(n10622), .A2(n10210), .ZN(n10611) );
  NAND2_X1 U13148 ( .A1(n10622), .A2(n10618), .ZN(n10614) );
  NAND2_X1 U13149 ( .A1(n10904), .A2(n10953), .ZN(n10595) );
  INV_X1 U13150 ( .A(n14172), .ZN(n10216) );
  NAND3_X1 U13151 ( .A1(n13385), .A2(n10216), .A3(n10215), .ZN(n17356) );
  NAND2_X1 U13152 ( .A1(n15130), .A2(n13462), .ZN(n15110) );
  AND2_X4 U13153 ( .A1(n10228), .A2(n14182), .ZN(n12012) );
  AND2_X2 U13154 ( .A1(n11782), .A2(n10228), .ZN(n11901) );
  OAI211_X2 U13155 ( .C1(n10230), .C2(n9866), .A(n9774), .B(n10229), .ZN(
        n11972) );
  AND2_X2 U13156 ( .A1(n12462), .A2(n9812), .ZN(n15213) );
  NAND3_X1 U13157 ( .A1(n15491), .A2(n10386), .A3(n12325), .ZN(n15485) );
  NOR2_X1 U13158 ( .A1(n15181), .A2(n10233), .ZN(n12629) );
  NOR2_X1 U13159 ( .A1(n15181), .A2(n10235), .ZN(n15156) );
  NAND2_X1 U13160 ( .A1(n10240), .A2(n9723), .ZN(n17139) );
  NAND2_X1 U13161 ( .A1(n14104), .A2(n10244), .ZN(n10243) );
  NAND2_X2 U13162 ( .A1(n10243), .A2(n10241), .ZN(n13194) );
  NAND2_X1 U13163 ( .A1(n17086), .A2(n10253), .ZN(n10249) );
  AND2_X1 U13164 ( .A1(n10258), .A2(n10257), .ZN(n13213) );
  NAND3_X1 U13165 ( .A1(n10261), .A2(n10260), .A3(n10259), .ZN(n14986) );
  AOI21_X1 U13166 ( .B1(n15915), .B2(n19676), .A(n10268), .ZN(n10267) );
  NAND2_X1 U13167 ( .A1(n15015), .A2(n10275), .ZN(n15023) );
  NAND2_X1 U13168 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10280) );
  NAND3_X1 U13169 ( .A1(n10281), .A2(n10279), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14996) );
  NAND3_X1 U13170 ( .A1(n10281), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14999) );
  NAND2_X2 U13171 ( .A1(n11600), .A2(n11599), .ZN(n18186) );
  INV_X2 U13172 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19488) );
  INV_X1 U13173 ( .A(n15999), .ZN(n10301) );
  OR2_X2 U13174 ( .A1(n15999), .A2(n10300), .ZN(n13556) );
  NAND3_X1 U13175 ( .A1(n14561), .A2(n11158), .A3(n9718), .ZN(n16200) );
  NAND2_X1 U13176 ( .A1(n13555), .A2(n10305), .ZN(n15926) );
  NAND2_X1 U13177 ( .A1(n16431), .A2(n10310), .ZN(n11566) );
  INV_X1 U13178 ( .A(n11566), .ZN(n11352) );
  NAND2_X1 U13179 ( .A1(n11262), .A2(n10311), .ZN(n14840) );
  NAND3_X2 U13180 ( .A1(n10317), .A2(n10316), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12858) );
  NAND2_X1 U13181 ( .A1(n16294), .A2(n9731), .ZN(n10324) );
  NAND2_X1 U13182 ( .A1(n16294), .A2(n16293), .ZN(n16292) );
  NAND2_X1 U13183 ( .A1(n16292), .A2(n12963), .ZN(n10322) );
  NAND2_X1 U13184 ( .A1(n16294), .A2(n10320), .ZN(n10319) );
  INV_X1 U13185 ( .A(n16293), .ZN(n10321) );
  NOR2_X2 U13186 ( .A1(n10330), .A2(n12946), .ZN(n16287) );
  AND2_X1 U13187 ( .A1(n10330), .A2(n12946), .ZN(n12947) );
  NOR2_X2 U13188 ( .A1(n12926), .A2(n12925), .ZN(n10330) );
  NAND2_X1 U13189 ( .A1(n14154), .A2(n12702), .ZN(n14302) );
  NAND2_X1 U13190 ( .A1(n16337), .A2(n10333), .ZN(n10332) );
  INV_X4 U13191 ( .A(n12906), .ZN(n10723) );
  NAND2_X2 U13192 ( .A1(n10339), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12906) );
  NAND2_X1 U13193 ( .A1(n11438), .A2(n10346), .ZN(n10342) );
  AOI21_X1 U13194 ( .B1(n10757), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10343), .ZN(n10347) );
  NAND3_X1 U13195 ( .A1(n10348), .A2(n10349), .A3(n10347), .ZN(n10777) );
  OAI21_X2 U13196 ( .B1(n16609), .B2(n16582), .A(n16607), .ZN(n16600) );
  AND2_X2 U13197 ( .A1(n13568), .A2(n9831), .ZN(n16485) );
  NAND2_X1 U13198 ( .A1(n10352), .A2(n10351), .ZN(n17382) );
  INV_X1 U13199 ( .A(n16948), .ZN(n10351) );
  NOR2_X1 U13200 ( .A1(n14475), .A2(n10353), .ZN(n14454) );
  NAND2_X1 U13201 ( .A1(n14663), .A2(n9724), .ZN(n15990) );
  NAND2_X1 U13202 ( .A1(n13559), .A2(n9815), .ZN(n11444) );
  AND2_X1 U13203 ( .A1(n13559), .A2(n9798), .ZN(n15919) );
  AND2_X1 U13204 ( .A1(n13559), .A2(n11431), .ZN(n11545) );
  INV_X1 U13205 ( .A(n11444), .ZN(n11443) );
  NAND2_X1 U13206 ( .A1(n14160), .A2(n10362), .ZN(n11504) );
  NAND4_X1 U13207 ( .A1(n10756), .A2(n10749), .A3(n9735), .A4(n10748), .ZN(
        n10767) );
  NAND2_X1 U13208 ( .A1(n10983), .A2(n9830), .ZN(n10365) );
  NAND3_X1 U13209 ( .A1(n10956), .A2(n16665), .A3(n10369), .ZN(n10368) );
  NAND3_X1 U13210 ( .A1(n11462), .A2(n10376), .A3(n10373), .ZN(n10372) );
  AND3_X2 U13211 ( .A1(n15527), .A2(n15705), .A3(n15538), .ZN(n15506) );
  NAND2_X1 U13212 ( .A1(n15506), .A2(n15505), .ZN(n10380) );
  NAND2_X1 U13213 ( .A1(n12000), .A2(n11951), .ZN(n10381) );
  NAND3_X1 U13214 ( .A1(n15680), .A2(n15681), .A3(n15679), .ZN(n15668) );
  NAND2_X1 U13215 ( .A1(n10518), .A2(n10517), .ZN(n10916) );
  OR2_X2 U13216 ( .A1(n13211), .A2(n14698), .ZN(n17101) );
  AND2_X1 U13217 ( .A1(n15154), .A2(n15081), .ZN(n15095) );
  INV_X1 U13218 ( .A(n11178), .ZN(n14602) );
  CLKBUF_X1 U13219 ( .A(n11453), .Z(n13009) );
  NOR2_X1 U13220 ( .A1(n13017), .A2(n10400), .ZN(n16532) );
  XNOR2_X1 U13221 ( .A(n11087), .B(n11088), .ZN(n16926) );
  NOR2_X2 U13222 ( .A1(n11937), .A2(n11940), .ZN(n11958) );
  NAND2_X1 U13223 ( .A1(n11937), .A2(n13874), .ZN(n11927) );
  AND3_X1 U13224 ( .A1(n11459), .A2(n11458), .A3(n11457), .ZN(n11460) );
  NAND2_X1 U13225 ( .A1(n12087), .A2(n20936), .ZN(n12293) );
  NAND2_X1 U13226 ( .A1(n11030), .A2(n10980), .ZN(n10518) );
  AOI22_X1 U13227 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10485) );
  INV_X1 U13228 ( .A(n18734), .ZN(n18703) );
  AND2_X1 U13229 ( .A1(n20653), .A2(n20818), .ZN(n20649) );
  OR2_X1 U13230 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n11755), .ZN(n10383) );
  OR2_X1 U13231 ( .A1(n11764), .A2(n11763), .ZN(P3_U2640) );
  INV_X1 U13232 ( .A(n18269), .ZN(n18276) );
  OR2_X1 U13233 ( .A1(n15120), .A2(n20770), .ZN(n10385) );
  AND2_X1 U13234 ( .A1(n15492), .A2(n15490), .ZN(n10386) );
  OR2_X1 U13235 ( .A1(n19808), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10387) );
  OR2_X1 U13236 ( .A1(n13571), .A2(n17400), .ZN(n10389) );
  AND2_X1 U13237 ( .A1(n11467), .A2(n20502), .ZN(n19796) );
  NAND2_X1 U13238 ( .A1(n11467), .A2(n20500), .ZN(n17400) );
  AND2_X1 U13239 ( .A1(n11529), .A2(n11528), .ZN(n10390) );
  INV_X2 U13240 ( .A(n14957), .ZN(n15497) );
  INV_X1 U13241 ( .A(n14840), .ZN(n11343) );
  NOR3_X1 U13242 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n10392) );
  AND2_X1 U13243 ( .A1(n11335), .A2(n11177), .ZN(n10394) );
  NOR2_X1 U13244 ( .A1(n16618), .A2(n16625), .ZN(n10395) );
  AND2_X1 U13245 ( .A1(n11126), .A2(n14523), .ZN(n10396) );
  AND3_X1 U13246 ( .A1(n13100), .A2(n13099), .A3(n13098), .ZN(n10398) );
  OR2_X1 U13247 ( .A1(n13016), .A2(n16538), .ZN(n10400) );
  AND4_X1 U13248 ( .A1(n14640), .A2(n12704), .A3(n14646), .A4(n14303), .ZN(
        n10401) );
  OR2_X1 U13249 ( .A1(n10980), .A2(n10596), .ZN(n10402) );
  AND4_X1 U13250 ( .A1(n12192), .A2(n15705), .A3(n14881), .A4(n15699), .ZN(
        n10403) );
  NAND2_X2 U13251 ( .A1(n15497), .A2(n14144), .ZN(n15501) );
  NAND2_X1 U13252 ( .A1(n10724), .A2(n10715), .ZN(n10404) );
  OR2_X1 U13253 ( .A1(n18700), .A2(n18956), .ZN(n10405) );
  AND2_X1 U13254 ( .A1(n10939), .A2(n10938), .ZN(n10406) );
  INV_X1 U13255 ( .A(n11518), .ZN(n11262) );
  INV_X2 U13256 ( .A(n21494), .ZN(n21439) );
  OR2_X1 U13257 ( .A1(n11561), .A2(n16549), .ZN(n10407) );
  INV_X1 U13258 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n16101) );
  INV_X1 U13259 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11114) );
  NOR2_X1 U13260 ( .A1(n21198), .A2(n21165), .ZN(n10408) );
  INV_X1 U13261 ( .A(n20773), .ZN(n12049) );
  AND3_X1 U13262 ( .A1(n10473), .A2(n10472), .A3(n10471), .ZN(n10409) );
  OR2_X1 U13263 ( .A1(n10980), .A2(n16101), .ZN(n10410) );
  AND2_X1 U13264 ( .A1(n12657), .A2(n16541), .ZN(n10411) );
  INV_X1 U13265 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12329) );
  INV_X1 U13266 ( .A(n12853), .ZN(n14449) );
  INV_X1 U13267 ( .A(n10722), .ZN(n12853) );
  NAND2_X1 U13268 ( .A1(n11342), .A2(n11341), .ZN(n10412) );
  INV_X2 U13269 ( .A(n18477), .ZN(n18484) );
  OR2_X1 U13270 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10413) );
  OR2_X1 U13271 ( .A1(n20032), .A2(n20333), .ZN(n20038) );
  INV_X1 U13272 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18253) );
  NAND2_X1 U13273 ( .A1(n11348), .A2(n11347), .ZN(n10414) );
  AND2_X1 U13274 ( .A1(n18714), .A2(n17504), .ZN(n10415) );
  INV_X1 U13275 ( .A(n12455), .ZN(n12426) );
  INV_X1 U13276 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19546) );
  OR2_X1 U13277 ( .A1(n18425), .A2(n18648), .ZN(n18455) );
  INV_X2 U13278 ( .A(n20674), .ZN(n20662) );
  OR2_X1 U13279 ( .A1(n19745), .A2(n19744), .ZN(n19747) );
  INV_X2 U13280 ( .A(n19747), .ZN(n19739) );
  OR2_X1 U13281 ( .A1(n10980), .A2(n10602), .ZN(n10416) );
  AND4_X1 U13282 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10417) );
  OR2_X1 U13283 ( .A1(n18488), .A2(n19503), .ZN(n18535) );
  INV_X2 U13284 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21306) );
  INV_X1 U13285 ( .A(n18589), .ZN(n11586) );
  INV_X1 U13286 ( .A(n12652), .ZN(n12653) );
  NAND3_X1 U13287 ( .A1(n11172), .A2(n11171), .A3(n11170), .ZN(n10418) );
  AND2_X1 U13288 ( .A1(n11335), .A2(n11173), .ZN(n10419) );
  NAND2_X2 U13289 ( .A1(n19639), .A2(n19515), .ZN(n10420) );
  AND2_X2 U13290 ( .A1(n19375), .A2(n19090), .ZN(n19409) );
  AND2_X1 U13291 ( .A1(n15025), .A2(n13572), .ZN(n10421) );
  INV_X1 U13292 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n12673) );
  OR2_X1 U13293 ( .A1(n20032), .A2(n20190), .ZN(n19947) );
  AND2_X1 U13294 ( .A1(n11513), .A2(n11512), .ZN(n10423) );
  INV_X1 U13295 ( .A(n11468), .ZN(n19748) );
  AND2_X1 U13296 ( .A1(n10805), .A2(n10804), .ZN(n10424) );
  AND3_X1 U13298 ( .A1(n10828), .A2(n10827), .A3(n10826), .ZN(n10425) );
  AND3_X1 U13299 ( .A1(n10815), .A2(n11002), .A3(n10814), .ZN(n10426) );
  AND2_X1 U13300 ( .A1(n10801), .A2(n10800), .ZN(n10427) );
  AND2_X1 U13301 ( .A1(n11963), .A2(n11962), .ZN(n10428) );
  OR2_X1 U13302 ( .A1(n12207), .A2(n12206), .ZN(n12195) );
  INV_X1 U13303 ( .A(n12218), .ZN(n12198) );
  OR2_X1 U13304 ( .A1(n12140), .A2(n12139), .ZN(n12158) );
  NAND2_X1 U13305 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11798) );
  AND2_X1 U13306 ( .A1(n19889), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10998) );
  AND2_X1 U13307 ( .A1(n10798), .A2(n10797), .ZN(n10816) );
  NAND2_X1 U13308 ( .A1(n10750), .A2(n10738), .ZN(n11055) );
  INV_X1 U13309 ( .A(n11942), .ZN(n11938) );
  INV_X1 U13310 ( .A(n11169), .ZN(n10882) );
  AND2_X1 U13311 ( .A1(n11133), .A2(n11131), .ZN(n10733) );
  AND2_X1 U13312 ( .A1(n11530), .A2(n16506), .ZN(n10616) );
  OR2_X1 U13313 ( .A1(n10852), .A2(n11323), .ZN(n10587) );
  NAND2_X1 U13314 ( .A1(n10741), .A2(n11133), .ZN(n11053) );
  INV_X1 U13315 ( .A(n11053), .ZN(n11054) );
  AOI22_X1 U13316 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12012), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11844) );
  INV_X1 U13317 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n21780) );
  INV_X1 U13318 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n21736) );
  NAND2_X1 U13319 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11917) );
  INV_X1 U13320 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U13321 ( .A1(n11943), .A2(n11959), .ZN(n12248) );
  INV_X1 U13322 ( .A(n12143), .ZN(n12144) );
  INV_X1 U13323 ( .A(n13468), .ZN(n13452) );
  OR2_X1 U13324 ( .A1(n12000), .A2(n11999), .ZN(n12005) );
  OR2_X1 U13325 ( .A1(n11834), .A2(n11833), .ZN(n12100) );
  AND2_X1 U13326 ( .A1(n10514), .A2(n10513), .ZN(n10996) );
  INV_X1 U13327 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11323) );
  INV_X2 U13328 ( .A(n12858), .ZN(n12986) );
  INV_X1 U13329 ( .A(n15966), .ZN(n11358) );
  NAND2_X1 U13330 ( .A1(n11086), .A2(n11085), .ZN(n11088) );
  NOR2_X1 U13331 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13196) );
  INV_X1 U13332 ( .A(n13113), .ZN(n13114) );
  AND4_X1 U13333 ( .A1(n11917), .A2(n11916), .A3(n11915), .A4(n11914), .ZN(
        n11918) );
  INV_X1 U13334 ( .A(n12513), .ZN(n12261) );
  INV_X1 U13335 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15239) );
  AND2_X1 U13336 ( .A1(n13437), .A2(n13436), .ZN(n15186) );
  AND2_X1 U13337 ( .A1(n13413), .A2(n13412), .ZN(n15332) );
  NAND2_X1 U13338 ( .A1(n12083), .A2(n14029), .ZN(n12126) );
  INV_X1 U13339 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14192) );
  OR2_X1 U13340 ( .A1(n17295), .A2(n13822), .ZN(n13826) );
  INV_X1 U13341 ( .A(n10996), .ZN(n11044) );
  INV_X1 U13342 ( .A(n12922), .ZN(n12903) );
  INV_X1 U13343 ( .A(n11519), .ZN(n11239) );
  NAND2_X1 U13344 ( .A1(n10488), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10489) );
  INV_X1 U13345 ( .A(n11536), .ZN(n10983) );
  AND2_X1 U13346 ( .A1(n16664), .A2(n16678), .ZN(n10955) );
  AND2_X1 U13347 ( .A1(n10903), .A2(n10902), .ZN(n11099) );
  NOR2_X1 U13348 ( .A1(n19494), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11739) );
  INV_X1 U13349 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18038) );
  INV_X1 U13350 ( .A(n13262), .ZN(n13264) );
  INV_X1 U13351 ( .A(n15320), .ZN(n13415) );
  NAND2_X1 U13352 ( .A1(n11936), .A2(n13823), .ZN(n11957) );
  AND2_X1 U13353 ( .A1(n12648), .A2(n15144), .ZN(n13671) );
  INV_X1 U13354 ( .A(n13666), .ZN(n14799) );
  NAND2_X1 U13355 ( .A1(n21306), .A2(n20830), .ZN(n14796) );
  NAND2_X1 U13356 ( .A1(n12333), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12422) );
  NOR2_X2 U13357 ( .A1(n20812), .A2(n21306), .ZN(n12455) );
  NAND2_X1 U13358 ( .A1(n15657), .A2(n15852), .ZN(n15640) );
  NOR2_X1 U13359 ( .A1(n17354), .A2(n17353), .ZN(n13392) );
  AND2_X1 U13360 ( .A1(n20896), .A2(n20926), .ZN(n20901) );
  INV_X1 U13361 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21066) );
  AND3_X1 U13362 ( .A1(n11837), .A2(n11836), .A3(n11835), .ZN(n12275) );
  OR2_X1 U13363 ( .A1(n11194), .A2(n11193), .ZN(n14541) );
  NAND2_X1 U13364 ( .A1(n12674), .A2(n12673), .ZN(n12688) );
  OR2_X1 U13365 ( .A1(n12942), .A2(n12948), .ZN(n12979) );
  OR2_X1 U13366 ( .A1(n12789), .A2(n12788), .ZN(n16336) );
  INV_X1 U13367 ( .A(n13756), .ZN(n14490) );
  AND2_X1 U13368 ( .A1(n11364), .A2(n11363), .ZN(n15924) );
  OR2_X1 U13369 ( .A1(n16028), .A2(n10642), .ZN(n16541) );
  OR2_X1 U13370 ( .A1(n14848), .A2(n19796), .ZN(n14849) );
  AND2_X1 U13371 ( .A1(n16855), .A2(n16813), .ZN(n16842) );
  AND3_X1 U13372 ( .A1(n11197), .A2(n11196), .A3(n11195), .ZN(n14518) );
  OR2_X1 U13373 ( .A1(n13238), .A2(n11745), .ZN(n13239) );
  OR2_X1 U13374 ( .A1(n11611), .A2(n11610), .ZN(n11612) );
  INV_X1 U13375 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n21584) );
  INV_X1 U13376 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14375) );
  INV_X1 U13377 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18084) );
  INV_X1 U13378 ( .A(n11663), .ZN(n18080) );
  INV_X1 U13379 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21564) );
  AND4_X1 U13380 ( .A1(n13141), .A2(n13140), .A3(n13139), .A4(n13138), .ZN(
        n13145) );
  NOR2_X1 U13381 ( .A1(n17598), .A2(n11585), .ZN(n18561) );
  AND2_X1 U13382 ( .A1(n13176), .A2(n13269), .ZN(n13190) );
  AND2_X1 U13383 ( .A1(n13746), .A2(n13744), .ZN(n13824) );
  INV_X1 U13384 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U13385 ( .A1(n13656), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13660) );
  OR2_X1 U13386 ( .A1(n21485), .A2(n14739), .ZN(n20561) );
  AND2_X1 U13387 ( .A1(n13445), .A2(n13444), .ZN(n15159) );
  NAND2_X1 U13388 ( .A1(n14140), .A2(n14139), .ZN(n14142) );
  INV_X1 U13389 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13595) );
  INV_X1 U13390 ( .A(n14796), .ZN(n14802) );
  INV_X1 U13391 ( .A(n15227), .ZN(n12479) );
  AND2_X1 U13392 ( .A1(n13486), .A2(n12251), .ZN(n13361) );
  INV_X1 U13393 ( .A(n20703), .ZN(n15577) );
  NAND2_X1 U13394 ( .A1(n15527), .A2(n15657), .ZN(n15530) );
  AND2_X1 U13395 ( .A1(n13423), .A2(n13422), .ZN(n15269) );
  INV_X1 U13396 ( .A(n15640), .ZN(n15643) );
  INV_X1 U13397 ( .A(n14186), .ZN(n14941) );
  OR2_X1 U13398 ( .A1(n20895), .A2(n21256), .ZN(n20788) );
  OR2_X1 U13399 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21037), .ZN(
        n21027) );
  NOR2_X1 U13400 ( .A1(n20778), .A2(n20945), .ZN(n21123) );
  AOI21_X1 U13401 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21677), .A(n20945), 
        .ZN(n21314) );
  AND2_X1 U13402 ( .A1(n17286), .A2(n17285), .ZN(n17298) );
  INV_X1 U13403 ( .A(n14991), .ZN(n14992) );
  NAND2_X1 U13404 ( .A1(n15039), .A2(n15038), .ZN(n19667) );
  INV_X1 U13405 ( .A(n19676), .ZN(n16270) );
  AND2_X1 U13406 ( .A1(n11041), .A2(n11040), .ZN(n13758) );
  NAND2_X1 U13407 ( .A1(n11461), .A2(n11460), .ZN(n14473) );
  NAND2_X1 U13408 ( .A1(n12694), .A2(n12693), .ZN(n14055) );
  INV_X1 U13409 ( .A(n16415), .ZN(n16461) );
  INV_X1 U13410 ( .A(n14590), .ZN(n11261) );
  INV_X1 U13411 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16530) );
  NOR2_X1 U13412 ( .A1(n16738), .A2(n13020), .ZN(n13024) );
  AND2_X1 U13413 ( .A1(n11350), .A2(n11349), .ZN(n16004) );
  NOR2_X1 U13414 ( .A1(n10665), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16562) );
  AND3_X1 U13415 ( .A1(n11338), .A2(n11337), .A3(n11336), .ZN(n14597) );
  INV_X1 U13416 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16937) );
  INV_X1 U13417 ( .A(n19788), .ZN(n17401) );
  AND2_X1 U13418 ( .A1(n20484), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20476) );
  INV_X1 U13419 ( .A(n19865), .ZN(n19861) );
  OR2_X1 U13420 ( .A1(n20032), .A2(n20257), .ZN(n20024) );
  OR2_X1 U13421 ( .A1(n20491), .A2(n20479), .ZN(n20125) );
  OR2_X1 U13422 ( .A1(n20491), .A2(n19957), .ZN(n20190) );
  NAND2_X1 U13423 ( .A1(n20298), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19847) );
  NAND2_X1 U13424 ( .A1(n17044), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14608) );
  INV_X1 U13425 ( .A(n19637), .ZN(n19629) );
  NOR2_X1 U13426 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  INV_X1 U13427 ( .A(n17511), .ZN(n17514) );
  AND2_X1 U13428 ( .A1(n18238), .A2(n17764), .ZN(n17746) );
  INV_X1 U13429 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17854) );
  NOR2_X1 U13430 ( .A1(n11613), .A2(n11612), .ZN(n11614) );
  INV_X1 U13431 ( .A(n18415), .ZN(n18346) );
  INV_X1 U13432 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14698) );
  AOI21_X1 U13433 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n9696), .A(n13547), .ZN(
        n13548) );
  INV_X1 U13434 ( .A(n18888), .ZN(n18644) );
  INV_X1 U13435 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18970) );
  AND2_X1 U13436 ( .A1(n13248), .A2(n13247), .ZN(n19464) );
  NAND2_X1 U13437 ( .A1(n19629), .A2(n13890), .ZN(n18889) );
  INV_X1 U13438 ( .A(n19245), .ZN(n19198) );
  AND2_X1 U13439 ( .A1(n19478), .A2(n19406), .ZN(n19345) );
  NOR2_X1 U13440 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19032), .ZN(n19375) );
  INV_X1 U13441 ( .A(n17368), .ZN(n21489) );
  INV_X1 U13442 ( .A(n15328), .ZN(n15274) );
  OR2_X1 U13443 ( .A1(n20612), .A2(n20610), .ZN(n15361) );
  NOR2_X2 U13444 ( .A1(n15056), .A2(n14737), .ZN(n20582) );
  AND2_X1 U13445 ( .A1(n20612), .A2(n20596), .ZN(n20586) );
  XNOR2_X1 U13446 ( .A(n13482), .B(n13481), .ZN(n14772) );
  INV_X1 U13447 ( .A(n20653), .ZN(n15404) );
  NAND2_X1 U13448 ( .A1(n14142), .A2(n14141), .ZN(n14957) );
  INV_X1 U13449 ( .A(n14296), .ZN(n20690) );
  NOR2_X1 U13450 ( .A1(n21497), .A2(n20792), .ZN(n20700) );
  AOI21_X1 U13451 ( .B1(n15551), .B2(n14802), .A(n12579), .ZN(n15144) );
  INV_X1 U13452 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13338) );
  OAI21_X1 U13453 ( .B1(n14726), .B2(n20760), .A(n13587), .ZN(n13588) );
  AND2_X1 U13454 ( .A1(n13449), .A2(n13448), .ZN(n15149) );
  NOR2_X1 U13455 ( .A1(n20733), .A2(n15851), .ZN(n17348) );
  NOR2_X1 U13456 ( .A1(n20743), .A2(n17328), .ZN(n17333) );
  INV_X1 U13457 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20734) );
  INV_X1 U13458 ( .A(n13858), .ZN(n21256) );
  OAI22_X1 U13459 ( .A1(n20789), .A2(n20788), .B1(n21126), .B2(n20940), .ZN(
        n20822) );
  OR2_X1 U13460 ( .A1(n20971), .A2(n20855), .ZN(n20974) );
  INV_X1 U13461 ( .A(n20905), .ZN(n20928) );
  INV_X1 U13462 ( .A(n20942), .ZN(n20963) );
  INV_X1 U13463 ( .A(n21028), .ZN(n20991) );
  OAI22_X1 U13464 ( .A1(n21006), .A2(n21005), .B1(n21004), .B2(n21254), .ZN(
        n21030) );
  INV_X1 U13465 ( .A(n21035), .ZN(n21060) );
  INV_X1 U13466 ( .A(n21050), .ZN(n21087) );
  INV_X1 U13467 ( .A(n20938), .ZN(n21197) );
  OAI22_X1 U13468 ( .A1(n21128), .A2(n21127), .B1(n21126), .B2(n21253), .ZN(
        n21159) );
  OAI22_X1 U13469 ( .A1(n21206), .A2(n21205), .B1(n21204), .B2(n21254), .ZN(
        n21221) );
  INV_X1 U13470 ( .A(n21262), .ZN(n21294) );
  NAND2_X1 U13471 ( .A1(n17370), .A2(n21306), .ZN(n17368) );
  INV_X1 U13472 ( .A(n21487), .ZN(n21378) );
  INV_X1 U13473 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21388) );
  AND2_X1 U13474 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21439), .ZN(n21423) );
  INV_X1 U13475 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16993) );
  OAI22_X1 U13476 ( .A1(n20503), .A2(n11115), .B1(n20501), .B2(n11052), .ZN(
        n11495) );
  NAND2_X1 U13477 ( .A1(n11443), .A2(n11442), .ZN(n14900) );
  INV_X1 U13478 ( .A(n17049), .ZN(n19681) );
  AND2_X1 U13479 ( .A1(n20521), .A2(n14984), .ZN(n19676) );
  AND2_X1 U13480 ( .A1(n13758), .A2(n17047), .ZN(n13721) );
  OR2_X1 U13481 ( .A1(n11334), .A2(n11333), .ZN(n14622) );
  OR2_X1 U13482 ( .A1(n11276), .A2(n11275), .ZN(n14554) );
  OR2_X1 U13483 ( .A1(n11215), .A2(n11214), .ZN(n14542) );
  OR2_X1 U13484 ( .A1(n14473), .A2(n13009), .ZN(n14448) );
  XNOR2_X1 U13485 ( .A(n13791), .B(n13790), .ZN(n20479) );
  NOR2_X1 U13486 ( .A1(n14924), .A2(n17029), .ZN(n16415) );
  INV_X1 U13487 ( .A(n16418), .ZN(n16466) );
  INV_X1 U13488 ( .A(n16462), .ZN(n19709) );
  AND2_X1 U13489 ( .A1(n13778), .A2(n13777), .ZN(n19745) );
  INV_X1 U13490 ( .A(n19696), .ZN(n19830) );
  INV_X1 U13491 ( .A(n13971), .ZN(n14024) );
  INV_X1 U13492 ( .A(n13328), .ZN(n13329) );
  AND2_X1 U13493 ( .A1(n9738), .A2(n14649), .ZN(n16832) );
  AND2_X1 U13494 ( .A1(n17388), .A2(n19778), .ZN(n19771) );
  INV_X1 U13495 ( .A(n17400), .ZN(n11071) );
  AND2_X1 U13496 ( .A1(n14434), .A2(n14208), .ZN(n17376) );
  AND2_X1 U13497 ( .A1(n11467), .A2(n11123), .ZN(n19792) );
  OAI21_X1 U13498 ( .B1(n17036), .B2(n17035), .A(n17034), .ZN(n19853) );
  NOR2_X1 U13499 ( .A1(n20219), .A2(n19919), .ZN(n19848) );
  INV_X1 U13500 ( .A(n19863), .ZN(n19883) );
  OAI21_X1 U13501 ( .B1(n19929), .B2(n19928), .A(n19927), .ZN(n19952) );
  INV_X1 U13502 ( .A(n19947), .ZN(n19932) );
  INV_X1 U13503 ( .A(n20024), .ZN(n20006) );
  NOR2_X1 U13504 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20067), .ZN(
        n20053) );
  INV_X1 U13505 ( .A(n20038), .ZN(n20086) );
  NAND2_X1 U13506 ( .A1(n20101), .A2(n20100), .ZN(n20117) );
  OAI21_X1 U13507 ( .B1(n20132), .B2(n20131), .A(n20130), .ZN(n20149) );
  AND2_X1 U13508 ( .A1(n20154), .A2(n20183), .ZN(n20177) );
  AOI21_X1 U13509 ( .B1(n20508), .B2(n20188), .A(n20187), .ZN(n20212) );
  AND2_X1 U13510 ( .A1(n20253), .A2(n20288), .ZN(n20294) );
  NOR2_X1 U13511 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20334), .ZN(
        n20321) );
  INV_X1 U13512 ( .A(n19991), .ZN(n20338) );
  INV_X1 U13513 ( .A(n20009), .ZN(n20357) );
  INV_X1 U13514 ( .A(n20018), .ZN(n20376) );
  INV_X1 U13515 ( .A(n20065), .ZN(n20333) );
  NAND2_X1 U13516 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20520) );
  INV_X1 U13517 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20394) );
  AND2_X1 U13518 ( .A1(n13242), .A2(n13241), .ZN(n19466) );
  NOR2_X1 U13519 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17724), .ZN(n17708) );
  INV_X1 U13520 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18091) );
  INV_X1 U13521 ( .A(n17852), .ZN(n17844) );
  NOR2_X1 U13522 ( .A1(n17597), .A2(n17963), .ZN(n17940) );
  INV_X1 U13523 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18050) );
  NOR2_X1 U13524 ( .A1(n18093), .A2(n18237), .ZN(n18173) );
  INV_X1 U13525 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18255) );
  OR4_X1 U13526 ( .A1(n17911), .A2(n17910), .A3(n17909), .A4(n17908), .ZN(
        n17916) );
  OR4_X1 U13527 ( .A1(n14407), .A2(n14406), .A3(n14405), .A4(n14404), .ZN(
        n17932) );
  NOR2_X1 U13528 ( .A1(n18452), .A2(n18352), .ZN(n18347) );
  AND2_X1 U13529 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18407), .ZN(n18394) );
  INV_X1 U13530 ( .A(n18694), .ZN(n18648) );
  INV_X1 U13531 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18425) );
  OR2_X1 U13532 ( .A1(n17082), .A2(n17081), .ZN(n17083) );
  AND2_X1 U13533 ( .A1(n18569), .A2(n13205), .ZN(n18551) );
  INV_X1 U13534 ( .A(n18691), .ZN(n18647) );
  INV_X1 U13535 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18853) );
  INV_X1 U13536 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18913) );
  NOR2_X1 U13537 ( .A1(n18715), .A2(n18947), .ZN(n18911) );
  AND2_X1 U13538 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18994), .ZN(
        n18945) );
  AND2_X1 U13539 ( .A1(n18951), .A2(n19465), .ZN(n19015) );
  INV_X1 U13540 ( .A(n19375), .ZN(n19312) );
  NAND2_X1 U13541 ( .A1(n18425), .A2(n19608), .ZN(n17869) );
  INV_X1 U13542 ( .A(n19130), .ZN(n19123) );
  NOR2_X1 U13543 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19487) );
  NOR2_X1 U13544 ( .A1(n19478), .A2(n19089), .ZN(n19154) );
  INV_X1 U13545 ( .A(n19215), .ZN(n19218) );
  INV_X1 U13546 ( .A(n19231), .ZN(n19239) );
  NOR2_X1 U13547 ( .A1(n19175), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19245) );
  INV_X1 U13548 ( .A(n19304), .ZN(n19308) );
  NOR2_X1 U13549 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n11737), .ZN(
        n19244) );
  INV_X1 U13550 ( .A(n19420), .ZN(n19380) );
  NOR2_X1 U13551 ( .A1(n19478), .A2(n19265), .ZN(n19347) );
  INV_X1 U13552 ( .A(n19342), .ZN(n19455) );
  NOR2_X1 U13553 ( .A1(n19515), .A2(n19512), .ZN(n19621) );
  INV_X1 U13554 ( .A(n19627), .ZN(n19529) );
  INV_X1 U13555 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19537) );
  INV_X1 U13556 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n17481) );
  NAND2_X1 U13557 ( .A1(n13730), .A2(n14038), .ZN(n14231) );
  OR3_X1 U13558 ( .A1(n20560), .A2(n21403), .A3(n21402), .ZN(n15328) );
  INV_X1 U13559 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21676) );
  INV_X1 U13560 ( .A(n20648), .ZN(n15395) );
  INV_X1 U13561 ( .A(n15623), .ZN(n15467) );
  OR2_X1 U13562 ( .A1(n15482), .A2(n15481), .ZN(n15684) );
  AND2_X1 U13563 ( .A1(n14228), .A2(n14227), .ZN(n20797) );
  OR2_X1 U13564 ( .A1(n20683), .A2(n14727), .ZN(n20654) );
  NAND2_X1 U13565 ( .A1(n21369), .A2(n17366), .ZN(n20674) );
  NAND2_X1 U13566 ( .A1(n14038), .A2(n14037), .ZN(n20683) );
  NOR2_X1 U13567 ( .A1(n14231), .A2(n14229), .ZN(n14294) );
  AOI21_X1 U13568 ( .B1(n15586), .B2(n15127), .A(n12265), .ZN(n12650) );
  OR2_X1 U13569 ( .A1(n20703), .A2(n14034), .ZN(n20714) );
  XNOR2_X1 U13570 ( .A(n15531), .B(n15717), .ZN(n15722) );
  INV_X1 U13571 ( .A(n20742), .ZN(n20760) );
  NAND2_X1 U13572 ( .A1(n13502), .A2(n13367), .ZN(n20753) );
  OAI21_X1 U13573 ( .B1(n17333), .B2(n20736), .A(n15850), .ZN(n20733) );
  INV_X1 U13574 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21474) );
  NAND2_X1 U13575 ( .A1(n13834), .A2(n13833), .ZN(n21457) );
  OR2_X1 U13576 ( .A1(n20897), .A2(n20938), .ZN(n20854) );
  OR2_X1 U13577 ( .A1(n20897), .A2(n20974), .ZN(n20883) );
  OR2_X1 U13578 ( .A1(n20897), .A2(n20889), .ZN(n20942) );
  NAND2_X1 U13579 ( .A1(n21034), .A2(n21197), .ZN(n20995) );
  NAND2_X1 U13580 ( .A1(n21034), .A2(n21252), .ZN(n21064) );
  NAND2_X1 U13581 ( .A1(n21164), .A2(n21197), .ZN(n21115) );
  NAND2_X1 U13582 ( .A1(n21164), .A2(n21226), .ZN(n21157) );
  NAND2_X1 U13583 ( .A1(n21164), .A2(n21252), .ZN(n21188) );
  NAND2_X1 U13584 ( .A1(n21164), .A2(n21163), .ZN(n21225) );
  NAND2_X1 U13585 ( .A1(n21311), .A2(n21226), .ZN(n21262) );
  NAND2_X1 U13586 ( .A1(n21311), .A2(n21252), .ZN(n21366) );
  INV_X1 U13587 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21660) );
  INV_X1 U13588 ( .A(n21448), .ZN(n21452) );
  NAND2_X1 U13589 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21487) );
  INV_X1 U13590 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21403) );
  NAND2_X1 U13591 ( .A1(n21439), .A2(n21388), .ZN(n21436) );
  INV_X1 U13592 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20512) );
  OR2_X1 U13593 ( .A1(n15042), .A2(n14980), .ZN(n16254) );
  AND2_X1 U13594 ( .A1(n13012), .A2(n13011), .ZN(n13013) );
  OR2_X1 U13595 ( .A1(n16451), .A2(n11133), .ZN(n16462) );
  OR2_X1 U13596 ( .A1(n16451), .A2(n14524), .ZN(n16468) );
  INV_X1 U13597 ( .A(n16451), .ZN(n14604) );
  AND2_X1 U13598 ( .A1(n16462), .A2(n16468), .ZN(n16475) );
  AND2_X1 U13599 ( .A1(n14925), .A2(n14924), .ZN(n19713) );
  NAND2_X1 U13600 ( .A1(n19745), .A2(n20511), .ZN(n13809) );
  INV_X1 U13601 ( .A(n19745), .ZN(n19742) );
  OR2_X1 U13602 ( .A1(n15032), .A2(n11002), .ZN(n15037) );
  NOR2_X1 U13603 ( .A1(n13330), .A2(n13329), .ZN(n13331) );
  NAND2_X1 U13604 ( .A1(n13728), .A2(n11507), .ZN(n17388) );
  XNOR2_X1 U13605 ( .A(n11562), .B(n10407), .ZN(n14922) );
  INV_X1 U13606 ( .A(n19796), .ZN(n16942) );
  INV_X1 U13607 ( .A(n20495), .ZN(n20498) );
  INV_X1 U13608 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19819) );
  AOI211_X2 U13609 ( .C1(n17030), .C2(n17026), .A(n17025), .B(n17024), .ZN(
        n19857) );
  NAND2_X1 U13610 ( .A1(n20123), .A2(n20059), .ZN(n19918) );
  AND2_X1 U13611 ( .A1(n19963), .A2(n19962), .ZN(n19972) );
  INV_X1 U13612 ( .A(n19968), .ZN(n19990) );
  NAND2_X1 U13613 ( .A1(n20059), .A2(n20250), .ZN(n20058) );
  NAND2_X1 U13614 ( .A1(n20065), .A2(n20059), .ZN(n20121) );
  INV_X1 U13615 ( .A(n20354), .ZN(n20271) );
  AOI22_X1 U13616 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19844), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19845), .ZN(n20308) );
  AOI221_X2 U13617 ( .B1(n20333), .B2(n20334), .C1(n20332), .C2(n20334), .A(
        n20331), .ZN(n20392) );
  INV_X1 U13618 ( .A(n20475), .ZN(n20393) );
  INV_X1 U13619 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20412) );
  INV_X1 U13620 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20437) );
  NAND2_X1 U13621 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20462), .ZN(n20458) );
  INV_X1 U13622 ( .A(n20462), .ZN(n20526) );
  INV_X1 U13623 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19625) );
  OR3_X1 U13624 ( .A1(n19566), .A2(n19563), .A3(n17682), .ZN(n17660) );
  INV_X1 U13625 ( .A(n17837), .ZN(n17823) );
  INV_X1 U13626 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17832) );
  AND2_X1 U13627 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17945), .ZN(n17939) );
  NOR2_X1 U13628 ( .A1(n17633), .A2(n17999), .ZN(n18015) );
  NAND2_X1 U13629 ( .A1(n18279), .A2(n18364), .ZN(n18269) );
  INV_X1 U13630 ( .A(n18276), .ZN(n18271) );
  INV_X1 U13631 ( .A(n18351), .ZN(n18363) );
  NAND2_X1 U13632 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18394), .ZN(n18392) );
  INV_X1 U13633 ( .A(n14692), .ZN(n18405) );
  AND2_X1 U13634 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18423), .ZN(n18418) );
  INV_X1 U13635 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18427) );
  INV_X1 U13636 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18444) );
  INV_X1 U13637 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18470) );
  OR2_X1 U13638 ( .A1(n19623), .A2(n18475), .ZN(n18477) );
  INV_X1 U13639 ( .A(n18533), .ZN(n18528) );
  INV_X1 U13640 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21610) );
  INV_X1 U13641 ( .A(n18790), .ZN(n18776) );
  INV_X1 U13642 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18887) );
  AOI22_X1 U13643 ( .A1(n17235), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n18895), .B2(n17234), .ZN(n17238) );
  INV_X1 U13644 ( .A(n19002), .ZN(n18976) );
  INV_X1 U13645 ( .A(n18951), .ZN(n19006) );
  INV_X1 U13646 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19018) );
  INV_X1 U13647 ( .A(n19015), .ZN(n17248) );
  INV_X1 U13648 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19494) );
  NAND2_X1 U13649 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19245), .ZN(
        n19282) );
  INV_X1 U13650 ( .A(n19433), .ZN(n19328) );
  NAND2_X1 U13651 ( .A1(n19409), .A2(BUF2_REG_23__SCAN_IN), .ZN(n19342) );
  INV_X1 U13652 ( .A(n19376), .ZN(n19413) );
  INV_X1 U13653 ( .A(n19296), .ZN(n19432) );
  NAND2_X1 U13654 ( .A1(n19483), .A2(n19346), .ZN(n19462) );
  INV_X1 U13655 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19608) );
  OAI21_X1 U13656 ( .B1(n19527), .B2(n17481), .A(n19523), .ZN(n19605) );
  INV_X1 U13657 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19543) );
  INV_X1 U13658 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19558) );
  OR2_X1 U13659 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n17481), .ZN(n19616) );
  INV_X1 U13660 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19049) );
  INV_X1 U13661 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19040) );
  INV_X1 U13662 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19062) );
  INV_X1 U13663 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19029) );
  INV_X1 U13664 ( .A(n17444), .ZN(n17433) );
  NAND2_X1 U13665 ( .A1(n13580), .A2(n10399), .ZN(P2_U2988) );
  OAI21_X1 U13666 ( .B1(n16785), .B2(n19785), .A(n13331), .ZN(P2_U2996) );
  OAI21_X1 U13667 ( .B1(n14922), .B2(n17400), .A(n11575), .ZN(P2_U3025) );
  NAND3_X1 U13668 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(n13704), .A3(n21445), .ZN(
        U214) );
  INV_X1 U13669 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10430) );
  OR2_X2 U13670 ( .A1(n12906), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12832) );
  OR2_X2 U13671 ( .A1(n12906), .A2(n10715), .ZN(n12808) );
  INV_X1 U13672 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10429) );
  OAI22_X1 U13673 ( .A1(n10430), .A2(n12832), .B1(n12808), .B2(n10429), .ZN(
        n10431) );
  INV_X1 U13674 ( .A(n10431), .ZN(n10441) );
  AND2_X4 U13675 ( .A1(n10445), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10724) );
  AOI22_X1 U13676 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10440) );
  BUF_X4 U13677 ( .A(n10724), .Z(n14480) );
  AND2_X2 U13678 ( .A1(n14480), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10840) );
  AND2_X2 U13679 ( .A1(n12911), .A2(n10715), .ZN(n10495) );
  INV_X1 U13680 ( .A(n10495), .ZN(n10851) );
  AOI22_X1 U13681 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10439) );
  INV_X1 U13682 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10436) );
  AND2_X1 U13683 ( .A1(n16991), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U13684 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10435) );
  AND2_X1 U13685 ( .A1(n14462), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10433) );
  AND2_X2 U13686 ( .A1(n12849), .A2(n10433), .ZN(n12842) );
  NAND2_X1 U13687 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10434) );
  OAI211_X1 U13688 ( .C1(n10559), .C2(n10436), .A(n10435), .B(n10434), .ZN(
        n10437) );
  INV_X1 U13689 ( .A(n10437), .ZN(n10438) );
  NAND4_X1 U13690 ( .A1(n10441), .A2(n10440), .A3(n10439), .A4(n10438), .ZN(
        n10451) );
  AND2_X4 U13691 ( .A1(n10445), .A2(n10317), .ZN(n10722) );
  AND2_X2 U13692 ( .A1(n12911), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10551) );
  AOI22_X1 U13693 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10519), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10449) );
  AND3_X4 U13694 ( .A1(n10443), .A2(n10442), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U13695 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10448) );
  INV_X2 U13696 ( .A(n9736), .ZN(n12828) );
  AOI22_X1 U13697 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12841), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10447) );
  AND2_X2 U13698 ( .A1(n9706), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10847) );
  NAND2_X1 U13699 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10446) );
  NAND4_X1 U13700 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10450) );
  INV_X1 U13701 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14164) );
  INV_X2 U13702 ( .A(n12858), .ZN(n12993) );
  AOI22_X1 U13703 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13704 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13705 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9710), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13706 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13707 ( .A1(n12993), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13708 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9710), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13709 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13710 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9706), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10456) );
  MUX2_X1 U13711 ( .A(n11159), .B(n14164), .S(n9700), .Z(n10931) );
  AOI22_X1 U13712 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10840), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13713 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10462) );
  INV_X2 U13714 ( .A(n10853), .ZN(n12841) );
  AOI22_X1 U13715 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12842), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U13716 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10460) );
  INV_X1 U13717 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10465) );
  INV_X1 U13718 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10788) );
  OAI22_X1 U13719 ( .A1(n10465), .A2(n10559), .B1(n12808), .B2(n10788), .ZN(
        n10466) );
  INV_X1 U13720 ( .A(n10466), .ZN(n10473) );
  INV_X2 U13721 ( .A(n10404), .ZN(n12834) );
  AOI22_X1 U13722 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10519), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10472) );
  INV_X1 U13723 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U13724 ( .A1(n12828), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13725 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10467) );
  OAI211_X1 U13726 ( .C1(n12832), .C2(n10469), .A(n10468), .B(n10467), .ZN(
        n10470) );
  INV_X1 U13727 ( .A(n10470), .ZN(n10471) );
  NAND2_X1 U13728 ( .A1(n11001), .A2(n10998), .ZN(n10476) );
  NAND2_X1 U13729 ( .A1(n20252), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10475) );
  NAND2_X1 U13730 ( .A1(n10476), .A2(n10475), .ZN(n10512) );
  XNOR2_X1 U13731 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13732 ( .A1(n10512), .A2(n10511), .ZN(n10513) );
  NAND2_X1 U13733 ( .A1(n20497), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10477) );
  NAND2_X1 U13734 ( .A1(n10513), .A2(n10477), .ZN(n11009) );
  INV_X1 U13735 ( .A(n11008), .ZN(n10478) );
  XNOR2_X1 U13736 ( .A(n11009), .B(n10478), .ZN(n11013) );
  AOI22_X1 U13737 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U13738 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9703), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13739 ( .A1(n12986), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13740 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10479) );
  NAND4_X1 U13741 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10483) );
  AOI22_X1 U13742 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13743 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9704), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13744 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13745 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10488) );
  MUX2_X1 U13746 ( .A(n11163), .B(n11013), .S(n14983), .Z(n11032) );
  INV_X1 U13747 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10491) );
  INV_X1 U13748 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10493) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10492) );
  OAI22_X1 U13750 ( .A1(n10493), .A2(n12832), .B1(n10559), .B2(n10492), .ZN(
        n10494) );
  INV_X1 U13751 ( .A(n10494), .ZN(n10504) );
  AOI22_X1 U13752 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10519), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10502) );
  INV_X1 U13754 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13755 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10498) );
  NAND2_X1 U13756 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10497) );
  OAI211_X1 U13757 ( .C1(n12808), .C2(n10499), .A(n10498), .B(n10497), .ZN(
        n10500) );
  INV_X1 U13758 ( .A(n10500), .ZN(n10501) );
  NAND4_X1 U13759 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10510) );
  AOI22_X1 U13760 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10840), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13761 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13762 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13763 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10505) );
  NAND4_X1 U13764 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10509) );
  NOR2_X1 U13765 ( .A1(n10510), .A2(n10509), .ZN(n11152) );
  INV_X1 U13766 ( .A(n11152), .ZN(n10516) );
  OR2_X1 U13767 ( .A1(n10512), .A2(n10511), .ZN(n10514) );
  NAND2_X1 U13768 ( .A1(n14983), .A2(n11044), .ZN(n10515) );
  OAI21_X1 U13769 ( .B1(n10516), .B2(n14983), .A(n10515), .ZN(n11030) );
  NOR2_X1 U13770 ( .A1(n10980), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10923) );
  INV_X1 U13771 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13792) );
  NAND2_X1 U13772 ( .A1(n10923), .A2(n13792), .ZN(n10539) );
  AOI22_X1 U13773 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13774 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13775 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10519), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13776 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13777 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12841), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U13778 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10520) );
  NAND4_X1 U13779 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10534) );
  INV_X1 U13780 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10526) );
  NAND2_X1 U13781 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10525) );
  NAND2_X1 U13782 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10524) );
  OAI211_X1 U13783 ( .C1(n10559), .C2(n10526), .A(n10525), .B(n10524), .ZN(
        n10527) );
  INV_X1 U13784 ( .A(n10527), .ZN(n10532) );
  INV_X1 U13785 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10529) );
  INV_X1 U13786 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10528) );
  OAI22_X1 U13787 ( .A1(n10529), .A2(n12832), .B1(n12808), .B2(n10528), .ZN(
        n10530) );
  INV_X1 U13788 ( .A(n10530), .ZN(n10531) );
  NAND3_X1 U13789 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n11142) );
  NAND2_X1 U13790 ( .A1(n11142), .A2(n10980), .ZN(n10538) );
  NOR2_X2 U13791 ( .A1(n10916), .A2(n10919), .ZN(n10912) );
  NAND2_X1 U13792 ( .A1(n10540), .A2(n10912), .ZN(n10930) );
  INV_X1 U13793 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10541) );
  INV_X1 U13794 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10871) );
  OAI22_X1 U13795 ( .A1(n10541), .A2(n12832), .B1(n12808), .B2(n10871), .ZN(
        n10542) );
  INV_X1 U13796 ( .A(n10542), .ZN(n10550) );
  AOI22_X1 U13797 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13798 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10548) );
  INV_X1 U13799 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U13800 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10544) );
  NAND2_X1 U13801 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10543) );
  OAI211_X1 U13802 ( .C1(n10559), .C2(n10545), .A(n10544), .B(n10543), .ZN(
        n10546) );
  INV_X1 U13803 ( .A(n10546), .ZN(n10547) );
  NAND4_X1 U13804 ( .A1(n10550), .A2(n10549), .A3(n10548), .A4(n10547), .ZN(
        n10557) );
  AOI22_X1 U13805 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10519), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13806 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13807 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n12841), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U13808 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10552) );
  NAND4_X1 U13809 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10556) );
  NOR2_X2 U13810 ( .A1(n10930), .A2(n10941), .ZN(n10905) );
  INV_X1 U13811 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10574) );
  INV_X1 U13812 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10887) );
  INV_X1 U13813 ( .A(n10839), .ZN(n10581) );
  INV_X1 U13814 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10886) );
  OAI22_X1 U13815 ( .A1(n10887), .A2(n12808), .B1(n10581), .B2(n10886), .ZN(
        n10558) );
  INV_X1 U13816 ( .A(n10558), .ZN(n10567) );
  INV_X1 U13817 ( .A(n10559), .ZN(n12835) );
  AOI22_X1 U13818 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13819 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10495), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10565) );
  INV_X1 U13820 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10562) );
  NAND2_X1 U13821 ( .A1(n12828), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10561) );
  NAND2_X1 U13822 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10560) );
  OAI211_X1 U13823 ( .C1(n12832), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        n10563) );
  INV_X1 U13824 ( .A(n10563), .ZN(n10564) );
  NAND4_X1 U13825 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10573) );
  AOI22_X1 U13826 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12724), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13828 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12842), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U13829 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10568) );
  NAND4_X1 U13830 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10572) );
  AND2_X2 U13831 ( .A1(n10905), .A2(n10906), .ZN(n10904) );
  INV_X1 U13832 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10576) );
  INV_X1 U13833 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10575) );
  OAI22_X1 U13834 ( .A1(n10576), .A2(n10559), .B1(n12808), .B2(n10575), .ZN(
        n10577) );
  INV_X1 U13835 ( .A(n10577), .ZN(n10586) );
  AOI22_X1 U13836 ( .A1(n11284), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13837 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10495), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10584) );
  INV_X1 U13838 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13839 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10579) );
  NAND2_X1 U13840 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10578) );
  OAI211_X1 U13841 ( .C1(n10581), .C2(n10580), .A(n10579), .B(n10578), .ZN(
        n10582) );
  INV_X1 U13842 ( .A(n10582), .ZN(n10583) );
  NAND4_X1 U13843 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10592) );
  AOI22_X1 U13844 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12724), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13845 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13846 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12841), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10588) );
  INV_X1 U13847 ( .A(n11209), .ZN(n10852) );
  NAND4_X1 U13848 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10591) );
  INV_X1 U13849 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10593) );
  MUX2_X1 U13850 ( .A(n10606), .B(n10593), .S(n19834), .Z(n10953) );
  NOR2_X1 U13851 ( .A1(n10980), .A2(n16157), .ZN(n10951) );
  INV_X1 U13852 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n16132) );
  INV_X1 U13853 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n14311) );
  NAND2_X1 U13854 ( .A1(n10672), .A2(n14311), .ZN(n10655) );
  NAND2_X1 U13855 ( .A1(n19834), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10653) );
  INV_X1 U13856 ( .A(n10643), .ZN(n10597) );
  NOR2_X1 U13857 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n10596) );
  NAND2_X1 U13858 ( .A1(n10597), .A2(n10402), .ZN(n10649) );
  INV_X1 U13859 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14666) );
  NOR2_X1 U13860 ( .A1(n10980), .A2(n14666), .ZN(n10636) );
  NOR2_X2 U13861 ( .A1(n10649), .A2(n10636), .ZN(n10630) );
  NAND2_X1 U13862 ( .A1(n9700), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10631) );
  INV_X1 U13863 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10598) );
  NOR2_X1 U13864 ( .A1(n10980), .A2(n10598), .ZN(n10657) );
  INV_X1 U13865 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10599) );
  NOR2_X1 U13866 ( .A1(n10980), .A2(n10599), .ZN(n10640) );
  INV_X1 U13867 ( .A(n10640), .ZN(n10600) );
  INV_X1 U13868 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13869 ( .A1(n10623), .A2(n10601), .ZN(n10617) );
  NAND2_X1 U13870 ( .A1(n10617), .A2(n10959), .ZN(n10622) );
  NAND2_X1 U13871 ( .A1(n19834), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10618) );
  INV_X1 U13872 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10602) );
  NOR2_X1 U13873 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_EBX_REG_26__SCAN_IN), 
        .ZN(n10603) );
  NAND2_X1 U13874 ( .A1(n15967), .A2(n10603), .ZN(n10690) );
  INV_X1 U13875 ( .A(n10687), .ZN(n14891) );
  INV_X1 U13876 ( .A(n15967), .ZN(n10613) );
  INV_X1 U13877 ( .A(n10608), .ZN(n15961) );
  AND2_X1 U13878 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10605) );
  NAND2_X1 U13879 ( .A1(n15961), .A2(n10605), .ZN(n10984) );
  INV_X1 U13880 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10607) );
  OAI21_X1 U13881 ( .B1(n10608), .B2(n10961), .A(n10607), .ZN(n10609) );
  INV_X1 U13882 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15979) );
  NOR2_X1 U13883 ( .A1(n10980), .A2(n15979), .ZN(n10610) );
  INV_X1 U13884 ( .A(n10959), .ZN(n10635) );
  AOI21_X1 U13885 ( .B1(n10611), .B2(n10610), .A(n10635), .ZN(n10612) );
  INV_X1 U13886 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13029) );
  NAND2_X1 U13887 ( .A1(n10620), .A2(n13029), .ZN(n13021) );
  XNOR2_X1 U13888 ( .A(n10614), .B(n10416), .ZN(n15998) );
  NAND2_X1 U13889 ( .A1(n15998), .A2(n11177), .ZN(n13018) );
  INV_X1 U13890 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16732) );
  NAND2_X1 U13891 ( .A1(n13018), .A2(n16732), .ZN(n10615) );
  NAND2_X1 U13892 ( .A1(n10959), .A2(n11177), .ZN(n10985) );
  NAND2_X1 U13893 ( .A1(n10985), .A2(n16717), .ZN(n16506) );
  NAND2_X1 U13894 ( .A1(n10617), .A2(n10211), .ZN(n10619) );
  NAND2_X1 U13895 ( .A1(n10614), .A2(n10619), .ZN(n16014) );
  NOR2_X1 U13896 ( .A1(n16538), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10662) );
  INV_X1 U13897 ( .A(n10620), .ZN(n10621) );
  INV_X1 U13898 ( .A(n10622), .ZN(n10625) );
  INV_X1 U13899 ( .A(n10623), .ZN(n10629) );
  NAND3_X1 U13900 ( .A1(n10629), .A2(n19834), .A3(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n10624) );
  NAND2_X1 U13901 ( .A1(n10625), .A2(n10624), .ZN(n16017) );
  INV_X1 U13902 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11564) );
  NOR2_X1 U13903 ( .A1(n10663), .A2(n11564), .ZN(n16549) );
  INV_X1 U13904 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n19666) );
  NOR2_X1 U13905 ( .A1(n10980), .A2(n19666), .ZN(n10627) );
  AOI21_X1 U13906 ( .B1(n10626), .B2(n10627), .A(n10635), .ZN(n10628) );
  INV_X1 U13907 ( .A(n10630), .ZN(n10632) );
  XNOR2_X1 U13908 ( .A(n10632), .B(n10631), .ZN(n16059) );
  AND2_X1 U13909 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10633) );
  NAND2_X1 U13910 ( .A1(n16059), .A2(n10633), .ZN(n14754) );
  INV_X1 U13911 ( .A(n10649), .ZN(n10634) );
  NAND2_X1 U13912 ( .A1(n10634), .A2(n14666), .ZN(n10638) );
  AOI21_X1 U13913 ( .B1(n10649), .B2(n10636), .A(n10635), .ZN(n10637) );
  AND2_X1 U13914 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10639) );
  NAND2_X1 U13915 ( .A1(n16073), .A2(n10639), .ZN(n14756) );
  NAND2_X1 U13916 ( .A1(n14754), .A2(n14756), .ZN(n16544) );
  NAND2_X1 U13917 ( .A1(n9741), .A2(n10640), .ZN(n10641) );
  NAND2_X1 U13918 ( .A1(n10626), .A2(n10641), .ZN(n16028) );
  NAND2_X1 U13919 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10642) );
  NAND2_X1 U13920 ( .A1(n19834), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10644) );
  MUX2_X1 U13921 ( .A(n9700), .B(n10644), .S(n10645), .Z(n10646) );
  OR2_X1 U13922 ( .A1(n10645), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10648) );
  AND2_X1 U13923 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10647) );
  NAND2_X1 U13924 ( .A1(n16092), .A2(n10647), .ZN(n16597) );
  NAND3_X1 U13925 ( .A1(n10648), .A2(n9700), .A3(P2_EBX_REG_15__SCAN_IN), .ZN(
        n10650) );
  AND2_X1 U13926 ( .A1(n10650), .A2(n10649), .ZN(n10670) );
  AND2_X1 U13927 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10651) );
  NAND2_X1 U13928 ( .A1(n10670), .A2(n10651), .ZN(n16584) );
  NAND2_X1 U13929 ( .A1(n16597), .A2(n16584), .ZN(n16545) );
  XNOR2_X1 U13930 ( .A(n10652), .B(n10410), .ZN(n16103) );
  NOR2_X1 U13931 ( .A1(n16545), .A2(n16542), .ZN(n12652) );
  INV_X1 U13932 ( .A(n10653), .ZN(n10654) );
  NAND2_X1 U13933 ( .A1(n10655), .A2(n10654), .ZN(n10656) );
  NAND2_X1 U13934 ( .A1(n10652), .A2(n10656), .ZN(n16106) );
  NAND2_X1 U13935 ( .A1(n10658), .A2(n10657), .ZN(n10659) );
  AND2_X1 U13936 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10660) );
  NAND2_X1 U13937 ( .A1(n16048), .A2(n10660), .ZN(n16543) );
  NAND4_X1 U13938 ( .A1(n16541), .A2(n12652), .A3(n16620), .A4(n16543), .ZN(
        n10661) );
  NOR4_X1 U13939 ( .A1(n16549), .A2(n11560), .A3(n16544), .A4(n10661), .ZN(
        n13015) );
  OAI211_X1 U13940 ( .C1(n10662), .C2(n13018), .A(n13022), .B(n13015), .ZN(
        n11531) );
  INV_X1 U13941 ( .A(n11531), .ZN(n10694) );
  INV_X1 U13942 ( .A(n10663), .ZN(n10664) );
  NOR2_X1 U13943 ( .A1(n10664), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11561) );
  INV_X1 U13944 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16758) );
  INV_X1 U13945 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U13946 ( .A1(n10666), .A2(n12664), .ZN(n12657) );
  NAND2_X1 U13947 ( .A1(n16092), .A2(n11177), .ZN(n10667) );
  INV_X1 U13948 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16817) );
  NAND2_X1 U13949 ( .A1(n10667), .A2(n16817), .ZN(n16598) );
  INV_X1 U13950 ( .A(n10668), .ZN(n10669) );
  INV_X1 U13951 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16829) );
  NAND2_X1 U13952 ( .A1(n10669), .A2(n16829), .ZN(n16606) );
  INV_X1 U13953 ( .A(n10670), .ZN(n16081) );
  INV_X1 U13954 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16799) );
  OAI21_X1 U13955 ( .B1(n16081), .B2(n10961), .A(n16799), .ZN(n16585) );
  INV_X1 U13956 ( .A(n10671), .ZN(n10675) );
  INV_X1 U13957 ( .A(n10672), .ZN(n10673) );
  NAND3_X1 U13958 ( .A1(n10673), .A2(n9699), .A3(P2_EBX_REG_11__SCAN_IN), .ZN(
        n10674) );
  NAND2_X1 U13959 ( .A1(n16125), .A2(n11177), .ZN(n10975) );
  INV_X1 U13960 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16863) );
  NAND2_X1 U13961 ( .A1(n10975), .A2(n16863), .ZN(n16634) );
  NAND2_X1 U13962 ( .A1(n16634), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10676) );
  OR2_X1 U13963 ( .A1(n16106), .A2(n10961), .ZN(n11555) );
  NAND2_X1 U13964 ( .A1(n10676), .A2(n11555), .ZN(n10677) );
  AND4_X1 U13965 ( .A1(n16598), .A2(n16606), .A3(n16585), .A4(n10677), .ZN(
        n10682) );
  NAND2_X1 U13966 ( .A1(n16048), .A2(n11177), .ZN(n10678) );
  INV_X1 U13967 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16776) );
  NAND2_X1 U13968 ( .A1(n10678), .A2(n16776), .ZN(n13314) );
  NAND2_X1 U13969 ( .A1(n16073), .A2(n11177), .ZN(n10679) );
  XNOR2_X1 U13970 ( .A(n10679), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12656) );
  NAND2_X1 U13971 ( .A1(n16059), .A2(n11177), .ZN(n10680) );
  NAND2_X1 U13972 ( .A1(n10680), .A2(n10038), .ZN(n14755) );
  NAND2_X1 U13973 ( .A1(n12656), .A2(n14755), .ZN(n11556) );
  INV_X1 U13974 ( .A(n11556), .ZN(n10681) );
  NAND4_X1 U13975 ( .A1(n12657), .A2(n10682), .A3(n13314), .A4(n10681), .ZN(
        n10683) );
  NAND2_X1 U13976 ( .A1(n19834), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10688) );
  INV_X1 U13977 ( .A(n10688), .ZN(n10689) );
  NAND2_X1 U13978 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NAND2_X1 U13979 ( .A1(n10981), .A2(n10691), .ZN(n15943) );
  NOR2_X1 U13980 ( .A1(n15943), .A2(n10961), .ZN(n11533) );
  INV_X1 U13981 ( .A(n11533), .ZN(n10693) );
  INV_X1 U13982 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10692) );
  INV_X1 U13983 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U13984 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9703), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13985 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13986 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10695) );
  NAND4_X1 U13987 ( .A1(n10698), .A2(n10697), .A3(n10696), .A4(n10695), .ZN(
        n10699) );
  NAND2_X1 U13988 ( .A1(n10699), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10706) );
  AOI22_X1 U13989 ( .A1(n12993), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13990 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9704), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13991 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13992 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13993 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10704) );
  NAND2_X1 U13994 ( .A1(n10704), .A2(n10715), .ZN(n10705) );
  AOI22_X1 U13995 ( .A1(n12993), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13996 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9704), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13997 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9710), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13998 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13999 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U14000 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9703), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U14001 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U14002 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10711) );
  INV_X1 U14003 ( .A(n11117), .ZN(n10753) );
  NAND2_X1 U14004 ( .A1(n11133), .A2(n11451), .ZN(n10730) );
  AOI22_X1 U14005 ( .A1(n12993), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U14006 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9704), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U14007 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10716) );
  NAND4_X1 U14008 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10720) );
  AOI22_X1 U14009 ( .A1(n12986), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U14010 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9703), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U14011 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U14012 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10725) );
  NAND4_X1 U14013 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10729) );
  AND2_X1 U14014 ( .A1(n10734), .A2(n11127), .ZN(n10735) );
  NAND2_X1 U14015 ( .A1(n11035), .A2(n10735), .ZN(n11120) );
  INV_X1 U14016 ( .A(n10747), .ZN(n10736) );
  NAND3_X1 U14017 ( .A1(n11120), .A2(n20511), .A3(n10736), .ZN(n10737) );
  INV_X1 U14018 ( .A(n11055), .ZN(n10740) );
  NAND2_X1 U14019 ( .A1(n10740), .A2(n10739), .ZN(n11060) );
  AND2_X1 U14020 ( .A1(n10761), .A2(n14979), .ZN(n10743) );
  NAND2_X1 U14021 ( .A1(n10762), .A2(n10743), .ZN(n10744) );
  AND2_X2 U14022 ( .A1(n19834), .A2(n14524), .ZN(n11126) );
  AOI22_X1 U14023 ( .A1(n14476), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n14511), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10748) );
  INV_X1 U14024 ( .A(n10750), .ZN(n10751) );
  NAND2_X1 U14025 ( .A1(n10751), .A2(n11131), .ZN(n11116) );
  INV_X1 U14026 ( .A(n11116), .ZN(n10754) );
  INV_X1 U14027 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10758) );
  INV_X1 U14028 ( .A(n14511), .ZN(n10760) );
  NAND2_X1 U14029 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10759) );
  NAND3_X1 U14030 ( .A1(n10762), .A2(n10761), .A3(n11455), .ZN(n10763) );
  INV_X1 U14031 ( .A(n14447), .ZN(n10765) );
  AOI22_X1 U14032 ( .A1(n10765), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n14511), .ZN(n10766) );
  OAI21_X1 U14033 ( .B1(n20497), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16993), 
        .ZN(n10768) );
  OAI21_X1 U14034 ( .B1(n20414), .B2(n11440), .A(n10769), .ZN(n10770) );
  BUF_X8 U14035 ( .A(n10757), .Z(n14898) );
  INV_X1 U14036 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U14037 ( .A1(n11438), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10771) );
  AOI22_X1 U14038 ( .A1(n10774), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n14511), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10775) );
  INV_X1 U14039 ( .A(n10781), .ZN(n10779) );
  AND2_X1 U14040 ( .A1(n10810), .A2(n10806), .ZN(n10780) );
  INV_X1 U14041 ( .A(n10782), .ZN(n10793) );
  AND2_X1 U14042 ( .A1(n10810), .A2(n10799), .ZN(n10783) );
  INV_X1 U14043 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10784) );
  OAI22_X1 U14044 ( .A1(n11246), .A2(n10867), .B1(n10868), .B2(n10784), .ZN(
        n10790) );
  BUF_X4 U14045 ( .A(n10785), .Z(n12681) );
  AND2_X1 U14046 ( .A1(n12681), .A2(n10799), .ZN(n10786) );
  AND2_X1 U14047 ( .A1(n12681), .A2(n10806), .ZN(n10787) );
  OAI22_X1 U14048 ( .A1(n10788), .A2(n10870), .B1(n10888), .B2(n20363), .ZN(
        n10789) );
  NOR2_X1 U14049 ( .A1(n10790), .A2(n10789), .ZN(n10798) );
  INV_X1 U14050 ( .A(n10792), .ZN(n10794) );
  NAND2_X1 U14051 ( .A1(n10794), .A2(n10793), .ZN(n10795) );
  NOR2_X1 U14052 ( .A1(n16966), .A2(n19788), .ZN(n10796) );
  AOI22_X1 U14054 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10864), .B1(
        n17033), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U14055 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19892), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U14056 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10877), .B1(
        n20061), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10800) );
  INV_X1 U14057 ( .A(n16966), .ZN(n10802) );
  NAND2_X1 U14058 ( .A1(n20099), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10805) );
  NAND2_X1 U14059 ( .A1(n10878), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10804) );
  AOI22_X1 U14061 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19926), .B1(
        n10876), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10815) );
  AND2_X1 U14062 ( .A1(n10810), .A2(n16966), .ZN(n10811) );
  AND2_X1 U14063 ( .A1(n12681), .A2(n16966), .ZN(n10812) );
  INV_X1 U14064 ( .A(n11163), .ZN(n10817) );
  NAND2_X1 U14065 ( .A1(n10817), .A2(n11051), .ZN(n10818) );
  AND2_X1 U14066 ( .A1(n20156), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10821) );
  INV_X1 U14067 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11203) );
  INV_X1 U14068 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10819) );
  OAI22_X1 U14069 ( .A1(n11203), .A2(n10867), .B1(n10868), .B2(n10819), .ZN(
        n10820) );
  NOR2_X1 U14070 ( .A1(n10821), .A2(n10820), .ZN(n10825) );
  AOI22_X1 U14071 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19892), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U14072 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10864), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U14073 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20061), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U14074 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17033), .B1(
        n19926), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U14075 ( .A1(n20099), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10827) );
  NAND2_X1 U14076 ( .A1(n10878), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10826) );
  INV_X1 U14077 ( .A(n10876), .ZN(n20036) );
  INV_X1 U14078 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11199) );
  INV_X1 U14079 ( .A(n10870), .ZN(n10829) );
  AOI21_X1 U14080 ( .B1(n10829), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n11051), .ZN(n10831) );
  INV_X1 U14081 ( .A(n10888), .ZN(n20329) );
  NAND2_X1 U14082 ( .A1(n20329), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10830) );
  OAI211_X1 U14083 ( .C1(n20036), .C2(n11199), .A(n10831), .B(n10830), .ZN(
        n10832) );
  INV_X1 U14084 ( .A(n10832), .ZN(n10833) );
  AOI22_X1 U14085 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U14086 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10837) );
  INV_X1 U14087 ( .A(n12808), .ZN(n12827) );
  NAND2_X1 U14088 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10836) );
  NAND2_X1 U14089 ( .A1(n11284), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10835) );
  NAND4_X1 U14090 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10846) );
  NAND2_X1 U14091 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U14092 ( .A1(n10840), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10843) );
  NAND2_X1 U14093 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U14094 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10841) );
  NAND4_X1 U14095 ( .A1(n10844), .A2(n10843), .A3(n10842), .A4(n10841), .ZN(
        n10845) );
  NOR2_X1 U14096 ( .A1(n10846), .A2(n10845), .ZN(n10860) );
  INV_X1 U14097 ( .A(n10847), .ZN(n11048) );
  INV_X1 U14098 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10849) );
  INV_X1 U14099 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21583) );
  OAI22_X1 U14100 ( .A1(n11048), .A2(n10849), .B1(n10848), .B2(n21583), .ZN(
        n10859) );
  INV_X1 U14101 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12706) );
  INV_X1 U14102 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10850) );
  OAI22_X1 U14103 ( .A1(n10851), .A2(n12706), .B1(n10404), .B2(n10850), .ZN(
        n10858) );
  INV_X1 U14104 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11182) );
  NOR2_X1 U14105 ( .A1(n10852), .A2(n11182), .ZN(n10856) );
  INV_X1 U14106 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10854) );
  INV_X1 U14107 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19971) );
  INV_X1 U14108 ( .A(n11137), .ZN(n10861) );
  NAND2_X1 U14109 ( .A1(n17396), .A2(n11142), .ZN(n11077) );
  NAND2_X1 U14110 ( .A1(n11077), .A2(n11152), .ZN(n10862) );
  AOI22_X1 U14111 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10864), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10875) );
  INV_X1 U14112 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21703) );
  INV_X1 U14113 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10869) );
  OAI22_X1 U14114 ( .A1(n21703), .A2(n20186), .B1(n10868), .B2(n10869), .ZN(
        n10873) );
  INV_X1 U14115 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12807) );
  OAI22_X1 U14116 ( .A1(n10871), .A2(n10870), .B1(n10888), .B2(n12807), .ZN(
        n10872) );
  NOR2_X1 U14117 ( .A1(n10873), .A2(n10872), .ZN(n10874) );
  AOI22_X1 U14118 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19926), .B1(
        n10876), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10881) );
  NAND2_X1 U14119 ( .A1(n20099), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10880) );
  NAND2_X1 U14120 ( .A1(n20225), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10879) );
  NAND2_X1 U14121 ( .A1(n10882), .A2(n11051), .ZN(n10883) );
  NAND2_X1 U14122 ( .A1(n10885), .A2(n10884), .ZN(n11098) );
  AOI22_X1 U14123 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10877), .B1(
        n20061), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U14124 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19892), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U14125 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20156), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10892) );
  OAI22_X1 U14126 ( .A1(n10887), .A2(n10870), .B1(n10868), .B2(n10886), .ZN(
        n10890) );
  INV_X1 U14127 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11282) );
  INV_X1 U14128 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12790) );
  OAI22_X1 U14129 ( .A1(n11282), .A2(n20186), .B1(n10888), .B2(n12790), .ZN(
        n10889) );
  NOR2_X1 U14130 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  NAND4_X1 U14131 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(
        n10900) );
  AOI22_X1 U14132 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19926), .B1(
        n10876), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U14133 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10864), .B1(
        n17033), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U14134 ( .A1(n20225), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10896) );
  NAND2_X1 U14135 ( .A1(n20099), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10895) );
  NAND4_X1 U14136 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10899) );
  INV_X1 U14137 ( .A(n11173), .ZN(n10901) );
  NAND2_X1 U14138 ( .A1(n10901), .A2(n11051), .ZN(n10902) );
  XNOR2_X1 U14139 ( .A(n11098), .B(n11099), .ZN(n11093) );
  NAND2_X1 U14140 ( .A1(n11093), .A2(n10961), .ZN(n10910) );
  INV_X1 U14141 ( .A(n10904), .ZN(n10954) );
  INV_X1 U14142 ( .A(n10905), .ZN(n10908) );
  INV_X1 U14143 ( .A(n10906), .ZN(n10907) );
  NAND2_X1 U14144 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  NAND2_X1 U14145 ( .A1(n10954), .A2(n10909), .ZN(n16195) );
  NAND2_X1 U14146 ( .A1(n10910), .A2(n16195), .ZN(n14861) );
  INV_X1 U14147 ( .A(n10912), .ZN(n10918) );
  INV_X1 U14148 ( .A(n10911), .ZN(n10913) );
  NAND2_X1 U14149 ( .A1(n10918), .A2(n10913), .ZN(n10914) );
  NAND2_X1 U14150 ( .A1(n9790), .A2(n10914), .ZN(n16234) );
  NAND2_X1 U14151 ( .A1(n10915), .A2(n16234), .ZN(n16927) );
  NAND2_X1 U14152 ( .A1(n10916), .A2(n10919), .ZN(n10917) );
  NAND2_X1 U14153 ( .A1(n10918), .A2(n10917), .ZN(n10928) );
  XNOR2_X1 U14154 ( .A(n10928), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19761) );
  INV_X1 U14155 ( .A(n10919), .ZN(n10922) );
  NAND2_X1 U14156 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10920) );
  NOR2_X1 U14157 ( .A1(n10980), .A2(n10920), .ZN(n10921) );
  OR2_X1 U14158 ( .A1(n10922), .A2(n10921), .ZN(n16258) );
  INV_X1 U14159 ( .A(n10923), .ZN(n10925) );
  NAND2_X1 U14160 ( .A1(n11137), .A2(n10980), .ZN(n10924) );
  NAND2_X1 U14161 ( .A1(n10925), .A2(n10924), .ZN(n17392) );
  INV_X1 U14162 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17395) );
  OR2_X1 U14163 ( .A1(n17392), .A2(n17395), .ZN(n17394) );
  OAI21_X1 U14164 ( .B1(n16258), .B2(n16963), .A(n17394), .ZN(n10927) );
  NAND2_X1 U14165 ( .A1(n16258), .A2(n16963), .ZN(n10926) );
  AND2_X1 U14166 ( .A1(n10927), .A2(n10926), .ZN(n19760) );
  NAND2_X1 U14167 ( .A1(n19761), .A2(n19760), .ZN(n19759) );
  INV_X1 U14168 ( .A(n10928), .ZN(n16250) );
  NAND2_X1 U14169 ( .A1(n16250), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10929) );
  AND2_X1 U14170 ( .A1(n19759), .A2(n10929), .ZN(n16930) );
  INV_X1 U14171 ( .A(n10931), .ZN(n10932) );
  NAND2_X1 U14172 ( .A1(n9790), .A2(n10932), .ZN(n10933) );
  NAND2_X1 U14173 ( .A1(n10930), .A2(n10933), .ZN(n16932) );
  AND2_X1 U14174 ( .A1(n16932), .A2(n16937), .ZN(n10935) );
  AOI21_X1 U14175 ( .B1(n16930), .B2(n16928), .A(n10935), .ZN(n10934) );
  INV_X1 U14176 ( .A(n16930), .ZN(n16946) );
  INV_X1 U14177 ( .A(n10935), .ZN(n10936) );
  NAND3_X1 U14178 ( .A1(n16946), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n10936), .ZN(n10939) );
  INV_X1 U14179 ( .A(n16932), .ZN(n10937) );
  NAND2_X1 U14180 ( .A1(n10937), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10938) );
  INV_X1 U14181 ( .A(n10941), .ZN(n10942) );
  XNOR2_X1 U14182 ( .A(n10930), .B(n10942), .ZN(n10943) );
  NAND2_X1 U14183 ( .A1(n10943), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10945) );
  INV_X1 U14184 ( .A(n10943), .ZN(n16211) );
  INV_X1 U14185 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16914) );
  NAND2_X1 U14186 ( .A1(n16211), .A2(n16914), .ZN(n10944) );
  AND2_X1 U14187 ( .A1(n10945), .A2(n10944), .ZN(n16919) );
  NAND2_X1 U14188 ( .A1(n16921), .A2(n16919), .ZN(n10949) );
  XNOR2_X1 U14189 ( .A(n11086), .B(n10946), .ZN(n11091) );
  OAI21_X1 U14190 ( .B1(n11091), .B2(n11177), .A(n16211), .ZN(n10947) );
  NAND2_X1 U14191 ( .A1(n10947), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10948) );
  NAND2_X1 U14192 ( .A1(n10949), .A2(n10948), .ZN(n16667) );
  NAND2_X1 U14193 ( .A1(n10595), .A2(n10951), .ZN(n10952) );
  NAND2_X1 U14194 ( .A1(n10950), .A2(n10952), .ZN(n16166) );
  NOR2_X1 U14195 ( .A1(n16166), .A2(n10961), .ZN(n10963) );
  NAND2_X1 U14196 ( .A1(n10963), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16664) );
  XNOR2_X1 U14197 ( .A(n10954), .B(n10953), .ZN(n10965) );
  NAND2_X1 U14198 ( .A1(n10965), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16678) );
  NAND2_X1 U14199 ( .A1(n19834), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10958) );
  INV_X1 U14200 ( .A(n10957), .ZN(n10967) );
  MUX2_X1 U14201 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n10958), .S(n10967), .Z(
        n10960) );
  NAND2_X1 U14202 ( .A1(n10960), .A2(n10959), .ZN(n16133) );
  OR2_X1 U14203 ( .A1(n16133), .A2(n10961), .ZN(n10962) );
  INV_X1 U14204 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14205 ( .A1(n10962), .A2(n11525), .ZN(n11498) );
  INV_X1 U14206 ( .A(n10963), .ZN(n10964) );
  NAND2_X1 U14207 ( .A1(n10964), .A2(n16886), .ZN(n16663) );
  INV_X1 U14208 ( .A(n10965), .ZN(n16178) );
  INV_X1 U14209 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16885) );
  NAND2_X1 U14210 ( .A1(n16178), .A2(n16885), .ZN(n16679) );
  AND2_X1 U14211 ( .A1(n16663), .A2(n16679), .ZN(n11499) );
  NAND2_X1 U14212 ( .A1(n19834), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10966) );
  MUX2_X1 U14213 ( .A(n9699), .B(n10966), .S(n10950), .Z(n10968) );
  NAND2_X1 U14214 ( .A1(n10968), .A2(n10967), .ZN(n16154) );
  INV_X1 U14215 ( .A(n16154), .ZN(n10969) );
  NAND2_X1 U14216 ( .A1(n10969), .A2(n11177), .ZN(n10970) );
  INV_X1 U14217 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14218 ( .A1(n10970), .A2(n11524), .ZN(n16645) );
  AND3_X1 U14219 ( .A1(n11498), .A2(n11499), .A3(n16645), .ZN(n10974) );
  INV_X1 U14220 ( .A(n10970), .ZN(n10971) );
  NAND2_X1 U14221 ( .A1(n10971), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16648) );
  NAND2_X1 U14222 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10972) );
  NAND2_X1 U14223 ( .A1(n16648), .A2(n11497), .ZN(n10973) );
  INV_X1 U14224 ( .A(n10975), .ZN(n10976) );
  NAND2_X1 U14225 ( .A1(n10976), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16635) );
  NAND2_X1 U14226 ( .A1(n16539), .A2(n10694), .ZN(n10977) );
  INV_X1 U14227 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15932) );
  NOR2_X1 U14228 ( .A1(n10980), .A2(n15932), .ZN(n10982) );
  AOI21_X1 U14229 ( .B1(n10982), .B2(n10981), .A(n10990), .ZN(n15936) );
  NAND2_X1 U14230 ( .A1(n15936), .A2(n11177), .ZN(n11536) );
  INV_X1 U14231 ( .A(n10984), .ZN(n10986) );
  NOR2_X1 U14232 ( .A1(n10985), .A2(n16717), .ZN(n16508) );
  NOR2_X1 U14233 ( .A1(n10986), .A2(n16508), .ZN(n11532) );
  NAND2_X1 U14234 ( .A1(n9699), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10989) );
  XNOR2_X1 U14235 ( .A(n10990), .B(n10989), .ZN(n10988) );
  INV_X1 U14236 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10987) );
  OAI21_X1 U14237 ( .B1(n10988), .B2(n10961), .A(n10987), .ZN(n16477) );
  INV_X1 U14238 ( .A(n10988), .ZN(n15923) );
  NAND3_X1 U14239 ( .A1(n15923), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11177), .ZN(n16478) );
  NAND2_X1 U14240 ( .A1(n14888), .A2(n16478), .ZN(n10995) );
  NAND2_X1 U14241 ( .A1(n19834), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10991) );
  XNOR2_X1 U14242 ( .A(n14889), .B(n10991), .ZN(n15915) );
  AOI21_X1 U14243 ( .B1(n15915), .B2(n11177), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14887) );
  AND2_X1 U14244 ( .A1(n11177), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10992) );
  NAND2_X1 U14245 ( .A1(n15915), .A2(n10992), .ZN(n14886) );
  INV_X1 U14246 ( .A(n14886), .ZN(n10993) );
  NAND2_X1 U14247 ( .A1(n11024), .A2(n11002), .ZN(n10997) );
  MUX2_X1 U14248 ( .A(n10997), .B(n14983), .S(n10996), .Z(n11007) );
  INV_X1 U14249 ( .A(n10998), .ZN(n11000) );
  NAND2_X1 U14250 ( .A1(n16991), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10999) );
  NAND2_X1 U14251 ( .A1(n11042), .A2(n11001), .ZN(n11029) );
  NAND2_X1 U14252 ( .A1(n14979), .A2(n11029), .ZN(n11004) );
  XNOR2_X1 U14253 ( .A(n11001), .B(n11000), .ZN(n11037) );
  OAI211_X1 U14254 ( .C1(n11002), .C2(n11042), .A(n20510), .B(n11037), .ZN(
        n11003) );
  OAI211_X1 U14255 ( .C1(n11005), .C2(n11044), .A(n11004), .B(n11003), .ZN(
        n11006) );
  NAND2_X1 U14256 ( .A1(n11007), .A2(n11006), .ZN(n11014) );
  NAND2_X1 U14257 ( .A1(n11009), .A2(n11008), .ZN(n11011) );
  NAND2_X1 U14258 ( .A1(n21570), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14259 ( .A1(n11011), .A2(n11010), .ZN(n11017) );
  INV_X1 U14260 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U14261 ( .A1(n11031), .A2(n11013), .ZN(n11036) );
  MUX2_X1 U14262 ( .A(n11014), .B(n14983), .S(n11036), .Z(n11015) );
  INV_X1 U14263 ( .A(n11015), .ZN(n11020) );
  NOR2_X1 U14264 ( .A1(n13772), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11016) );
  NAND2_X1 U14265 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13772), .ZN(
        n11018) );
  NOR2_X1 U14266 ( .A1(n11020), .A2(n11023), .ZN(n11021) );
  MUX2_X1 U14267 ( .A(n11021), .B(n13772), .S(n17044), .Z(n11026) );
  OAI21_X1 U14268 ( .B1(n11026), .B2(n14498), .A(n10741), .ZN(n11028) );
  INV_X1 U14269 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20395) );
  NOR2_X4 U14270 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20394), .ZN(n20462) );
  INV_X1 U14271 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21644) );
  NAND2_X1 U14272 ( .A1(n21644), .A2(n20394), .ZN(n20407) );
  NAND2_X1 U14273 ( .A1(n11022), .A2(n14445), .ZN(n11027) );
  NOR2_X1 U14274 ( .A1(n14605), .A2(n11051), .ZN(n13775) );
  MUX2_X1 U14275 ( .A(n11028), .B(n11027), .S(n13775), .Z(n11069) );
  NAND2_X1 U14276 ( .A1(n11030), .A2(n11029), .ZN(n11033) );
  NAND3_X1 U14277 ( .A1(n11033), .A2(n11032), .A3(n11031), .ZN(n11034) );
  NAND2_X1 U14278 ( .A1(n11034), .A2(n11040), .ZN(n20503) );
  AND2_X1 U14279 ( .A1(n11051), .A2(n14498), .ZN(n11056) );
  NAND2_X1 U14280 ( .A1(n14499), .A2(n11056), .ZN(n11115) );
  INV_X1 U14281 ( .A(n11036), .ZN(n11046) );
  INV_X1 U14282 ( .A(n11037), .ZN(n11038) );
  NOR2_X1 U14283 ( .A1(n11044), .A2(n11038), .ZN(n11039) );
  NAND2_X1 U14284 ( .A1(n11046), .A2(n11039), .ZN(n11041) );
  INV_X1 U14285 ( .A(n11042), .ZN(n11043) );
  NOR2_X1 U14286 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  AOI21_X1 U14287 ( .B1(n11046), .B2(n11045), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n11050) );
  AOI21_X1 U14288 ( .B1(n14475), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13770) );
  NAND2_X1 U14289 ( .A1(n11048), .A2(n13770), .ZN(n11049) );
  INV_X1 U14290 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13766) );
  AOI21_X1 U14291 ( .B1(n11049), .B2(n13766), .A(n16993), .ZN(n16975) );
  NAND2_X1 U14292 ( .A1(n14499), .A2(n11002), .ZN(n11052) );
  OAI21_X1 U14293 ( .B1(n11054), .B2(n11022), .A(n13718), .ZN(n11063) );
  NAND2_X1 U14294 ( .A1(n11055), .A2(n14524), .ZN(n11057) );
  NAND2_X1 U14295 ( .A1(n11057), .A2(n11056), .ZN(n11450) );
  AOI21_X1 U14296 ( .B1(n11051), .B2(n10741), .A(n14498), .ZN(n11058) );
  OAI21_X1 U14297 ( .B1(n11058), .B2(n19846), .A(n10734), .ZN(n11059) );
  AND4_X1 U14298 ( .A1(n11450), .A2(n11060), .A3(n10752), .A4(n11059), .ZN(
        n11062) );
  NAND3_X1 U14299 ( .A1(n10747), .A2(n13758), .A3(n14445), .ZN(n11061) );
  MUX2_X1 U14300 ( .A(n10747), .B(n11022), .S(n11051), .Z(n11065) );
  INV_X1 U14301 ( .A(n13758), .ZN(n14492) );
  NOR2_X1 U14302 ( .A1(n14492), .A2(n20509), .ZN(n11064) );
  NAND2_X1 U14303 ( .A1(n11065), .A2(n11064), .ZN(n11066) );
  NAND2_X1 U14304 ( .A1(n13760), .A2(n11066), .ZN(n11067) );
  NOR2_X1 U14305 ( .A1(n11495), .A2(n11067), .ZN(n11068) );
  NAND2_X1 U14306 ( .A1(n11069), .A2(n11068), .ZN(n11070) );
  AND2_X1 U14307 ( .A1(n14499), .A2(n14979), .ZN(n20500) );
  INV_X1 U14308 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11464) );
  INV_X1 U14309 ( .A(n17396), .ZN(n11072) );
  NAND2_X1 U14310 ( .A1(n11072), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17398) );
  INV_X1 U14311 ( .A(n11142), .ZN(n11073) );
  XNOR2_X1 U14312 ( .A(n11137), .B(n11073), .ZN(n11074) );
  NOR2_X1 U14313 ( .A1(n17398), .A2(n11074), .ZN(n11076) );
  AOI21_X1 U14314 ( .B1(n17398), .B2(n11074), .A(n11076), .ZN(n11075) );
  INV_X1 U14315 ( .A(n11075), .ZN(n13733) );
  NOR2_X1 U14316 ( .A1(n16963), .A2(n13733), .ZN(n13732) );
  NOR2_X1 U14317 ( .A1(n11076), .A2(n13732), .ZN(n11079) );
  XNOR2_X1 U14318 ( .A(n11464), .B(n11079), .ZN(n19766) );
  INV_X1 U14319 ( .A(n19766), .ZN(n11078) );
  XNOR2_X1 U14320 ( .A(n11152), .B(n11077), .ZN(n19764) );
  NAND2_X1 U14321 ( .A1(n11078), .A2(n19764), .ZN(n19768) );
  OR2_X1 U14322 ( .A1(n11079), .A2(n11464), .ZN(n11080) );
  NAND2_X1 U14323 ( .A1(n19768), .A2(n11080), .ZN(n11081) );
  XNOR2_X1 U14324 ( .A(n11081), .B(n16928), .ZN(n16948) );
  NAND2_X1 U14325 ( .A1(n11081), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11082) );
  INV_X1 U14326 ( .A(n11159), .ZN(n11083) );
  NAND2_X1 U14327 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  INV_X1 U14328 ( .A(n11087), .ZN(n11089) );
  NAND2_X1 U14329 ( .A1(n11089), .A2(n11088), .ZN(n11090) );
  INV_X1 U14330 ( .A(n11091), .ZN(n11092) );
  INV_X1 U14331 ( .A(n11094), .ZN(n11095) );
  INV_X1 U14332 ( .A(n11099), .ZN(n11096) );
  NAND2_X1 U14333 ( .A1(n9765), .A2(n11096), .ZN(n14858) );
  INV_X1 U14334 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11097) );
  INV_X1 U14335 ( .A(n11098), .ZN(n11100) );
  NAND2_X1 U14336 ( .A1(n11100), .A2(n11099), .ZN(n11101) );
  NAND2_X1 U14337 ( .A1(n16657), .A2(n16885), .ZN(n11102) );
  INV_X1 U14338 ( .A(n11101), .ZN(n11105) );
  NAND2_X1 U14339 ( .A1(n11105), .A2(n11177), .ZN(n16660) );
  NAND2_X1 U14340 ( .A1(n16660), .A2(n16886), .ZN(n11104) );
  AND2_X1 U14341 ( .A1(n11102), .A2(n11104), .ZN(n11103) );
  INV_X1 U14342 ( .A(n16657), .ZN(n16658) );
  NAND3_X1 U14343 ( .A1(n11104), .A2(n16658), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11107) );
  NAND3_X1 U14344 ( .A1(n11105), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11177), .ZN(n11106) );
  NAND2_X1 U14345 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16730) );
  NOR2_X1 U14346 ( .A1(n16730), .A2(n13029), .ZN(n11487) );
  AND2_X1 U14347 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16818) );
  AND2_X1 U14348 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11109) );
  NAND3_X1 U14349 ( .A1(n16818), .A2(n16813), .A3(n11109), .ZN(n14845) );
  NAND3_X1 U14350 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11110) );
  NOR2_X1 U14351 ( .A1(n14845), .A2(n11110), .ZN(n16773) );
  NAND2_X1 U14352 ( .A1(n12662), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16760) );
  NAND2_X1 U14353 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11111) );
  NOR2_X1 U14354 ( .A1(n16760), .A2(n11111), .ZN(n11563) );
  AND2_X1 U14355 ( .A1(n11487), .A2(n11563), .ZN(n13014) );
  NAND2_X1 U14356 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16705) );
  INV_X1 U14357 ( .A(n16705), .ZN(n11112) );
  AND2_X1 U14358 ( .A1(n13014), .A2(n11112), .ZN(n11113) );
  AND2_X2 U14359 ( .A1(n14760), .A2(n11113), .ZN(n13568) );
  AND2_X1 U14360 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11478) );
  INV_X1 U14361 ( .A(n11478), .ZN(n14968) );
  INV_X1 U14362 ( .A(n11115), .ZN(n20502) );
  MUX2_X1 U14363 ( .A(n11116), .B(n11133), .S(n11451), .Z(n11119) );
  NAND2_X1 U14364 ( .A1(n13726), .A2(n11117), .ZN(n11118) );
  INV_X1 U14365 ( .A(n11120), .ZN(n11121) );
  NAND2_X1 U14366 ( .A1(n14467), .A2(n11121), .ZN(n14491) );
  NAND2_X1 U14367 ( .A1(n14514), .A2(n13718), .ZN(n14493) );
  NAND2_X1 U14368 ( .A1(n14493), .A2(n11002), .ZN(n11122) );
  NAND2_X1 U14369 ( .A1(n14491), .A2(n11122), .ZN(n11123) );
  NOR2_X1 U14370 ( .A1(n9996), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11125) );
  NOR2_X1 U14371 ( .A1(n14524), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11340) );
  AOI222_X1 U14372 ( .A1(n14962), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n14961), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n11138), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11365) );
  AOI21_X1 U14373 ( .B1(n11127), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U14374 ( .A1(n19846), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11128) );
  OAI211_X1 U14375 ( .C1(n11140), .C2(n10758), .A(n11129), .B(n11128), .ZN(
        n14534) );
  NAND2_X1 U14376 ( .A1(n11131), .A2(n11130), .ZN(n11465) );
  INV_X1 U14377 ( .A(n11133), .ZN(n11134) );
  NAND2_X1 U14378 ( .A1(n11134), .A2(n11138), .ZN(n11150) );
  NAND2_X1 U14379 ( .A1(n14524), .A2(n12673), .ZN(n11135) );
  NAND2_X1 U14380 ( .A1(n19889), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16974) );
  NAND2_X1 U14381 ( .A1(n11135), .A2(n16974), .ZN(n11136) );
  NAND2_X1 U14382 ( .A1(n14534), .A2(n14535), .ZN(n11145) );
  AOI22_X1 U14383 ( .A1(n11340), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11139) );
  OAI21_X1 U14384 ( .B1(n11140), .B2(n20412), .A(n11139), .ZN(n11146) );
  XNOR2_X1 U14385 ( .A(n11145), .B(n11146), .ZN(n14564) );
  NAND2_X1 U14386 ( .A1(n11133), .A2(n14524), .ZN(n11141) );
  MUX2_X1 U14387 ( .A(n11141), .B(n20252), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11144) );
  NAND2_X1 U14388 ( .A1(n11335), .A2(n11142), .ZN(n11143) );
  AND2_X1 U14389 ( .A1(n11144), .A2(n11143), .ZN(n14563) );
  NAND2_X1 U14390 ( .A1(n14564), .A2(n14563), .ZN(n14562) );
  INV_X1 U14391 ( .A(n11146), .ZN(n11147) );
  NAND2_X1 U14392 ( .A1(n11145), .A2(n11147), .ZN(n11148) );
  NAND2_X1 U14393 ( .A1(n14562), .A2(n11148), .ZN(n11157) );
  NAND2_X1 U14394 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11151) );
  OAI211_X1 U14395 ( .C1(n11149), .C2(n11152), .A(n11151), .B(n11150), .ZN(
        n11155) );
  XNOR2_X1 U14396 ( .A(n11157), .B(n11155), .ZN(n14559) );
  NAND2_X1 U14397 ( .A1(n14962), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11154) );
  AOI22_X1 U14398 ( .A1(n14961), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11153) );
  AND2_X1 U14399 ( .A1(n11154), .A2(n11153), .ZN(n14558) );
  NAND2_X1 U14400 ( .A1(n14559), .A2(n14558), .ZN(n14561) );
  INV_X1 U14401 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U14402 ( .A1(n11157), .A2(n11156), .ZN(n11158) );
  NAND2_X1 U14403 ( .A1(n11335), .A2(n11159), .ZN(n11162) );
  AOI22_X1 U14404 ( .A1(n14961), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14405 ( .A1(n14962), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11160) );
  AND3_X1 U14406 ( .A1(n11162), .A2(n11161), .A3(n11160), .ZN(n16214) );
  NAND2_X1 U14407 ( .A1(n11335), .A2(n11163), .ZN(n11168) );
  AOI22_X1 U14408 ( .A1(n11138), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11165) );
  NAND2_X1 U14409 ( .A1(n14961), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11164) );
  AND2_X1 U14410 ( .A1(n11165), .A2(n11164), .ZN(n11167) );
  NAND2_X1 U14411 ( .A1(n14962), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11166) );
  NAND2_X1 U14412 ( .A1(n11335), .A2(n11169), .ZN(n11172) );
  AOI22_X1 U14413 ( .A1(n14961), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U14414 ( .A1(n14962), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11170) );
  AOI21_X1 U14415 ( .B1(n11174), .B2(n10418), .A(n10419), .ZN(n11175) );
  INV_X1 U14416 ( .A(n11175), .ZN(n14593) );
  INV_X1 U14417 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20420) );
  AOI22_X1 U14418 ( .A1(n14961), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11176) );
  OAI21_X1 U14419 ( .B1(n11140), .B2(n20420), .A(n11176), .ZN(n14594) );
  AOI21_X1 U14420 ( .B1(n14593), .B2(n14594), .A(n10394), .ZN(n11178) );
  AOI22_X1 U14421 ( .A1(n14961), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11179) );
  OAI21_X1 U14422 ( .B1(n11140), .B2(n21760), .A(n11179), .ZN(n14601) );
  NAND2_X1 U14423 ( .A1(n14602), .A2(n14601), .ZN(n14517) );
  AOI22_X1 U14424 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11187) );
  NAND2_X1 U14425 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11181) );
  NAND2_X1 U14426 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11180) );
  OAI211_X1 U14427 ( .C1(n10559), .C2(n11182), .A(n11181), .B(n11180), .ZN(
        n11183) );
  INV_X1 U14428 ( .A(n11183), .ZN(n11186) );
  AOI22_X1 U14429 ( .A1(n11284), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14430 ( .A1(n12724), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11184) );
  NAND4_X1 U14431 ( .A1(n11187), .A2(n11186), .A3(n11185), .A4(n11184), .ZN(
        n11194) );
  AOI22_X1 U14432 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14433 ( .A1(n11209), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14434 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11190) );
  NAND2_X1 U14435 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11189) );
  NAND4_X1 U14436 ( .A1(n11192), .A2(n11191), .A3(n11190), .A4(n11189), .ZN(
        n11193) );
  NAND2_X1 U14437 ( .A1(n11335), .A2(n14541), .ZN(n11197) );
  AOI22_X1 U14438 ( .A1(n14961), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U14439 ( .A1(n14962), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11195) );
  INV_X1 U14440 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11198) );
  OAI22_X1 U14441 ( .A1(n11199), .A2(n12832), .B1(n12808), .B2(n11198), .ZN(
        n11200) );
  INV_X1 U14442 ( .A(n11200), .ZN(n11208) );
  AOI22_X1 U14443 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14444 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12724), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14445 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11202) );
  NAND2_X1 U14446 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11201) );
  OAI211_X1 U14447 ( .C1(n10559), .C2(n11203), .A(n11202), .B(n11201), .ZN(
        n11204) );
  INV_X1 U14448 ( .A(n11204), .ZN(n11205) );
  NAND4_X1 U14449 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n11215) );
  AOI22_X1 U14450 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14451 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14452 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U14453 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11210) );
  NAND4_X1 U14454 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n11214) );
  INV_X1 U14455 ( .A(n14542), .ZN(n11218) );
  AOI22_X1 U14456 ( .A1(n14961), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11138), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U14457 ( .A1(n14962), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11216) );
  OAI211_X1 U14458 ( .C1(n11149), .C2(n11218), .A(n11217), .B(n11216), .ZN(
        n14599) );
  NAND2_X1 U14459 ( .A1(n14516), .A2(n14599), .ZN(n11517) );
  INV_X1 U14460 ( .A(n11517), .ZN(n11240) );
  INV_X1 U14461 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11220) );
  INV_X1 U14462 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11219) );
  OAI22_X1 U14463 ( .A1(n11220), .A2(n12832), .B1(n10559), .B2(n11219), .ZN(
        n11221) );
  INV_X1 U14464 ( .A(n11221), .ZN(n11229) );
  AOI22_X1 U14465 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10840), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11227) );
  INV_X1 U14467 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14468 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14469 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11222) );
  OAI211_X1 U14470 ( .C1(n12808), .C2(n11224), .A(n11223), .B(n11222), .ZN(
        n11225) );
  INV_X1 U14471 ( .A(n11225), .ZN(n11226) );
  NAND4_X1 U14472 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11235) );
  AOI22_X1 U14473 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10519), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14474 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12841), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U14476 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11230) );
  NAND4_X1 U14477 ( .A1(n11233), .A2(n11232), .A3(n11231), .A4(n11230), .ZN(
        n11234) );
  NAND2_X1 U14478 ( .A1(n11335), .A2(n14303), .ZN(n11238) );
  AOI22_X1 U14479 ( .A1(n14961), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U14480 ( .A1(n14962), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11236) );
  NAND2_X1 U14481 ( .A1(n11240), .A2(n11239), .ZN(n11518) );
  INV_X1 U14482 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11242) );
  INV_X1 U14483 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11241) );
  OAI22_X1 U14484 ( .A1(n11242), .A2(n12832), .B1(n12808), .B2(n11241), .ZN(
        n11243) );
  INV_X1 U14485 ( .A(n11243), .ZN(n11251) );
  AOI22_X1 U14486 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14487 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12724), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U14488 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11245) );
  NAND2_X1 U14489 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11244) );
  OAI211_X1 U14490 ( .C1(n10559), .C2(n11246), .A(n11245), .B(n11244), .ZN(
        n11247) );
  INV_X1 U14491 ( .A(n11247), .ZN(n11248) );
  NAND4_X1 U14492 ( .A1(n11251), .A2(n11250), .A3(n11249), .A4(n11248), .ZN(
        n11257) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14494 ( .A1(n11209), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14495 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U14496 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11252) );
  NAND4_X1 U14497 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n11256) );
  OR2_X1 U14498 ( .A1(n11257), .A2(n11256), .ZN(n14307) );
  NAND2_X1 U14499 ( .A1(n11335), .A2(n14307), .ZN(n11260) );
  AOI22_X1 U14500 ( .A1(n14961), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11259) );
  NAND2_X1 U14501 ( .A1(n14962), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11258) );
  INV_X1 U14502 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11263) );
  INV_X1 U14503 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21502) );
  OAI22_X1 U14504 ( .A1(n11263), .A2(n10559), .B1(n12808), .B2(n21502), .ZN(
        n11264) );
  INV_X1 U14505 ( .A(n11264), .ZN(n11270) );
  AOI22_X1 U14506 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10496), .B1(
        n12842), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11266) );
  NAND2_X1 U14507 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11265) );
  AND2_X1 U14508 ( .A1(n11266), .A2(n11265), .ZN(n11269) );
  AOI22_X1 U14509 ( .A1(n11284), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14510 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12834), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11267) );
  NAND4_X1 U14511 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11276) );
  AOI22_X1 U14512 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14513 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U14515 ( .A1(n11209), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11271) );
  NAND4_X1 U14516 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11275) );
  NAND2_X1 U14517 ( .A1(n11335), .A2(n14554), .ZN(n11279) );
  AOI22_X1 U14518 ( .A1(n14961), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11278) );
  NAND2_X1 U14519 ( .A1(n14962), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11277) );
  AOI22_X1 U14520 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12827), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U14521 ( .A1(n12828), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11281) );
  NAND2_X1 U14522 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11280) );
  OAI211_X1 U14523 ( .C1(n10559), .C2(n11282), .A(n11281), .B(n11280), .ZN(
        n11283) );
  INV_X1 U14524 ( .A(n11283), .ZN(n11287) );
  AOI22_X1 U14525 ( .A1(n11284), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14526 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10495), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11285) );
  NAND4_X1 U14527 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n11294) );
  AOI22_X1 U14528 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10551), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14529 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12841), .B1(
        n12842), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U14531 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11289) );
  NAND4_X1 U14532 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11293) );
  NOR2_X1 U14533 ( .A1(n11294), .A2(n11293), .ZN(n12703) );
  AOI22_X1 U14534 ( .A1(n14961), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U14535 ( .A1(n14962), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11295) );
  OAI211_X1 U14536 ( .C1(n11149), .C2(n12703), .A(n11296), .B(n11295), .ZN(
        n14528) );
  INV_X1 U14537 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11298) );
  INV_X1 U14538 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11297) );
  OAI22_X1 U14539 ( .A1(n11298), .A2(n12832), .B1(n12808), .B2(n11297), .ZN(
        n11299) );
  INV_X1 U14540 ( .A(n11299), .ZN(n11306) );
  AOI22_X1 U14541 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11305) );
  BUF_X1 U14542 ( .A(n10840), .Z(n12724) );
  AOI22_X1 U14543 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12724), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11304) );
  NAND2_X1 U14544 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11301) );
  NAND2_X1 U14545 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11300) );
  OAI211_X1 U14546 ( .C1(n10559), .C2(n21703), .A(n11301), .B(n11300), .ZN(
        n11302) );
  INV_X1 U14547 ( .A(n11302), .ZN(n11303) );
  NAND4_X1 U14548 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(
        n11312) );
  AOI22_X1 U14549 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14550 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14551 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U14552 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11307) );
  NAND4_X1 U14553 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11311) );
  OR2_X1 U14554 ( .A1(n11312), .A2(n11311), .ZN(n14646) );
  INV_X1 U14555 ( .A(n14646), .ZN(n14638) );
  AOI22_X1 U14556 ( .A1(n14961), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14557 ( .A1(n14962), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11313) );
  OAI211_X1 U14558 ( .C1(n11149), .C2(n14638), .A(n11314), .B(n11313), .ZN(
        n14582) );
  AND2_X1 U14559 ( .A1(n14528), .A2(n14582), .ZN(n11315) );
  INV_X1 U14560 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U14561 ( .A1(n14961), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11316) );
  OAI21_X1 U14562 ( .B1(n11140), .B2(n20439), .A(n11316), .ZN(n14842) );
  AOI22_X1 U14563 ( .A1(n14961), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11317) );
  OAI21_X1 U14564 ( .B1(n11140), .B2(n20437), .A(n11317), .ZN(n16062) );
  INV_X1 U14565 ( .A(n16062), .ZN(n11339) );
  INV_X1 U14566 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11319) );
  INV_X1 U14567 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11318) );
  OAI22_X1 U14568 ( .A1(n11319), .A2(n12832), .B1(n12808), .B2(n11318), .ZN(
        n11320) );
  INV_X1 U14569 ( .A(n11320), .ZN(n11328) );
  AOI22_X1 U14570 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14571 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11326) );
  NAND2_X1 U14572 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U14573 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11321) );
  OAI211_X1 U14574 ( .C1(n10559), .C2(n11323), .A(n11322), .B(n11321), .ZN(
        n11324) );
  INV_X1 U14575 ( .A(n11324), .ZN(n11325) );
  NAND4_X1 U14576 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11334) );
  AOI22_X1 U14577 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14578 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14579 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U14580 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11329) );
  NAND4_X1 U14581 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11333) );
  NAND2_X1 U14582 ( .A1(n11335), .A2(n14622), .ZN(n11338) );
  AOI22_X1 U14583 ( .A1(n14961), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U14584 ( .A1(n14962), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11336) );
  NOR2_X1 U14585 ( .A1(n11339), .A2(n14597), .ZN(n14841) );
  NAND2_X1 U14586 ( .A1(n14962), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14587 ( .A1(n14961), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14588 ( .A1(n14962), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14589 ( .A1(n14961), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11344) );
  INV_X1 U14590 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U14591 ( .A1(n14961), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11346) );
  OAI21_X1 U14592 ( .B1(n11140), .B2(n19665), .A(n11346), .ZN(n16430) );
  NAND2_X1 U14593 ( .A1(n14962), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14594 ( .A1(n14961), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U14595 ( .A1(n14962), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14596 ( .A1(n14961), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11349) );
  INV_X1 U14597 ( .A(n16004), .ZN(n11351) );
  NAND2_X1 U14598 ( .A1(n11352), .A2(n11351), .ZN(n15999) );
  NAND2_X1 U14599 ( .A1(n14962), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14600 ( .A1(n14961), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11353) );
  INV_X1 U14601 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15985) );
  AOI22_X1 U14602 ( .A1(n14961), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11355) );
  OAI21_X1 U14603 ( .B1(n11140), .B2(n15985), .A(n11355), .ZN(n13033) );
  NAND2_X1 U14604 ( .A1(n14962), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14605 ( .A1(n14961), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11356) );
  AND2_X1 U14606 ( .A1(n11357), .A2(n11356), .ZN(n15966) );
  NAND2_X1 U14607 ( .A1(n14962), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14608 ( .A1(n14961), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11359) );
  INV_X1 U14609 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20455) );
  AOI22_X1 U14610 ( .A1(n14961), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11361) );
  OAI21_X1 U14611 ( .B1(n11140), .B2(n20455), .A(n11361), .ZN(n15938) );
  INV_X1 U14612 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20456) );
  AOI22_X1 U14613 ( .A1(n14961), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11362) );
  OAI21_X1 U14614 ( .B1(n11140), .B2(n20456), .A(n11362), .ZN(n11541) );
  NAND2_X1 U14615 ( .A1(n14962), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14616 ( .A1(n14961), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11138), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U14617 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11370) );
  INV_X1 U14618 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11367) );
  OAI22_X1 U14619 ( .A1(n10345), .A2(n14164), .B1(n16993), .B2(n11367), .ZN(
        n11368) );
  AOI21_X1 U14620 ( .B1(n11420), .B2(P2_REIP_REG_4__SCAN_IN), .A(n11368), .ZN(
        n11369) );
  NAND2_X1 U14621 ( .A1(n11370), .A2(n11369), .ZN(n14162) );
  NAND2_X1 U14622 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11374) );
  INV_X1 U14623 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11371) );
  OAI22_X1 U14624 ( .A1(n10345), .A2(n11371), .B1(n16993), .B2(n16201), .ZN(
        n11372) );
  AOI21_X1 U14625 ( .B1(n11420), .B2(P2_REIP_REG_5__SCAN_IN), .A(n11372), .ZN(
        n11373) );
  NAND2_X1 U14626 ( .A1(n11374), .A2(n11373), .ZN(n14207) );
  NAND2_X1 U14627 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11377) );
  INV_X1 U14628 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16158) );
  OAI22_X1 U14629 ( .A1(n10345), .A2(n16157), .B1(n16993), .B2(n16158), .ZN(
        n11375) );
  AOI21_X1 U14630 ( .B1(n11420), .B2(P2_REIP_REG_8__SCAN_IN), .A(n11375), .ZN(
        n11376) );
  NAND2_X1 U14631 ( .A1(n11377), .A2(n11376), .ZN(n14652) );
  AOI22_X1 U14632 ( .A1(n11438), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11378) );
  AOI21_X1 U14633 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11379), .ZN(n14317) );
  AOI22_X1 U14634 ( .A1(n11438), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11380) );
  OAI21_X1 U14635 ( .B1(n11440), .B2(n20420), .A(n11380), .ZN(n11381) );
  AOI21_X1 U14636 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11381), .ZN(n14435) );
  NOR2_X1 U14637 ( .A1(n14317), .A2(n14435), .ZN(n14315) );
  AND2_X1 U14638 ( .A1(n14652), .A2(n14315), .ZN(n11382) );
  INV_X1 U14639 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20424) );
  AOI22_X1 U14640 ( .A1(n11438), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11383) );
  OAI21_X1 U14641 ( .B1(n11440), .B2(n20424), .A(n11383), .ZN(n11384) );
  AOI21_X1 U14642 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11384), .ZN(n14545) );
  INV_X1 U14643 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20426) );
  AOI22_X1 U14644 ( .A1(n11438), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11385) );
  AOI21_X1 U14645 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11386), .ZN(n11505) );
  INV_X1 U14646 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20428) );
  AOI22_X1 U14647 ( .A1(n11438), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11387) );
  OAI21_X1 U14648 ( .B1(n11440), .B2(n20428), .A(n11387), .ZN(n11388) );
  AOI21_X1 U14649 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11388), .ZN(n14308) );
  NAND2_X1 U14650 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11390) );
  INV_X1 U14651 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20430) );
  AOI22_X1 U14652 ( .A1(n11438), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11389) );
  NAND2_X1 U14653 ( .A1(n11390), .A2(n9758), .ZN(n14549) );
  NAND2_X1 U14654 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11394) );
  INV_X1 U14655 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n21718) );
  AOI22_X1 U14656 ( .A1(n14895), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11391) );
  OAI21_X1 U14657 ( .B1(n11440), .B2(n21718), .A(n11391), .ZN(n11392) );
  INV_X1 U14658 ( .A(n11392), .ZN(n11393) );
  NAND2_X1 U14659 ( .A1(n11394), .A2(n11393), .ZN(n14648) );
  INV_X1 U14660 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20435) );
  AOI22_X1 U14661 ( .A1(n14895), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11395) );
  OAI21_X1 U14662 ( .B1(n11440), .B2(n20435), .A(n11395), .ZN(n11396) );
  AOI21_X1 U14663 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11396), .ZN(n14618) );
  INV_X1 U14664 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20433) );
  AOI22_X1 U14665 ( .A1(n14895), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11397) );
  AOI21_X1 U14666 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11398), .ZN(n14635) );
  OR2_X1 U14667 ( .A1(n14618), .A2(n14635), .ZN(n11399) );
  NAND2_X1 U14668 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11401) );
  AOI22_X1 U14669 ( .A1(n14895), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11400) );
  NAND2_X1 U14670 ( .A1(n11401), .A2(n9799), .ZN(n14664) );
  NAND2_X1 U14671 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11405) );
  AOI22_X1 U14672 ( .A1(n14895), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11402) );
  OAI21_X1 U14673 ( .B1(n11440), .B2(n20439), .A(n11402), .ZN(n11403) );
  INV_X1 U14674 ( .A(n11403), .ZN(n11404) );
  NAND2_X1 U14675 ( .A1(n11405), .A2(n11404), .ZN(n14762) );
  NAND2_X1 U14676 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11407) );
  AOI22_X1 U14677 ( .A1(n14895), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11406) );
  NAND2_X1 U14678 ( .A1(n11407), .A2(n9756), .ZN(n16334) );
  INV_X1 U14679 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U14680 ( .A1(n14895), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11408) );
  OAI21_X1 U14681 ( .B1(n11440), .B2(n20442), .A(n11408), .ZN(n11409) );
  AOI21_X1 U14682 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11409), .ZN(n12667) );
  INV_X1 U14683 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U14684 ( .A1(n14895), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11410) );
  AOI21_X1 U14685 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11411), .ZN(n13320) );
  NOR2_X1 U14686 ( .A1(n12667), .A2(n13320), .ZN(n12665) );
  AND2_X1 U14687 ( .A1(n16334), .A2(n12665), .ZN(n11412) );
  INV_X1 U14688 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20444) );
  AOI22_X1 U14689 ( .A1(n14895), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11413) );
  OAI21_X1 U14690 ( .B1(n11440), .B2(n20444), .A(n11413), .ZN(n11414) );
  AOI21_X1 U14691 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11414), .ZN(n11569) );
  INV_X1 U14692 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20446) );
  AOI22_X1 U14693 ( .A1(n11438), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11415) );
  AOI21_X1 U14694 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11416), .ZN(n16006) );
  INV_X1 U14695 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20448) );
  AOI22_X1 U14696 ( .A1(n11438), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11417) );
  OAI21_X1 U14697 ( .B1(n11440), .B2(n20448), .A(n11417), .ZN(n11418) );
  AOI21_X1 U14698 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11418), .ZN(n15991) );
  NAND2_X1 U14699 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11422) );
  OAI22_X1 U14700 ( .A1(n10345), .A2(n15979), .B1(n16993), .B2(n10278), .ZN(
        n11419) );
  AOI21_X1 U14701 ( .B1(n11420), .B2(P2_REIP_REG_24__SCAN_IN), .A(n11419), 
        .ZN(n11421) );
  NAND2_X1 U14702 ( .A1(n11422), .A2(n11421), .ZN(n13027) );
  NAND2_X1 U14703 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11426) );
  INV_X1 U14704 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20451) );
  AOI22_X1 U14705 ( .A1(n11438), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11423) );
  OAI21_X1 U14706 ( .B1(n11440), .B2(n20451), .A(n11423), .ZN(n11424) );
  INV_X1 U14707 ( .A(n11424), .ZN(n11425) );
  NAND2_X1 U14708 ( .A1(n11426), .A2(n11425), .ZN(n15964) );
  INV_X1 U14709 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20452) );
  AOI22_X1 U14710 ( .A1(n11438), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11427) );
  OAI21_X1 U14711 ( .B1(n11440), .B2(n20452), .A(n11427), .ZN(n11428) );
  AOI21_X1 U14712 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11428), .ZN(n13561) );
  AOI22_X1 U14713 ( .A1(n11438), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11429) );
  AOI21_X1 U14714 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11430), .ZN(n15940) );
  INV_X1 U14715 ( .A(n15940), .ZN(n11431) );
  NAND2_X1 U14716 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11435) );
  AOI22_X1 U14717 ( .A1(n11438), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11432) );
  OAI21_X1 U14718 ( .B1(n11440), .B2(n20456), .A(n11432), .ZN(n11433) );
  INV_X1 U14719 ( .A(n11433), .ZN(n11434) );
  NAND2_X1 U14720 ( .A1(n11435), .A2(n11434), .ZN(n11546) );
  NAND2_X1 U14721 ( .A1(n14898), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11437) );
  INV_X1 U14722 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20459) );
  AOI22_X1 U14723 ( .A1(n11438), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11436) );
  NAND2_X1 U14724 ( .A1(n11437), .A2(n9800), .ZN(n15918) );
  INV_X1 U14725 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14726 ( .A1(n11438), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11439) );
  OAI21_X1 U14727 ( .B1(n11440), .B2(n11480), .A(n11439), .ZN(n11441) );
  AOI21_X1 U14728 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11441), .ZN(n11445) );
  INV_X1 U14729 ( .A(n11445), .ZN(n11442) );
  NAND2_X1 U14730 ( .A1(n11444), .A2(n11445), .ZN(n11446) );
  NAND2_X1 U14731 ( .A1(n14900), .A2(n11446), .ZN(n15917) );
  NAND2_X1 U14732 ( .A1(n14476), .A2(n11051), .ZN(n11447) );
  NAND2_X1 U14733 ( .A1(n11447), .A2(n14447), .ZN(n11448) );
  NAND2_X2 U14734 ( .A1(n11467), .A2(n11448), .ZN(n19803) );
  NAND2_X1 U14735 ( .A1(n11449), .A2(n11002), .ZN(n14459) );
  NAND2_X1 U14736 ( .A1(n14459), .A2(n11450), .ZN(n11452) );
  NAND2_X1 U14737 ( .A1(n11452), .A2(n11451), .ZN(n11461) );
  OAI211_X1 U14738 ( .C1(n13768), .C2(n13009), .A(n11455), .B(n11454), .ZN(
        n11459) );
  INV_X1 U14739 ( .A(n13726), .ZN(n13725) );
  NAND2_X1 U14740 ( .A1(n10752), .A2(n10739), .ZN(n11456) );
  AOI22_X1 U14741 ( .A1(n13725), .A2(n11456), .B1(n11022), .B2(n14498), .ZN(
        n11458) );
  OR2_X1 U14742 ( .A1(n14473), .A2(n11462), .ZN(n11463) );
  NAND2_X1 U14743 ( .A1(n11467), .A2(n11463), .ZN(n19808) );
  NOR2_X1 U14744 ( .A1(n17395), .A2(n16963), .ZN(n19807) );
  INV_X1 U14745 ( .A(n19807), .ZN(n16969) );
  NOR2_X1 U14746 ( .A1(n11464), .A2(n16969), .ZN(n19797) );
  NOR2_X1 U14747 ( .A1(n19808), .A2(n19797), .ZN(n19794) );
  NOR2_X1 U14748 ( .A1(n11465), .A2(n11022), .ZN(n11466) );
  NAND2_X1 U14749 ( .A1(n11467), .A2(n13756), .ZN(n19801) );
  NOR2_X1 U14750 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19807), .ZN(
        n19798) );
  INV_X1 U14751 ( .A(n19798), .ZN(n11483) );
  INV_X1 U14752 ( .A(n11467), .ZN(n11469) );
  NAND2_X1 U14753 ( .A1(n20484), .A2(n16993), .ZN(n13722) );
  OR2_X2 U14754 ( .A1(n13722), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U14755 ( .A1(n11469), .A2(n11468), .ZN(n19806) );
  OAI21_X1 U14756 ( .B1(n19801), .B2(n11483), .A(n19806), .ZN(n11470) );
  NOR2_X1 U14757 ( .A1(n19794), .A2(n11470), .ZN(n16952) );
  AND2_X2 U14758 ( .A1(n19801), .A2(n19808), .ZN(n17406) );
  INV_X1 U14759 ( .A(n17406), .ZN(n16970) );
  NAND2_X1 U14760 ( .A1(n16970), .A2(n16928), .ZN(n11471) );
  NOR2_X1 U14761 ( .A1(n16914), .A2(n16937), .ZN(n16913) );
  NAND2_X1 U14762 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16913), .ZN(
        n11472) );
  NAND2_X1 U14763 ( .A1(n16970), .A2(n11472), .ZN(n11473) );
  NAND2_X1 U14764 ( .A1(n16936), .A2(n11473), .ZN(n16902) );
  AND2_X1 U14765 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11481) );
  NOR2_X1 U14766 ( .A1(n17406), .A2(n11481), .ZN(n11474) );
  NOR2_X1 U14767 ( .A1(n17406), .A2(n11563), .ZN(n11475) );
  OR2_X1 U14768 ( .A1(n16872), .A2(n11475), .ZN(n16745) );
  NOR2_X1 U14769 ( .A1(n17406), .A2(n11487), .ZN(n11476) );
  NAND2_X1 U14770 ( .A1(n16936), .A2(n17406), .ZN(n16811) );
  NAND2_X1 U14771 ( .A1(n16811), .A2(n16705), .ZN(n11477) );
  NAND2_X1 U14772 ( .A1(n16719), .A2(n11477), .ZN(n16709) );
  AOI21_X1 U14773 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11478), .A(
        n17406), .ZN(n11479) );
  NOR2_X1 U14774 ( .A1(n16709), .A2(n11479), .ZN(n14967) );
  INV_X1 U14775 ( .A(n14967), .ZN(n11490) );
  NOR2_X1 U14776 ( .A1(n11468), .A2(n11480), .ZN(n14909) );
  INV_X1 U14777 ( .A(n11481), .ZN(n11486) );
  INV_X1 U14778 ( .A(n19797), .ZN(n11482) );
  NAND2_X1 U14779 ( .A1(n19801), .A2(n11482), .ZN(n11484) );
  NAND2_X1 U14780 ( .A1(n11484), .A2(n11483), .ZN(n16950) );
  NOR3_X1 U14781 ( .A1(n17406), .A2(n16928), .A3(n16950), .ZN(n16912) );
  NAND2_X1 U14782 ( .A1(n16913), .A2(n16912), .ZN(n14863) );
  NAND2_X1 U14783 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16884), .ZN(
        n11485) );
  NOR2_X2 U14784 ( .A1(n11486), .A2(n11485), .ZN(n16772) );
  NAND2_X1 U14785 ( .A1(n11563), .A2(n16772), .ZN(n16747) );
  INV_X1 U14786 ( .A(n11487), .ZN(n11488) );
  OR2_X1 U14787 ( .A1(n16747), .A2(n11488), .ZN(n16718) );
  NOR3_X1 U14788 ( .A1(n16693), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14968), .ZN(n11489) );
  AOI211_X1 U14789 ( .C1(n11490), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14909), .B(n11489), .ZN(n11491) );
  OAI21_X1 U14790 ( .B1(n15917), .B2(n19803), .A(n11491), .ZN(n11492) );
  AOI21_X1 U14791 ( .B1(n19792), .B2(n15908), .A(n11492), .ZN(n11493) );
  AND2_X1 U14793 ( .A1(n14498), .A2(n17047), .ZN(n11494) );
  INV_X1 U14794 ( .A(n13728), .ZN(n11496) );
  NAND2_X1 U14795 ( .A1(n11515), .A2(n19781), .ZN(n11514) );
  NAND2_X1 U14796 ( .A1(n11498), .A2(n11497), .ZN(n11503) );
  NAND2_X1 U14797 ( .A1(n11500), .A2(n11499), .ZN(n16647) );
  INV_X1 U14798 ( .A(n16645), .ZN(n11501) );
  NAND2_X1 U14799 ( .A1(n16644), .A2(n16648), .ZN(n11502) );
  XOR2_X1 U14800 ( .A(n11503), .B(n11502), .Z(n11516) );
  NAND2_X1 U14801 ( .A1(n11504), .A2(n11505), .ZN(n11506) );
  NOR2_X1 U14802 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17009) );
  OR2_X1 U14803 ( .A1(n20484), .A2(n17009), .ZN(n16986) );
  NAND2_X1 U14804 ( .A1(n16986), .A2(n17044), .ZN(n11507) );
  AND2_X1 U14805 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16984) );
  NAND2_X1 U14806 ( .A1(n20512), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15029) );
  NAND2_X1 U14807 ( .A1(n14608), .A2(n15029), .ZN(n19778) );
  NAND2_X1 U14808 ( .A1(n15001), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15004) );
  AND2_X1 U14809 ( .A1(n9733), .A2(n11508), .ZN(n11509) );
  OR2_X1 U14810 ( .A1(n11509), .A2(n14994), .ZN(n16130) );
  NOR2_X1 U14811 ( .A1(n11468), .A2(n20426), .ZN(n11520) );
  AOI21_X1 U14812 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n11520), .ZN(n11510) );
  OAI21_X1 U14813 ( .B1(n19758), .B2(n16130), .A(n11510), .ZN(n11511) );
  AOI21_X1 U14814 ( .B1(n16142), .B2(n19787), .A(n11511), .ZN(n11512) );
  NAND2_X1 U14815 ( .A1(n11514), .A2(n10423), .ZN(P2_U3004) );
  AOI21_X1 U14816 ( .B1(n11519), .B2(n11517), .A(n11262), .ZN(n14532) );
  INV_X1 U14817 ( .A(n16855), .ZN(n11523) );
  NAND2_X1 U14818 ( .A1(n16142), .A2(n16967), .ZN(n11522) );
  INV_X1 U14819 ( .A(n11520), .ZN(n11521) );
  OAI211_X1 U14820 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n11523), .A(
        n11522), .B(n11521), .ZN(n11527) );
  OAI21_X1 U14821 ( .B1(n16872), .B2(n11524), .A(n16811), .ZN(n16862) );
  NOR2_X1 U14822 ( .A1(n16862), .A2(n11525), .ZN(n11526) );
  AOI211_X1 U14823 ( .C1(n19792), .C2(n14532), .A(n11527), .B(n11526), .ZN(
        n11528) );
  XNOR2_X1 U14824 ( .A(n11534), .B(n10693), .ZN(n16498) );
  AND2_X1 U14825 ( .A1(n11534), .A2(n11533), .ZN(n11535) );
  AOI21_X1 U14826 ( .B1(n16498), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11535), .ZN(n11538) );
  XOR2_X1 U14827 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n11536), .Z(
        n11537) );
  XNOR2_X1 U14828 ( .A(n11538), .B(n11537), .ZN(n16497) );
  OR2_X1 U14829 ( .A1(n11540), .A2(n11541), .ZN(n11542) );
  NAND2_X1 U14830 ( .A1(n11539), .A2(n11542), .ZN(n16373) );
  INV_X1 U14831 ( .A(n16811), .ZN(n11544) );
  INV_X1 U14832 ( .A(n16709), .ZN(n11543) );
  OAI21_X1 U14833 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11544), .A(
        n11543), .ZN(n16695) );
  NAND2_X1 U14834 ( .A1(n19748), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16491) );
  OAI21_X1 U14835 ( .B1(n16693), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16491), .ZN(n11549) );
  NOR2_X1 U14836 ( .A1(n11545), .A2(n11546), .ZN(n11547) );
  OR2_X2 U14837 ( .A1(n15919), .A2(n11547), .ZN(n15933) );
  NOR2_X1 U14838 ( .A1(n15933), .A2(n19803), .ZN(n11548) );
  AOI211_X2 U14839 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16695), .A(
        n11549), .B(n11548), .ZN(n11550) );
  OAI21_X1 U14840 ( .B1(n16958), .B2(n16373), .A(n11550), .ZN(n11551) );
  OAI21_X1 U14841 ( .B1(n16497), .B2(n17400), .A(n11552), .ZN(P2_U3018) );
  AND2_X1 U14842 ( .A1(n16635), .A2(n16620), .ZN(n11554) );
  INV_X1 U14843 ( .A(n16634), .ZN(n16622) );
  AND2_X1 U14844 ( .A1(n16620), .A2(n16622), .ZN(n16618) );
  NAND2_X1 U14845 ( .A1(n11555), .A2(n10204), .ZN(n16621) );
  INV_X1 U14846 ( .A(n16621), .ZN(n16625) );
  INV_X1 U14847 ( .A(n16606), .ZN(n16582) );
  OR2_X1 U14848 ( .A1(n16582), .A2(n9780), .ZN(n12651) );
  OR2_X1 U14849 ( .A1(n12651), .A2(n11556), .ZN(n11557) );
  INV_X1 U14850 ( .A(n16544), .ZN(n11558) );
  NAND3_X1 U14851 ( .A1(n16541), .A2(n11558), .A3(n16543), .ZN(n11559) );
  NAND2_X1 U14852 ( .A1(n14760), .A2(n12662), .ZN(n13317) );
  INV_X1 U14853 ( .A(n11565), .ZN(n11567) );
  OAI21_X1 U14854 ( .B1(n11567), .B2(n10414), .A(n11566), .ZN(n16429) );
  INV_X1 U14855 ( .A(n11568), .ZN(n11570) );
  OAI21_X1 U14856 ( .B1(n11570), .B2(n10356), .A(n9754), .ZN(n16333) );
  INV_X1 U14857 ( .A(n16333), .ZN(n16025) );
  NOR2_X1 U14858 ( .A1(n11468), .A2(n20444), .ZN(n14916) );
  INV_X1 U14859 ( .A(n16772), .ZN(n16868) );
  NOR3_X1 U14860 ( .A1(n16760), .A2(n16758), .A3(n16868), .ZN(n11571) );
  MUX2_X1 U14861 ( .A(n11571), .B(n16745), .S(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(n11572) );
  AOI211_X1 U14862 ( .C1(n16025), .C2(n16967), .A(n14916), .B(n11572), .ZN(
        n11573) );
  OAI21_X1 U14863 ( .B1(n16958), .B2(n16429), .A(n11573), .ZN(n11574) );
  INV_X1 U14864 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17505) );
  NAND2_X1 U14865 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17151), .ZN(
        n17143) );
  NAND2_X1 U14866 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17743) );
  INV_X1 U14867 ( .A(n17743), .ZN(n18754) );
  NAND3_X1 U14868 ( .A1(n18720), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17689) );
  NAND2_X1 U14869 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18652) );
  NAND2_X1 U14870 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18629) );
  NAND2_X1 U14871 ( .A1(n18616), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18592) );
  NAND2_X1 U14872 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18594) );
  NAND2_X1 U14873 ( .A1(n18566), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18539) );
  NAND2_X1 U14874 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18542) );
  NAND2_X1 U14875 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14700) );
  XNOR2_X1 U14876 ( .A(n17505), .B(n11591), .ZN(n17504) );
  OR2_X1 U14877 ( .A1(n11577), .A2(n17860), .ZN(n11587) );
  INV_X1 U14878 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17106) );
  NOR2_X1 U14879 ( .A1(n11587), .A2(n17106), .ZN(n11590) );
  AND2_X1 U14880 ( .A1(n11587), .A2(n17106), .ZN(n11578) );
  NOR2_X1 U14881 ( .A1(n11590), .A2(n11578), .ZN(n17538) );
  INV_X1 U14882 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17598) );
  INV_X1 U14883 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17618) );
  INV_X1 U14884 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17132) );
  NAND2_X1 U14885 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17133), .ZN(
        n17650) );
  INV_X1 U14886 ( .A(n17131), .ZN(n17124) );
  NOR2_X1 U14887 ( .A1(n18629), .A2(n17124), .ZN(n18590) );
  INV_X1 U14888 ( .A(n18590), .ZN(n17627) );
  NOR2_X1 U14889 ( .A1(n17618), .A2(n17627), .ZN(n11584) );
  NAND2_X1 U14890 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11584), .ZN(
        n11585) );
  NAND2_X1 U14891 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18561), .ZN(
        n11582) );
  NOR2_X1 U14892 ( .A1(n18542), .A2(n11582), .ZN(n14694) );
  OAI21_X1 U14893 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n14694), .A(
        n11587), .ZN(n11579) );
  INV_X1 U14894 ( .A(n11579), .ZN(n17550) );
  INV_X1 U14895 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18557) );
  NOR2_X1 U14896 ( .A1(n18557), .A2(n11582), .ZN(n11581) );
  INV_X1 U14897 ( .A(n14694), .ZN(n11580) );
  OAI21_X1 U14898 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n11581), .A(
        n11580), .ZN(n18544) );
  INV_X1 U14899 ( .A(n18544), .ZN(n17561) );
  AOI21_X1 U14900 ( .B1(n18557), .B2(n11582), .A(n11581), .ZN(n18555) );
  OAI21_X1 U14901 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18561), .A(
        n11582), .ZN(n18562) );
  INV_X1 U14902 ( .A(n18562), .ZN(n17582) );
  AOI21_X1 U14903 ( .B1(n17618), .B2(n17627), .A(n11584), .ZN(n18621) );
  INV_X1 U14904 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18664) );
  NOR2_X1 U14905 ( .A1(n17860), .A2(n18646), .ZN(n18649) );
  INV_X1 U14906 ( .A(n18649), .ZN(n17690) );
  NOR2_X1 U14907 ( .A1(n18664), .A2(n17690), .ZN(n17672) );
  NAND2_X1 U14908 ( .A1(n17854), .A2(n17672), .ZN(n17666) );
  INV_X1 U14909 ( .A(n17666), .ZN(n17667) );
  XNOR2_X2 U14910 ( .A(n11583), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11593) );
  OAI21_X1 U14911 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11584), .A(
        n11585), .ZN(n18602) );
  INV_X1 U14912 ( .A(n18602), .ZN(n17607) );
  AOI21_X1 U14913 ( .B1(n17598), .B2(n11585), .A(n18561), .ZN(n18589) );
  NOR2_X1 U14914 ( .A1(n17580), .A2(n17820), .ZN(n17573) );
  NOR2_X1 U14915 ( .A1(n18555), .A2(n17573), .ZN(n17572) );
  NOR2_X1 U14916 ( .A1(n17572), .A2(n17820), .ZN(n17560) );
  NOR2_X1 U14917 ( .A1(n17561), .A2(n17560), .ZN(n17559) );
  NOR2_X1 U14918 ( .A1(n17559), .A2(n17820), .ZN(n17549) );
  NOR2_X1 U14919 ( .A1(n17550), .A2(n17549), .ZN(n17548) );
  NOR2_X1 U14920 ( .A1(n17548), .A2(n17820), .ZN(n17537) );
  NOR2_X1 U14921 ( .A1(n17538), .A2(n17537), .ZN(n17536) );
  OR2_X1 U14922 ( .A1(n17536), .A2(n17820), .ZN(n17526) );
  INV_X1 U14923 ( .A(n11587), .ZN(n11589) );
  INV_X1 U14924 ( .A(n14700), .ZN(n11588) );
  NAND2_X1 U14925 ( .A1(n11589), .A2(n11588), .ZN(n17089) );
  OAI21_X1 U14926 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11590), .A(
        n17089), .ZN(n14703) );
  INV_X1 U14927 ( .A(n14703), .ZN(n17530) );
  NAND2_X1 U14928 ( .A1(n17526), .A2(n14703), .ZN(n17527) );
  AOI21_X1 U14929 ( .B1(n17089), .B2(n10088), .A(n11591), .ZN(n17515) );
  INV_X1 U14930 ( .A(n17515), .ZN(n11592) );
  NAND2_X1 U14931 ( .A1(n17511), .A2(n11592), .ZN(n17512) );
  NAND3_X1 U14932 ( .A1(n19515), .A2(n19512), .A3(n19625), .ZN(n19513) );
  NOR2_X2 U14933 ( .A1(n18425), .A2(n19513), .ZN(n17837) );
  NAND2_X1 U14934 ( .A1(n11593), .A2(n17837), .ZN(n17853) );
  NOR3_X1 U14935 ( .A1(n17504), .A2(n17503), .A3(n17853), .ZN(n11764) );
  INV_X1 U14936 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18223) );
  AND2_X2 U14937 ( .A1(n13907), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11609) );
  AOI22_X1 U14938 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11596) );
  NAND2_X2 U14939 ( .A1(n14675), .A2(n11598), .ZN(n18224) );
  INV_X1 U14940 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11594) );
  OAI211_X1 U14941 ( .C1(n18223), .C2(n9702), .A(n11596), .B(n11595), .ZN(
        n11597) );
  INV_X1 U14942 ( .A(n11597), .ZN(n11615) );
  NAND2_X1 U14943 ( .A1(n11609), .A2(n11600), .ZN(n13055) );
  AOI22_X1 U14944 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11605) );
  AND2_X2 U14945 ( .A1(n11608), .A2(n11599), .ZN(n17890) );
  AOI22_X1 U14946 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18152), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11604) );
  INV_X2 U14947 ( .A(n18085), .ZN(n18207) );
  AOI22_X1 U14948 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11603) );
  NOR2_X1 U14949 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14950 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14951 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11613) );
  AND2_X2 U14952 ( .A1(n11606), .A2(n13906), .ZN(n13086) );
  INV_X1 U14953 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18062) );
  AND2_X2 U14954 ( .A1(n13884), .A2(n11607), .ZN(n13047) );
  INV_X1 U14955 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18061) );
  OAI22_X1 U14956 ( .A1(n13142), .A2(n18062), .B1(n18198), .B2(n18061), .ZN(
        n11611) );
  INV_X1 U14957 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14373) );
  OAI22_X1 U14958 ( .A1(n18203), .A2(n14373), .B1(n9745), .B2(n14375), .ZN(
        n11610) );
  INV_X2 U14959 ( .A(n13055), .ZN(n11663) );
  INV_X2 U14960 ( .A(n11663), .ZN(n18141) );
  NAND2_X1 U14961 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U14962 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11616) );
  OAI211_X1 U14963 ( .C1(n18038), .C2(n18141), .A(n11617), .B(n11616), .ZN(
        n11618) );
  INV_X1 U14964 ( .A(n11618), .ZN(n11622) );
  AOI22_X1 U14965 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14966 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11620) );
  INV_X1 U14967 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18197) );
  NAND4_X1 U14968 ( .A1(n11622), .A2(n11621), .A3(n11620), .A4(n11619), .ZN(
        n11628) );
  AOI22_X1 U14969 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14970 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14971 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14972 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14973 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11627) );
  NAND2_X1 U14974 ( .A1(n19035), .A2(n18490), .ZN(n13892) );
  INV_X1 U14975 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18081) );
  INV_X1 U14976 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11629) );
  OR2_X1 U14977 ( .A1(n18224), .A2(n11629), .ZN(n11632) );
  NAND2_X1 U14978 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U14979 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11630) );
  INV_X2 U14980 ( .A(n9745), .ZN(n18194) );
  NAND2_X1 U14981 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U14982 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11636) );
  NAND2_X1 U14983 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14984 ( .A1(n9701), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14985 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11641) );
  INV_X2 U14986 ( .A(n18203), .ZN(n18134) );
  NAND2_X1 U14987 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U14988 ( .A1(n13086), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U14989 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14990 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U14991 ( .A1(n9707), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U14992 ( .A1(n13929), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14993 ( .A1(n18222), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11642) );
  INV_X1 U14994 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U14995 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11651) );
  NAND2_X1 U14996 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11650) );
  OAI211_X1 U14997 ( .C1(n14345), .C2(n18141), .A(n11651), .B(n11650), .ZN(
        n11652) );
  INV_X1 U14998 ( .A(n11652), .ZN(n11656) );
  AOI22_X1 U14999 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U15000 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11654) );
  OR2_X1 U15001 ( .A1(n18224), .A2(n21780), .ZN(n11653) );
  NAND4_X1 U15002 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11662) );
  AOI22_X1 U15003 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U15004 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U15005 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U15006 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U15007 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11661) );
  INV_X1 U15008 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U15009 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11665) );
  NAND2_X1 U15010 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11664) );
  OAI211_X1 U15011 ( .C1(n11666), .C2(n18141), .A(n11665), .B(n11664), .ZN(
        n11667) );
  INV_X1 U15012 ( .A(n11667), .ZN(n11671) );
  AOI22_X1 U15013 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U15014 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11669) );
  INV_X1 U15015 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17969) );
  OR2_X1 U15016 ( .A1(n18224), .A2(n17969), .ZN(n11668) );
  NAND4_X1 U15017 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n11677) );
  AOI22_X1 U15018 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18207), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U15019 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13086), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U15020 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U15021 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11672) );
  NAND4_X1 U15022 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(
        n11676) );
  INV_X1 U15023 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18025) );
  NAND2_X1 U15024 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11679) );
  NAND2_X1 U15025 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11678) );
  OAI211_X1 U15026 ( .C1(n18025), .C2(n18080), .A(n11679), .B(n11678), .ZN(
        n11680) );
  INV_X1 U15027 ( .A(n11680), .ZN(n11685) );
  AOI22_X1 U15028 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U15029 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11683) );
  INV_X1 U15030 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11681) );
  OR2_X1 U15031 ( .A1(n18224), .A2(n11681), .ZN(n11682) );
  NAND4_X1 U15032 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11691) );
  AOI22_X1 U15033 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18207), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U15034 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U15035 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U15036 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U15037 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11690) );
  AOI22_X1 U15038 ( .A1(n13086), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17886), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U15039 ( .A1(n9701), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11696) );
  INV_X1 U15040 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U15041 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18152), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11692) );
  OAI21_X1 U15042 ( .B1(n14388), .B2(n11693), .A(n11692), .ZN(n11694) );
  AOI21_X1 U15043 ( .B1(n18180), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11694), .ZN(n11695) );
  AOI22_X1 U15044 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U15045 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18207), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U15046 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U15047 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11663), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U15048 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11704) );
  NAND2_X1 U15049 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11703) );
  OAI211_X1 U15050 ( .C1(n21736), .C2(n18141), .A(n11704), .B(n11703), .ZN(
        n11705) );
  INV_X1 U15051 ( .A(n11705), .ZN(n11710) );
  AOI22_X1 U15052 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U15053 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11708) );
  INV_X1 U15054 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11706) );
  OR2_X1 U15055 ( .A1(n18224), .A2(n11706), .ZN(n11707) );
  NAND4_X1 U15056 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11717) );
  AOI22_X1 U15057 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U15058 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U15059 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U15060 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11712) );
  NAND4_X1 U15061 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  NAND2_X1 U15062 ( .A1(n19035), .A2(n18364), .ZN(n11730) );
  NAND2_X1 U15063 ( .A1(n18428), .A2(n19626), .ZN(n13288) );
  INV_X1 U15064 ( .A(n14218), .ZN(n13885) );
  AND2_X1 U15065 ( .A1(n18364), .A2(n13885), .ZN(n11718) );
  NOR2_X1 U15066 ( .A1(n13288), .A2(n11718), .ZN(n13226) );
  INV_X1 U15067 ( .A(n13226), .ZN(n11719) );
  OAI21_X1 U15068 ( .B1(n13289), .B2(n11720), .A(n11719), .ZN(n11726) );
  AOI22_X1 U15069 ( .A1(n19046), .A2(n11730), .B1(n19051), .B2(n14218), .ZN(
        n11725) );
  NAND2_X1 U15070 ( .A1(n19042), .A2(n13892), .ZN(n13221) );
  AOI21_X1 U15071 ( .B1(n18364), .B2(n11722), .A(n19051), .ZN(n11721) );
  AOI21_X1 U15072 ( .B1(n11722), .B2(n13221), .A(n11721), .ZN(n11724) );
  NAND2_X1 U15073 ( .A1(n19058), .A2(n13223), .ZN(n13910) );
  NOR2_X1 U15074 ( .A1(n19058), .A2(n18286), .ZN(n13222) );
  INV_X1 U15075 ( .A(n13222), .ZN(n11729) );
  NAND4_X1 U15076 ( .A1(n19042), .A2(n19035), .A3(n13910), .A4(n11729), .ZN(
        n11723) );
  NAND2_X1 U15077 ( .A1(n19046), .A2(n19042), .ZN(n13909) );
  NOR2_X1 U15078 ( .A1(n11730), .A2(n14214), .ZN(n11731) );
  AND2_X1 U15079 ( .A1(n11731), .A2(n19626), .ZN(n11732) );
  OR2_X2 U15080 ( .A1(n13284), .A2(n11732), .ZN(n13886) );
  MUX2_X1 U15081 ( .A(n19478), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13236) );
  NAND2_X1 U15082 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19477), .ZN(
        n13229) );
  INV_X1 U15083 ( .A(n13229), .ZN(n11748) );
  NAND2_X1 U15084 ( .A1(n13236), .A2(n11748), .ZN(n11746) );
  NAND2_X1 U15085 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19478), .ZN(
        n11733) );
  NAND2_X1 U15086 ( .A1(n11746), .A2(n11733), .ZN(n11744) );
  MUX2_X1 U15087 ( .A(n19028), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11743) );
  NOR2_X1 U15088 ( .A1(n13907), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11734) );
  AOI21_X1 U15089 ( .B1(n11744), .B2(n11743), .A(n11734), .ZN(n11735) );
  AOI21_X1 U15090 ( .B1(n11735), .B2(n19488), .A(n11739), .ZN(n11738) );
  OR2_X1 U15091 ( .A1(n11735), .A2(n19488), .ZN(n11740) );
  NAND2_X1 U15092 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11740), .ZN(
        n11736) );
  AOI22_X1 U15093 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19494), .B1(
        n11738), .B2(n11736), .ZN(n13240) );
  INV_X1 U15094 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11737) );
  OR2_X1 U15095 ( .A1(n11738), .A2(n11737), .ZN(n11742) );
  NAND2_X1 U15096 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  NAND2_X1 U15097 ( .A1(n11742), .A2(n11741), .ZN(n13238) );
  XNOR2_X1 U15098 ( .A(n11744), .B(n11743), .ZN(n11745) );
  INV_X1 U15099 ( .A(n13239), .ZN(n11747) );
  OAI211_X1 U15100 ( .C1(n13236), .C2(n11748), .A(n11747), .B(n11746), .ZN(
        n11749) );
  NAND2_X1 U15101 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18490), .ZN(n11750) );
  AOI211_X4 U15102 ( .C1(n19625), .C2(n19627), .A(n19640), .B(n11750), .ZN(
        n17829) );
  INV_X1 U15103 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18238) );
  NAND2_X1 U15104 ( .A1(n17833), .A2(n18255), .ZN(n17828) );
  NOR2_X1 U15105 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17828), .ZN(n17801) );
  NAND2_X1 U15106 ( .A1(n17801), .A2(n18091), .ZN(n17796) );
  NOR2_X1 U15107 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17796), .ZN(n17779) );
  INV_X1 U15108 ( .A(n17779), .ZN(n17765) );
  NOR2_X1 U15109 ( .A1(n17765), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17764) );
  INV_X1 U15110 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17740) );
  NAND2_X1 U15111 ( .A1(n17746), .A2(n17740), .ZN(n17728) );
  NAND2_X1 U15112 ( .A1(n17727), .A2(n21783), .ZN(n17724) );
  NAND2_X1 U15113 ( .A1(n17708), .A2(n18129), .ZN(n17705) );
  INV_X1 U15114 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17678) );
  NAND2_X1 U15115 ( .A1(n17683), .A2(n17678), .ZN(n17676) );
  NAND2_X1 U15116 ( .A1(n17661), .A2(n18050), .ZN(n17654) );
  INV_X1 U15117 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17633) );
  NAND2_X1 U15118 ( .A1(n17639), .A2(n17633), .ZN(n17631) );
  INV_X1 U15119 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17979) );
  NAND2_X1 U15120 ( .A1(n17617), .A2(n17979), .ZN(n17611) );
  INV_X1 U15121 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17586) );
  NAND2_X1 U15122 ( .A1(n17593), .A2(n17586), .ZN(n17585) );
  INV_X1 U15123 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17874) );
  NAND2_X1 U15124 ( .A1(n17571), .A2(n17874), .ZN(n17563) );
  INV_X1 U15125 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17543) );
  NAND2_X1 U15126 ( .A1(n17547), .A2(n17543), .ZN(n17542) );
  INV_X1 U15127 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17875) );
  NAND2_X1 U15128 ( .A1(n17525), .A2(n17875), .ZN(n17502) );
  NOR2_X1 U15129 ( .A1(n17864), .A2(n17502), .ZN(n17508) );
  INV_X1 U15130 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17880) );
  NAND2_X1 U15131 ( .A1(n17508), .A2(n17880), .ZN(n11762) );
  INV_X1 U15132 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19588) );
  INV_X1 U15133 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n17483) );
  NAND2_X2 U15134 ( .A1(n19635), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19593) );
  NAND2_X1 U15135 ( .A1(n17481), .A2(n19537), .ZN(n19522) );
  AOI211_X1 U15136 ( .C1(n19624), .C2(n19626), .A(n19529), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n11754) );
  INV_X1 U15137 ( .A(n11754), .ZN(n19502) );
  NAND2_X1 U15138 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17524) );
  NAND2_X1 U15139 ( .A1(n18425), .A2(n19512), .ZN(n14680) );
  INV_X1 U15140 ( .A(n14680), .ZN(n19630) );
  NAND3_X1 U15141 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .A3(n19630), .ZN(n11751) );
  AND3_X1 U15142 ( .A1(n10420), .A2(n17823), .A3(n11751), .ZN(n11752) );
  INV_X1 U15143 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19583) );
  INV_X1 U15144 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19580) );
  INV_X1 U15145 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19576) );
  INV_X1 U15146 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21741) );
  INV_X1 U15147 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19551) );
  NAND3_X1 U15148 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17818) );
  NOR2_X1 U15149 ( .A1(n19543), .A2(n17818), .ZN(n17791) );
  NAND2_X1 U15150 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17791), .ZN(n17783) );
  NOR2_X1 U15151 ( .A1(n19546), .A2(n17783), .ZN(n17766) );
  NAND2_X1 U15152 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17766), .ZN(n17754) );
  NOR2_X1 U15153 ( .A1(n19551), .A2(n17754), .ZN(n17730) );
  NAND4_X1 U15154 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17730), .A3(
        P3_REIP_REG_9__SCAN_IN), .A4(P3_REIP_REG_10__SCAN_IN), .ZN(n17714) );
  NOR2_X1 U15155 ( .A1(n19558), .A2(n17714), .ZN(n17614) );
  NAND3_X1 U15156 ( .A1(n17614), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .ZN(n17625) );
  NAND3_X1 U15157 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_17__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n17626) );
  NAND2_X1 U15158 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17636) );
  NOR4_X1 U15159 ( .A1(n21741), .A2(n17625), .A3(n17626), .A4(n17636), .ZN(
        n17592) );
  NAND2_X1 U15160 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17592), .ZN(n17596) );
  NOR2_X1 U15161 ( .A1(n19576), .A2(n17596), .ZN(n17578) );
  NAND2_X1 U15162 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17578), .ZN(n17558) );
  NOR2_X1 U15163 ( .A1(n19580), .A2(n17558), .ZN(n17564) );
  NAND2_X1 U15164 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17564), .ZN(n17557) );
  NOR2_X1 U15165 ( .A1(n19583), .A2(n17557), .ZN(n11753) );
  OR2_X1 U15166 ( .A1(n17857), .A2(n11753), .ZN(n17556) );
  NAND2_X1 U15167 ( .A1(n17868), .A2(n17556), .ZN(n17553) );
  AOI221_X1 U15168 ( .B1(n19588), .B2(n17846), .C1(n17524), .C2(n17846), .A(
        n17553), .ZN(n17523) );
  NAND2_X1 U15169 ( .A1(n17846), .A2(n11753), .ZN(n17539) );
  NOR2_X1 U15170 ( .A1(n17539), .A2(n17524), .ZN(n17518) );
  NAND2_X1 U15171 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17518), .ZN(n11755) );
  INV_X1 U15172 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19591) );
  AOI21_X1 U15173 ( .B1(n17523), .B2(n10383), .A(n19591), .ZN(n11760) );
  AOI211_X4 U15174 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18490), .A(n11754), .B(
        n19640), .ZN(n17804) );
  INV_X1 U15175 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21720) );
  NOR3_X1 U15176 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21720), .A3(n11755), 
        .ZN(n11756) );
  AOI21_X1 U15177 ( .B1(n17804), .B2(P3_EBX_REG_31__SCAN_IN), .A(n11756), .ZN(
        n11758) );
  INV_X1 U15178 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17067) );
  OR2_X1 U15179 ( .A1(n17852), .A2(n17067), .ZN(n11757) );
  NAND2_X1 U15180 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  NAND2_X1 U15181 ( .A1(n11762), .A2(n11761), .ZN(n11763) );
  INV_X1 U15182 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11765) );
  AND2_X2 U15183 ( .A1(n11765), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15184 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11769) );
  NAND2_X1 U15185 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11768) );
  NAND2_X1 U15186 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11767) );
  AND2_X2 U15187 ( .A1(n13841), .A2(n14182), .ZN(n11913) );
  NAND2_X1 U15188 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11766) );
  INV_X1 U15189 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11770) );
  NAND2_X1 U15190 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U15191 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U15192 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11772) );
  NAND2_X1 U15193 ( .A1(n12011), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11771) );
  NAND2_X1 U15194 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U15195 ( .A1(n12012), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U15196 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11776) );
  NAND3_X1 U15197 ( .A1(n11778), .A2(n11777), .A3(n11776), .ZN(n11779) );
  AND2_X2 U15198 ( .A1(n11781), .A2(n11782), .ZN(n11975) );
  NAND2_X1 U15199 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U15200 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U15201 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U15202 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U15203 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U15204 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11793) );
  NAND2_X1 U15205 ( .A1(n12012), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U15206 ( .A1(n11912), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U15207 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U15208 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U15209 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U15210 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U15211 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U15212 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11800) );
  NAND2_X1 U15213 ( .A1(n12011), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U15214 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U15215 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U15216 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U15217 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11803) );
  INV_X1 U15218 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11811) );
  OR2_X1 U15219 ( .A1(n12222), .A2(n11811), .ZN(n11837) );
  INV_X1 U15220 ( .A(n11887), .ZN(n12035) );
  AOI22_X1 U15221 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U15222 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U15223 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U15224 ( .A1(n14775), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U15225 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11823) );
  AOI22_X1 U15226 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U15227 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U15228 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U15229 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U15230 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11822) );
  INV_X1 U15231 ( .A(n12173), .ZN(n12169) );
  NAND2_X1 U15232 ( .A1(n11992), .A2(n12169), .ZN(n11836) );
  AOI22_X1 U15233 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U15234 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U15235 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U15236 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U15237 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11834) );
  AOI22_X1 U15238 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U15239 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U15240 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U15241 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11829) );
  NAND4_X1 U15242 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n11833) );
  NAND2_X1 U15243 ( .A1(n10019), .A2(n12100), .ZN(n11835) );
  INV_X1 U15244 ( .A(n12275), .ZN(n11994) );
  AND2_X1 U15245 ( .A1(n11912), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11839) );
  NOR2_X1 U15246 ( .A1(n11839), .A2(n11838), .ZN(n11843) );
  AOI22_X1 U15247 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U15248 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15249 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U15250 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U15251 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15252 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11896), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11845) );
  INV_X1 U15253 ( .A(n12266), .ZN(n11859) );
  AOI22_X1 U15254 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U15255 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14776), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U15256 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12012), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15257 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15258 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U15259 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U15260 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11912), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U15261 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11854) );
  NAND2_X1 U15262 ( .A1(n11859), .A2(n11925), .ZN(n11965) );
  AOI22_X1 U15263 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U15264 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12636), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11863) );
  AOI21_X1 U15265 ( .B1(n11912), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n11861), .ZN(n11862) );
  NAND3_X1 U15266 ( .A1(n9768), .A2(n11863), .A3(n11862), .ZN(n11869) );
  AOI22_X1 U15267 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U15268 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U15269 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11864) );
  NAND4_X1 U15270 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11868) );
  AOI22_X1 U15271 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12636), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15272 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U15273 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U15274 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11881) );
  AOI22_X1 U15275 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14776), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15276 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11896), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15277 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U15278 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U15279 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11880) );
  AOI22_X1 U15280 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U15281 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U15282 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U15283 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15284 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U15285 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12012), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U15286 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U15287 ( .A1(n12249), .A2(n20808), .ZN(n12102) );
  INV_X1 U15288 ( .A(n11936), .ZN(n11922) );
  NAND2_X1 U15289 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U15290 ( .A1(n11975), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11899) );
  NAND2_X1 U15291 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U15292 ( .A1(n11896), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11897) );
  NAND2_X1 U15293 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15294 ( .A1(n12011), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11904) );
  NAND2_X1 U15295 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11903) );
  NAND2_X1 U15296 ( .A1(n12012), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11902) );
  NAND2_X1 U15297 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U15298 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11910) );
  NAND2_X1 U15299 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U15300 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U15301 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15302 ( .A1(n11912), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11915) );
  NAND2_X1 U15303 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U15304 ( .A1(n12266), .A2(n14143), .ZN(n11923) );
  NOR2_X1 U15305 ( .A1(n11927), .A2(n11940), .ZN(n11924) );
  NAND4_X1 U15306 ( .A1(n11959), .A2(n11924), .A3(n13369), .A4(n11942), .ZN(
        n13366) );
  NAND2_X1 U15307 ( .A1(n14143), .A2(n11936), .ZN(n12200) );
  INV_X1 U15308 ( .A(n12200), .ZN(n11930) );
  INV_X1 U15309 ( .A(n11927), .ZN(n11929) );
  NOR2_X1 U15310 ( .A1(n11940), .A2(n12266), .ZN(n11928) );
  NAND3_X1 U15311 ( .A1(n11930), .A2(n11929), .A3(n11928), .ZN(n13742) );
  NAND2_X1 U15312 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21385) );
  OAI21_X1 U15313 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n21385), .ZN(n13340) );
  INV_X1 U15314 ( .A(n13340), .ZN(n11932) );
  NAND2_X1 U15315 ( .A1(n13730), .A2(n11932), .ZN(n11933) );
  INV_X2 U15316 ( .A(n11949), .ZN(n13823) );
  NAND2_X1 U15317 ( .A1(n20796), .A2(n20776), .ZN(n11941) );
  OAI211_X1 U15318 ( .C1(n13874), .C2(n11957), .A(n13484), .B(n11941), .ZN(
        n11961) );
  INV_X1 U15319 ( .A(n20800), .ZN(n13370) );
  NOR2_X1 U15320 ( .A1(n11961), .A2(n13370), .ZN(n11946) );
  INV_X1 U15321 ( .A(n12266), .ZN(n12282) );
  INV_X1 U15322 ( .A(n12248), .ZN(n11944) );
  NAND2_X1 U15323 ( .A1(n11944), .A2(n13874), .ZN(n13346) );
  NAND2_X1 U15324 ( .A1(n13346), .A2(n11945), .ZN(n11954) );
  NAND2_X1 U15325 ( .A1(n13487), .A2(n20796), .ZN(n11947) );
  NAND2_X1 U15326 ( .A1(n21302), .A2(n21677), .ZN(n21198) );
  NAND2_X1 U15327 ( .A1(n21198), .A2(n21166), .ZN(n21120) );
  NAND2_X1 U15328 ( .A1(n21370), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11998) );
  OAI21_X1 U15329 ( .B1(n12264), .B2(n21120), .A(n11998), .ZN(n11950) );
  INV_X1 U15330 ( .A(n11950), .ZN(n11951) );
  INV_X1 U15331 ( .A(n21370), .ZN(n11952) );
  MUX2_X1 U15332 ( .A(n11952), .B(n12264), .S(n21677), .Z(n11953) );
  NAND2_X1 U15333 ( .A1(n14727), .A2(n20792), .ZN(n15352) );
  INV_X1 U15334 ( .A(n14944), .ZN(n11955) );
  NOR2_X1 U15335 ( .A1(n11955), .A2(n21369), .ZN(n11956) );
  AND2_X1 U15336 ( .A1(n15352), .A2(n11956), .ZN(n11963) );
  NAND2_X1 U15337 ( .A1(n11958), .A2(n12282), .ZN(n13495) );
  OAI21_X1 U15338 ( .B1(n11957), .B2(n11959), .A(n13495), .ZN(n11960) );
  NOR2_X1 U15339 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  NAND3_X1 U15340 ( .A1(n15351), .A2(n11965), .A3(n20800), .ZN(n11966) );
  NAND2_X1 U15341 ( .A1(n11964), .A2(n11966), .ZN(n11967) );
  OAI211_X1 U15342 ( .C1(n11954), .C2(n13823), .A(n10428), .B(n11967), .ZN(
        n11970) );
  NAND2_X1 U15343 ( .A1(n11992), .A2(n12100), .ZN(n11969) );
  INV_X1 U15344 ( .A(n11970), .ZN(n11971) );
  XNOR2_X1 U15345 ( .A(n11972), .B(n11971), .ZN(n12284) );
  NAND2_X1 U15346 ( .A1(n12284), .A2(n21369), .ZN(n11988) );
  AOI22_X1 U15348 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15349 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13615), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15350 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15351 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11976) );
  NAND4_X1 U15352 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11985) );
  AOI22_X1 U15353 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15354 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13632), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15355 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11906), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15356 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11912), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11980) );
  NAND4_X1 U15357 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11984) );
  XNOR2_X1 U15358 ( .A(n12101), .B(n12173), .ZN(n11986) );
  NAND2_X1 U15359 ( .A1(n11986), .A2(n11992), .ZN(n11987) );
  NAND2_X1 U15360 ( .A1(n11988), .A2(n11987), .ZN(n12106) );
  AOI21_X1 U15361 ( .B1(n13874), .B2(n12173), .A(n21369), .ZN(n11990) );
  NAND2_X1 U15362 ( .A1(n14727), .A2(n12107), .ZN(n11989) );
  NAND2_X1 U15363 ( .A1(n11992), .A2(n12173), .ZN(n11993) );
  NAND2_X1 U15364 ( .A1(n12099), .A2(n11995), .ZN(n12273) );
  AND2_X1 U15365 ( .A1(n11997), .A2(n11998), .ZN(n11999) );
  NAND2_X1 U15366 ( .A1(n12007), .A2(n12005), .ZN(n12003) );
  XNOR2_X1 U15367 ( .A(n21166), .B(n21066), .ZN(n20785) );
  NOR2_X1 U15368 ( .A1(n20785), .A2(n12264), .ZN(n12001) );
  NAND2_X1 U15369 ( .A1(n21370), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U15370 ( .A1(n12006), .A2(n12004), .ZN(n12002) );
  NAND4_X1 U15371 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(
        n12008) );
  INV_X1 U15372 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21706) );
  AOI22_X1 U15373 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15374 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15375 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15376 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12013) );
  NAND4_X1 U15377 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12022) );
  AOI22_X1 U15378 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15379 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15380 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15381 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12017) );
  NAND4_X1 U15382 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n12021) );
  INV_X1 U15383 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12023) );
  INV_X1 U15384 ( .A(n12082), .ZN(n12050) );
  NAND2_X1 U15385 ( .A1(n12027), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12032) );
  OAI21_X1 U15386 ( .B1(n21166), .B2(n21066), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12029) );
  INV_X1 U15387 ( .A(n21166), .ZN(n21300) );
  NAND2_X1 U15388 ( .A1(n21474), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20997) );
  INV_X1 U15389 ( .A(n20997), .ZN(n12028) );
  NAND2_X1 U15390 ( .A1(n21300), .A2(n12028), .ZN(n21035) );
  NAND2_X1 U15391 ( .A1(n12029), .A2(n21035), .ZN(n21067) );
  INV_X1 U15392 ( .A(n12264), .ZN(n12030) );
  AOI22_X1 U15393 ( .A1(n21067), .A2(n12030), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21370), .ZN(n12031) );
  AOI22_X1 U15394 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15395 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15396 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15397 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12036) );
  NAND4_X1 U15398 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12045) );
  AOI22_X1 U15399 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15400 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15401 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15402 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12040) );
  NAND4_X1 U15403 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12044) );
  NAND2_X1 U15404 ( .A1(n12246), .A2(n12088), .ZN(n12046) );
  OAI21_X1 U15405 ( .B1(n12047), .B2(n12222), .A(n12046), .ZN(n12048) );
  NAND2_X2 U15406 ( .A1(n12050), .A2(n12049), .ZN(n12087) );
  AOI22_X1 U15407 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15408 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15409 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15410 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12051) );
  NAND4_X1 U15411 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12060) );
  AOI22_X1 U15412 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15413 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15414 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15415 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U15416 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12059) );
  NAND2_X1 U15417 ( .A1(n12246), .A2(n12090), .ZN(n12063) );
  INV_X1 U15418 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12061) );
  NAND2_X1 U15419 ( .A1(n12234), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12076) );
  AOI22_X1 U15420 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15421 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15422 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15423 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12065) );
  NAND4_X1 U15424 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12074) );
  AOI22_X1 U15425 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15426 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15427 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15428 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12069) );
  NAND4_X1 U15429 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12073) );
  NAND2_X1 U15430 ( .A1(n12246), .A2(n12159), .ZN(n12075) );
  NAND2_X1 U15431 ( .A1(n12100), .A2(n12107), .ZN(n12095) );
  NAND2_X1 U15432 ( .A1(n12095), .A2(n12094), .ZN(n12089) );
  AND2_X1 U15433 ( .A1(n12088), .A2(n12090), .ZN(n12079) );
  NAND2_X1 U15434 ( .A1(n12089), .A2(n12079), .ZN(n12161) );
  XNOR2_X1 U15435 ( .A(n12161), .B(n12159), .ZN(n12080) );
  INV_X1 U15436 ( .A(n11957), .ZN(n12174) );
  NAND2_X1 U15437 ( .A1(n12080), .A2(n12174), .ZN(n12081) );
  INV_X1 U15438 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17326) );
  NAND2_X1 U15439 ( .A1(n12082), .A2(n20773), .ZN(n20936) );
  INV_X1 U15440 ( .A(n12293), .ZN(n12083) );
  INV_X1 U15441 ( .A(n12088), .ZN(n12084) );
  XNOR2_X1 U15442 ( .A(n12089), .B(n12084), .ZN(n12085) );
  NAND2_X1 U15443 ( .A1(n12085), .A2(n12174), .ZN(n12124) );
  XNOR2_X1 U15444 ( .A(n12087), .B(n12086), .ZN(n12309) );
  NAND2_X1 U15445 ( .A1(n12089), .A2(n12088), .ZN(n12091) );
  XNOR2_X1 U15446 ( .A(n12091), .B(n12090), .ZN(n12092) );
  NAND2_X1 U15447 ( .A1(n12092), .A2(n12174), .ZN(n12093) );
  NAND3_X1 U15448 ( .A1(n14574), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U15449 ( .A1(n15905), .A2(n14029), .ZN(n12098) );
  XNOR2_X1 U15450 ( .A(n12095), .B(n12094), .ZN(n12096) );
  AND2_X1 U15451 ( .A1(n14727), .A2(n20800), .ZN(n12108) );
  AOI21_X1 U15452 ( .B1(n12096), .B2(n12174), .A(n12108), .ZN(n12097) );
  NAND2_X1 U15453 ( .A1(n12098), .A2(n12097), .ZN(n14630) );
  OR2_X1 U15454 ( .A1(n12099), .A2(n13823), .ZN(n12105) );
  XNOR2_X1 U15455 ( .A(n12101), .B(n12100), .ZN(n12103) );
  AOI21_X1 U15456 ( .B1(n12103), .B2(n12174), .A(n12102), .ZN(n12104) );
  AND2_X1 U15457 ( .A1(n12105), .A2(n12104), .ZN(n14669) );
  INV_X1 U15458 ( .A(n12106), .ZN(n12113) );
  OR2_X1 U15459 ( .A1(n11957), .A2(n12107), .ZN(n12110) );
  INV_X1 U15460 ( .A(n12108), .ZN(n12109) );
  NAND2_X1 U15461 ( .A1(n12110), .A2(n12109), .ZN(n14028) );
  NOR2_X1 U15462 ( .A1(n12281), .A2(n14028), .ZN(n12112) );
  OAI21_X1 U15463 ( .B1(n14028), .B2(n14029), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12111) );
  AOI21_X1 U15464 ( .B1(n12113), .B2(n12112), .A(n12111), .ZN(n12116) );
  OR2_X1 U15465 ( .A1(n12114), .A2(n14028), .ZN(n12115) );
  NAND2_X1 U15466 ( .A1(n12116), .A2(n12115), .ZN(n14030) );
  INV_X1 U15467 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20767) );
  NAND2_X1 U15468 ( .A1(n14669), .A2(n12117), .ZN(n12119) );
  NAND2_X1 U15469 ( .A1(n14030), .A2(n20767), .ZN(n12118) );
  NAND2_X1 U15470 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  XNOR2_X1 U15471 ( .A(n12120), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14629) );
  INV_X1 U15472 ( .A(n12120), .ZN(n12121) );
  NAND2_X1 U15473 ( .A1(n12121), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12122) );
  INV_X1 U15474 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12123) );
  AND2_X1 U15475 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  NAND2_X1 U15476 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  NAND2_X1 U15477 ( .A1(n12129), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U15478 ( .A1(n12234), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12142) );
  AOI22_X1 U15479 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15480 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15481 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15482 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12131) );
  NAND4_X1 U15483 ( .A1(n12134), .A2(n12133), .A3(n12132), .A4(n12131), .ZN(
        n12140) );
  AOI22_X1 U15484 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15485 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15486 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15487 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U15488 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12139) );
  NAND2_X1 U15489 ( .A1(n12246), .A2(n12158), .ZN(n12141) );
  NAND2_X1 U15490 ( .A1(n12302), .A2(n12143), .ZN(n12319) );
  NAND3_X1 U15491 ( .A1(n12319), .A2(n14029), .A3(n12171), .ZN(n12149) );
  INV_X1 U15492 ( .A(n12161), .ZN(n12145) );
  NAND2_X1 U15493 ( .A1(n12145), .A2(n12159), .ZN(n12146) );
  XNOR2_X1 U15494 ( .A(n12146), .B(n12158), .ZN(n12147) );
  NAND2_X1 U15495 ( .A1(n12147), .A2(n12174), .ZN(n12148) );
  NAND2_X1 U15496 ( .A1(n12149), .A2(n12148), .ZN(n12153) );
  INV_X1 U15497 ( .A(n12153), .ZN(n12151) );
  INV_X1 U15498 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12150) );
  NAND2_X1 U15499 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  NAND2_X1 U15500 ( .A1(n12153), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12154) );
  INV_X1 U15501 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12156) );
  NAND2_X1 U15502 ( .A1(n12246), .A2(n12173), .ZN(n12155) );
  XNOR2_X1 U15503 ( .A(n12171), .B(n12157), .ZN(n12326) );
  NAND2_X1 U15504 ( .A1(n12326), .A2(n14029), .ZN(n12164) );
  NAND2_X1 U15505 ( .A1(n12159), .A2(n12158), .ZN(n12160) );
  OR2_X1 U15506 ( .A1(n12161), .A2(n12160), .ZN(n12172) );
  XNOR2_X1 U15507 ( .A(n12172), .B(n12173), .ZN(n12162) );
  NAND2_X1 U15508 ( .A1(n12162), .A2(n12174), .ZN(n12163) );
  NAND2_X1 U15509 ( .A1(n12164), .A2(n12163), .ZN(n12167) );
  INV_X1 U15510 ( .A(n12167), .ZN(n12166) );
  INV_X1 U15511 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U15512 ( .A1(n12166), .A2(n12165), .ZN(n17309) );
  NAND2_X1 U15513 ( .A1(n12167), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17308) );
  NOR2_X1 U15514 ( .A1(n13344), .A2(n12169), .ZN(n12170) );
  INV_X4 U15515 ( .A(n12190), .ZN(n15641) );
  INV_X1 U15516 ( .A(n12172), .ZN(n12175) );
  NAND3_X1 U15517 ( .A1(n12175), .A2(n12174), .A3(n12173), .ZN(n12176) );
  NAND2_X1 U15518 ( .A1(n15641), .A2(n12176), .ZN(n15689) );
  INV_X4 U15519 ( .A(n12190), .ZN(n15657) );
  INV_X1 U15520 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15592) );
  INV_X1 U15521 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15833) );
  XNOR2_X1 U15522 ( .A(n15641), .B(n15833), .ZN(n15644) );
  NAND2_X1 U15523 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12177) );
  AND2_X1 U15524 ( .A1(n15657), .A2(n12177), .ZN(n15635) );
  INV_X1 U15525 ( .A(n15635), .ZN(n12178) );
  INV_X1 U15526 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15852) );
  INV_X1 U15527 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15820) );
  NAND2_X1 U15528 ( .A1(n15657), .A2(n15820), .ZN(n15596) );
  AND2_X1 U15529 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15804) );
  NAND2_X1 U15530 ( .A1(n15804), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12179) );
  NAND2_X1 U15531 ( .A1(n15657), .A2(n12179), .ZN(n12180) );
  NAND2_X1 U15532 ( .A1(n15596), .A2(n12180), .ZN(n12181) );
  NOR2_X1 U15533 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12182) );
  OR2_X1 U15534 ( .A1(n15657), .A2(n12182), .ZN(n12183) );
  INV_X1 U15535 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U15536 ( .A1(n15657), .A2(n15793), .ZN(n12184) );
  NOR2_X1 U15537 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12185) );
  INV_X1 U15538 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15806) );
  NAND2_X1 U15539 ( .A1(n15613), .A2(n15617), .ZN(n15597) );
  INV_X1 U15540 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15666) );
  INV_X1 U15541 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15861) );
  NAND2_X1 U15542 ( .A1(n15666), .A2(n15861), .ZN(n15636) );
  NOR2_X1 U15543 ( .A1(n15636), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12186) );
  NOR2_X1 U15544 ( .A1(n15641), .A2(n12186), .ZN(n15593) );
  NOR2_X1 U15545 ( .A1(n15597), .A2(n15593), .ZN(n12187) );
  XNOR2_X1 U15546 ( .A(n15641), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15584) );
  AND2_X1 U15547 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U15548 ( .A1(n15758), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15743) );
  NOR2_X1 U15549 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12189) );
  INV_X1 U15550 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15752) );
  NAND2_X1 U15551 ( .A1(n15556), .A2(n15752), .ZN(n12191) );
  INV_X1 U15552 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14824) );
  INV_X1 U15553 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13508) );
  INV_X1 U15554 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13335) );
  NAND2_X1 U15555 ( .A1(n21302), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12194) );
  NAND2_X1 U15556 ( .A1(n11997), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12193) );
  NAND2_X1 U15557 ( .A1(n12194), .A2(n12193), .ZN(n12207) );
  NAND2_X1 U15558 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21677), .ZN(
        n12206) );
  NAND2_X1 U15559 ( .A1(n21066), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U15560 ( .A1(n13852), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12196) );
  NAND2_X1 U15561 ( .A1(n12199), .A2(n12196), .ZN(n12217) );
  INV_X1 U15562 ( .A(n12217), .ZN(n12197) );
  NAND2_X1 U15563 ( .A1(n12198), .A2(n12197), .ZN(n12219) );
  NAND2_X1 U15564 ( .A1(n12219), .A2(n12199), .ZN(n12231) );
  XNOR2_X1 U15565 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12230) );
  AOI222_X1 U15566 ( .A1(n12228), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12228), .B2(n12312), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n12312), .ZN(n13352) );
  NAND2_X1 U15567 ( .A1(n13352), .A2(n12240), .ZN(n12245) );
  NAND2_X1 U15568 ( .A1(n12200), .A2(n13823), .ZN(n12225) );
  INV_X1 U15569 ( .A(n12206), .ZN(n12201) );
  AOI21_X1 U15570 ( .B1(n9866), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12201), .ZN(n12202) );
  OAI211_X1 U15571 ( .C1(n14727), .C2(n13487), .A(n12225), .B(n12202), .ZN(
        n12205) );
  INV_X1 U15572 ( .A(n12240), .ZN(n12242) );
  NAND2_X1 U15573 ( .A1(n12246), .A2(n12202), .ZN(n12203) );
  NAND2_X1 U15574 ( .A1(n12242), .A2(n12203), .ZN(n12204) );
  XNOR2_X1 U15575 ( .A(n12207), .B(n12206), .ZN(n13349) );
  INV_X1 U15576 ( .A(n13349), .ZN(n12211) );
  NAND2_X1 U15577 ( .A1(n12246), .A2(n20792), .ZN(n12208) );
  NAND2_X1 U15578 ( .A1(n14143), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12209) );
  OAI211_X1 U15579 ( .C1(n12222), .C2(n12211), .A(n12208), .B(n12209), .ZN(
        n12213) );
  NAND2_X1 U15580 ( .A1(n12209), .A2(n20792), .ZN(n12210) );
  NOR2_X1 U15581 ( .A1(n12210), .A2(n12246), .ZN(n12212) );
  OAI22_X1 U15582 ( .A1(n12214), .A2(n12213), .B1(n12212), .B2(n12211), .ZN(
        n12216) );
  NAND2_X1 U15583 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  NAND2_X1 U15584 ( .A1(n12216), .A2(n12215), .ZN(n12224) );
  NAND2_X1 U15585 ( .A1(n12218), .A2(n12217), .ZN(n12220) );
  NAND2_X1 U15586 ( .A1(n12220), .A2(n12219), .ZN(n13350) );
  NAND2_X1 U15587 ( .A1(n12246), .A2(n12226), .ZN(n12221) );
  OAI211_X1 U15588 ( .C1(n12226), .C2(n12222), .A(n12225), .B(n12221), .ZN(
        n12223) );
  NAND2_X1 U15589 ( .A1(n12224), .A2(n12223), .ZN(n12238) );
  INV_X1 U15590 ( .A(n12225), .ZN(n12227) );
  NAND3_X1 U15591 ( .A1(n12227), .A2(n12226), .A3(n12246), .ZN(n12237) );
  AND2_X1 U15592 ( .A1(n12312), .A2(n12228), .ZN(n12229) );
  NAND2_X1 U15593 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12229), .ZN(
        n13351) );
  NOR2_X1 U15594 ( .A1(n12231), .A2(n12230), .ZN(n12232) );
  OR2_X1 U15595 ( .A1(n12233), .A2(n12232), .ZN(n13348) );
  INV_X1 U15596 ( .A(n13348), .ZN(n12235) );
  AOI21_X1 U15597 ( .B1(n13351), .B2(n12235), .A(n12234), .ZN(n12236) );
  AOI21_X1 U15598 ( .B1(n12238), .B2(n12237), .A(n12236), .ZN(n12244) );
  NOR2_X1 U15599 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12312), .ZN(n12239) );
  AOI21_X1 U15600 ( .B1(n12240), .B2(n13348), .A(n12239), .ZN(n12241) );
  OAI21_X1 U15601 ( .B1(n13351), .B2(n12242), .A(n12241), .ZN(n12243) );
  NAND2_X1 U15602 ( .A1(n13352), .A2(n12246), .ZN(n12247) );
  INV_X1 U15603 ( .A(n13359), .ZN(n14038) );
  NAND2_X1 U15604 ( .A1(n12249), .A2(n20800), .ZN(n12250) );
  NAND2_X1 U15605 ( .A1(n11945), .A2(n14727), .ZN(n12251) );
  NAND2_X1 U15606 ( .A1(n21304), .A2(n12264), .ZN(n21486) );
  NAND2_X1 U15607 ( .A1(n21486), .A2(n21369), .ZN(n12252) );
  NAND2_X1 U15608 ( .A1(n21369), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17287) );
  NAND2_X1 U15609 ( .A1(n20830), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12253) );
  AND2_X1 U15610 ( .A1(n17287), .A2(n12253), .ZN(n14034) );
  NAND2_X1 U15611 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12294) );
  INV_X1 U15612 ( .A(n12294), .ZN(n12254) );
  NAND2_X1 U15613 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12254), .ZN(
        n12314) );
  NAND2_X1 U15614 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12255) );
  NOR2_X2 U15615 ( .A1(n12314), .A2(n12255), .ZN(n12321) );
  NAND2_X1 U15616 ( .A1(n12321), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12327) );
  NAND2_X1 U15617 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12256) );
  OR2_X2 U15618 ( .A1(n12375), .A2(n12256), .ZN(n12391) );
  NOR2_X2 U15619 ( .A1(n12391), .A2(n12390), .ZN(n12333) );
  NAND2_X1 U15620 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12257) );
  OR2_X2 U15621 ( .A1(n12422), .A2(n12257), .ZN(n12430) );
  INV_X1 U15622 ( .A(n12446), .ZN(n12259) );
  OR2_X2 U15623 ( .A1(n12463), .A2(n15239), .ZN(n12480) );
  OR2_X2 U15624 ( .A1(n12530), .A2(n12529), .ZN(n12547) );
  INV_X1 U15625 ( .A(n12547), .ZN(n12262) );
  INV_X1 U15626 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12613) );
  OR2_X2 U15627 ( .A1(n12580), .A2(n12613), .ZN(n13596) );
  XNOR2_X1 U15628 ( .A(n13596), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15127) );
  NAND2_X1 U15629 ( .A1(n20718), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15732) );
  OAI21_X1 U15630 ( .B1(n15577), .B2(n13595), .A(n15732), .ZN(n12265) );
  NAND2_X1 U15631 ( .A1(n15905), .A2(n12455), .ZN(n12271) );
  NAND2_X1 U15632 ( .A1(n12297), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12269) );
  NOR2_X2 U15633 ( .A1(n20818), .A2(n21306), .ZN(n12320) );
  INV_X1 U15634 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14627) );
  XNOR2_X1 U15635 ( .A(n14627), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20624) );
  OAI21_X1 U15636 ( .B1(n20624), .B2(n14796), .A(n12492), .ZN(n12267) );
  AOI21_X1 U15637 ( .B1(n12320), .B2(P1_EAX_REG_2__SCAN_IN), .A(n12267), .ZN(
        n12268) );
  AND2_X1 U15638 ( .A1(n12269), .A2(n12268), .ZN(n12270) );
  NAND2_X1 U15639 ( .A1(n12271), .A2(n12270), .ZN(n12272) );
  NAND2_X1 U15640 ( .A1(n14803), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12292) );
  NAND2_X1 U15641 ( .A1(n12272), .A2(n12292), .ZN(n14169) );
  INV_X1 U15642 ( .A(n14169), .ZN(n12291) );
  NAND2_X1 U15643 ( .A1(n20971), .A2(n12455), .ZN(n12280) );
  AOI22_X1 U15644 ( .A1(n12320), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21306), .ZN(n12278) );
  NAND2_X1 U15645 ( .A1(n12297), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12277) );
  AND2_X1 U15646 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NAND2_X1 U15647 ( .A1(n12280), .A2(n12279), .ZN(n14061) );
  NAND2_X1 U15648 ( .A1(n20855), .A2(n12282), .ZN(n12283) );
  NAND2_X1 U15649 ( .A1(n12283), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13879) );
  INV_X1 U15650 ( .A(n12297), .ZN(n12313) );
  NAND2_X1 U15651 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U15652 ( .A1(n12320), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12285) );
  OAI211_X1 U15653 ( .C1(n12313), .C2(n9866), .A(n12286), .B(n12285), .ZN(
        n12287) );
  AOI21_X1 U15654 ( .B1(n20893), .B2(n12455), .A(n12287), .ZN(n12288) );
  OR2_X1 U15655 ( .A1(n13879), .A2(n12288), .ZN(n13880) );
  INV_X1 U15656 ( .A(n12288), .ZN(n13881) );
  OR2_X1 U15657 ( .A1(n13881), .A2(n14796), .ZN(n12289) );
  NAND2_X1 U15658 ( .A1(n13880), .A2(n12289), .ZN(n14060) );
  NAND2_X1 U15659 ( .A1(n14061), .A2(n14060), .ZN(n14168) );
  NAND2_X1 U15660 ( .A1(n12291), .A2(n12290), .ZN(n14166) );
  INV_X1 U15661 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U15662 ( .A1(n14577), .A2(n12294), .ZN(n12295) );
  AND2_X1 U15663 ( .A1(n12295), .A2(n12314), .ZN(n20607) );
  OAI22_X1 U15664 ( .A1(n20607), .A2(n14796), .B1(n14577), .B2(n12492), .ZN(
        n12296) );
  AOI21_X1 U15665 ( .B1(n12320), .B2(P1_EAX_REG_3__SCAN_IN), .A(n12296), .ZN(
        n12299) );
  NAND2_X1 U15666 ( .A1(n12297), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12298) );
  OAI211_X1 U15667 ( .C1(n21463), .C2(n12426), .A(n12299), .B(n12298), .ZN(
        n14439) );
  AND2_X1 U15668 ( .A1(n12300), .A2(n12455), .ZN(n12301) );
  NAND2_X1 U15669 ( .A1(n12302), .A2(n12301), .ZN(n12308) );
  INV_X1 U15670 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20589) );
  INV_X1 U15671 ( .A(n12314), .ZN(n12303) );
  AOI21_X1 U15672 ( .B1(n12303), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12304) );
  OR2_X1 U15673 ( .A1(n12304), .A2(n12321), .ZN(n20587) );
  NAND2_X1 U15674 ( .A1(n20587), .A2(n14802), .ZN(n12305) );
  OAI21_X1 U15675 ( .B1(n12492), .B2(n20589), .A(n12305), .ZN(n12306) );
  AOI21_X1 U15676 ( .B1(n12320), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12306), .ZN(
        n12307) );
  NAND2_X1 U15677 ( .A1(n12308), .A2(n12307), .ZN(n15492) );
  INV_X1 U15678 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15679 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12311) );
  NAND2_X1 U15680 ( .A1(n12320), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12310) );
  OAI211_X1 U15681 ( .C1(n12313), .C2(n12312), .A(n12311), .B(n12310), .ZN(
        n12317) );
  INV_X1 U15682 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12315) );
  XNOR2_X1 U15683 ( .A(n12315), .B(n12314), .ZN(n20713) );
  AND2_X1 U15684 ( .A1(n20713), .A2(n14802), .ZN(n12316) );
  AOI21_X1 U15685 ( .B1(n12317), .B2(n14796), .A(n12316), .ZN(n12318) );
  INV_X1 U15686 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n15488) );
  OR2_X1 U15687 ( .A1(n12321), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12322) );
  NAND2_X1 U15688 ( .A1(n12327), .A2(n12322), .ZN(n20580) );
  AOI22_X1 U15689 ( .A1(n20580), .A2(n14802), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n14803), .ZN(n12323) );
  OAI21_X1 U15690 ( .B1(n14797), .B2(n15488), .A(n12323), .ZN(n12324) );
  AOI21_X1 U15691 ( .B1(n12319), .B2(n12455), .A(n12324), .ZN(n15400) );
  INV_X1 U15692 ( .A(n15400), .ZN(n12325) );
  INV_X1 U15693 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U15694 ( .A1(n12327), .A2(n12329), .ZN(n12328) );
  NAND2_X1 U15695 ( .A1(n12375), .A2(n12328), .ZN(n20565) );
  NOR2_X1 U15696 ( .A1(n12492), .A2(n12329), .ZN(n12330) );
  AOI21_X1 U15697 ( .B1(n20565), .B2(n14802), .A(n12330), .ZN(n12331) );
  OAI21_X1 U15698 ( .B1(n14797), .B2(n14260), .A(n12331), .ZN(n12332) );
  INV_X1 U15699 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U15700 ( .A1(n12320), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12337) );
  INV_X1 U15701 ( .A(n12333), .ZN(n12334) );
  NAND2_X1 U15702 ( .A1(n12334), .A2(n12338), .ZN(n12335) );
  NAND2_X1 U15703 ( .A1(n12422), .A2(n12335), .ZN(n15662) );
  NAND2_X1 U15704 ( .A1(n15662), .A2(n14802), .ZN(n12336) );
  OAI211_X1 U15705 ( .C1(n12492), .C2(n12338), .A(n12337), .B(n12336), .ZN(
        n15282) );
  AOI22_X1 U15706 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15707 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13615), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15708 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15709 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12339) );
  NAND4_X1 U15710 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12348) );
  AOI22_X1 U15711 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15712 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15713 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15714 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12343) );
  NAND4_X1 U15715 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12347) );
  OR2_X1 U15716 ( .A1(n12348), .A2(n12347), .ZN(n12349) );
  AND2_X1 U15717 ( .A1(n12455), .A2(n12349), .ZN(n15281) );
  OR2_X1 U15718 ( .A1(n15282), .A2(n15281), .ZN(n12396) );
  AOI22_X1 U15719 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12548), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15720 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13615), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15721 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15722 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12350) );
  NAND4_X1 U15723 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12359) );
  AOI22_X1 U15724 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15725 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15726 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15727 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n14774), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12354) );
  NAND4_X1 U15728 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12358) );
  OAI21_X1 U15729 ( .B1(n12359), .B2(n12358), .A(n12455), .ZN(n12364) );
  NAND2_X1 U15730 ( .A1(n12320), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12363) );
  INV_X1 U15731 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12360) );
  XNOR2_X1 U15732 ( .A(n12375), .B(n12360), .ZN(n15691) );
  NAND2_X1 U15733 ( .A1(n15691), .A2(n14802), .ZN(n12362) );
  NAND2_X1 U15734 ( .A1(n14803), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12361) );
  NAND4_X1 U15735 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n15343) );
  AOI22_X1 U15736 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15737 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15738 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15739 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12365) );
  NAND4_X1 U15740 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12374) );
  AOI22_X1 U15741 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15742 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15743 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15744 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15745 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  NOR2_X1 U15746 ( .A1(n12374), .A2(n12373), .ZN(n12379) );
  INV_X1 U15747 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21679) );
  OAI21_X1 U15748 ( .B1(n12375), .B2(n12360), .A(n21679), .ZN(n12376) );
  NAND2_X1 U15749 ( .A1(n12376), .A2(n12391), .ZN(n20557) );
  AOI22_X1 U15750 ( .A1(n20557), .A2(n14802), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n14803), .ZN(n12378) );
  NAND2_X1 U15751 ( .A1(n12320), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12377) );
  OAI211_X1 U15752 ( .C1(n12426), .C2(n12379), .A(n12378), .B(n12377), .ZN(
        n15479) );
  AOI22_X1 U15753 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15754 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15755 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15756 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15757 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12389) );
  AOI22_X1 U15758 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15759 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15760 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15761 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12384) );
  NAND4_X1 U15762 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12388) );
  OAI21_X1 U15763 ( .B1(n12389), .B2(n12388), .A(n12455), .ZN(n12395) );
  NAND2_X1 U15764 ( .A1(n12320), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12394) );
  XNOR2_X1 U15765 ( .A(n12391), .B(n12390), .ZN(n15673) );
  NAND2_X1 U15766 ( .A1(n15673), .A2(n14802), .ZN(n12393) );
  NAND2_X1 U15767 ( .A1(n14803), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12392) );
  NAND4_X1 U15768 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n15330) );
  AND4_X1 U15769 ( .A1(n12396), .A2(n15343), .A3(n15479), .A4(n15330), .ZN(
        n12428) );
  AOI22_X1 U15770 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15771 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13615), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15772 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15773 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12397) );
  NAND4_X1 U15774 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12406) );
  AOI22_X1 U15775 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15776 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15777 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15778 ( .A1(n14775), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12401) );
  NAND4_X1 U15779 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n12401), .ZN(
        n12405) );
  NOR2_X1 U15780 ( .A1(n12406), .A2(n12405), .ZN(n12411) );
  INV_X1 U15781 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15307) );
  OR2_X1 U15782 ( .A1(n12422), .A2(n15307), .ZN(n12408) );
  INV_X1 U15783 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12407) );
  XNOR2_X1 U15784 ( .A(n12408), .B(n12407), .ZN(n15633) );
  NAND2_X1 U15785 ( .A1(n15633), .A2(n14802), .ZN(n12410) );
  AOI22_X1 U15786 ( .A1(n12320), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n14803), .ZN(n12409) );
  OAI211_X1 U15787 ( .C1(n12411), .C2(n12426), .A(n12410), .B(n12409), .ZN(
        n15286) );
  AOI22_X1 U15788 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15789 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15790 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15791 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15792 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12421) );
  AOI22_X1 U15793 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15794 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15795 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15796 ( .A1(n14775), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12416) );
  NAND4_X1 U15797 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n12416), .ZN(
        n12420) );
  NOR2_X1 U15798 ( .A1(n12421), .A2(n12420), .ZN(n12427) );
  XNOR2_X1 U15799 ( .A(n12422), .B(n15307), .ZN(n15653) );
  NAND2_X1 U15800 ( .A1(n15653), .A2(n14802), .ZN(n12425) );
  NOR2_X1 U15801 ( .A1(n12492), .A2(n15307), .ZN(n12423) );
  AOI21_X1 U15802 ( .B1(n12320), .B2(P1_EAX_REG_12__SCAN_IN), .A(n12423), .ZN(
        n12424) );
  OAI211_X1 U15803 ( .C1(n12427), .C2(n12426), .A(n12425), .B(n12424), .ZN(
        n15284) );
  AND3_X1 U15804 ( .A1(n12428), .A2(n15286), .A3(n15284), .ZN(n12429) );
  INV_X1 U15805 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15271) );
  XNOR2_X1 U15806 ( .A(n12430), .B(n15271), .ZN(n15629) );
  NAND2_X1 U15807 ( .A1(n15629), .A2(n14802), .ZN(n12445) );
  AOI22_X1 U15808 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15809 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15810 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15811 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12431) );
  NAND4_X1 U15812 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12440) );
  AOI22_X1 U15813 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15814 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15815 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15816 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15817 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  OAI21_X1 U15818 ( .B1(n12440), .B2(n12439), .A(n12455), .ZN(n12443) );
  NAND2_X1 U15819 ( .A1(n12320), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U15820 ( .A1(n14803), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12441) );
  AND3_X1 U15821 ( .A1(n12443), .A2(n12442), .A3(n12441), .ZN(n12444) );
  NAND2_X1 U15822 ( .A1(n12445), .A2(n12444), .ZN(n15265) );
  NAND2_X1 U15823 ( .A1(n15264), .A2(n15265), .ZN(n15250) );
  INV_X1 U15824 ( .A(n15250), .ZN(n12462) );
  INV_X1 U15825 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15258) );
  XNOR2_X1 U15826 ( .A(n12446), .B(n15258), .ZN(n15621) );
  INV_X1 U15827 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20661) );
  AOI22_X1 U15828 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15829 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15830 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15831 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12447) );
  NAND4_X1 U15832 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12457) );
  AOI22_X1 U15833 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15834 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15835 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15836 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12451) );
  NAND4_X1 U15837 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12456) );
  OAI21_X1 U15838 ( .B1(n12457), .B2(n12456), .A(n12455), .ZN(n12459) );
  NAND2_X1 U15839 ( .A1(n14803), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12458) );
  OAI211_X1 U15840 ( .C1(n14797), .C2(n20661), .A(n12459), .B(n12458), .ZN(
        n12460) );
  AOI21_X1 U15841 ( .B1(n15621), .B2(n14802), .A(n12460), .ZN(n15251) );
  NAND2_X1 U15842 ( .A1(n12463), .A2(n15239), .ZN(n12464) );
  NAND2_X1 U15843 ( .A1(n12480), .A2(n12464), .ZN(n15608) );
  AOI22_X1 U15844 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11817), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15845 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15846 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15847 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13633), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12465) );
  NAND4_X1 U15848 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(
        n12474) );
  AOI22_X1 U15849 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n13632), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15850 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15851 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n14784), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15852 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12469) );
  NAND4_X1 U15853 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12469), .ZN(
        n12473) );
  NOR2_X1 U15854 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  NOR2_X1 U15855 ( .A1(n13666), .A2(n12475), .ZN(n12478) );
  INV_X1 U15856 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U15857 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12476) );
  OAI211_X1 U15858 ( .C1(n14797), .C2(n15459), .A(n14796), .B(n12476), .ZN(
        n12477) );
  OAI22_X1 U15859 ( .A1(n15608), .A2(n14796), .B1(n12478), .B2(n12477), .ZN(
        n15227) );
  INV_X1 U15860 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21646) );
  NAND2_X1 U15861 ( .A1(n12480), .A2(n21646), .ZN(n12481) );
  NAND2_X1 U15862 ( .A1(n12497), .A2(n12481), .ZN(n15602) );
  AOI22_X1 U15863 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15864 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15865 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15866 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12482) );
  NAND4_X1 U15867 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n12491) );
  AOI22_X1 U15868 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15869 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15870 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15871 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U15872 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n12490) );
  NOR2_X1 U15873 ( .A1(n12491), .A2(n12490), .ZN(n12495) );
  NOR2_X1 U15874 ( .A1(n12492), .A2(n21646), .ZN(n12493) );
  AOI21_X1 U15875 ( .B1(n12320), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12493), .ZN(
        n12494) );
  OAI21_X1 U15876 ( .B1(n13666), .B2(n12495), .A(n12494), .ZN(n12496) );
  AOI21_X1 U15877 ( .B1(n15602), .B2(n14802), .A(n12496), .ZN(n15214) );
  NAND2_X1 U15878 ( .A1(n12497), .A2(n15204), .ZN(n12498) );
  AND2_X1 U15879 ( .A1(n12513), .A2(n12498), .ZN(n15585) );
  AOI22_X1 U15880 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15881 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15882 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15883 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15884 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12508) );
  AOI22_X1 U15885 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15886 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15887 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15888 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12503) );
  NAND4_X1 U15889 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12507) );
  OR2_X1 U15890 ( .A1(n12508), .A2(n12507), .ZN(n12511) );
  INV_X1 U15891 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U15892 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12509) );
  OAI211_X1 U15893 ( .C1(n14797), .C2(n15451), .A(n14796), .B(n12509), .ZN(
        n12510) );
  AOI21_X1 U15894 ( .B1(n14799), .B2(n12511), .A(n12510), .ZN(n12512) );
  AOI21_X1 U15895 ( .B1(n15585), .B2(n14802), .A(n12512), .ZN(n15202) );
  NAND2_X1 U15896 ( .A1(n15213), .A2(n15202), .ZN(n15181) );
  XNOR2_X1 U15897 ( .A(n12513), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15581) );
  NAND2_X1 U15898 ( .A1(n15581), .A2(n14802), .ZN(n12528) );
  AOI22_X1 U15899 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15900 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U15901 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15902 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12514) );
  NAND4_X1 U15903 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n12514), .ZN(
        n12523) );
  AOI22_X1 U15904 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U15905 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15906 ( .A1(n14775), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15907 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12518) );
  NAND4_X1 U15908 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        n12522) );
  NOR2_X1 U15909 ( .A1(n12523), .A2(n12522), .ZN(n12526) );
  INV_X1 U15910 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15576) );
  AOI21_X1 U15911 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15576), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12524) );
  AOI21_X1 U15912 ( .B1(n12320), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12524), .ZN(
        n12525) );
  OAI21_X1 U15913 ( .B1(n13666), .B2(n12526), .A(n12525), .ZN(n12527) );
  NAND2_X1 U15914 ( .A1(n12528), .A2(n12527), .ZN(n15182) );
  NAND2_X1 U15915 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  NAND2_X1 U15916 ( .A1(n12547), .A2(n12531), .ZN(n15570) );
  AOI22_X1 U15917 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12535) );
  AOI22_X1 U15918 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15919 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15920 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12532) );
  NAND4_X1 U15921 ( .A1(n12535), .A2(n12534), .A3(n12533), .A4(n12532), .ZN(
        n12541) );
  AOI22_X1 U15922 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15923 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15924 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15925 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12536) );
  NAND4_X1 U15926 ( .A1(n12539), .A2(n12538), .A3(n12537), .A4(n12536), .ZN(
        n12540) );
  NOR2_X1 U15927 ( .A1(n12541), .A2(n12540), .ZN(n12542) );
  NOR2_X1 U15928 ( .A1(n13666), .A2(n12542), .ZN(n12545) );
  INV_X1 U15929 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15443) );
  NAND2_X1 U15930 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12543) );
  OAI211_X1 U15931 ( .C1(n14797), .C2(n15443), .A(n14796), .B(n12543), .ZN(
        n12544) );
  OAI22_X1 U15932 ( .A1(n15570), .A2(n14796), .B1(n12545), .B2(n12544), .ZN(
        n15171) );
  XNOR2_X1 U15933 ( .A(n12547), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15564) );
  AOI22_X1 U15934 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15935 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15936 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15937 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12550) );
  NAND4_X1 U15938 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12559) );
  AOI22_X1 U15939 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15940 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15941 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15942 ( .A1(n11812), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12554) );
  NAND4_X1 U15943 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12558) );
  OR2_X1 U15944 ( .A1(n12559), .A2(n12558), .ZN(n12562) );
  INV_X1 U15945 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U15946 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12560) );
  OAI211_X1 U15947 ( .C1(n14797), .C2(n15439), .A(n14796), .B(n12560), .ZN(
        n12561) );
  AOI21_X1 U15948 ( .B1(n14799), .B2(n12562), .A(n12561), .ZN(n12563) );
  AOI21_X1 U15949 ( .B1(n15564), .B2(n14802), .A(n12563), .ZN(n15155) );
  NAND2_X1 U15950 ( .A1(n12564), .A2(n15549), .ZN(n12565) );
  AOI22_X1 U15951 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15952 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15953 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15954 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12566) );
  NAND4_X1 U15955 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12575) );
  AOI22_X1 U15956 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15957 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15958 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15959 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12570) );
  NAND4_X1 U15960 ( .A1(n12573), .A2(n12572), .A3(n12571), .A4(n12570), .ZN(
        n12574) );
  OR2_X1 U15961 ( .A1(n12575), .A2(n12574), .ZN(n12578) );
  INV_X1 U15962 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15435) );
  OAI21_X1 U15963 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20830), .A(
        n21306), .ZN(n12576) );
  OAI21_X1 U15964 ( .B1(n14797), .B2(n15435), .A(n12576), .ZN(n12577) );
  AOI21_X1 U15965 ( .B1(n14799), .B2(n12578), .A(n12577), .ZN(n12579) );
  NAND2_X1 U15966 ( .A1(n12580), .A2(n12613), .ZN(n12581) );
  NAND2_X1 U15967 ( .A1(n13596), .A2(n12581), .ZN(n14730) );
  OR2_X1 U15968 ( .A1(n14730), .A2(n14796), .ZN(n12618) );
  AOI22_X1 U15969 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15970 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13615), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15971 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15972 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12582) );
  NAND4_X1 U15973 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12591) );
  AOI22_X1 U15974 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15975 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15976 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15977 ( .A1(n14775), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U15978 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12590) );
  NOR2_X1 U15979 ( .A1(n12591), .A2(n12590), .ZN(n12620) );
  AOI22_X1 U15980 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15981 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13609), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15982 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15983 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15984 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12602) );
  AOI22_X1 U15985 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n14774), .B1(
        n13615), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15986 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15987 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15988 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12597) );
  NAND4_X1 U15989 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12601) );
  NOR2_X1 U15990 ( .A1(n12602), .A2(n12601), .ZN(n12621) );
  NOR2_X1 U15991 ( .A1(n12620), .A2(n12621), .ZN(n12631) );
  AOI22_X1 U15992 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15993 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15994 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15995 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12603) );
  NAND4_X1 U15996 ( .A1(n12606), .A2(n12605), .A3(n12604), .A4(n12603), .ZN(
        n12612) );
  AOI22_X1 U15997 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15998 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12609) );
  INV_X1 U15999 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21787) );
  AOI22_X1 U16000 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U16001 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12607) );
  NAND4_X1 U16002 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n12611) );
  OR2_X1 U16003 ( .A1(n12612), .A2(n12611), .ZN(n12630) );
  XNOR2_X1 U16004 ( .A(n12631), .B(n12630), .ZN(n12616) );
  AOI21_X1 U16005 ( .B1(n12613), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12614) );
  AOI21_X1 U16006 ( .B1(n12320), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12614), .ZN(
        n12615) );
  OAI21_X1 U16007 ( .B1(n12616), .B2(n13666), .A(n12615), .ZN(n12617) );
  NAND2_X1 U16008 ( .A1(n12618), .A2(n12617), .ZN(n14709) );
  XNOR2_X1 U16009 ( .A(n12619), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15140) );
  NAND2_X1 U16010 ( .A1(n15140), .A2(n14802), .ZN(n12628) );
  XOR2_X1 U16011 ( .A(n12621), .B(n12620), .Z(n12622) );
  NAND2_X1 U16012 ( .A1(n12622), .A2(n14799), .ZN(n12626) );
  NAND2_X1 U16013 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12623) );
  NAND2_X1 U16014 ( .A1(n14796), .A2(n12623), .ZN(n12624) );
  AOI21_X1 U16015 ( .B1(n12320), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12624), .ZN(
        n12625) );
  NAND2_X1 U16016 ( .A1(n12626), .A2(n12625), .ZN(n12627) );
  NAND2_X1 U16017 ( .A1(n12628), .A2(n12627), .ZN(n14833) );
  NOR2_X1 U16018 ( .A1(n14709), .A2(n14833), .ZN(n12647) );
  NAND2_X1 U16019 ( .A1(n12631), .A2(n12630), .ZN(n13607) );
  AOI22_X1 U16020 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U16021 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U16022 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U16023 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12632) );
  NAND4_X1 U16024 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12642) );
  AOI22_X1 U16025 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U16026 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U16027 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U16028 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12637) );
  NAND4_X1 U16029 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12641) );
  NOR2_X1 U16030 ( .A1(n12642), .A2(n12641), .ZN(n13608) );
  XOR2_X1 U16031 ( .A(n13607), .B(n13608), .Z(n12645) );
  INV_X1 U16032 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15427) );
  NAND2_X1 U16033 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12643) );
  OAI211_X1 U16034 ( .C1(n14797), .C2(n15427), .A(n14796), .B(n12643), .ZN(
        n12644) );
  AOI21_X1 U16035 ( .B1(n12645), .B2(n14799), .A(n12644), .ZN(n12646) );
  AOI21_X1 U16036 ( .B1(n15127), .B2(n14802), .A(n12646), .ZN(n12649) );
  AND2_X1 U16037 ( .A1(n12649), .A2(n12647), .ZN(n12648) );
  NAND2_X1 U16038 ( .A1(n15154), .A2(n13671), .ZN(n15108) );
  OAI21_X1 U16039 ( .B1(n14711), .B2(n12649), .A(n15108), .ZN(n15120) );
  AND2_X1 U16040 ( .A1(n21369), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14725) );
  NAND2_X1 U16041 ( .A1(n14725), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n17364) );
  OAI211_X1 U16042 ( .C1(n15738), .C2(n20537), .A(n12650), .B(n10385), .ZN(
        P1_U2974) );
  INV_X1 U16043 ( .A(n12656), .ZN(n16572) );
  XNOR2_X1 U16044 ( .A(n12658), .B(n10411), .ZN(n14940) );
  AOI21_X1 U16045 ( .B1(n12659), .B2(n16040), .A(n16431), .ZN(n16027) );
  INV_X1 U16046 ( .A(n12662), .ZN(n12660) );
  OAI21_X1 U16047 ( .B1(n16872), .B2(n12660), .A(n16811), .ZN(n16777) );
  NOR2_X1 U16048 ( .A1(n11468), .A2(n20442), .ZN(n14935) );
  INV_X1 U16049 ( .A(n14935), .ZN(n12663) );
  AND2_X1 U16050 ( .A1(n16772), .A2(n12664), .ZN(n12661) );
  NAND2_X1 U16051 ( .A1(n12662), .A2(n12661), .ZN(n16759) );
  OAI211_X1 U16052 ( .C1(n16777), .C2(n12664), .A(n12663), .B(n16759), .ZN(
        n12669) );
  INV_X1 U16053 ( .A(n12666), .ZN(n14761) );
  OR2_X1 U16054 ( .A1(n14761), .A2(n13320), .ZN(n13318) );
  AND2_X1 U16055 ( .A1(n12666), .A2(n12665), .ZN(n16335) );
  AOI21_X1 U16056 ( .B1(n12667), .B2(n13318), .A(n16335), .ZN(n16038) );
  INV_X1 U16057 ( .A(n16038), .ZN(n16346) );
  NOR2_X1 U16058 ( .A1(n16346), .A2(n19803), .ZN(n12668) );
  AOI211_X1 U16059 ( .C1(n16027), .C2(n19792), .A(n12669), .B(n12668), .ZN(
        n12670) );
  INV_X1 U16060 ( .A(n12670), .ZN(n12671) );
  OAI21_X1 U16061 ( .B1(n14940), .B2(n17400), .A(n12672), .ZN(P2_U3027) );
  NAND2_X1 U16062 ( .A1(n14523), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12674) );
  OAI21_X1 U16063 ( .B1(n19920), .B2(n20497), .A(n21570), .ZN(n12675) );
  NAND2_X1 U16064 ( .A1(n20184), .A2(n20288), .ZN(n20328) );
  AND3_X1 U16065 ( .A1(n12675), .A2(n20328), .A3(n20484), .ZN(n20218) );
  AOI21_X1 U16066 ( .B1(n12688), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20218), .ZN(n12676) );
  INV_X1 U16067 ( .A(n12697), .ZN(n12677) );
  NAND2_X1 U16068 ( .A1(n12677), .A2(n12678), .ZN(n12680) );
  INV_X1 U16069 ( .A(n12678), .ZN(n12679) );
  NAND2_X1 U16070 ( .A1(n12697), .A2(n12679), .ZN(n14157) );
  NAND2_X1 U16071 ( .A1(n12681), .A2(n12691), .ZN(n12683) );
  XNOR2_X1 U16072 ( .A(n19920), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19958) );
  AOI22_X1 U16073 ( .A1(n12688), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20484), .B2(n19958), .ZN(n12682) );
  NAND2_X1 U16074 ( .A1(n12683), .A2(n12682), .ZN(n12685) );
  AOI22_X1 U16075 ( .A1(n12688), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20484), .B2(n19889), .ZN(n12686) );
  NAND2_X1 U16076 ( .A1(n12688), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12689) );
  NAND2_X1 U16077 ( .A1(n20252), .A2(n19889), .ZN(n20219) );
  NAND3_X1 U16078 ( .A1(n20484), .A2(n20219), .A3(n19920), .ZN(n20290) );
  NAND2_X1 U16079 ( .A1(n12689), .A2(n20290), .ZN(n12690) );
  NAND2_X1 U16080 ( .A1(n13791), .A2(n13790), .ZN(n12694) );
  INV_X1 U16081 ( .A(n13814), .ZN(n16998) );
  NAND2_X1 U16082 ( .A1(n16998), .A2(n12692), .ZN(n12693) );
  NAND2_X1 U16083 ( .A1(n14523), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12696) );
  NAND2_X1 U16084 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12698) );
  NAND2_X1 U16085 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U16086 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12699) );
  NOR2_X1 U16087 ( .A1(n14314), .A2(n12699), .ZN(n12700) );
  NAND3_X1 U16088 ( .A1(n14541), .A2(n12700), .A3(n14542), .ZN(n12701) );
  NOR2_X1 U16089 ( .A1(n14153), .A2(n12701), .ZN(n12702) );
  INV_X1 U16090 ( .A(n12703), .ZN(n14640) );
  AND2_X1 U16091 ( .A1(n14554), .A2(n14307), .ZN(n12704) );
  INV_X1 U16092 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12705) );
  OAI22_X1 U16093 ( .A1(n12832), .A2(n12706), .B1(n12808), .B2(n12705), .ZN(
        n12707) );
  INV_X1 U16094 ( .A(n12707), .ZN(n12715) );
  AOI22_X1 U16095 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U16096 ( .A1(n10840), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12713) );
  INV_X1 U16097 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U16098 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12709) );
  NAND2_X1 U16099 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12708) );
  OAI211_X1 U16100 ( .C1(n10559), .C2(n12710), .A(n12709), .B(n12708), .ZN(
        n12711) );
  INV_X1 U16101 ( .A(n12711), .ZN(n12712) );
  NAND4_X1 U16102 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12712), .ZN(
        n12721) );
  AOI22_X1 U16103 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U16104 ( .A1(n11209), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U16105 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12828), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U16106 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12716) );
  NAND4_X1 U16107 ( .A1(n12719), .A2(n12718), .A3(n12717), .A4(n12716), .ZN(
        n12720) );
  OR2_X1 U16108 ( .A1(n12721), .A2(n12720), .ZN(n14661) );
  INV_X1 U16109 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12722) );
  OAI22_X1 U16110 ( .A1(n12722), .A2(n12832), .B1(n12808), .B2(n20350), .ZN(
        n12723) );
  INV_X1 U16111 ( .A(n12723), .ZN(n12732) );
  AOI22_X1 U16112 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U16113 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12724), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12730) );
  INV_X1 U16114 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U16115 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12726) );
  NAND2_X1 U16116 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12725) );
  OAI211_X1 U16117 ( .C1(n10559), .C2(n12727), .A(n12726), .B(n12725), .ZN(
        n12728) );
  INV_X1 U16118 ( .A(n12728), .ZN(n12729) );
  NAND4_X1 U16119 ( .A1(n12732), .A2(n12731), .A3(n12730), .A4(n12729), .ZN(
        n12738) );
  AOI22_X1 U16120 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U16121 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U16122 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U16123 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12733) );
  NAND4_X1 U16124 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12737) );
  OR2_X1 U16125 ( .A1(n12738), .A2(n12737), .ZN(n16347) );
  INV_X1 U16126 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12740) );
  INV_X1 U16127 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12739) );
  OAI22_X1 U16128 ( .A1(n12740), .A2(n12832), .B1(n12808), .B2(n12739), .ZN(
        n12741) );
  INV_X1 U16129 ( .A(n12741), .ZN(n12749) );
  AOI22_X1 U16130 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U16131 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12747) );
  INV_X1 U16132 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U16133 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12743) );
  NAND2_X1 U16134 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12742) );
  OAI211_X1 U16135 ( .C1(n10559), .C2(n12744), .A(n12743), .B(n12742), .ZN(
        n12745) );
  INV_X1 U16136 ( .A(n12745), .ZN(n12746) );
  NAND4_X1 U16137 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12755) );
  AOI22_X1 U16138 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U16139 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U16140 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U16141 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12750) );
  NAND4_X1 U16142 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12754) );
  OR2_X1 U16143 ( .A1(n12755), .A2(n12754), .ZN(n16349) );
  NAND4_X1 U16144 ( .A1(n14622), .A2(n14661), .A3(n16347), .A4(n16349), .ZN(
        n12756) );
  NOR2_X2 U16145 ( .A1(n14619), .A2(n12756), .ZN(n16343) );
  INV_X1 U16146 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12757) );
  OAI22_X1 U16147 ( .A1(n12757), .A2(n12832), .B1(n12808), .B2(n20363), .ZN(
        n12758) );
  INV_X1 U16148 ( .A(n12758), .ZN(n12766) );
  AOI22_X1 U16149 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U16150 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12764) );
  INV_X1 U16151 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U16152 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12760) );
  NAND2_X1 U16153 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12759) );
  OAI211_X1 U16154 ( .C1(n10559), .C2(n12761), .A(n12760), .B(n12759), .ZN(
        n12762) );
  INV_X1 U16155 ( .A(n12762), .ZN(n12763) );
  NAND4_X1 U16156 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12772) );
  AOI22_X1 U16157 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16158 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16159 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U16160 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12767) );
  NAND4_X1 U16161 ( .A1(n12770), .A2(n12769), .A3(n12768), .A4(n12767), .ZN(
        n12771) );
  OR2_X1 U16162 ( .A1(n12772), .A2(n12771), .ZN(n16342) );
  INV_X1 U16163 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12774) );
  INV_X1 U16164 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12773) );
  OAI22_X1 U16165 ( .A1(n12774), .A2(n12832), .B1(n12808), .B2(n12773), .ZN(
        n12775) );
  INV_X1 U16166 ( .A(n12775), .ZN(n12783) );
  AOI22_X1 U16167 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U16168 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12781) );
  INV_X1 U16169 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12778) );
  NAND2_X1 U16170 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12777) );
  NAND2_X1 U16171 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12776) );
  OAI211_X1 U16172 ( .C1(n10559), .C2(n12778), .A(n12777), .B(n12776), .ZN(
        n12779) );
  INV_X1 U16173 ( .A(n12779), .ZN(n12780) );
  NAND4_X1 U16174 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        n12789) );
  AOI22_X1 U16175 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16176 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U16177 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U16178 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12784) );
  NAND4_X1 U16179 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12788) );
  INV_X1 U16180 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12791) );
  OAI22_X1 U16181 ( .A1(n12791), .A2(n12832), .B1(n12808), .B2(n12790), .ZN(
        n12792) );
  INV_X1 U16182 ( .A(n12792), .ZN(n12800) );
  AOI22_X1 U16183 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16184 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12724), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12798) );
  INV_X1 U16185 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12795) );
  NAND2_X1 U16186 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12794) );
  NAND2_X1 U16187 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12793) );
  OAI211_X1 U16188 ( .C1(n10559), .C2(n12795), .A(n12794), .B(n12793), .ZN(
        n12796) );
  INV_X1 U16189 ( .A(n12796), .ZN(n12797) );
  NAND4_X1 U16190 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12806) );
  AOI22_X1 U16191 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U16192 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16193 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12802) );
  NAND2_X1 U16194 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12801) );
  NAND4_X1 U16195 ( .A1(n12804), .A2(n12803), .A3(n12802), .A4(n12801), .ZN(
        n12805) );
  NOR2_X1 U16196 ( .A1(n12806), .A2(n12805), .ZN(n16326) );
  INV_X1 U16197 ( .A(n16326), .ZN(n12825) );
  INV_X1 U16198 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12809) );
  OAI22_X1 U16199 ( .A1(n12809), .A2(n12832), .B1(n12808), .B2(n12807), .ZN(
        n12810) );
  INV_X1 U16200 ( .A(n12810), .ZN(n12818) );
  AOI22_X1 U16201 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16202 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12816) );
  INV_X1 U16203 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U16204 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12812) );
  NAND2_X1 U16205 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12811) );
  OAI211_X1 U16206 ( .C1(n10559), .C2(n12813), .A(n12812), .B(n12811), .ZN(
        n12814) );
  INV_X1 U16207 ( .A(n12814), .ZN(n12815) );
  NAND4_X1 U16208 ( .A1(n12818), .A2(n12817), .A3(n12816), .A4(n12815), .ZN(
        n12824) );
  AOI22_X1 U16209 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U16210 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16211 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12828), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U16212 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12819) );
  NAND4_X1 U16213 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12823) );
  OR2_X1 U16214 ( .A1(n12824), .A2(n12823), .ZN(n16330) );
  AND2_X1 U16215 ( .A1(n12825), .A2(n16330), .ZN(n12826) );
  AOI22_X1 U16216 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12827), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12839) );
  INV_X1 U16217 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U16218 ( .A1(n12828), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12830) );
  NAND2_X1 U16219 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12829) );
  OAI211_X1 U16220 ( .C1(n12832), .C2(n12831), .A(n12830), .B(n12829), .ZN(
        n12833) );
  INV_X1 U16221 ( .A(n12833), .ZN(n12838) );
  AOI22_X1 U16222 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16223 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10840), .B1(
        n10495), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12836) );
  NAND4_X1 U16224 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        n12848) );
  AOI22_X1 U16225 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10551), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U16226 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11209), .B1(
        n12840), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U16227 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12842), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U16228 ( .A1(n10847), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12843) );
  NAND4_X1 U16229 ( .A1(n12846), .A2(n12845), .A3(n12844), .A4(n12843), .ZN(
        n12847) );
  OR2_X1 U16230 ( .A1(n12848), .A2(n12847), .ZN(n12882) );
  AOI22_X1 U16231 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9711), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12857) );
  AND2_X1 U16232 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12850) );
  OR2_X1 U16233 ( .A1(n12850), .A2(n12849), .ZN(n12997) );
  INV_X1 U16234 ( .A(n12997), .ZN(n14474) );
  NAND2_X1 U16235 ( .A1(n12989), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12852) );
  NAND2_X1 U16236 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12851) );
  AND3_X1 U16237 ( .A1(n14474), .A2(n12852), .A3(n12851), .ZN(n12856) );
  AOI22_X1 U16238 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16239 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12854) );
  NAND4_X1 U16240 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n12854), .ZN(
        n12866) );
  AOI22_X1 U16241 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9709), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16242 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12996), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U16243 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12862) );
  NAND2_X1 U16244 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12860) );
  NAND2_X1 U16245 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12859) );
  AND3_X1 U16246 ( .A1(n12860), .A2(n12997), .A3(n12859), .ZN(n12861) );
  NAND4_X1 U16247 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n12861), .ZN(
        n12865) );
  NAND2_X1 U16248 ( .A1(n12882), .A2(n16312), .ZN(n12887) );
  AOI22_X1 U16249 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9709), .B1(n9711), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12872) );
  AOI22_X1 U16250 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9704), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U16251 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12911), .B1(
        n14449), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12870) );
  NAND2_X1 U16252 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12868) );
  NAND2_X1 U16253 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12867) );
  AND3_X1 U16254 ( .A1(n12868), .A2(n12867), .A3(n12997), .ZN(n12869) );
  NAND4_X1 U16255 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n12869), .ZN(
        n12880) );
  AOI22_X1 U16256 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12878) );
  NAND2_X1 U16257 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12874) );
  NAND2_X1 U16258 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12873) );
  AND3_X1 U16259 ( .A1(n14474), .A2(n12874), .A3(n12873), .ZN(n12877) );
  AOI22_X1 U16260 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9703), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U16261 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12875) );
  NAND4_X1 U16262 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        n12879) );
  NAND2_X1 U16263 ( .A1(n12880), .A2(n12879), .ZN(n12886) );
  XNOR2_X1 U16264 ( .A(n12887), .B(n12886), .ZN(n12881) );
  NOR2_X1 U16265 ( .A1(n12881), .A2(n14153), .ZN(n16316) );
  NAND2_X1 U16266 ( .A1(n11002), .A2(n16312), .ZN(n12883) );
  XNOR2_X1 U16267 ( .A(n12883), .B(n12882), .ZN(n16313) );
  NAND2_X1 U16268 ( .A1(n16316), .A2(n16313), .ZN(n12885) );
  NOR2_X1 U16269 ( .A1(n11002), .A2(n12886), .ZN(n16315) );
  NAND3_X1 U16270 ( .A1(n16313), .A2(n16312), .A3(n16315), .ZN(n12884) );
  NOR2_X1 U16271 ( .A1(n12887), .A2(n12886), .ZN(n12902) );
  AOI22_X1 U16272 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U16273 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12889) );
  NAND2_X1 U16274 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12888) );
  AND3_X1 U16275 ( .A1(n14474), .A2(n12889), .A3(n12888), .ZN(n12892) );
  AOI22_X1 U16276 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16277 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12890) );
  NAND4_X1 U16278 ( .A1(n12893), .A2(n12892), .A3(n12891), .A4(n12890), .ZN(
        n12901) );
  AOI22_X1 U16279 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12986), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16280 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9706), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16281 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12897) );
  NAND2_X1 U16282 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12895) );
  NAND2_X1 U16283 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12894) );
  AND3_X1 U16284 ( .A1(n12895), .A2(n12894), .A3(n12997), .ZN(n12896) );
  NAND4_X1 U16285 ( .A1(n12899), .A2(n12898), .A3(n12897), .A4(n12896), .ZN(
        n12900) );
  AND2_X1 U16286 ( .A1(n12901), .A2(n12900), .ZN(n12920) );
  NAND2_X1 U16287 ( .A1(n12902), .A2(n12920), .ZN(n12941) );
  OAI211_X1 U16288 ( .C1(n12902), .C2(n12920), .A(n12943), .B(n12941), .ZN(
        n12922) );
  AOI22_X1 U16289 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12986), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12910) );
  NAND2_X1 U16290 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12905) );
  NAND2_X1 U16291 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12904) );
  AND3_X1 U16292 ( .A1(n14474), .A2(n12905), .A3(n12904), .ZN(n12909) );
  INV_X1 U16293 ( .A(n12906), .ZN(n12970) );
  AOI22_X1 U16294 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16295 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12907) );
  NAND4_X1 U16296 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n12907), .ZN(
        n12919) );
  AOI22_X1 U16297 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16298 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9706), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16299 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12915) );
  NAND2_X1 U16300 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12913) );
  NAND2_X1 U16301 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12912) );
  AND3_X1 U16302 ( .A1(n12913), .A2(n12912), .A3(n12997), .ZN(n12914) );
  NAND4_X1 U16303 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n12918) );
  NAND2_X1 U16304 ( .A1(n12919), .A2(n12918), .ZN(n16299) );
  NAND2_X1 U16305 ( .A1(n11051), .A2(n12920), .ZN(n16308) );
  INV_X1 U16306 ( .A(n12921), .ZN(n12923) );
  XNOR2_X1 U16307 ( .A(n12941), .B(n16299), .ZN(n12924) );
  NOR2_X1 U16308 ( .A1(n12924), .A2(n14153), .ZN(n16301) );
  AOI22_X1 U16309 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9709), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U16310 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16311 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16312 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U16313 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12927) );
  AND3_X1 U16314 ( .A1(n12928), .A2(n12927), .A3(n12997), .ZN(n12929) );
  NAND4_X1 U16315 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12940) );
  AOI22_X1 U16316 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12938) );
  NAND2_X1 U16317 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12934) );
  NAND2_X1 U16318 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12933) );
  AND3_X1 U16319 ( .A1(n14474), .A2(n12934), .A3(n12933), .ZN(n12937) );
  AOI22_X1 U16320 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9706), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16321 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12935) );
  NAND4_X1 U16322 ( .A1(n12938), .A2(n12937), .A3(n12936), .A4(n12935), .ZN(
        n12939) );
  NAND2_X1 U16323 ( .A1(n12940), .A2(n12939), .ZN(n12948) );
  INV_X1 U16324 ( .A(n12948), .ZN(n12945) );
  OR2_X1 U16325 ( .A1(n12941), .A2(n16299), .ZN(n12942) );
  INV_X1 U16326 ( .A(n12942), .ZN(n12944) );
  OAI211_X1 U16327 ( .C1(n12945), .C2(n12944), .A(n12979), .B(n12943), .ZN(
        n12946) );
  NOR2_X2 U16328 ( .A1(n12947), .A2(n16287), .ZN(n16294) );
  NOR2_X1 U16329 ( .A1(n11002), .A2(n12948), .ZN(n16293) );
  INV_X1 U16330 ( .A(n16287), .ZN(n12963) );
  AOI22_X1 U16331 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12986), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U16332 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16333 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12952) );
  NAND2_X1 U16334 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12950) );
  NAND2_X1 U16335 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12949) );
  AND3_X1 U16336 ( .A1(n12950), .A2(n12949), .A3(n12997), .ZN(n12951) );
  NAND4_X1 U16337 ( .A1(n12954), .A2(n12953), .A3(n12952), .A4(n12951), .ZN(
        n12962) );
  AOI22_X1 U16338 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12960) );
  NAND2_X1 U16339 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12956) );
  NAND2_X1 U16340 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12955) );
  AND3_X1 U16341 ( .A1(n14474), .A2(n12956), .A3(n12955), .ZN(n12959) );
  AOI22_X1 U16342 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9704), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U16343 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12957) );
  NAND4_X1 U16344 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n12961) );
  NAND2_X1 U16345 ( .A1(n12962), .A2(n12961), .ZN(n16288) );
  AOI22_X1 U16346 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12986), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12969) );
  NAND2_X1 U16347 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12965) );
  NAND2_X1 U16348 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12964) );
  AND3_X1 U16349 ( .A1(n14474), .A2(n12965), .A3(n12964), .ZN(n12968) );
  AOI22_X1 U16350 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9706), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16351 ( .A1(n12989), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16352 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12978) );
  AOI22_X1 U16353 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U16354 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12996), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U16355 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U16356 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12972) );
  NAND2_X1 U16357 ( .A1(n9703), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12971) );
  AND3_X1 U16358 ( .A1(n12972), .A2(n12997), .A3(n12971), .ZN(n12973) );
  NAND4_X1 U16359 ( .A1(n12976), .A2(n12975), .A3(n12974), .A4(n12973), .ZN(
        n12977) );
  NAND2_X1 U16360 ( .A1(n12978), .A2(n12977), .ZN(n12983) );
  INV_X1 U16361 ( .A(n12979), .ZN(n16286) );
  INV_X1 U16362 ( .A(n16288), .ZN(n12980) );
  AND2_X1 U16363 ( .A1(n11127), .A2(n12980), .ZN(n12981) );
  NAND2_X1 U16364 ( .A1(n16286), .A2(n12981), .ZN(n12982) );
  NOR2_X1 U16365 ( .A1(n12982), .A2(n12983), .ZN(n12984) );
  AOI21_X1 U16366 ( .B1(n12983), .B2(n12982), .A(n12984), .ZN(n16281) );
  INV_X1 U16367 ( .A(n12984), .ZN(n12985) );
  AOI22_X1 U16368 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16369 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U16370 ( .A1(n12988), .A2(n12987), .ZN(n13004) );
  INV_X1 U16371 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12992) );
  AOI21_X1 U16372 ( .B1(n12996), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12997), .ZN(n12991) );
  AOI22_X1 U16373 ( .A1(n12989), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12990) );
  OAI211_X1 U16374 ( .C1(n12853), .C2(n12992), .A(n12991), .B(n12990), .ZN(
        n13003) );
  AOI22_X1 U16375 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16376 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9704), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U16377 ( .A1(n12995), .A2(n12994), .ZN(n13002) );
  AOI22_X1 U16378 ( .A1(n14449), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12989), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U16379 ( .A1(n12996), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12999) );
  NAND2_X1 U16380 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12998) );
  NAND4_X1 U16381 ( .A1(n13000), .A2(n12999), .A3(n12998), .A4(n12997), .ZN(
        n13001) );
  OAI22_X1 U16382 ( .A1(n13004), .A2(n13003), .B1(n13002), .B2(n13001), .ZN(
        n13005) );
  INV_X1 U16383 ( .A(n13005), .ZN(n13006) );
  INV_X1 U16384 ( .A(n14491), .ZN(n13008) );
  NAND2_X1 U16385 ( .A1(n14605), .A2(n13008), .ZN(n13761) );
  INV_X1 U16386 ( .A(n17047), .ZN(n13010) );
  INV_X1 U16387 ( .A(n15917), .ZN(n14912) );
  NAND2_X1 U16388 ( .A1(n14912), .A2(n16350), .ZN(n13012) );
  NAND2_X1 U16389 ( .A1(n16360), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13011) );
  OAI21_X1 U16390 ( .B1(n14932), .B2(n16353), .A(n13013), .ZN(P2_U2857) );
  OAI21_X1 U16391 ( .B1(n16526), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16514), .ZN(n16525) );
  INV_X1 U16392 ( .A(n13015), .ZN(n13016) );
  XNOR2_X1 U16393 ( .A(n13018), .B(n16732), .ZN(n16531) );
  NOR2_X1 U16394 ( .A1(n16532), .A2(n16531), .ZN(n16738) );
  INV_X1 U16395 ( .A(n13018), .ZN(n13019) );
  AND2_X1 U16396 ( .A1(n13019), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13020) );
  AND2_X1 U16397 ( .A1(n13022), .A2(n13021), .ZN(n13023) );
  NAND2_X1 U16398 ( .A1(n16523), .A2(n11071), .ZN(n13037) );
  NOR2_X1 U16399 ( .A1(n13026), .A2(n13027), .ZN(n13028) );
  OR2_X1 U16400 ( .A1(n13025), .A2(n13028), .ZN(n16521) );
  OR2_X1 U16401 ( .A1(n11468), .A2(n15985), .ZN(n16517) );
  OR2_X1 U16402 ( .A1(n16747), .A2(n16730), .ZN(n13030) );
  MUX2_X1 U16403 ( .A(n16719), .B(n13030), .S(n13029), .Z(n13031) );
  OAI211_X1 U16404 ( .C1(n16521), .C2(n19803), .A(n16517), .B(n13031), .ZN(
        n13035) );
  OAI21_X1 U16405 ( .B1(n16000), .B2(n13033), .A(n13032), .ZN(n16403) );
  NOR2_X1 U16406 ( .A1(n16403), .A2(n16958), .ZN(n13034) );
  NOR2_X1 U16407 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  OAI211_X1 U16408 ( .C1(n16942), .C2(n16525), .A(n13037), .B(n13036), .ZN(
        P2_U3022) );
  INV_X1 U16409 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13310) );
  INV_X1 U16410 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U16411 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13039) );
  NAND2_X1 U16412 ( .A1(n18216), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13038) );
  OAI211_X1 U16413 ( .C1(n14403), .C2(n18080), .A(n13039), .B(n13038), .ZN(
        n13040) );
  INV_X1 U16414 ( .A(n13040), .ZN(n13046) );
  AOI22_X1 U16415 ( .A1(n13105), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16416 ( .A1(n13929), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13044) );
  INV_X1 U16417 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13042) );
  OR2_X1 U16418 ( .A1(n18224), .A2(n13042), .ZN(n13043) );
  NAND4_X1 U16419 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13053) );
  AOI22_X1 U16420 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U16421 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13086), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16422 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13049) );
  INV_X2 U16423 ( .A(n9745), .ZN(n18230) );
  AOI22_X1 U16424 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13048) );
  NAND4_X1 U16425 ( .A1(n13051), .A2(n13050), .A3(n13049), .A4(n13048), .ZN(
        n13052) );
  OR2_X2 U16426 ( .A1(n13053), .A2(n13052), .ZN(n14300) );
  INV_X1 U16427 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13054) );
  OR2_X1 U16428 ( .A1(n18224), .A2(n13054), .ZN(n13059) );
  INV_X1 U16429 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18202) );
  OR2_X1 U16430 ( .A1(n13055), .A2(n18202), .ZN(n13058) );
  NAND2_X1 U16431 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13057) );
  NAND2_X1 U16432 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13056) );
  AND4_X1 U16433 ( .A1(n13059), .A2(n13058), .A3(n13057), .A4(n13056), .ZN(
        n13076) );
  NAND2_X1 U16434 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13063) );
  NAND2_X1 U16435 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13062) );
  NAND2_X1 U16436 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13061) );
  NAND2_X1 U16437 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13060) );
  NAND2_X1 U16438 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13067) );
  NAND2_X1 U16439 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13066) );
  NAND2_X1 U16440 ( .A1(n13086), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13065) );
  NAND2_X1 U16441 ( .A1(n13047), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13064) );
  NAND2_X1 U16442 ( .A1(n13105), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13072) );
  NAND2_X1 U16443 ( .A1(n13068), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13071) );
  NAND2_X1 U16444 ( .A1(n13929), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13070) );
  NAND2_X1 U16445 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13069) );
  NAND4_X4 U16446 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13249) );
  NAND2_X2 U16447 ( .A1(n14300), .A2(n13249), .ZN(n13116) );
  OAI21_X2 U16448 ( .B1(n14300), .B2(n13249), .A(n13116), .ZN(n13094) );
  XNOR2_X1 U16449 ( .A(n13249), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17176) );
  NAND2_X1 U16450 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13078) );
  NAND2_X1 U16451 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13077) );
  OAI211_X1 U16452 ( .C1(n14359), .C2(n18223), .A(n13078), .B(n13077), .ZN(
        n13079) );
  INV_X1 U16453 ( .A(n13079), .ZN(n13085) );
  AOI22_X1 U16454 ( .A1(n13068), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16455 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13083) );
  INV_X1 U16456 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13081) );
  OR2_X1 U16457 ( .A1(n18224), .A2(n13081), .ZN(n13082) );
  AOI22_X1 U16458 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13105), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16459 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13086), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16460 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16461 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13088) );
  AND2_X1 U16462 ( .A1(n14223), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17177) );
  NAND2_X1 U16463 ( .A1(n17176), .A2(n17177), .ZN(n13093) );
  INV_X1 U16464 ( .A(n13249), .ZN(n14222) );
  NAND2_X1 U16465 ( .A1(n14222), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13092) );
  NAND2_X1 U16466 ( .A1(n13093), .A2(n13092), .ZN(n14099) );
  NAND2_X1 U16467 ( .A1(n14098), .A2(n14099), .ZN(n13097) );
  INV_X1 U16468 ( .A(n13094), .ZN(n13095) );
  NAND2_X1 U16469 ( .A1(n13095), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13096) );
  NAND2_X1 U16470 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13100) );
  NAND2_X1 U16471 ( .A1(n13929), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13099) );
  NAND2_X1 U16472 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13098) );
  AOI22_X1 U16473 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16474 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13103) );
  INV_X1 U16475 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13101) );
  OR2_X1 U16476 ( .A1(n18224), .A2(n13101), .ZN(n13102) );
  NAND4_X1 U16477 ( .A1(n10398), .A2(n13104), .A3(n13103), .A4(n13102), .ZN(
        n13111) );
  AOI22_X1 U16478 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16479 ( .A1(n13086), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13108) );
  AOI22_X1 U16480 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13105), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16481 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13106) );
  NAND4_X1 U16482 ( .A1(n13109), .A2(n13108), .A3(n13107), .A4(n13106), .ZN(
        n13110) );
  INV_X1 U16483 ( .A(n13255), .ZN(n18420) );
  XNOR2_X1 U16484 ( .A(n18420), .B(n13116), .ZN(n13113) );
  NAND2_X1 U16485 ( .A1(n13112), .A2(n13114), .ZN(n13115) );
  INV_X1 U16486 ( .A(n13116), .ZN(n13117) );
  NAND2_X1 U16487 ( .A1(n13117), .A2(n13255), .ZN(n13136) );
  INV_X1 U16488 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14417) );
  NAND2_X1 U16489 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13119) );
  NAND2_X1 U16490 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13118) );
  OAI211_X1 U16491 ( .C1(n14417), .C2(n18141), .A(n13119), .B(n13118), .ZN(
        n13120) );
  INV_X1 U16492 ( .A(n13120), .ZN(n13125) );
  AOI22_X1 U16493 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13068), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16494 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13123) );
  INV_X1 U16495 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13121) );
  OR2_X1 U16496 ( .A1(n18224), .A2(n13121), .ZN(n13122) );
  NAND4_X1 U16497 ( .A1(n13125), .A2(n13124), .A3(n13123), .A4(n13122), .ZN(
        n13131) );
  AOI22_X1 U16498 ( .A1(n13087), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16499 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13086), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16500 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13127) );
  AOI22_X1 U16501 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13126) );
  NAND4_X1 U16502 ( .A1(n13129), .A2(n13128), .A3(n13127), .A4(n13126), .ZN(
        n13130) );
  XNOR2_X1 U16503 ( .A(n13136), .B(n18416), .ZN(n13132) );
  XNOR2_X1 U16504 ( .A(n13132), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18783) );
  INV_X1 U16505 ( .A(n13132), .ZN(n13133) );
  NAND2_X1 U16506 ( .A1(n13133), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13134) );
  NAND2_X2 U16507 ( .A1(n13135), .A2(n13134), .ZN(n13154) );
  INV_X1 U16508 ( .A(n13136), .ZN(n13137) );
  NAND2_X1 U16509 ( .A1(n13137), .A2(n13259), .ZN(n13156) );
  INV_X1 U16510 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17968) );
  OR2_X1 U16511 ( .A1(n18224), .A2(n17968), .ZN(n13141) );
  NAND2_X1 U16512 ( .A1(n18222), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13140) );
  NAND2_X1 U16513 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13139) );
  NAND2_X1 U16514 ( .A1(n9701), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13138) );
  AOI22_X1 U16515 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18194), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U16516 ( .A1(n14395), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13143) );
  NAND3_X1 U16517 ( .A1(n13145), .A2(n13144), .A3(n13143), .ZN(n13151) );
  AOI22_X1 U16518 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13149) );
  AOI22_X1 U16519 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13148) );
  AOI22_X1 U16520 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16521 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13146) );
  NAND4_X1 U16522 ( .A1(n13149), .A2(n13148), .A3(n13147), .A4(n13146), .ZN(
        n13150) );
  INV_X1 U16523 ( .A(n13250), .ZN(n18412) );
  XNOR2_X1 U16524 ( .A(n13156), .B(n18412), .ZN(n13152) );
  XNOR2_X2 U16525 ( .A(n13154), .B(n13152), .ZN(n14104) );
  INV_X1 U16526 ( .A(n13152), .ZN(n13153) );
  NAND2_X1 U16527 ( .A1(n13154), .A2(n13153), .ZN(n13155) );
  INV_X1 U16528 ( .A(n13156), .ZN(n13157) );
  NAND2_X1 U16529 ( .A1(n13157), .A2(n13250), .ZN(n13175) );
  INV_X1 U16530 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17906) );
  NAND2_X1 U16531 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13159) );
  NAND2_X1 U16532 ( .A1(n18216), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13158) );
  OAI211_X1 U16533 ( .C1(n17906), .C2(n18141), .A(n13159), .B(n13158), .ZN(
        n13160) );
  INV_X1 U16534 ( .A(n13160), .ZN(n13165) );
  AOI22_X1 U16535 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U16536 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13163) );
  INV_X1 U16537 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13161) );
  OR2_X1 U16538 ( .A1(n18224), .A2(n13161), .ZN(n13162) );
  NAND4_X1 U16539 ( .A1(n13165), .A2(n13164), .A3(n13163), .A4(n13162), .ZN(
        n13171) );
  AOI22_X1 U16540 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13169) );
  AOI22_X1 U16541 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16542 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U16543 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13166) );
  NAND4_X1 U16544 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        n13170) );
  XNOR2_X1 U16545 ( .A(n13175), .B(n18409), .ZN(n13172) );
  XNOR2_X1 U16546 ( .A(n13172), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14079) );
  INV_X1 U16547 ( .A(n13172), .ZN(n13173) );
  NAND2_X1 U16548 ( .A1(n13173), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13174) );
  INV_X1 U16549 ( .A(n13175), .ZN(n13176) );
  INV_X1 U16550 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21625) );
  NAND2_X1 U16551 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13178) );
  NAND2_X1 U16552 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13177) );
  OAI211_X1 U16553 ( .C1(n21625), .C2(n18141), .A(n13178), .B(n13177), .ZN(
        n13179) );
  INV_X1 U16554 ( .A(n13179), .ZN(n13183) );
  AOI22_X1 U16555 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16556 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13181) );
  OR2_X1 U16557 ( .A1(n18224), .A2(n18084), .ZN(n13180) );
  NAND4_X1 U16558 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13189) );
  AOI22_X1 U16559 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U16560 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U16561 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U16562 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13184) );
  NAND4_X1 U16563 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13188) );
  INV_X1 U16564 ( .A(n13190), .ZN(n13534) );
  NAND2_X1 U16565 ( .A1(n13534), .A2(n18405), .ZN(n13191) );
  NAND2_X1 U16566 ( .A1(n18734), .A2(n13191), .ZN(n13192) );
  INV_X1 U16567 ( .A(n13192), .ZN(n13193) );
  NAND2_X1 U16568 ( .A1(n13194), .A2(n13193), .ZN(n13195) );
  NAND2_X1 U16569 ( .A1(n18734), .A2(n13196), .ZN(n13197) );
  NOR2_X1 U16570 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13198) );
  INV_X1 U16571 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13199) );
  INV_X1 U16572 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18991) );
  NOR2_X1 U16573 ( .A1(n18991), .A2(n18970), .ZN(n18958) );
  NAND2_X1 U16574 ( .A1(n18958), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18715) );
  NAND2_X1 U16575 ( .A1(n18911), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18917) );
  OR2_X2 U16576 ( .A1(n18956), .A2(n18644), .ZN(n18899) );
  NOR2_X1 U16577 ( .A1(n18734), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13201) );
  AOI21_X1 U16578 ( .B1(n18899), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n13201), .ZN(n13202) );
  INV_X1 U16579 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17239) );
  NAND2_X1 U16580 ( .A1(n17129), .A2(n17239), .ZN(n13203) );
  NAND2_X1 U16581 ( .A1(n13204), .A2(n18899), .ZN(n18643) );
  INV_X1 U16582 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18587) );
  NOR2_X1 U16583 ( .A1(n18887), .A2(n18853), .ZN(n18867) );
  NAND2_X1 U16584 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18867), .ZN(
        n18843) );
  NOR2_X1 U16585 ( .A1(n18587), .A2(n18843), .ZN(n18842) );
  AND2_X1 U16586 ( .A1(n18842), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18569) );
  AND2_X1 U16587 ( .A1(n17229), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13205) );
  NAND2_X1 U16588 ( .A1(n18643), .A2(n18551), .ZN(n13208) );
  NAND2_X1 U16589 ( .A1(n18734), .A2(n18587), .ZN(n18636) );
  NOR2_X1 U16590 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18636), .ZN(
        n13206) );
  NAND2_X1 U16591 ( .A1(n13206), .A2(n18853), .ZN(n18609) );
  NOR2_X1 U16592 ( .A1(n18609), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18582) );
  INV_X1 U16593 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18857) );
  INV_X1 U16594 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18796) );
  NAND3_X1 U16595 ( .A1(n18582), .A2(n18857), .A3(n18796), .ZN(n13207) );
  INV_X1 U16596 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18830) );
  NAND2_X1 U16597 ( .A1(n18643), .A2(n17229), .ZN(n18607) );
  NAND2_X1 U16598 ( .A1(n18568), .A2(n18607), .ZN(n18637) );
  AND2_X1 U16599 ( .A1(n18569), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13209) );
  NAND2_X1 U16600 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17214) );
  OAI21_X1 U16601 ( .B1(n18547), .B2(n17214), .A(n18703), .ZN(n13210) );
  OAI21_X2 U16602 ( .B1(n17110), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13210), .ZN(n13211) );
  OR2_X1 U16603 ( .A1(n18734), .A2(n21581), .ZN(n13526) );
  NAND2_X1 U16604 ( .A1(n13211), .A2(n14698), .ZN(n13524) );
  NAND2_X1 U16605 ( .A1(n18734), .A2(n21581), .ZN(n13525) );
  OR2_X2 U16606 ( .A1(n13524), .A2(n13525), .ZN(n13212) );
  OAI21_X2 U16607 ( .B1(n17101), .B2(n13526), .A(n13212), .ZN(n17086) );
  INV_X1 U16608 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13306) );
  NAND2_X1 U16609 ( .A1(n18734), .A2(n13310), .ZN(n13215) );
  AOI21_X1 U16610 ( .B1(n13213), .B2(n17072), .A(n13215), .ZN(n13214) );
  INV_X1 U16611 ( .A(n13214), .ZN(n13220) );
  OAI21_X1 U16612 ( .B1(n18703), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13216) );
  OAI211_X1 U16613 ( .C1(n17072), .C2(n18703), .A(n13216), .B(n13215), .ZN(
        n13217) );
  AOI21_X1 U16614 ( .B1(n17073), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13217), .ZN(n13218) );
  INV_X1 U16615 ( .A(n13218), .ZN(n13219) );
  NAND3_X1 U16616 ( .A1(n9775), .A2(n13220), .A3(n13219), .ZN(n17071) );
  INV_X1 U16617 ( .A(n13283), .ZN(n13291) );
  NOR3_X1 U16618 ( .A1(n13222), .A2(n13291), .A3(n13221), .ZN(n13225) );
  NAND2_X1 U16619 ( .A1(n13223), .A2(n13885), .ZN(n13224) );
  NAND2_X1 U16620 ( .A1(n9797), .A2(n13248), .ZN(n13227) );
  AOI21_X1 U16621 ( .B1(n13228), .B2(n13227), .A(n13226), .ZN(n13894) );
  OAI21_X1 U16622 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19477), .A(
        n13229), .ZN(n13234) );
  NOR2_X1 U16623 ( .A1(n13239), .A2(n13234), .ZN(n14687) );
  NOR2_X1 U16624 ( .A1(n19626), .A2(n13230), .ZN(n13233) );
  NAND2_X1 U16625 ( .A1(n13233), .A2(n13231), .ZN(n13246) );
  OAI21_X1 U16626 ( .B1(n19042), .B2(n18490), .A(n19624), .ZN(n13232) );
  OAI21_X1 U16627 ( .B1(n13233), .B2(n13232), .A(n19627), .ZN(n19472) );
  OAI22_X1 U16628 ( .A1(n14687), .A2(n13246), .B1(n13289), .B2(n19472), .ZN(
        n13243) );
  INV_X1 U16629 ( .A(n13234), .ZN(n13235) );
  NAND2_X1 U16630 ( .A1(n13236), .A2(n13235), .ZN(n13237) );
  OR2_X1 U16631 ( .A1(n13238), .A2(n13237), .ZN(n13242) );
  AND2_X1 U16632 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  AOI22_X1 U16633 ( .A1(n13243), .A2(n19469), .B1(n13289), .B2(n19466), .ZN(
        n13244) );
  NAND2_X1 U16634 ( .A1(n13894), .A2(n13244), .ZN(n13245) );
  INV_X1 U16635 ( .A(n13246), .ZN(n13247) );
  INV_X1 U16636 ( .A(n14300), .ZN(n13251) );
  NAND2_X1 U16637 ( .A1(n13254), .A2(n13251), .ZN(n13256) );
  NAND2_X1 U16638 ( .A1(n13256), .A2(n13255), .ZN(n13260) );
  NOR2_X1 U16639 ( .A1(n18416), .A2(n13260), .ZN(n13266) );
  NAND2_X1 U16640 ( .A1(n13266), .A2(n13250), .ZN(n13270) );
  NOR2_X1 U16641 ( .A1(n18409), .A2(n13270), .ZN(n13274) );
  NAND2_X1 U16642 ( .A1(n13274), .A2(n14692), .ZN(n13275) );
  XNOR2_X1 U16643 ( .A(n13254), .B(n13251), .ZN(n13252) );
  NOR2_X1 U16644 ( .A1(n14223), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17175) );
  INV_X1 U16645 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U16646 ( .B1(n13256), .B2(n13255), .A(n13260), .ZN(n13257) );
  XNOR2_X1 U16647 ( .A(n14130), .B(n13257), .ZN(n14132) );
  NOR2_X1 U16648 ( .A1(n14133), .A2(n14132), .ZN(n14131) );
  NOR2_X1 U16649 ( .A1(n14130), .A2(n13257), .ZN(n13258) );
  XOR2_X1 U16650 ( .A(n13260), .B(n13259), .Z(n13263) );
  NOR2_X1 U16651 ( .A1(n13264), .A2(n13263), .ZN(n13265) );
  XNOR2_X1 U16652 ( .A(n13266), .B(n18412), .ZN(n13267) );
  XNOR2_X1 U16653 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13267), .ZN(
        n14109) );
  AND2_X1 U16654 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13267), .ZN(
        n13268) );
  NOR2_X1 U16655 ( .A1(n14108), .A2(n13268), .ZN(n13272) );
  XOR2_X1 U16656 ( .A(n13270), .B(n13269), .Z(n13271) );
  NOR2_X1 U16657 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  XNOR2_X1 U16658 ( .A(n13272), .B(n13271), .ZN(n14075) );
  INV_X1 U16659 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14086) );
  NOR2_X1 U16660 ( .A1(n14075), .A2(n14086), .ZN(n14074) );
  NOR2_X1 U16661 ( .A1(n13273), .A2(n14074), .ZN(n13276) );
  XNOR2_X1 U16662 ( .A(n13274), .B(n14692), .ZN(n13277) );
  NAND2_X1 U16663 ( .A1(n13276), .A2(n13277), .ZN(n14116) );
  NAND2_X1 U16664 ( .A1(n14116), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13279) );
  NOR2_X1 U16665 ( .A1(n13275), .A2(n13279), .ZN(n13281) );
  INV_X1 U16666 ( .A(n13275), .ZN(n13280) );
  OR2_X1 U16667 ( .A1(n13277), .A2(n13276), .ZN(n14117) );
  OAI21_X1 U16668 ( .B1(n13280), .B2(n13279), .A(n14117), .ZN(n13278) );
  AOI21_X1 U16669 ( .B1(n13280), .B2(n13279), .A(n13278), .ZN(n17141) );
  INV_X1 U16670 ( .A(n18911), .ZN(n18660) );
  INV_X1 U16671 ( .A(n18551), .ZN(n17113) );
  AND2_X1 U16672 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13304) );
  INV_X1 U16673 ( .A(n13886), .ZN(n13282) );
  NAND2_X2 U16674 ( .A1(n13282), .A2(n13887), .ZN(n18981) );
  NOR3_X1 U16675 ( .A1(n13284), .A2(n13283), .A3(n19626), .ZN(n13287) );
  INV_X1 U16676 ( .A(n13285), .ZN(n13286) );
  OAI21_X2 U16677 ( .B1(n13909), .B2(n13886), .A(n13908), .ZN(n18978) );
  NAND2_X1 U16678 ( .A1(n13892), .A2(n13288), .ZN(n19637) );
  INV_X1 U16679 ( .A(n13289), .ZN(n13290) );
  INV_X1 U16680 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21598) );
  INV_X1 U16681 ( .A(n18899), .ZN(n13292) );
  NAND2_X1 U16682 ( .A1(n18551), .A2(n13292), .ZN(n18824) );
  NOR2_X1 U16683 ( .A1(n18830), .A2(n18824), .ZN(n18538) );
  NAND2_X1 U16684 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18538), .ZN(
        n18537) );
  NOR2_X1 U16685 ( .A1(n21598), .A2(n18537), .ZN(n17210) );
  NAND2_X1 U16686 ( .A1(n17210), .A2(n13304), .ZN(n17096) );
  AND2_X1 U16687 ( .A1(n18951), .A2(n18996), .ZN(n18926) );
  INV_X1 U16688 ( .A(n18926), .ZN(n18820) );
  INV_X1 U16689 ( .A(n18569), .ZN(n18573) );
  AOI21_X1 U16690 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14077) );
  INV_X1 U16691 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14120) );
  INV_X1 U16692 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14106) );
  NOR3_X1 U16693 ( .A1(n14106), .A2(n14130), .A3(n19018), .ZN(n14081) );
  NAND2_X1 U16694 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14081), .ZN(
        n14119) );
  OR2_X1 U16695 ( .A1(n14120), .A2(n14119), .ZN(n18980) );
  NOR2_X1 U16696 ( .A1(n18993), .A2(n18980), .ZN(n13294) );
  INV_X1 U16697 ( .A(n13294), .ZN(n13293) );
  NOR2_X1 U16698 ( .A1(n14077), .A2(n13293), .ZN(n18912) );
  NAND3_X1 U16699 ( .A1(n17229), .A2(n18888), .A3(n18912), .ZN(n17232) );
  INV_X1 U16700 ( .A(n17232), .ZN(n18847) );
  NAND2_X1 U16701 ( .A1(n10299), .A2(n18847), .ZN(n13540) );
  AOI21_X1 U16702 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18978), .A(
        n18981), .ZN(n14090) );
  INV_X1 U16703 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14103) );
  NOR2_X1 U16704 ( .A1(n14103), .A2(n13253), .ZN(n14076) );
  NAND2_X1 U16705 ( .A1(n14076), .A2(n13294), .ZN(n18916) );
  NOR2_X1 U16706 ( .A1(n18644), .A2(n18916), .ZN(n18846) );
  NAND3_X1 U16707 ( .A1(n17229), .A2(n18569), .A3(n18846), .ZN(n17215) );
  OAI22_X1 U16708 ( .A1(n18573), .A2(n13540), .B1(n14090), .B2(n17215), .ZN(
        n18809) );
  INV_X1 U16709 ( .A(n17214), .ZN(n13298) );
  NAND2_X1 U16710 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18808) );
  INV_X1 U16711 ( .A(n18808), .ZN(n18810) );
  NAND2_X1 U16712 ( .A1(n13298), .A2(n18810), .ZN(n13300) );
  INV_X1 U16713 ( .A(n13300), .ZN(n17220) );
  AND2_X1 U16714 ( .A1(n17220), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13295) );
  AND2_X1 U16715 ( .A1(n18951), .A2(n13295), .ZN(n13545) );
  NAND3_X1 U16716 ( .A1(n18809), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n13545), .ZN(n13296) );
  OAI21_X1 U16717 ( .B1(n17096), .B2(n18820), .A(n13296), .ZN(n13297) );
  INV_X1 U16718 ( .A(n17204), .ZN(n13312) );
  NAND3_X1 U16719 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n13310), .ZN(n17063) );
  INV_X1 U16720 ( .A(n17063), .ZN(n13311) );
  NOR2_X1 U16721 ( .A1(n18573), .A2(n17232), .ZN(n18825) );
  NAND3_X1 U16722 ( .A1(n13298), .A2(n18825), .A3(n18810), .ZN(n13299) );
  NAND2_X1 U16723 ( .A1(n10299), .A2(n13299), .ZN(n17216) );
  AND2_X1 U16724 ( .A1(n18998), .A2(n17216), .ZN(n13303) );
  OAI22_X1 U16725 ( .A1(n18978), .A2(n18981), .B1(n17215), .B2(n13300), .ZN(
        n13302) );
  NAND2_X1 U16726 ( .A1(n18978), .A2(n10151), .ZN(n14072) );
  INV_X1 U16727 ( .A(n14072), .ZN(n17228) );
  AOI21_X1 U16728 ( .B1(n18978), .B2(n14698), .A(n17228), .ZN(n13301) );
  AND2_X1 U16729 ( .A1(n13302), .A2(n13301), .ZN(n17202) );
  NAND2_X1 U16730 ( .A1(n13303), .A2(n17202), .ZN(n13528) );
  AND2_X1 U16731 ( .A1(n18951), .A2(n18892), .ZN(n19010) );
  AND2_X1 U16732 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n13304), .ZN(
        n13305) );
  AOI22_X1 U16733 ( .A1(n13528), .A2(n10420), .B1(n19010), .B2(n10165), .ZN(
        n17191) );
  OAI21_X1 U16734 ( .B1(n13306), .B2(n17187), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17051) );
  NAND2_X1 U16735 ( .A1(n9696), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n17059) );
  AND2_X1 U16736 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13306), .ZN(
        n13308) );
  NAND2_X1 U16737 ( .A1(n17210), .A2(n13305), .ZN(n17189) );
  OAI21_X1 U16738 ( .B1(n13306), .B2(n17189), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17062) );
  INV_X1 U16739 ( .A(n17062), .ZN(n13307) );
  AOI22_X1 U16740 ( .A1(n19010), .A2(n13308), .B1(n18926), .B2(n13307), .ZN(
        n13309) );
  OAI21_X1 U16741 ( .B1(n17071), .B2(n18976), .A(n13313), .ZN(P3_U2831) );
  NAND2_X1 U16742 ( .A1(n13314), .A2(n16543), .ZN(n13315) );
  XNOR2_X1 U16743 ( .A(n13316), .B(n13315), .ZN(n16785) );
  NOR2_X1 U16744 ( .A1(n16770), .A2(n16690), .ZN(n13330) );
  INV_X1 U16745 ( .A(n13318), .ZN(n13319) );
  AOI21_X1 U16746 ( .B1(n13320), .B2(n14761), .A(n13319), .ZN(n16779) );
  NAND2_X1 U16747 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n15013), .ZN(
        n15012) );
  INV_X1 U16748 ( .A(n15012), .ZN(n13321) );
  INV_X1 U16749 ( .A(n14763), .ZN(n13323) );
  INV_X1 U16750 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13322) );
  NAND2_X1 U16751 ( .A1(n13323), .A2(n13322), .ZN(n13324) );
  NAND2_X1 U16752 ( .A1(n9725), .A2(n13324), .ZN(n16045) );
  NOR2_X1 U16753 ( .A1(n11468), .A2(n13325), .ZN(n16771) );
  AOI21_X1 U16754 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16771), .ZN(n13326) );
  OAI21_X1 U16755 ( .B1(n19758), .B2(n16045), .A(n13326), .ZN(n13327) );
  AOI21_X1 U16756 ( .B1(n16779), .B2(n19787), .A(n13327), .ZN(n13328) );
  AND2_X1 U16757 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13497) );
  NAND2_X1 U16758 ( .A1(n13497), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15513) );
  NAND2_X1 U16759 ( .A1(n13336), .A2(n15513), .ZN(n13333) );
  NAND2_X1 U16760 ( .A1(n13334), .A2(n13333), .ZN(n15527) );
  NAND3_X1 U16761 ( .A1(n13335), .A2(n14824), .A3(n13508), .ZN(n15515) );
  OAI21_X2 U16762 ( .B1(n13336), .B2(n15515), .A(n12192), .ZN(n15538) );
  NOR2_X1 U16763 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15705) );
  INV_X1 U16764 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14881) );
  INV_X1 U16765 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15699) );
  AND2_X1 U16766 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15706) );
  NAND4_X1 U16767 ( .A1(n15657), .A2(n15706), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13337) );
  NOR2_X1 U16768 ( .A1(n20812), .A2(n20804), .ZN(n13339) );
  NAND2_X1 U16769 ( .A1(n13486), .A2(n13339), .ZN(n13820) );
  INV_X1 U16770 ( .A(n17306), .ZN(n17290) );
  OAI21_X1 U16771 ( .B1(n20792), .B2(n17290), .A(n21487), .ZN(n14731) );
  INV_X1 U16772 ( .A(n14146), .ZN(n13341) );
  OAI211_X1 U16773 ( .C1(n13820), .C2(n14731), .A(n20776), .B(n13341), .ZN(
        n13342) );
  NAND2_X1 U16774 ( .A1(n13342), .A2(n12249), .ZN(n13358) );
  OR2_X1 U16775 ( .A1(n13744), .A2(n13361), .ZN(n13347) );
  NOR2_X1 U16776 ( .A1(n13344), .A2(n20812), .ZN(n13498) );
  NOR2_X1 U16777 ( .A1(n13498), .A2(n14727), .ZN(n13345) );
  NAND2_X1 U16778 ( .A1(n13346), .A2(n13345), .ZN(n13494) );
  NOR3_X1 U16779 ( .A1(n13350), .A2(n13349), .A3(n13348), .ZN(n13353) );
  OAI21_X1 U16780 ( .B1(n13353), .B2(n13352), .A(n13351), .ZN(n13746) );
  NAND2_X1 U16781 ( .A1(n20792), .A2(n17306), .ZN(n13354) );
  NAND4_X1 U16782 ( .A1(n13746), .A2(n20796), .A3(n21487), .A4(n13354), .ZN(
        n13355) );
  NAND3_X1 U16783 ( .A1(n13356), .A2(n13828), .A3(n13355), .ZN(n13357) );
  NAND2_X1 U16784 ( .A1(n13361), .A2(n11926), .ZN(n13844) );
  INV_X1 U16785 ( .A(n13844), .ZN(n13362) );
  NOR2_X1 U16786 ( .A1(n13362), .A2(n17277), .ZN(n13741) );
  NAND2_X1 U16787 ( .A1(n13744), .A2(n13823), .ZN(n13838) );
  INV_X1 U16788 ( .A(n13363), .ZN(n13364) );
  NAND2_X1 U16789 ( .A1(n13364), .A2(n20804), .ZN(n13365) );
  NAND4_X1 U16790 ( .A1(n13366), .A2(n13741), .A3(n13838), .A4(n13365), .ZN(
        n13367) );
  NAND2_X1 U16791 ( .A1(n13400), .A2(n20767), .ZN(n13372) );
  INV_X1 U16792 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U16793 ( .A1(n14064), .A2(n15355), .ZN(n13371) );
  NAND3_X1 U16794 ( .A1(n13372), .A2(n13375), .A3(n13371), .ZN(n13373) );
  NAND2_X1 U16795 ( .A1(n13400), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13377) );
  INV_X1 U16796 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13883) );
  NAND2_X1 U16797 ( .A1(n13375), .A2(n13883), .ZN(n13376) );
  NAND2_X1 U16798 ( .A1(n13377), .A2(n13376), .ZN(n13871) );
  XNOR2_X1 U16799 ( .A(n13378), .B(n13871), .ZN(n14065) );
  NAND2_X1 U16800 ( .A1(n14065), .A2(n14064), .ZN(n14063) );
  NAND2_X1 U16801 ( .A1(n14063), .A2(n13378), .ZN(n14172) );
  OR2_X1 U16802 ( .A1(n13470), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13383) );
  INV_X1 U16803 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20751) );
  NAND2_X1 U16804 ( .A1(n13400), .A2(n20751), .ZN(n13381) );
  INV_X1 U16805 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13379) );
  NAND2_X1 U16806 ( .A1(n14064), .A2(n13379), .ZN(n13380) );
  NAND3_X1 U16807 ( .A1(n13381), .A2(n13375), .A3(n13380), .ZN(n13382) );
  AND2_X1 U16808 ( .A1(n13383), .A2(n13382), .ZN(n14171) );
  MUX2_X1 U16809 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13384) );
  OAI21_X1 U16810 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13870), .A(
        n13384), .ZN(n14442) );
  INV_X1 U16811 ( .A(n14442), .ZN(n13385) );
  MUX2_X1 U16812 ( .A(n13470), .B(n13400), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13388) );
  INV_X1 U16813 ( .A(n13400), .ZN(n13395) );
  NAND2_X1 U16814 ( .A1(n13395), .A2(n13819), .ZN(n13402) );
  NAND2_X1 U16815 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13819), .ZN(
        n13386) );
  AND2_X1 U16816 ( .A1(n13402), .A2(n13386), .ZN(n13387) );
  INV_X1 U16817 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20652) );
  NAND2_X1 U16818 ( .A1(n14064), .A2(n20652), .ZN(n13390) );
  NAND2_X1 U16819 ( .A1(n13375), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13389) );
  NAND3_X1 U16820 ( .A1(n13390), .A2(n13400), .A3(n13389), .ZN(n13391) );
  OAI21_X1 U16821 ( .B1(n13468), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13391), .ZN(
        n17353) );
  MUX2_X1 U16822 ( .A(n13470), .B(n13400), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13394) );
  NAND2_X1 U16823 ( .A1(n13819), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13393) );
  INV_X1 U16824 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20646) );
  NAND2_X1 U16825 ( .A1(n13452), .A2(n20646), .ZN(n13399) );
  NAND2_X1 U16826 ( .A1(n14064), .A2(n20646), .ZN(n13397) );
  NAND2_X1 U16827 ( .A1(n13375), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13396) );
  NAND3_X1 U16828 ( .A1(n13397), .A2(n13400), .A3(n13396), .ZN(n13398) );
  MUX2_X1 U16829 ( .A(n13470), .B(n13400), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13404) );
  NAND2_X1 U16830 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13819), .ZN(
        n13401) );
  AND2_X1 U16831 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  NAND2_X1 U16832 ( .A1(n13404), .A2(n13403), .ZN(n15879) );
  INV_X1 U16833 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20642) );
  NAND2_X1 U16834 ( .A1(n13452), .A2(n20642), .ZN(n13408) );
  NAND2_X1 U16835 ( .A1(n14064), .A2(n20642), .ZN(n13406) );
  NAND2_X1 U16836 ( .A1(n13375), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13405) );
  NAND3_X1 U16837 ( .A1(n13406), .A2(n13400), .A3(n13405), .ZN(n13407) );
  AND2_X1 U16838 ( .A1(n13408), .A2(n13407), .ZN(n15878) );
  AND2_X1 U16839 ( .A1(n15879), .A2(n15878), .ZN(n13409) );
  OR2_X1 U16840 ( .A1(n13470), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13413) );
  NAND2_X1 U16841 ( .A1(n13400), .A2(n15666), .ZN(n13411) );
  INV_X1 U16842 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15394) );
  NAND2_X1 U16843 ( .A1(n14064), .A2(n15394), .ZN(n13410) );
  NAND3_X1 U16844 ( .A1(n13411), .A2(n13375), .A3(n13410), .ZN(n13412) );
  MUX2_X1 U16845 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13414) );
  OAI21_X1 U16846 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13870), .A(
        n13414), .ZN(n15320) );
  MUX2_X1 U16847 ( .A(n13470), .B(n13400), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13417) );
  NAND2_X1 U16848 ( .A1(n13819), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13416) );
  NAND2_X1 U16849 ( .A1(n13417), .A2(n13416), .ZN(n15304) );
  NAND2_X1 U16850 ( .A1(n10397), .A2(n15304), .ZN(n15306) );
  MUX2_X1 U16851 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13418) );
  OAI21_X1 U16852 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13870), .A(
        n13418), .ZN(n15287) );
  OR2_X1 U16853 ( .A1(n13470), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n13423) );
  NAND2_X1 U16854 ( .A1(n13400), .A2(n15820), .ZN(n13421) );
  INV_X1 U16855 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13419) );
  NAND2_X1 U16856 ( .A1(n14064), .A2(n13419), .ZN(n13420) );
  NAND3_X1 U16857 ( .A1(n13421), .A2(n13368), .A3(n13420), .ZN(n13422) );
  INV_X1 U16858 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n13424) );
  NAND2_X1 U16859 ( .A1(n14064), .A2(n13424), .ZN(n13426) );
  NAND2_X1 U16860 ( .A1(n13375), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13425) );
  NAND3_X1 U16861 ( .A1(n13426), .A2(n13400), .A3(n13425), .ZN(n13427) );
  OAI21_X1 U16862 ( .B1(n13468), .B2(P1_EBX_REG_15__SCAN_IN), .A(n13427), .ZN(
        n15256) );
  OR2_X1 U16863 ( .A1(n13470), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n13431) );
  INV_X1 U16864 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15805) );
  NAND2_X1 U16865 ( .A1(n13400), .A2(n15805), .ZN(n13429) );
  INV_X1 U16866 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U16867 ( .A1(n14064), .A2(n15387), .ZN(n13428) );
  NAND3_X1 U16868 ( .A1(n13429), .A2(n13375), .A3(n13428), .ZN(n13430) );
  NAND2_X1 U16869 ( .A1(n13431), .A2(n13430), .ZN(n15235) );
  MUX2_X1 U16870 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13433) );
  OR2_X1 U16871 ( .A1(n13870), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13432) );
  NAND2_X1 U16872 ( .A1(n13452), .A2(n21676), .ZN(n13437) );
  NAND2_X1 U16873 ( .A1(n14064), .A2(n21676), .ZN(n13435) );
  NAND2_X1 U16874 ( .A1(n13375), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13434) );
  NAND3_X1 U16875 ( .A1(n13435), .A2(n13400), .A3(n13434), .ZN(n13436) );
  OR2_X1 U16876 ( .A1(n13470), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n13442) );
  INV_X1 U16877 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13438) );
  NAND2_X1 U16878 ( .A1(n13400), .A2(n13438), .ZN(n13440) );
  INV_X1 U16879 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U16880 ( .A1(n14064), .A2(n15385), .ZN(n13439) );
  NAND3_X1 U16881 ( .A1(n13440), .A2(n13375), .A3(n13439), .ZN(n13441) );
  NAND2_X1 U16882 ( .A1(n13442), .A2(n13441), .ZN(n15185) );
  NAND2_X1 U16883 ( .A1(n15186), .A2(n15185), .ZN(n13443) );
  MUX2_X1 U16884 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13445) );
  OR2_X1 U16885 ( .A1(n13870), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13444) );
  MUX2_X1 U16886 ( .A(n13470), .B(n13400), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13447) );
  NAND2_X1 U16887 ( .A1(n13819), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13446) );
  NAND2_X1 U16888 ( .A1(n13447), .A2(n13446), .ZN(n15172) );
  MUX2_X1 U16889 ( .A(n13470), .B(n13400), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13449) );
  NAND2_X1 U16890 ( .A1(n13819), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13448) );
  MUX2_X1 U16891 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13450) );
  OAI21_X1 U16892 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13870), .A(
        n13450), .ZN(n14826) );
  NOR2_X1 U16893 ( .A1(n15149), .A2(n14826), .ZN(n13451) );
  INV_X1 U16894 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n13453) );
  NAND2_X1 U16895 ( .A1(n13452), .A2(n13453), .ZN(n13457) );
  NAND2_X1 U16896 ( .A1(n14064), .A2(n13453), .ZN(n13455) );
  NAND2_X1 U16897 ( .A1(n13368), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13454) );
  NAND3_X1 U16898 ( .A1(n13455), .A2(n13400), .A3(n13454), .ZN(n13456) );
  AND2_X1 U16899 ( .A1(n13457), .A2(n13456), .ZN(n15128) );
  OR2_X1 U16900 ( .A1(n13470), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U16901 ( .A1(n13400), .A2(n13508), .ZN(n13459) );
  INV_X1 U16902 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14745) );
  NAND2_X1 U16903 ( .A1(n14064), .A2(n14745), .ZN(n13458) );
  NAND3_X1 U16904 ( .A1(n13459), .A2(n13375), .A3(n13458), .ZN(n13460) );
  NAND2_X1 U16905 ( .A1(n13461), .A2(n13460), .ZN(n15129) );
  AND2_X1 U16906 ( .A1(n15128), .A2(n15129), .ZN(n13462) );
  OR2_X1 U16907 ( .A1(n13470), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13467) );
  INV_X1 U16908 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21717) );
  NAND2_X1 U16909 ( .A1(n13400), .A2(n21717), .ZN(n13465) );
  INV_X1 U16910 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U16911 ( .A1(n14064), .A2(n13463), .ZN(n13464) );
  NAND3_X1 U16912 ( .A1(n13465), .A2(n13375), .A3(n13464), .ZN(n13466) );
  AND2_X1 U16913 ( .A1(n13467), .A2(n13466), .ZN(n15112) );
  MUX2_X1 U16914 ( .A(n13468), .B(n13375), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13469) );
  OAI21_X1 U16915 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13870), .A(
        n13469), .ZN(n15103) );
  OR2_X1 U16916 ( .A1(n13470), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13475) );
  INV_X1 U16917 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15519) );
  NAND2_X1 U16918 ( .A1(n13400), .A2(n15519), .ZN(n13473) );
  INV_X1 U16919 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U16920 ( .A1(n14064), .A2(n13471), .ZN(n13472) );
  NAND3_X1 U16921 ( .A1(n13473), .A2(n13375), .A3(n13472), .ZN(n13474) );
  NAND2_X1 U16922 ( .A1(n13475), .A2(n13474), .ZN(n15084) );
  INV_X1 U16923 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13476) );
  NAND2_X1 U16924 ( .A1(n14064), .A2(n13476), .ZN(n13478) );
  OR2_X1 U16925 ( .A1(n13870), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13477) );
  NAND2_X1 U16926 ( .A1(n13477), .A2(n13478), .ZN(n15061) );
  MUX2_X1 U16927 ( .A(n13478), .B(n15061), .S(n13375), .Z(n14876) );
  AOI22_X1 U16928 ( .A1(n13870), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13819), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15063) );
  NAND2_X1 U16929 ( .A1(n15062), .A2(n15063), .ZN(n13479) );
  AOI22_X1 U16930 ( .A1(n13870), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13819), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13481) );
  OAI21_X1 U16931 ( .B1(n13363), .B2(n20804), .A(n17288), .ZN(n13483) );
  INV_X1 U16932 ( .A(n13870), .ZN(n13485) );
  OR2_X1 U16933 ( .A1(n13486), .A2(n13485), .ZN(n13492) );
  OR2_X1 U16934 ( .A1(n11958), .A2(n13487), .ZN(n13490) );
  INV_X1 U16935 ( .A(n15352), .ZN(n13489) );
  NAND2_X1 U16936 ( .A1(n14146), .A2(n14727), .ZN(n13488) );
  AOI22_X1 U16937 ( .A1(n13490), .A2(n13489), .B1(n13488), .B2(n20796), .ZN(
        n13491) );
  NAND2_X1 U16938 ( .A1(n11964), .A2(n11926), .ZN(n13493) );
  AND3_X1 U16939 ( .A1(n13499), .A2(n13494), .A3(n13493), .ZN(n13839) );
  OAI211_X1 U16940 ( .C1(n13484), .C2(n20776), .A(n13839), .B(n13495), .ZN(
        n13496) );
  NAND2_X1 U16941 ( .A1(n13502), .A2(n13496), .ZN(n15781) );
  INV_X1 U16942 ( .A(n15781), .ZN(n15894) );
  INV_X1 U16943 ( .A(n13497), .ZN(n13519) );
  INV_X1 U16944 ( .A(n20736), .ZN(n15840) );
  INV_X1 U16945 ( .A(n15743), .ZN(n13500) );
  NAND2_X1 U16946 ( .A1(n13500), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13518) );
  AND2_X1 U16947 ( .A1(n13744), .A2(n20792), .ZN(n14186) );
  NAND2_X1 U16948 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17323) );
  NOR2_X1 U16949 ( .A1(n17323), .A2(n12150), .ZN(n15867) );
  AND2_X1 U16950 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13501) );
  NAND2_X1 U16951 ( .A1(n15867), .A2(n13501), .ZN(n15838) );
  OR2_X1 U16952 ( .A1(n15838), .A2(n15861), .ZN(n15839) );
  NOR2_X1 U16953 ( .A1(n15839), .A2(n15852), .ZN(n13504) );
  INV_X1 U16954 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20716) );
  NOR2_X1 U16955 ( .A1(n20716), .A2(n12123), .ZN(n20715) );
  NAND2_X1 U16956 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20715), .ZN(
        n15851) );
  NAND2_X1 U16957 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17328) );
  NOR2_X1 U16958 ( .A1(n15851), .A2(n17328), .ZN(n15837) );
  NAND2_X1 U16959 ( .A1(n13504), .A2(n15837), .ZN(n15777) );
  NAND2_X1 U16960 ( .A1(n20735), .A2(n15777), .ZN(n13505) );
  OR2_X1 U16961 ( .A1(n13502), .A2(n20718), .ZN(n15895) );
  OR2_X1 U16962 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15781), .ZN(
        n13503) );
  AOI21_X1 U16963 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20720) );
  NOR2_X1 U16964 ( .A1(n15851), .A2(n20720), .ZN(n15842) );
  NAND2_X1 U16965 ( .A1(n15842), .A2(n13504), .ZN(n13511) );
  NAND2_X1 U16966 ( .A1(n20736), .A2(n13511), .ZN(n15784) );
  AND3_X1 U16967 ( .A1(n13505), .A2(n20750), .A3(n15784), .ZN(n13507) );
  AND2_X1 U16968 ( .A1(n15804), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15786) );
  NAND2_X1 U16969 ( .A1(n15786), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13517) );
  OR3_X1 U16970 ( .A1(n15833), .A2(n15820), .A3(n13517), .ZN(n13506) );
  AOI21_X1 U16971 ( .B1(n15894), .B2(n13519), .A(n13583), .ZN(n13510) );
  NAND2_X1 U16972 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13520) );
  INV_X1 U16973 ( .A(n15779), .ZN(n15896) );
  AOI22_X1 U16974 ( .A1(n15896), .A2(n15513), .B1(n20736), .B2(n13508), .ZN(
        n13509) );
  AOI211_X1 U16975 ( .C1(n13510), .C2(n17334), .A(n13338), .B(n15697), .ZN(
        n13523) );
  INV_X1 U16976 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21438) );
  NOR2_X1 U16977 ( .A1(n20576), .A2(n21438), .ZN(n15054) );
  INV_X1 U16978 ( .A(n13511), .ZN(n13512) );
  NAND2_X1 U16979 ( .A1(n20736), .A2(n13512), .ZN(n13515) );
  NOR2_X1 U16980 ( .A1(n15777), .A2(n20734), .ZN(n15780) );
  INV_X1 U16981 ( .A(n15780), .ZN(n13513) );
  OR2_X1 U16982 ( .A1(n15781), .A2(n13513), .ZN(n13514) );
  OAI21_X1 U16983 ( .B1(n15777), .B2(n15779), .A(n15785), .ZN(n15832) );
  AND2_X1 U16984 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13516) );
  NAND2_X1 U16985 ( .A1(n15832), .A2(n13516), .ZN(n15815) );
  NOR2_X1 U16986 ( .A1(n14820), .A2(n13519), .ZN(n15723) );
  INV_X1 U16987 ( .A(n13520), .ZN(n13521) );
  NAND3_X1 U16988 ( .A1(n15714), .A2(n15706), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15698) );
  NOR3_X1 U16989 ( .A1(n15698), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15699), .ZN(n13522) );
  INV_X1 U16990 ( .A(n17087), .ZN(n17052) );
  NAND2_X1 U16991 ( .A1(n17101), .A2(n18703), .ZN(n14686) );
  NAND2_X1 U16992 ( .A1(n13526), .A2(n13525), .ZN(n14685) );
  AOI21_X2 U16993 ( .B1(n14686), .B2(n13524), .A(n14685), .ZN(n14708) );
  OAI211_X1 U16994 ( .C1(n17101), .C2(n13534), .A(n19464), .B(n14692), .ZN(
        n13527) );
  NOR2_X1 U16995 ( .A1(n14708), .A2(n13527), .ZN(n13532) );
  NAND2_X1 U16996 ( .A1(n17096), .A2(n18996), .ZN(n13530) );
  INV_X1 U16997 ( .A(n13528), .ZN(n13529) );
  INV_X1 U16998 ( .A(n18981), .ZN(n18845) );
  NAND2_X1 U16999 ( .A1(n18845), .A2(n18889), .ZN(n18968) );
  NAND2_X1 U17000 ( .A1(n18968), .A2(n14698), .ZN(n17198) );
  NAND3_X1 U17001 ( .A1(n13530), .A2(n13529), .A3(n17198), .ZN(n13531) );
  NOR3_X1 U17002 ( .A1(n13533), .A2(n9696), .A3(n21581), .ZN(n13551) );
  INV_X1 U17003 ( .A(n13524), .ZN(n13536) );
  NOR3_X1 U17004 ( .A1(n14708), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n13534), .ZN(n13535) );
  AOI21_X1 U17005 ( .B1(n13536), .B2(n14685), .A(n13535), .ZN(n13549) );
  INV_X1 U17006 ( .A(n19465), .ZN(n18933) );
  OR2_X1 U17007 ( .A1(n13537), .A2(n18933), .ZN(n13539) );
  INV_X1 U17008 ( .A(n18996), .ZN(n18931) );
  OR2_X1 U17009 ( .A1(n18956), .A2(n18931), .ZN(n13538) );
  NAND2_X1 U17010 ( .A1(n13539), .A2(n13538), .ZN(n18944) );
  AND2_X1 U17011 ( .A1(n18888), .A2(n17229), .ZN(n13544) );
  NAND2_X1 U17012 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18846), .ZN(
        n17227) );
  NOR3_X1 U17013 ( .A1(n17239), .A2(n14090), .A3(n17227), .ZN(n13542) );
  INV_X1 U17014 ( .A(n13540), .ZN(n13541) );
  OR2_X1 U17015 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  AOI21_X1 U17016 ( .B1(n18944), .B2(n13544), .A(n13543), .ZN(n18841) );
  OR2_X1 U17017 ( .A1(n18841), .A2(n18573), .ZN(n18797) );
  NAND2_X1 U17018 ( .A1(n13545), .A2(n21581), .ZN(n13546) );
  NOR2_X1 U17019 ( .A1(n18797), .A2(n13546), .ZN(n13547) );
  AOI21_X1 U17020 ( .B1(n9739), .B2(n16506), .A(n16508), .ZN(n13554) );
  INV_X1 U17021 ( .A(n13552), .ZN(n13553) );
  XNOR2_X1 U17022 ( .A(n13554), .B(n13553), .ZN(n13571) );
  AND2_X1 U17023 ( .A1(n13556), .A2(n13557), .ZN(n13558) );
  NOR2_X1 U17024 ( .A1(n13555), .A2(n13558), .ZN(n16390) );
  INV_X1 U17025 ( .A(n13559), .ZN(n15941) );
  NAND2_X1 U17026 ( .A1(n13560), .A2(n13561), .ZN(n13562) );
  NAND2_X1 U17027 ( .A1(n15941), .A2(n13562), .ZN(n16304) );
  INV_X1 U17028 ( .A(n16719), .ZN(n13565) );
  OAI21_X1 U17029 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16705), .ZN(n13563) );
  OR2_X1 U17030 ( .A1(n11468), .A2(n20452), .ZN(n13573) );
  OAI21_X1 U17031 ( .B1(n16718), .B2(n13563), .A(n13573), .ZN(n13564) );
  AOI21_X1 U17032 ( .B1(n13565), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13564), .ZN(n13566) );
  OAI21_X1 U17033 ( .B1(n16304), .B2(n19803), .A(n13566), .ZN(n13567) );
  AOI21_X1 U17034 ( .B1(n16390), .B2(n19792), .A(n13567), .ZN(n13570) );
  INV_X1 U17035 ( .A(n13568), .ZN(n16500) );
  NAND3_X1 U17036 ( .A1(n10389), .A2(n13570), .A3(n13569), .ZN(P2_U3020) );
  NOR2_X1 U17037 ( .A1(n13571), .A2(n19785), .ZN(n13579) );
  INV_X1 U17038 ( .A(n16304), .ZN(n13576) );
  INV_X1 U17039 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15956) );
  INV_X1 U17040 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U17041 ( .A1(n15023), .A2(n15956), .ZN(n13572) );
  NAND2_X1 U17042 ( .A1(n19771), .A2(n10421), .ZN(n13574) );
  OAI211_X1 U17043 ( .C1(n17388), .C2(n15956), .A(n13574), .B(n13573), .ZN(
        n13575) );
  INV_X1 U17044 ( .A(n13577), .ZN(n13578) );
  NAND2_X1 U17045 ( .A1(n14713), .A2(n20738), .ZN(n13590) );
  XNOR2_X1 U17046 ( .A(n15130), .B(n15129), .ZN(n14726) );
  NAND2_X1 U17047 ( .A1(n15779), .A2(n20734), .ZN(n20756) );
  NAND2_X1 U17048 ( .A1(n20735), .A2(n20756), .ZN(n20743) );
  INV_X1 U17049 ( .A(n13583), .ZN(n13584) );
  OAI21_X1 U17050 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20743), .A(
        n13584), .ZN(n13586) );
  INV_X1 U17051 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21426) );
  NOR2_X1 U17052 ( .A1(n20576), .A2(n21426), .ZN(n14715) );
  NOR3_X1 U17053 ( .A1(n14820), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14824), .ZN(n13585) );
  AOI211_X1 U17054 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n13586), .A(
        n14715), .B(n13585), .ZN(n13587) );
  INV_X1 U17055 ( .A(n13588), .ZN(n13589) );
  NAND2_X1 U17056 ( .A1(n13590), .A2(n13589), .ZN(P1_U3007) );
  INV_X1 U17057 ( .A(n15706), .ZN(n15502) );
  NAND2_X1 U17058 ( .A1(n15528), .A2(n15706), .ZN(n13591) );
  OAI21_X1 U17059 ( .B1(n15506), .B2(n15641), .A(n13591), .ZN(n13594) );
  NOR2_X1 U17060 ( .A1(n15641), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15505) );
  INV_X1 U17061 ( .A(n15505), .ZN(n13592) );
  NAND2_X1 U17062 ( .A1(n15657), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15503) );
  NAND2_X1 U17063 ( .A1(n13592), .A2(n15503), .ZN(n13593) );
  XNOR2_X1 U17064 ( .A(n13594), .B(n13593), .ZN(n14885) );
  NOR2_X2 U17065 ( .A1(n13596), .A2(n13595), .ZN(n13656) );
  INV_X1 U17066 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15534) );
  OR2_X2 U17067 ( .A1(n13660), .A2(n15534), .ZN(n13674) );
  OR2_X2 U17068 ( .A1(n13674), .A2(n13673), .ZN(n13676) );
  XNOR2_X1 U17069 ( .A(n14723), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15078) );
  INV_X1 U17070 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U17071 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U17072 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U17073 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U17074 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13597) );
  NAND4_X1 U17075 ( .A1(n13600), .A2(n13599), .A3(n13598), .A4(n13597), .ZN(
        n13606) );
  AOI22_X1 U17076 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U17077 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13603) );
  AOI22_X1 U17078 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13602) );
  AOI22_X1 U17079 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13601) );
  NAND4_X1 U17080 ( .A1(n13604), .A2(n13603), .A3(n13602), .A4(n13601), .ZN(
        n13605) );
  NOR2_X1 U17081 ( .A1(n13606), .A2(n13605), .ZN(n13648) );
  NOR2_X1 U17082 ( .A1(n13608), .A2(n13607), .ZN(n13662) );
  AOI22_X1 U17083 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U17084 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U17085 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U17086 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13611) );
  NAND4_X1 U17087 ( .A1(n13614), .A2(n13613), .A3(n13612), .A4(n13611), .ZN(
        n13621) );
  AOI22_X1 U17088 ( .A1(n13615), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U17089 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U17090 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U17091 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13616) );
  NAND4_X1 U17092 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13620) );
  OR2_X1 U17093 ( .A1(n13621), .A2(n13620), .ZN(n13661) );
  NAND2_X1 U17094 ( .A1(n13662), .A2(n13661), .ZN(n13649) );
  NOR2_X1 U17095 ( .A1(n13648), .A2(n13649), .ZN(n13679) );
  AOI22_X1 U17096 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13625) );
  AOI22_X1 U17097 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U17098 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U17099 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11912), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13622) );
  NAND4_X1 U17100 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n13631) );
  AOI22_X1 U17101 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14774), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13629) );
  AOI22_X1 U17102 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U17103 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13627) );
  AOI22_X1 U17104 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13626) );
  NAND4_X1 U17105 ( .A1(n13629), .A2(n13628), .A3(n13627), .A4(n13626), .ZN(
        n13630) );
  OR2_X1 U17106 ( .A1(n13631), .A2(n13630), .ZN(n13677) );
  NAND2_X1 U17107 ( .A1(n13679), .A2(n13677), .ZN(n14791) );
  AOI22_X1 U17108 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13637) );
  AOI22_X1 U17109 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13633), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U17110 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13635) );
  AOI22_X1 U17111 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11912), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13634) );
  NAND4_X1 U17112 ( .A1(n13637), .A2(n13636), .A3(n13635), .A4(n13634), .ZN(
        n13643) );
  AOI22_X1 U17113 ( .A1(n14782), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13641) );
  AOI22_X1 U17114 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U17115 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13639) );
  AOI22_X1 U17116 ( .A1(n14775), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13638) );
  NAND4_X1 U17117 ( .A1(n13641), .A2(n13640), .A3(n13639), .A4(n13638), .ZN(
        n13642) );
  NOR2_X1 U17118 ( .A1(n13643), .A2(n13642), .ZN(n14792) );
  XOR2_X1 U17119 ( .A(n14791), .B(n14792), .Z(n13644) );
  NAND2_X1 U17120 ( .A1(n13644), .A2(n14799), .ZN(n13646) );
  OAI21_X1 U17121 ( .B1(n20830), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n21306), .ZN(n13645) );
  OAI211_X1 U17122 ( .C1(n14797), .C2(n15408), .A(n13646), .B(n13645), .ZN(
        n13647) );
  OAI21_X1 U17123 ( .B1(n15078), .B2(n14796), .A(n13647), .ZN(n13687) );
  XNOR2_X1 U17124 ( .A(n13660), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15532) );
  NAND2_X1 U17125 ( .A1(n15532), .A2(n14802), .ZN(n13655) );
  XOR2_X1 U17126 ( .A(n13649), .B(n13648), .Z(n13650) );
  NAND2_X1 U17127 ( .A1(n13650), .A2(n14799), .ZN(n13653) );
  AOI21_X1 U17128 ( .B1(n15534), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13651) );
  AOI21_X1 U17129 ( .B1(n12320), .B2(P1_EAX_REG_27__SCAN_IN), .A(n13651), .ZN(
        n13652) );
  NAND2_X1 U17130 ( .A1(n13653), .A2(n13652), .ZN(n13654) );
  NAND2_X1 U17131 ( .A1(n13655), .A2(n13654), .ZN(n15096) );
  INV_X1 U17132 ( .A(n15096), .ZN(n13672) );
  INV_X1 U17133 ( .A(n13656), .ZN(n13658) );
  INV_X1 U17134 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13657) );
  NAND2_X1 U17135 ( .A1(n13658), .A2(n13657), .ZN(n13659) );
  NAND2_X1 U17136 ( .A1(n13660), .A2(n13659), .ZN(n15542) );
  OR2_X1 U17137 ( .A1(n15542), .A2(n14796), .ZN(n13669) );
  XNOR2_X1 U17138 ( .A(n13662), .B(n13661), .ZN(n13667) );
  NAND2_X1 U17139 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13663) );
  NAND2_X1 U17140 ( .A1(n14796), .A2(n13663), .ZN(n13664) );
  AOI21_X1 U17141 ( .B1(n12320), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13664), .ZN(
        n13665) );
  OAI21_X1 U17142 ( .B1(n13667), .B2(n13666), .A(n13665), .ZN(n13668) );
  NAND2_X1 U17143 ( .A1(n13669), .A2(n13668), .ZN(n15109) );
  INV_X1 U17144 ( .A(n15109), .ZN(n13670) );
  NAND2_X1 U17145 ( .A1(n13674), .A2(n13673), .ZN(n13675) );
  AND2_X1 U17146 ( .A1(n13676), .A2(n13675), .ZN(n15521) );
  INV_X1 U17147 ( .A(n13677), .ZN(n13678) );
  XNOR2_X1 U17148 ( .A(n13679), .B(n13678), .ZN(n13682) );
  INV_X1 U17149 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15413) );
  NAND2_X1 U17150 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13680) );
  OAI211_X1 U17151 ( .C1(n14797), .C2(n15413), .A(n14796), .B(n13680), .ZN(
        n13681) );
  AOI21_X1 U17152 ( .B1(n13682), .B2(n14799), .A(n13681), .ZN(n13683) );
  AOI21_X1 U17153 ( .B1(n15521), .B2(n14802), .A(n13683), .ZN(n15083) );
  NAND2_X1 U17154 ( .A1(n15154), .A2(n13684), .ZN(n15082) );
  INV_X1 U17155 ( .A(n13684), .ZN(n13685) );
  NOR2_X1 U17156 ( .A1(n13687), .A2(n13685), .ZN(n13686) );
  AOI21_X1 U17157 ( .B1(n13687), .B2(n15082), .A(n14951), .ZN(n15072) );
  INV_X1 U17158 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21434) );
  NOR2_X1 U17159 ( .A1(n20576), .A2(n21434), .ZN(n14878) );
  AOI21_X1 U17160 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14878), .ZN(n13688) );
  OAI21_X1 U17161 ( .B1(n15078), .B2(n20714), .A(n13688), .ZN(n13689) );
  AOI21_X1 U17162 ( .B1(n15072), .B2(n20709), .A(n13689), .ZN(n13690) );
  OAI21_X1 U17163 ( .B1(n14885), .B2(n20537), .A(n13690), .ZN(P1_U2970) );
  NOR2_X1 U17164 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n20499), .ZN(n13692) );
  NOR4_X1 U17165 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13691) );
  NAND4_X1 U17166 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13692), .A3(n13691), .A4(
        n21773), .ZN(n13714) );
  NOR2_X4 U17167 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13714), .ZN(n17471)
         );
  INV_X2 U17168 ( .A(n17471), .ZN(U215) );
  NOR2_X1 U17169 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21511) );
  NOR3_X1 U17170 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13695) );
  NOR4_X1 U17171 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13694) );
  NOR4_X1 U17172 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13693) );
  AND4_X1 U17173 ( .A1(n21511), .A2(n13695), .A3(n13694), .A4(n13693), .ZN(
        n13701) );
  NOR4_X1 U17174 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_16__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13699) );
  NOR4_X1 U17175 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13698) );
  NOR4_X1 U17176 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13697) );
  NOR4_X1 U17177 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n13696) );
  AND4_X1 U17178 ( .A1(n13699), .A2(n13698), .A3(n13697), .A4(n13696), .ZN(
        n13700) );
  NAND2_X1 U17179 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  NAND4_X1 U17180 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(n21789), .A3(n21549), .A4(
        n21567), .ZN(n13703) );
  NOR4_X1 U17181 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13708) );
  NOR4_X1 U17182 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13707) );
  NOR4_X1 U17183 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13706) );
  NOR4_X1 U17184 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13705) );
  NAND4_X1 U17185 ( .A1(n13708), .A2(n13707), .A3(n13706), .A4(n13705), .ZN(
        n13713) );
  NOR2_X1 U17186 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21512) );
  NOR3_X1 U17187 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n13711) );
  NOR4_X1 U17188 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13710) );
  NOR4_X1 U17189 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13709) );
  NAND4_X1 U17190 ( .A1(n21512), .A2(n13711), .A3(n13710), .A4(n13709), .ZN(
        n13712) );
  NOR3_X1 U17191 ( .A1(n20520), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n17044), 
        .ZN(n17041) );
  INV_X1 U17192 ( .A(n16978), .ZN(n13715) );
  NAND2_X1 U17193 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13715), .ZN(n14611) );
  INV_X1 U17194 ( .A(n14611), .ZN(n16980) );
  NOR2_X1 U17195 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13717) );
  NOR3_X1 U17196 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n13716) );
  NOR4_X1 U17197 ( .A1(n17041), .A2(n16980), .A3(n13717), .A4(n13716), .ZN(
        P2_U3178) );
  NAND2_X1 U17198 ( .A1(n13774), .A2(n13721), .ZN(n16279) );
  INV_X1 U17199 ( .A(n16279), .ZN(n13720) );
  INV_X1 U17200 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20528) );
  INV_X1 U17201 ( .A(n13721), .ZN(n13719) );
  OAI211_X1 U17202 ( .C1(n13720), .C2(n20528), .A(n13722), .B(n15032), .ZN(
        P2_U2814) );
  INV_X1 U17203 ( .A(n15042), .ZN(n20521) );
  INV_X1 U17204 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19644) );
  OAI22_X1 U17205 ( .A1(n20521), .A2(n19644), .B1(n17044), .B2(n13722), .ZN(
        P2_U2816) );
  INV_X1 U17206 ( .A(n13722), .ZN(n13723) );
  OAI21_X1 U17207 ( .B1(n13723), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n15042), 
        .ZN(n13724) );
  OAI21_X1 U17208 ( .B1(n13725), .B2(n15042), .A(n13724), .ZN(P2_U3612) );
  AND2_X1 U17209 ( .A1(n13726), .A2(n20520), .ZN(n13757) );
  NOR2_X1 U17210 ( .A1(n13757), .A2(n14445), .ZN(n13727) );
  NAND3_X1 U17211 ( .A1(n14493), .A2(n13758), .A3(n13727), .ZN(n14504) );
  NAND2_X1 U17212 ( .A1(n14504), .A2(n17047), .ZN(n20507) );
  INV_X1 U17213 ( .A(n20507), .ZN(n13729) );
  OAI21_X1 U17214 ( .B1(n13729), .B2(n13766), .A(n13728), .ZN(P2_U2819) );
  NAND2_X1 U17215 ( .A1(n13824), .A2(n14141), .ZN(n13753) );
  AND2_X1 U17216 ( .A1(n9694), .A2(n17370), .ZN(n20530) );
  AOI21_X1 U17217 ( .B1(n13753), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n20530), 
        .ZN(n13731) );
  NAND2_X1 U17218 ( .A1(n14231), .A2(n13731), .ZN(P1_U2801) );
  INV_X1 U17219 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16264) );
  AOI21_X1 U17220 ( .B1(n13733), .B2(n16963), .A(n13732), .ZN(n16968) );
  NOR2_X1 U17221 ( .A1(n11468), .A2(n20412), .ZN(n16965) );
  XNOR2_X1 U17222 ( .A(n17394), .B(n16963), .ZN(n13734) );
  XNOR2_X1 U17223 ( .A(n13734), .B(n16258), .ZN(n16962) );
  OAI22_X1 U17224 ( .A1(n19785), .A2(n16962), .B1(n17388), .B2(n16264), .ZN(
        n13735) );
  AOI211_X1 U17225 ( .C1(n19781), .C2(n16968), .A(n16965), .B(n13735), .ZN(
        n13737) );
  NAND2_X1 U17226 ( .A1(n16966), .A2(n19787), .ZN(n13736) );
  OAI211_X1 U17227 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19758), .A(
        n13737), .B(n13736), .ZN(P2_U3013) );
  NAND2_X1 U17228 ( .A1(n17295), .A2(n15351), .ZN(n13739) );
  OR2_X1 U17229 ( .A1(n13824), .A2(n13730), .ZN(n13738) );
  NAND2_X1 U17230 ( .A1(n13739), .A2(n13738), .ZN(n20532) );
  NAND3_X1 U17231 ( .A1(n15351), .A2(n13819), .A3(n17306), .ZN(n13740) );
  AND2_X1 U17232 ( .A1(n13740), .A2(n21487), .ZN(n21488) );
  NOR2_X1 U17233 ( .A1(n20532), .A2(n21488), .ZN(n17278) );
  OR2_X1 U17234 ( .A1(n17278), .A2(n20531), .ZN(n13750) );
  INV_X1 U17235 ( .A(n13750), .ZN(n20539) );
  INV_X1 U17236 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13752) );
  INV_X1 U17237 ( .A(n13873), .ZN(n13845) );
  AND2_X1 U17238 ( .A1(n13742), .A2(n13741), .ZN(n13743) );
  MUX2_X1 U17239 ( .A(n13845), .B(n13743), .S(n17295), .Z(n13748) );
  INV_X1 U17240 ( .A(n13744), .ZN(n13745) );
  OR2_X1 U17241 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  NAND2_X1 U17242 ( .A1(n13748), .A2(n13747), .ZN(n13749) );
  NAND2_X1 U17243 ( .A1(n13749), .A2(n20818), .ZN(n17280) );
  OR2_X1 U17244 ( .A1(n13750), .A2(n17280), .ZN(n13751) );
  OAI21_X1 U17245 ( .B1(n20539), .B2(n13752), .A(n13751), .ZN(P1_U3484) );
  NOR2_X1 U17246 ( .A1(n11926), .A2(n11939), .ZN(n13755) );
  NOR3_X1 U17247 ( .A1(n21485), .A2(n20530), .A3(P1_READREQUEST_REG_SCAN_IN), 
        .ZN(n13754) );
  AOI21_X1 U17248 ( .B1(n13755), .B2(n21485), .A(n13754), .ZN(P1_U3487) );
  NAND3_X1 U17249 ( .A1(n14493), .A2(n13758), .A3(n13757), .ZN(n13759) );
  NAND2_X1 U17250 ( .A1(n13761), .A2(n13760), .ZN(n13762) );
  NOR2_X1 U17251 ( .A1(n14521), .A2(n13762), .ZN(n13764) );
  NAND3_X1 U17252 ( .A1(n13775), .A2(n13774), .A3(n14445), .ZN(n13763) );
  NAND2_X1 U17253 ( .A1(n17044), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13765) );
  AND2_X1 U17254 ( .A1(n13765), .A2(n14611), .ZN(n14515) );
  AOI21_X1 U17255 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n13766), .A(n14515), 
        .ZN(n13767) );
  INV_X1 U17256 ( .A(n17020), .ZN(n13773) );
  AND2_X1 U17257 ( .A1(n13769), .A2(n13768), .ZN(n14501) );
  INV_X1 U17258 ( .A(n13770), .ZN(n14500) );
  NAND4_X1 U17259 ( .A1(n13773), .A2(n14501), .A3(n14500), .A4(n17009), .ZN(
        n13771) );
  OAI21_X1 U17260 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(P2_U3595) );
  INV_X1 U17261 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13780) );
  NAND3_X1 U17262 ( .A1(n13775), .A2(n17047), .A3(n13774), .ZN(n13776) );
  NAND2_X1 U17263 ( .A1(n13776), .A2(n15037), .ZN(n13778) );
  INV_X1 U17264 ( .A(n20513), .ZN(n13777) );
  NOR2_X4 U17265 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16978), .ZN(n19744) );
  AOI22_X1 U17266 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n19739), .B1(n19744), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13779) );
  OAI21_X1 U17267 ( .B1(n13780), .B2(n13809), .A(n13779), .ZN(P2_U2926) );
  INV_X1 U17268 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U17269 ( .A1(n19744), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13781) );
  OAI21_X1 U17270 ( .B1(n14012), .B2(n13809), .A(n13781), .ZN(P2_U2935) );
  INV_X1 U17271 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U17272 ( .A1(n19744), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13782) );
  OAI21_X1 U17273 ( .B1(n13783), .B2(n13809), .A(n13782), .ZN(P2_U2932) );
  INV_X1 U17274 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13785) );
  AOI22_X1 U17275 ( .A1(n19744), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13784) );
  OAI21_X1 U17276 ( .B1(n13785), .B2(n13809), .A(n13784), .ZN(P2_U2934) );
  INV_X1 U17277 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U17278 ( .A1(n19744), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13786) );
  OAI21_X1 U17279 ( .B1(n13787), .B2(n13809), .A(n13786), .ZN(P2_U2930) );
  INV_X1 U17280 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U17281 ( .A1(n19744), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13788) );
  OAI21_X1 U17282 ( .B1(n13789), .B2(n13809), .A(n13788), .ZN(P2_U2933) );
  NOR2_X1 U17283 ( .A1(n16350), .A2(n13792), .ZN(n13793) );
  AOI21_X1 U17284 ( .B1(n16350), .B2(n16966), .A(n13793), .ZN(n13794) );
  OAI21_X1 U17285 ( .B1(n19957), .B2(n16353), .A(n13794), .ZN(P2_U2886) );
  INV_X1 U17286 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U17287 ( .A1(n19744), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13795) );
  OAI21_X1 U17288 ( .B1(n13967), .B2(n13809), .A(n13795), .ZN(P2_U2921) );
  INV_X1 U17289 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13797) );
  AOI22_X1 U17290 ( .A1(n19744), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13796) );
  OAI21_X1 U17291 ( .B1(n13797), .B2(n13809), .A(n13796), .ZN(P2_U2931) );
  INV_X1 U17292 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U17293 ( .A1(n19744), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13798) );
  OAI21_X1 U17294 ( .B1(n14023), .B2(n13809), .A(n13798), .ZN(P2_U2925) );
  INV_X1 U17295 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U17296 ( .A1(n19744), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13799) );
  OAI21_X1 U17297 ( .B1(n13800), .B2(n13809), .A(n13799), .ZN(P2_U2923) );
  INV_X1 U17298 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U17299 ( .A1(n19744), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U17300 ( .B1(n13802), .B2(n13809), .A(n13801), .ZN(P2_U2929) );
  INV_X1 U17301 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U17302 ( .A1(n19744), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13803) );
  OAI21_X1 U17303 ( .B1(n13804), .B2(n13809), .A(n13803), .ZN(P2_U2928) );
  INV_X1 U17304 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14027) );
  AOI22_X1 U17305 ( .A1(n19744), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13805) );
  OAI21_X1 U17306 ( .B1(n14027), .B2(n13809), .A(n13805), .ZN(P2_U2927) );
  INV_X1 U17307 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U17308 ( .A1(n19744), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13806) );
  OAI21_X1 U17309 ( .B1(n13807), .B2(n13809), .A(n13806), .ZN(P2_U2922) );
  INV_X1 U17310 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U17311 ( .A1(n19744), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13808) );
  OAI21_X1 U17312 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(P2_U2924) );
  AOI21_X1 U17313 ( .B1(n11127), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13811) );
  AND2_X1 U17314 ( .A1(n13812), .A2(n13811), .ZN(n13813) );
  NOR2_X1 U17315 ( .A1(n16360), .A2(n17401), .ZN(n13815) );
  AOI21_X1 U17316 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n16360), .A(n13815), .ZN(
        n13816) );
  OAI21_X1 U17317 ( .B1(n16353), .B2(n20090), .A(n13816), .ZN(P2_U2887) );
  INV_X1 U17318 ( .A(n13820), .ZN(n13817) );
  OAI211_X1 U17319 ( .C1(n14186), .C2(n13817), .A(n17290), .B(n21487), .ZN(
        n13818) );
  MUX2_X1 U17320 ( .A(n13818), .B(n13845), .S(n17295), .Z(n13830) );
  NAND3_X1 U17321 ( .A1(n13824), .A2(n13823), .A3(n21487), .ZN(n13825) );
  OR2_X1 U17322 ( .A1(n15352), .A2(n20796), .ZN(n13827) );
  AND2_X1 U17323 ( .A1(n13828), .A2(n13827), .ZN(n13829) );
  NAND3_X1 U17324 ( .A1(n13830), .A2(n14140), .A3(n13829), .ZN(n17265) );
  NAND2_X1 U17325 ( .A1(n17265), .A2(n14141), .ZN(n13834) );
  INV_X1 U17326 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20538) );
  NAND2_X1 U17327 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17366), .ZN(n17372) );
  OR2_X1 U17328 ( .A1(n20538), .A2(n17372), .ZN(n13832) );
  NAND2_X1 U17329 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21369), .ZN(n13831) );
  AND2_X1 U17330 ( .A1(n13832), .A2(n13831), .ZN(n13833) );
  NAND2_X1 U17331 ( .A1(n21457), .A2(n14944), .ZN(n21459) );
  INV_X1 U17332 ( .A(n21459), .ZN(n14947) );
  INV_X1 U17333 ( .A(n13838), .ZN(n14198) );
  INV_X1 U17334 ( .A(n20939), .ZN(n21201) );
  OR2_X1 U17335 ( .A1(n12026), .A2(n21201), .ZN(n13835) );
  XNOR2_X1 U17336 ( .A(n13835), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20599) );
  NAND3_X1 U17337 ( .A1(n14947), .A2(n14198), .A3(n20599), .ZN(n13836) );
  OAI21_X1 U17338 ( .B1(n12312), .B2(n21457), .A(n13836), .ZN(P1_U3468) );
  AND2_X1 U17339 ( .A1(n13484), .A2(n20808), .ZN(n13837) );
  AND2_X1 U17340 ( .A1(n13838), .A2(n13837), .ZN(n13840) );
  NAND2_X1 U17341 ( .A1(n13840), .A2(n13839), .ZN(n14191) );
  INV_X1 U17342 ( .A(n13841), .ZN(n13842) );
  NAND2_X1 U17343 ( .A1(n13842), .A2(n13852), .ZN(n14178) );
  NAND2_X1 U17344 ( .A1(n13841), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14176) );
  NAND2_X1 U17345 ( .A1(n14178), .A2(n14176), .ZN(n13847) );
  INV_X1 U17346 ( .A(n13847), .ZN(n13854) );
  NAND2_X1 U17347 ( .A1(n11958), .A2(n13854), .ZN(n13850) );
  INV_X1 U17348 ( .A(n14191), .ZN(n14945) );
  OR2_X1 U17349 ( .A1(n13843), .A2(n14945), .ZN(n13849) );
  NAND2_X1 U17350 ( .A1(n13845), .A2(n13844), .ZN(n14180) );
  XNOR2_X1 U17351 ( .A(n11997), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13846) );
  AOI22_X1 U17352 ( .A1(n14180), .A2(n13847), .B1(n14186), .B2(n13846), .ZN(
        n13848) );
  OAI211_X1 U17353 ( .C1(n14191), .C2(n13850), .A(n13849), .B(n13848), .ZN(
        n14193) );
  INV_X1 U17354 ( .A(n14193), .ZN(n13856) );
  INV_X1 U17355 ( .A(n21457), .ZN(n14942) );
  NOR2_X1 U17356 ( .A1(n14942), .A2(n21454), .ZN(n14948) );
  NOR2_X1 U17357 ( .A1(n17370), .A2(n20734), .ZN(n13865) );
  AOI22_X1 U17358 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20767), .B2(n13338), .ZN(
        n13863) );
  NAND3_X1 U17359 ( .A1(n21457), .A2(n13865), .A3(n13863), .ZN(n13851) );
  OAI21_X1 U17360 ( .B1(n21457), .B2(n13852), .A(n13851), .ZN(n13853) );
  AOI21_X1 U17361 ( .B1(n14948), .B2(n13854), .A(n13853), .ZN(n13855) );
  OAI21_X1 U17362 ( .B1(n13856), .B2(n21459), .A(n13855), .ZN(P1_U3472) );
  OR2_X1 U17363 ( .A1(n13858), .A2(n14945), .ZN(n13862) );
  NOR2_X1 U17364 ( .A1(n13859), .A2(n13841), .ZN(n13868) );
  AOI22_X1 U17365 ( .A1(n14186), .A2(n11997), .B1(n13868), .B2(n13860), .ZN(
        n13861) );
  AND2_X1 U17366 ( .A1(n13862), .A2(n13861), .ZN(n17264) );
  INV_X1 U17367 ( .A(n13863), .ZN(n13864) );
  NAND3_X1 U17368 ( .A1(n21457), .A2(n13865), .A3(n13864), .ZN(n13866) );
  OAI21_X1 U17369 ( .B1(n21457), .B2(n11997), .A(n13866), .ZN(n13867) );
  AOI21_X1 U17370 ( .B1(n14948), .B2(n13868), .A(n13867), .ZN(n13869) );
  OAI21_X1 U17371 ( .B1(n17264), .B2(n21459), .A(n13869), .ZN(P1_U3473) );
  OR2_X1 U17372 ( .A1(n13870), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13872) );
  NAND2_X1 U17373 ( .A1(n13872), .A2(n13871), .ZN(n15891) );
  NAND2_X1 U17374 ( .A1(n17295), .A2(n13873), .ZN(n13877) );
  AND4_X1 U17375 ( .A1(n14956), .A2(n14143), .A3(n13874), .A4(n20812), .ZN(
        n13875) );
  NAND2_X1 U17376 ( .A1(n14138), .A2(n14064), .ZN(n13876) );
  NAND2_X1 U17377 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  INV_X1 U17378 ( .A(n13879), .ZN(n13882) );
  OAI21_X1 U17379 ( .B1(n13882), .B2(n13881), .A(n13880), .ZN(n15367) );
  INV_X2 U17380 ( .A(n20649), .ZN(n15399) );
  OAI222_X1 U17381 ( .A1(n15891), .A2(n15395), .B1(n13883), .B2(n20653), .C1(
        n15367), .C2(n15399), .ZN(P1_U2872) );
  NOR2_X1 U17382 ( .A1(n13884), .A2(n13906), .ZN(n17849) );
  INV_X1 U17383 ( .A(n18978), .ZN(n18961) );
  NAND2_X1 U17384 ( .A1(n18961), .A2(n13885), .ZN(n13901) );
  AOI21_X1 U17385 ( .B1(n18978), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13886), .ZN(n13912) );
  NAND2_X1 U17386 ( .A1(n13912), .A2(n13887), .ZN(n13927) );
  AOI22_X1 U17387 ( .A1(n17849), .A2(n13901), .B1(n13927), .B2(n13888), .ZN(
        n19481) );
  INV_X1 U17388 ( .A(n19481), .ZN(n13889) );
  INV_X1 U17389 ( .A(n17869), .ZN(n13932) );
  AOI22_X1 U17390 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13253), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13310), .ZN(n13917) );
  NOR2_X1 U17391 ( .A1(n18425), .A2(n10151), .ZN(n13919) );
  AOI222_X1 U17392 ( .A1(n13889), .A2(n13932), .B1(n13917), .B2(n13919), .C1(
        n19506), .C2(n17849), .ZN(n13900) );
  NAND2_X1 U17393 ( .A1(n19466), .A2(n13890), .ZN(n14212) );
  INV_X1 U17394 ( .A(n19469), .ZN(n14688) );
  NAND3_X1 U17395 ( .A1(n19473), .A2(n18426), .A3(n19627), .ZN(n13893) );
  AND3_X1 U17396 ( .A1(n13894), .A2(n14212), .A3(n13893), .ZN(n13895) );
  NAND2_X1 U17397 ( .A1(n14216), .A2(n13895), .ZN(n19490) );
  NAND2_X1 U17398 ( .A1(n19490), .A2(n19509), .ZN(n13898) );
  INV_X1 U17399 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19021) );
  NAND2_X1 U17400 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19621), .ZN(n19606) );
  NOR2_X1 U17401 ( .A1(n19021), .A2(n19606), .ZN(n13896) );
  NOR2_X1 U17402 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19608), .ZN(n19034) );
  NOR2_X1 U17403 ( .A1(n13896), .A2(n19034), .ZN(n13897) );
  NAND2_X1 U17404 ( .A1(n14677), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13899) );
  OAI21_X1 U17405 ( .B1(n13900), .B2(n14677), .A(n13899), .ZN(P3_U3289) );
  MUX2_X1 U17406 ( .A(n13901), .B(n18981), .S(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n19479) );
  INV_X1 U17407 ( .A(n19506), .ZN(n13902) );
  OAI22_X1 U17408 ( .A1(n13902), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18425), .ZN(n13903) );
  AOI21_X1 U17409 ( .B1(n19479), .B2(n13932), .A(n13903), .ZN(n13905) );
  NAND2_X1 U17410 ( .A1(n14677), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13904) );
  OAI21_X1 U17411 ( .B1(n13905), .B2(n14677), .A(n13904), .ZN(P3_U3290) );
  INV_X1 U17412 ( .A(n13906), .ZN(n13911) );
  NAND2_X1 U17413 ( .A1(n13911), .A2(n13907), .ZN(n13925) );
  NAND2_X1 U17414 ( .A1(n13926), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13930) );
  AND2_X1 U17415 ( .A1(n13925), .A2(n13930), .ZN(n17835) );
  OAI21_X1 U17416 ( .B1(n13910), .B2(n13909), .A(n13908), .ZN(n13923) );
  NAND3_X1 U17417 ( .A1(n13923), .A2(n13911), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13916) );
  INV_X1 U17418 ( .A(n13912), .ZN(n13914) );
  OAI211_X1 U17419 ( .C1(n14676), .C2(n13914), .A(n10413), .B(n13913), .ZN(
        n13915) );
  OAI211_X1 U17420 ( .C1(n18889), .C2(n17835), .A(n13916), .B(n13915), .ZN(
        n19476) );
  INV_X1 U17421 ( .A(n13917), .ZN(n13918) );
  AOI222_X1 U17422 ( .A1(n19476), .A2(n13932), .B1(n13919), .B2(n13918), .C1(
        n19506), .C2(n17835), .ZN(n13921) );
  NAND2_X1 U17423 ( .A1(n14677), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13920) );
  OAI21_X1 U17424 ( .B1(n13921), .B2(n14677), .A(n13920), .ZN(P3_U3288) );
  OAI21_X1 U17425 ( .B1(n18845), .B2(n13926), .A(n13925), .ZN(n13922) );
  AOI21_X1 U17426 ( .B1(n13923), .B2(n13930), .A(n13922), .ZN(n19489) );
  NOR2_X1 U17427 ( .A1(n19489), .A2(n17869), .ZN(n13924) );
  NOR2_X1 U17428 ( .A1(n13924), .A2(n14677), .ZN(n13934) );
  AOI22_X1 U17429 ( .A1(n13927), .A2(n13926), .B1(n10299), .B2(n13925), .ZN(
        n13928) );
  NOR2_X1 U17430 ( .A1(n13928), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n19492) );
  NAND2_X1 U17431 ( .A1(n13930), .A2(n19488), .ZN(n13931) );
  AND2_X1 U17432 ( .A1(n14359), .A2(n13931), .ZN(n17827) );
  AOI22_X1 U17433 ( .A1(n19492), .A2(n13932), .B1(n17827), .B2(n19506), .ZN(
        n13933) );
  OAI22_X1 U17434 ( .A1(n13934), .A2(n19488), .B1(n13933), .B2(n14677), .ZN(
        P3_U3285) );
  INV_X1 U17435 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13939) );
  INV_X1 U17436 ( .A(n13935), .ZN(n13936) );
  INV_X1 U17437 ( .A(n14019), .ZN(n13938) );
  AOI22_X1 U17438 ( .A1(n17029), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17027), .ZN(n14598) );
  INV_X1 U17439 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13937) );
  OAI222_X1 U17440 ( .A1(n13939), .A2(n13971), .B1(n13938), .B2(n14598), .C1(
        n13937), .C2(n15037), .ZN(P2_U2982) );
  AOI22_X1 U17441 ( .A1(n13968), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n15049), .ZN(n13943) );
  NAND2_X1 U17442 ( .A1(n14016), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13942) );
  INV_X1 U17443 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13940) );
  OR2_X1 U17444 ( .A1(n17027), .A2(n13940), .ZN(n13941) );
  NAND2_X1 U17445 ( .A1(n13942), .A2(n13941), .ZN(n19849) );
  NAND2_X1 U17446 ( .A1(n14019), .A2(n19849), .ZN(n14008) );
  NAND2_X1 U17447 ( .A1(n13943), .A2(n14008), .ZN(P2_U2974) );
  AOI22_X1 U17448 ( .A1(n13968), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n15049), .ZN(n13947) );
  INV_X1 U17449 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13944) );
  OR2_X1 U17450 ( .A1(n17027), .A2(n13944), .ZN(n13946) );
  NAND2_X1 U17451 ( .A1(n17027), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13945) );
  AND2_X1 U17452 ( .A1(n13946), .A2(n13945), .ZN(n19696) );
  NAND2_X1 U17453 ( .A1(n14019), .A2(n19830), .ZN(n14000) );
  NAND2_X1 U17454 ( .A1(n13947), .A2(n14000), .ZN(P2_U2971) );
  AOI22_X1 U17455 ( .A1(n13968), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n15049), .ZN(n13950) );
  NAND2_X1 U17456 ( .A1(n17027), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13949) );
  INV_X1 U17457 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17440) );
  OR2_X1 U17458 ( .A1(n17027), .A2(n17440), .ZN(n13948) );
  NAND2_X1 U17459 ( .A1(n13949), .A2(n13948), .ZN(n17037) );
  NAND2_X1 U17460 ( .A1(n14019), .A2(n17037), .ZN(n13992) );
  NAND2_X1 U17461 ( .A1(n13950), .A2(n13992), .ZN(P2_U2969) );
  AOI22_X1 U17462 ( .A1(n13968), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n15049), .ZN(n13951) );
  AOI22_X1 U17463 ( .A1(n17029), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17027), .ZN(n19714) );
  INV_X1 U17464 ( .A(n19714), .ZN(n19820) );
  NAND2_X1 U17465 ( .A1(n14019), .A2(n19820), .ZN(n14004) );
  NAND2_X1 U17466 ( .A1(n13951), .A2(n14004), .ZN(P2_U2968) );
  AOI22_X1 U17467 ( .A1(n13968), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n15049), .ZN(n13953) );
  AOI22_X1 U17468 ( .A1(n17029), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17027), .ZN(n13952) );
  INV_X1 U17469 ( .A(n13952), .ZN(n19835) );
  NAND2_X1 U17470 ( .A1(n14019), .A2(n19835), .ZN(n14002) );
  NAND2_X1 U17471 ( .A1(n13953), .A2(n14002), .ZN(P2_U2972) );
  AOI22_X1 U17472 ( .A1(n13968), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n15049), .ZN(n13954) );
  AOI22_X1 U17473 ( .A1(n17029), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17027), .ZN(n19703) );
  INV_X1 U17474 ( .A(n19703), .ZN(n19825) );
  NAND2_X1 U17475 ( .A1(n14019), .A2(n19825), .ZN(n13998) );
  NAND2_X1 U17476 ( .A1(n13954), .A2(n13998), .ZN(P2_U2970) );
  AOI22_X1 U17477 ( .A1(n13968), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n15049), .ZN(n13958) );
  NAND2_X1 U17478 ( .A1(n14016), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13957) );
  INV_X1 U17479 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13955) );
  OR2_X1 U17480 ( .A1(n17027), .A2(n13955), .ZN(n13956) );
  NAND2_X1 U17481 ( .A1(n13957), .A2(n13956), .ZN(n19840) );
  NAND2_X1 U17482 ( .A1(n14019), .A2(n19840), .ZN(n14006) );
  NAND2_X1 U17483 ( .A1(n13958), .A2(n14006), .ZN(P2_U2973) );
  AOI22_X1 U17484 ( .A1(n13968), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n15049), .ZN(n13962) );
  INV_X1 U17485 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13959) );
  OR2_X1 U17486 ( .A1(n17027), .A2(n13959), .ZN(n13961) );
  NAND2_X1 U17487 ( .A1(n14016), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13960) );
  NAND2_X1 U17488 ( .A1(n13961), .A2(n13960), .ZN(n16393) );
  NAND2_X1 U17489 ( .A1(n14019), .A2(n16393), .ZN(n13986) );
  NAND2_X1 U17490 ( .A1(n13962), .A2(n13986), .ZN(P2_U2976) );
  NAND2_X1 U17491 ( .A1(n13968), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13966) );
  INV_X1 U17492 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13963) );
  OR2_X1 U17493 ( .A1(n17027), .A2(n13963), .ZN(n13965) );
  NAND2_X1 U17494 ( .A1(n14016), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13964) );
  NAND2_X1 U17495 ( .A1(n13965), .A2(n13964), .ZN(n14926) );
  NAND2_X1 U17496 ( .A1(n14019), .A2(n14926), .ZN(n13969) );
  OAI211_X1 U17497 ( .C1(n13967), .C2(n15037), .A(n13966), .B(n13969), .ZN(
        P2_U2966) );
  INV_X1 U17498 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19718) );
  NAND2_X1 U17499 ( .A1(n13968), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13970) );
  OAI211_X1 U17500 ( .C1(n19718), .C2(n15037), .A(n13970), .B(n13969), .ZN(
        P2_U2981) );
  AOI22_X1 U17501 ( .A1(n14024), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n15049), .ZN(n13975) );
  NAND2_X1 U17502 ( .A1(n17027), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13974) );
  INV_X1 U17503 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13972) );
  OR2_X1 U17504 ( .A1(n17027), .A2(n13972), .ZN(n13973) );
  NAND2_X1 U17505 ( .A1(n13974), .A2(n13973), .ZN(n19814) );
  NAND2_X1 U17506 ( .A1(n14019), .A2(n19814), .ZN(n14010) );
  NAND2_X1 U17507 ( .A1(n13975), .A2(n14010), .ZN(P2_U2967) );
  AOI22_X1 U17508 ( .A1(n14024), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n15049), .ZN(n13979) );
  INV_X1 U17509 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n13976) );
  OR2_X1 U17510 ( .A1(n17027), .A2(n13976), .ZN(n13978) );
  NAND2_X1 U17511 ( .A1(n14016), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13977) );
  NAND2_X1 U17512 ( .A1(n13978), .A2(n13977), .ZN(n16370) );
  NAND2_X1 U17513 ( .A1(n14019), .A2(n16370), .ZN(n13980) );
  NAND2_X1 U17514 ( .A1(n13979), .A2(n13980), .ZN(P2_U2979) );
  AOI22_X1 U17515 ( .A1(n14024), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n15049), .ZN(n13981) );
  NAND2_X1 U17516 ( .A1(n13981), .A2(n13980), .ZN(P2_U2964) );
  AOI22_X1 U17517 ( .A1(n14024), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n15049), .ZN(n13985) );
  INV_X1 U17518 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13982) );
  OR2_X1 U17519 ( .A1(n17027), .A2(n13982), .ZN(n13984) );
  NAND2_X1 U17520 ( .A1(n14016), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13983) );
  NAND2_X1 U17521 ( .A1(n13984), .A2(n13983), .ZN(n16363) );
  NAND2_X1 U17522 ( .A1(n14019), .A2(n16363), .ZN(n13994) );
  NAND2_X1 U17523 ( .A1(n13985), .A2(n13994), .ZN(P2_U2965) );
  AOI22_X1 U17524 ( .A1(n14024), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n15049), .ZN(n13987) );
  NAND2_X1 U17525 ( .A1(n13987), .A2(n13986), .ZN(P2_U2961) );
  AOI22_X1 U17526 ( .A1(n14024), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n15049), .ZN(n13991) );
  INV_X1 U17527 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13988) );
  OR2_X1 U17528 ( .A1(n17027), .A2(n13988), .ZN(n13990) );
  NAND2_X1 U17529 ( .A1(n14016), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13989) );
  NAND2_X1 U17530 ( .A1(n13990), .A2(n13989), .ZN(n16378) );
  NAND2_X1 U17531 ( .A1(n14019), .A2(n16378), .ZN(n13996) );
  NAND2_X1 U17532 ( .A1(n13991), .A2(n13996), .ZN(P2_U2978) );
  AOI22_X1 U17533 ( .A1(n14024), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n15049), .ZN(n13993) );
  NAND2_X1 U17534 ( .A1(n13993), .A2(n13992), .ZN(P2_U2954) );
  AOI22_X1 U17535 ( .A1(n14024), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n15049), .ZN(n13995) );
  NAND2_X1 U17536 ( .A1(n13995), .A2(n13994), .ZN(P2_U2980) );
  AOI22_X1 U17537 ( .A1(n14024), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n15049), .ZN(n13997) );
  NAND2_X1 U17538 ( .A1(n13997), .A2(n13996), .ZN(P2_U2963) );
  AOI22_X1 U17539 ( .A1(n14024), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n15049), .ZN(n13999) );
  NAND2_X1 U17540 ( .A1(n13999), .A2(n13998), .ZN(P2_U2955) );
  AOI22_X1 U17541 ( .A1(n14024), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n15049), .ZN(n14001) );
  NAND2_X1 U17542 ( .A1(n14001), .A2(n14000), .ZN(P2_U2956) );
  AOI22_X1 U17543 ( .A1(n14024), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n15049), .ZN(n14003) );
  NAND2_X1 U17544 ( .A1(n14003), .A2(n14002), .ZN(P2_U2957) );
  AOI22_X1 U17545 ( .A1(n14024), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n15049), .ZN(n14005) );
  NAND2_X1 U17546 ( .A1(n14005), .A2(n14004), .ZN(P2_U2953) );
  AOI22_X1 U17547 ( .A1(n14024), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n15049), .ZN(n14007) );
  NAND2_X1 U17548 ( .A1(n14007), .A2(n14006), .ZN(P2_U2958) );
  AOI22_X1 U17549 ( .A1(n14024), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n15049), .ZN(n14009) );
  NAND2_X1 U17550 ( .A1(n14009), .A2(n14008), .ZN(P2_U2959) );
  NAND2_X1 U17551 ( .A1(n14024), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14011) );
  OAI211_X1 U17552 ( .C1(n14012), .C2(n15037), .A(n14011), .B(n14010), .ZN(
        P2_U2952) );
  INV_X1 U17553 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19726) );
  NAND2_X1 U17554 ( .A1(n14024), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14015) );
  INV_X1 U17555 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17430) );
  OR2_X1 U17556 ( .A1(n17027), .A2(n17430), .ZN(n14014) );
  NAND2_X1 U17557 ( .A1(n14016), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U17558 ( .A1(n14014), .A2(n14013), .ZN(n16385) );
  NAND2_X1 U17559 ( .A1(n14019), .A2(n16385), .ZN(n14021) );
  OAI211_X1 U17560 ( .C1(n19726), .C2(n15037), .A(n14015), .B(n14021), .ZN(
        P2_U2977) );
  INV_X1 U17561 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19730) );
  NAND2_X1 U17562 ( .A1(n14024), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n14020) );
  INV_X1 U17563 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n21711) );
  OR2_X1 U17564 ( .A1(n17027), .A2(n21711), .ZN(n14018) );
  NAND2_X1 U17565 ( .A1(n14016), .A2(BUF2_REG_8__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U17566 ( .A1(n14018), .A2(n14017), .ZN(n16401) );
  NAND2_X1 U17567 ( .A1(n14019), .A2(n16401), .ZN(n14025) );
  OAI211_X1 U17568 ( .C1(n19730), .C2(n15037), .A(n14020), .B(n14025), .ZN(
        P2_U2975) );
  NAND2_X1 U17569 ( .A1(n14024), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14022) );
  OAI211_X1 U17570 ( .C1(n14023), .C2(n15037), .A(n14022), .B(n14021), .ZN(
        P2_U2962) );
  NAND2_X1 U17571 ( .A1(n14024), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14026) );
  OAI211_X1 U17572 ( .C1(n14027), .C2(n15037), .A(n14026), .B(n14025), .ZN(
        P2_U2960) );
  AOI211_X1 U17573 ( .C1(n20774), .C2(n14029), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n14028), .ZN(n14031) );
  INV_X1 U17574 ( .A(n14030), .ZN(n14668) );
  NOR2_X1 U17575 ( .A1(n14031), .A2(n14668), .ZN(n15890) );
  INV_X1 U17576 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14032) );
  NOR2_X1 U17577 ( .A1(n20576), .A2(n14032), .ZN(n15892) );
  INV_X1 U17578 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14033) );
  AOI21_X1 U17579 ( .B1(n15577), .B2(n14034), .A(n14033), .ZN(n14035) );
  AOI211_X1 U17580 ( .C1(n15890), .C2(n20710), .A(n15892), .B(n14035), .ZN(
        n14036) );
  OAI21_X1 U17581 ( .B1(n20770), .B2(n15367), .A(n14036), .ZN(P1_U2999) );
  INV_X1 U17582 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U17583 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20662), .B1(n20681), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14040) );
  OAI21_X1 U17584 ( .B1(n14041), .B2(n20654), .A(n14040), .ZN(P1_U2910) );
  AOI22_X1 U17585 ( .A1(n20662), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14042) );
  OAI21_X1 U17586 ( .B1(n15435), .B2(n20654), .A(n14042), .ZN(P1_U2914) );
  AOI22_X1 U17587 ( .A1(n20662), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14043) );
  OAI21_X1 U17588 ( .B1(n15443), .B2(n20654), .A(n14043), .ZN(P1_U2916) );
  INV_X1 U17589 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14718) );
  AOI22_X1 U17590 ( .A1(n20662), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14044) );
  OAI21_X1 U17591 ( .B1(n14718), .B2(n20654), .A(n14044), .ZN(P1_U2912) );
  INV_X1 U17592 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U17593 ( .A1(n20662), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14045) );
  OAI21_X1 U17594 ( .B1(n14046), .B2(n20654), .A(n14045), .ZN(P1_U2919) );
  AOI22_X1 U17595 ( .A1(n20662), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14047) );
  OAI21_X1 U17596 ( .B1(n15413), .B2(n20654), .A(n14047), .ZN(P1_U2908) );
  INV_X1 U17597 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U17598 ( .A1(n20662), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14048) );
  OAI21_X1 U17599 ( .B1(n14049), .B2(n20654), .A(n14048), .ZN(P1_U2917) );
  INV_X1 U17600 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17601 ( .A1(n20662), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14050) );
  OAI21_X1 U17602 ( .B1(n14241), .B2(n20654), .A(n14050), .ZN(P1_U2909) );
  INV_X1 U17603 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U17604 ( .A1(n20662), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14051) );
  OAI21_X1 U17605 ( .B1(n14236), .B2(n20654), .A(n14051), .ZN(P1_U2906) );
  AOI22_X1 U17606 ( .A1(n20662), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14052) );
  OAI21_X1 U17607 ( .B1(n15439), .B2(n20654), .A(n14052), .ZN(P1_U2915) );
  INV_X1 U17608 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17609 ( .A1(n20662), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14053) );
  OAI21_X1 U17610 ( .B1(n14054), .B2(n20654), .A(n14053), .ZN(P1_U2913) );
  XNOR2_X2 U17611 ( .A(n14057), .B(n14056), .ZN(n20491) );
  INV_X1 U17612 ( .A(n20491), .ZN(n17015) );
  INV_X1 U17613 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14058) );
  MUX2_X1 U17614 ( .A(n19802), .B(n14058), .S(n16360), .Z(n14059) );
  OAI21_X1 U17615 ( .B1(n17015), .B2(n16353), .A(n14059), .ZN(P2_U2885) );
  OR2_X1 U17616 ( .A1(n14061), .A2(n14060), .ZN(n14062) );
  NAND2_X1 U17617 ( .A1(n14168), .A2(n14062), .ZN(n15360) );
  OAI21_X1 U17618 ( .B1(n14065), .B2(n14064), .A(n14063), .ZN(n20758) );
  AOI22_X1 U17619 ( .A1(n20648), .A2(n20758), .B1(n15404), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n14066) );
  OAI21_X1 U17620 ( .B1(n15360), .B2(n15399), .A(n14066), .ZN(P1_U2871) );
  MUX2_X1 U17621 ( .A(n10100), .B(n10491), .S(n16360), .Z(n14071) );
  OAI21_X1 U17622 ( .B1(n20124), .B2(n16353), .A(n14071), .ZN(P2_U2884) );
  INV_X1 U17623 ( .A(n19010), .ZN(n18999) );
  NAND2_X1 U17624 ( .A1(n10299), .A2(n14077), .ZN(n14095) );
  OAI211_X1 U17625 ( .C1(n18822), .C2(n14076), .A(n14072), .B(n14095), .ZN(
        n14127) );
  AOI21_X1 U17626 ( .B1(n18951), .B2(n14127), .A(n19008), .ZN(n14073) );
  OAI21_X1 U17627 ( .B1(n14081), .B2(n18999), .A(n14073), .ZN(n14105) );
  INV_X1 U17628 ( .A(n14105), .ZN(n14085) );
  AOI21_X1 U17629 ( .B1(n14086), .B2(n14075), .A(n14074), .ZN(n18769) );
  NAND2_X1 U17630 ( .A1(n18769), .A2(n19015), .ZN(n14084) );
  INV_X1 U17631 ( .A(n14076), .ZN(n18982) );
  OAI22_X1 U17632 ( .A1(n14077), .A2(n18889), .B1(n14090), .B2(n18982), .ZN(
        n14128) );
  INV_X1 U17633 ( .A(n14128), .ZN(n17233) );
  NOR3_X1 U17634 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17233), .A3(
        n19006), .ZN(n14082) );
  INV_X1 U17635 ( .A(n17252), .ZN(n19012) );
  XNOR2_X1 U17636 ( .A(n14078), .B(n14079), .ZN(n18766) );
  OAI22_X1 U17637 ( .A1(n19012), .A2(n18766), .B1(n10420), .B2(n19546), .ZN(
        n14080) );
  AOI21_X1 U17638 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(n14083) );
  OAI211_X1 U17639 ( .C1(n14086), .C2(n14085), .A(n14084), .B(n14083), .ZN(
        P3_U2856) );
  AOI21_X1 U17640 ( .B1(n14088), .B2(n14087), .A(n9823), .ZN(n14089) );
  INV_X1 U17641 ( .A(n14089), .ZN(n17170) );
  OR2_X1 U17642 ( .A1(n13253), .A2(n14090), .ZN(n14094) );
  NAND2_X1 U17643 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14091) );
  OAI22_X1 U17644 ( .A1(n18822), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18889), .B2(n14091), .ZN(n14092) );
  NOR2_X1 U17645 ( .A1(n17228), .A2(n14092), .ZN(n14093) );
  MUX2_X1 U17646 ( .A(n14094), .B(n14093), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n14096) );
  OAI211_X1 U17647 ( .C1(n18933), .C2(n17170), .A(n14096), .B(n14095), .ZN(
        n14097) );
  NAND2_X1 U17648 ( .A1(n14097), .A2(n18951), .ZN(n14102) );
  XOR2_X1 U17649 ( .A(n14098), .B(n14099), .Z(n17173) );
  NAND2_X1 U17650 ( .A1(n9696), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n17167) );
  INV_X1 U17651 ( .A(n17167), .ZN(n14100) );
  AOI21_X1 U17652 ( .B1(n17252), .B2(n17173), .A(n14100), .ZN(n14101) );
  OAI211_X1 U17653 ( .C1(n18998), .C2(n14103), .A(n14102), .B(n14101), .ZN(
        P3_U2860) );
  XNOR2_X1 U17654 ( .A(n14104), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18774) );
  NAND3_X1 U17655 ( .A1(n18951), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n14128), .ZN(n19019) );
  NOR2_X1 U17656 ( .A1(n19018), .A2(n19019), .ZN(n14107) );
  INV_X1 U17657 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n21593) );
  NOR2_X1 U17658 ( .A1(n10420), .A2(n21593), .ZN(n18778) );
  AOI221_X1 U17659 ( .B1(n14107), .B2(n14106), .C1(n14105), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18778), .ZN(n14111) );
  AOI21_X1 U17660 ( .B1(n9822), .B2(n14109), .A(n14108), .ZN(n18779) );
  NAND2_X1 U17661 ( .A1(n18779), .A2(n19015), .ZN(n14110) );
  OAI211_X1 U17662 ( .C1(n18774), .C2(n19012), .A(n14111), .B(n14110), .ZN(
        P3_U2857) );
  NOR2_X1 U17663 ( .A1(n17175), .A2(n17177), .ZN(n17186) );
  NOR2_X1 U17664 ( .A1(n10299), .A2(n18978), .ZN(n18910) );
  NOR3_X1 U17665 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18910), .A3(
        n19006), .ZN(n17253) );
  AOI21_X1 U17666 ( .B1(n18845), .B2(n18951), .A(n10151), .ZN(n14112) );
  OAI21_X1 U17667 ( .B1(n17253), .B2(n14112), .A(n10420), .ZN(n14115) );
  INV_X1 U17668 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n14113) );
  NOR2_X1 U17669 ( .A1(n10420), .A2(n14113), .ZN(n17182) );
  AOI21_X1 U17670 ( .B1(n17252), .B2(n17186), .A(n17182), .ZN(n14114) );
  OAI211_X1 U17671 ( .C1(n17186), .C2(n17248), .A(n14115), .B(n14114), .ZN(
        P3_U2862) );
  NAND2_X1 U17672 ( .A1(n14117), .A2(n14116), .ZN(n14118) );
  XNOR2_X1 U17673 ( .A(n14118), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17155) );
  INV_X1 U17674 ( .A(n17155), .ZN(n14126) );
  AOI21_X1 U17675 ( .B1(n18892), .B2(n18980), .A(n14127), .ZN(n19000) );
  AOI221_X1 U17676 ( .B1(n17233), .B2(n14120), .C1(n14119), .C2(n14120), .A(
        n19000), .ZN(n14122) );
  INV_X1 U17677 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19548) );
  NOR2_X1 U17678 ( .A1(n10420), .A2(n19548), .ZN(n17152) );
  AND2_X1 U17679 ( .A1(n19008), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14121) );
  AOI211_X1 U17680 ( .C1(n14122), .C2(n18951), .A(n17152), .B(n14121), .ZN(
        n14125) );
  XOR2_X1 U17681 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n14123), .Z(
        n17154) );
  NAND2_X1 U17682 ( .A1(n17154), .A2(n17252), .ZN(n14124) );
  OAI211_X1 U17683 ( .C1(n14126), .C2(n17248), .A(n14125), .B(n14124), .ZN(
        P3_U2855) );
  NAND2_X1 U17684 ( .A1(n9696), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n17158) );
  OR2_X1 U17685 ( .A1(n14130), .A2(n14127), .ZN(n19009) );
  OAI211_X1 U17686 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n14128), .A(
        n18951), .B(n19009), .ZN(n14129) );
  OAI211_X1 U17687 ( .C1(n18998), .C2(n14130), .A(n17158), .B(n14129), .ZN(
        n14137) );
  AOI21_X1 U17688 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n17165) );
  INV_X1 U17689 ( .A(n17165), .ZN(n14135) );
  XNOR2_X1 U17690 ( .A(n14134), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17159) );
  OAI22_X1 U17691 ( .A1(n17248), .A2(n14135), .B1(n19012), .B2(n17159), .ZN(
        n14136) );
  OR2_X1 U17692 ( .A1(n14137), .A2(n14136), .ZN(P3_U2859) );
  NAND2_X1 U17693 ( .A1(n14138), .A2(n11926), .ZN(n14139) );
  AND2_X1 U17694 ( .A1(n14143), .A2(n20818), .ZN(n14145) );
  AND2_X1 U17695 ( .A1(n15497), .A2(n14146), .ZN(n14720) );
  NAND2_X1 U17696 ( .A1(n20769), .A2(DATAI_0_), .ZN(n14149) );
  NAND2_X1 U17697 ( .A1(n20771), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14148) );
  AND2_X1 U17698 ( .A1(n14149), .A2(n14148), .ZN(n20783) );
  INV_X1 U17699 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20684) );
  OAI222_X1 U17700 ( .A1(n15501), .A2(n15367), .B1(n15499), .B2(n20783), .C1(
        n15497), .C2(n20684), .ZN(P1_U2904) );
  NAND2_X1 U17701 ( .A1(n20769), .A2(DATAI_1_), .ZN(n14151) );
  NAND2_X1 U17702 ( .A1(n20771), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14150) );
  AND2_X1 U17703 ( .A1(n14151), .A2(n14150), .ZN(n20793) );
  OAI222_X1 U17704 ( .A1(n15501), .A2(n15360), .B1(n15499), .B2(n20793), .C1(
        n15497), .C2(n14280), .ZN(P1_U2903) );
  INV_X1 U17705 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14152) );
  NOR2_X1 U17706 ( .A1(n14153), .A2(n14152), .ZN(n14155) );
  NAND2_X1 U17707 ( .A1(n14154), .A2(n14155), .ZN(n14429) );
  INV_X1 U17708 ( .A(n14155), .ZN(n14156) );
  NAND3_X1 U17709 ( .A1(n14158), .A2(n14157), .A3(n14156), .ZN(n14159) );
  NAND2_X1 U17710 ( .A1(n14429), .A2(n14159), .ZN(n19691) );
  NOR2_X1 U17711 ( .A1(n14161), .A2(n14162), .ZN(n14163) );
  OR2_X1 U17712 ( .A1(n14160), .A2(n14163), .ZN(n19753) );
  MUX2_X1 U17713 ( .A(n19753), .B(n14164), .S(n16360), .Z(n14165) );
  OAI21_X1 U17714 ( .B1(n19691), .B2(n16353), .A(n14165), .ZN(P2_U2883) );
  INV_X1 U17715 ( .A(n14166), .ZN(n14167) );
  AOI21_X1 U17716 ( .B1(n14169), .B2(n14168), .A(n14167), .ZN(n20634) );
  INV_X1 U17717 ( .A(n20634), .ZN(n14634) );
  AND2_X1 U17718 ( .A1(n14172), .A2(n14171), .ZN(n14173) );
  OR2_X1 U17719 ( .A1(n14170), .A2(n14173), .ZN(n20637) );
  INV_X1 U17720 ( .A(n20637), .ZN(n20741) );
  AOI22_X1 U17721 ( .A1(n20648), .A2(n20741), .B1(n15404), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14174) );
  OAI21_X1 U17722 ( .B1(n14634), .B2(n15399), .A(n14174), .ZN(P1_U2870) );
  NAND2_X1 U17723 ( .A1(n14176), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14177) );
  NAND2_X1 U17724 ( .A1(n12035), .A2(n14177), .ZN(n21453) );
  NAND2_X1 U17725 ( .A1(n11958), .A2(n21453), .ZN(n14189) );
  XNOR2_X1 U17726 ( .A(n14178), .B(n14192), .ZN(n14179) );
  NAND2_X1 U17727 ( .A1(n14180), .A2(n14179), .ZN(n14188) );
  INV_X1 U17728 ( .A(n14181), .ZN(n14185) );
  INV_X1 U17729 ( .A(n14182), .ZN(n14183) );
  MUX2_X1 U17730 ( .A(n14183), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n11997), .Z(n14184) );
  NAND3_X1 U17731 ( .A1(n14186), .A2(n14185), .A3(n14184), .ZN(n14187) );
  OAI211_X1 U17732 ( .C1(n14191), .C2(n14189), .A(n14188), .B(n14187), .ZN(
        n14190) );
  AOI21_X1 U17733 ( .B1(n21464), .B2(n14191), .A(n14190), .ZN(n21460) );
  MUX2_X1 U17734 ( .A(n14192), .B(n21460), .S(n17265), .Z(n17273) );
  NOR2_X1 U17735 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n17370), .ZN(n14194) );
  INV_X1 U17736 ( .A(n14194), .ZN(n14199) );
  OAI22_X1 U17737 ( .A1(n17273), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n14192), 
        .B2(n14199), .ZN(n14197) );
  MUX2_X1 U17738 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14193), .S(
        n17265), .Z(n17272) );
  AOI22_X1 U17739 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14194), .B1(
        n17272), .B2(n17370), .ZN(n14195) );
  INV_X1 U17740 ( .A(n14195), .ZN(n14196) );
  NAND2_X1 U17741 ( .A1(n14197), .A2(n14196), .ZN(n17284) );
  NAND3_X1 U17742 ( .A1(n20599), .A2(n17370), .A3(n14198), .ZN(n14202) );
  OAI21_X1 U17743 ( .B1(n17265), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n14199), 
        .ZN(n14200) );
  NAND2_X1 U17744 ( .A1(n14200), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14201) );
  AND2_X1 U17745 ( .A1(n14202), .A2(n14201), .ZN(n17282) );
  OAI21_X1 U17746 ( .B1(n17284), .B2(n13859), .A(n17282), .ZN(n15900) );
  NOR2_X1 U17747 ( .A1(n15900), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14203) );
  INV_X1 U17748 ( .A(n21475), .ZN(n21472) );
  NOR2_X1 U17749 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n17370), .ZN(n21465) );
  INV_X1 U17750 ( .A(n21465), .ZN(n15902) );
  INV_X1 U17751 ( .A(n20971), .ZN(n21171) );
  NAND2_X1 U17752 ( .A1(n20971), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21038) );
  NAND2_X1 U17753 ( .A1(n21038), .A2(n9694), .ZN(n20898) );
  AOI21_X1 U17754 ( .B1(n21171), .B2(n20830), .A(n20898), .ZN(n14204) );
  AOI21_X1 U17755 ( .B1(n15902), .B2(n21256), .A(n14204), .ZN(n14206) );
  NAND2_X1 U17756 ( .A1(n21472), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14205) );
  OAI21_X1 U17757 ( .B1(n21472), .B2(n14206), .A(n14205), .ZN(P1_U3477) );
  XOR2_X1 U17758 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14429), .Z(n14211)
         );
  INV_X1 U17759 ( .A(n14316), .ZN(n14434) );
  OR2_X1 U17760 ( .A1(n14160), .A2(n14207), .ZN(n14208) );
  NOR2_X1 U17761 ( .A1(n16350), .A2(n11371), .ZN(n14209) );
  AOI21_X1 U17762 ( .B1(n17376), .B2(n16350), .A(n14209), .ZN(n14210) );
  OAI21_X1 U17763 ( .B1(n14211), .B2(n16353), .A(n14210), .ZN(P2_U2882) );
  NAND2_X1 U17764 ( .A1(n19065), .A2(n19051), .ZN(n14213) );
  NAND3_X1 U17765 ( .A1(n19035), .A2(n19626), .A3(n14322), .ZN(n14215) );
  NAND2_X1 U17766 ( .A1(n14216), .A2(n14215), .ZN(n14217) );
  NOR2_X1 U17767 ( .A1(n14218), .A2(n18415), .ZN(n18390) );
  NAND2_X1 U17768 ( .A1(n18390), .A2(BUF2_REG_1__SCAN_IN), .ZN(n14221) );
  AND2_X1 U17769 ( .A1(n18282), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n14219) );
  NAND2_X1 U17770 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n18281) );
  NAND2_X1 U17771 ( .A1(n18282), .A2(n19065), .ZN(n18372) );
  NOR2_X1 U17772 ( .A1(n18281), .A2(n18372), .ZN(n18419) );
  INV_X1 U17773 ( .A(n18419), .ZN(n18403) );
  OAI211_X1 U17774 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n14219), .A(n18415), .B(
        n18403), .ZN(n14220) );
  OAI211_X1 U17775 ( .C1(n14222), .C2(n18421), .A(n14221), .B(n14220), .ZN(
        P3_U2734) );
  NAND2_X1 U17776 ( .A1(n18390), .A2(BUF2_REG_0__SCAN_IN), .ZN(n14226) );
  INV_X1 U17777 ( .A(n18282), .ZN(n14224) );
  AOI22_X1 U17778 ( .A1(n14224), .A2(P3_EAX_REG_0__SCAN_IN), .B1(n14223), .B2(
        n18399), .ZN(n14225) );
  OAI211_X1 U17779 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(n18372), .A(n14226), .B(
        n14225), .ZN(P3_U2735) );
  NAND2_X1 U17780 ( .A1(n20769), .A2(DATAI_2_), .ZN(n14228) );
  NAND2_X1 U17781 ( .A1(n20771), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14227) );
  INV_X1 U17782 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20679) );
  OAI222_X1 U17783 ( .A1(n15501), .A2(n14634), .B1(n15499), .B2(n20797), .C1(
        n15497), .C2(n20679), .ZN(P1_U2902) );
  NAND2_X1 U17784 ( .A1(n20792), .A2(n21487), .ZN(n14230) );
  NAND2_X1 U17785 ( .A1(n20769), .A2(DATAI_14_), .ZN(n14233) );
  NAND2_X1 U17786 ( .A1(n20771), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14232) );
  AND2_X1 U17787 ( .A1(n14233), .A2(n14232), .ZN(n15469) );
  INV_X1 U17788 ( .A(n15469), .ZN(n14234) );
  NAND2_X1 U17789 ( .A1(n20690), .A2(n14234), .ZN(n20701) );
  NAND2_X1 U17790 ( .A1(n21497), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14235) );
  OAI211_X1 U17791 ( .C1(n21499), .C2(n14236), .A(n20701), .B(n14235), .ZN(
        P1_U2951) );
  NAND2_X1 U17792 ( .A1(n20769), .A2(DATAI_11_), .ZN(n14238) );
  NAND2_X1 U17793 ( .A1(n20771), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14237) );
  AND2_X1 U17794 ( .A1(n14238), .A2(n14237), .ZN(n15476) );
  INV_X1 U17795 ( .A(n15476), .ZN(n14239) );
  NAND2_X1 U17796 ( .A1(n20690), .A2(n14239), .ZN(n20694) );
  NAND2_X1 U17797 ( .A1(n21497), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14240) );
  OAI211_X1 U17798 ( .C1(n21499), .C2(n14241), .A(n20694), .B(n14240), .ZN(
        P1_U2948) );
  NAND2_X1 U17799 ( .A1(n20769), .A2(DATAI_12_), .ZN(n14243) );
  NAND2_X1 U17800 ( .A1(n20771), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14242) );
  AND2_X1 U17801 ( .A1(n14243), .A2(n14242), .ZN(n15473) );
  INV_X1 U17802 ( .A(n15473), .ZN(n14244) );
  NAND2_X1 U17803 ( .A1(n20690), .A2(n14244), .ZN(n20696) );
  NAND2_X1 U17804 ( .A1(n21497), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14245) );
  OAI211_X1 U17805 ( .C1(n21499), .C2(n15413), .A(n20696), .B(n14245), .ZN(
        P1_U2949) );
  INV_X1 U17806 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14248) );
  INV_X1 U17807 ( .A(DATAI_10_), .ZN(n14246) );
  MUX2_X1 U17808 ( .A(n14246), .B(n17430), .S(n20771), .Z(n15478) );
  NOR2_X1 U17809 ( .A1(n14296), .A2(n15478), .ZN(n21496) );
  AOI21_X1 U17810 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n21497), .A(n21496), 
        .ZN(n14247) );
  OAI21_X1 U17811 ( .B1(n14248), .B2(n21499), .A(n14247), .ZN(P1_U2962) );
  INV_X1 U17812 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n14252) );
  NAND2_X1 U17813 ( .A1(n20769), .A2(DATAI_4_), .ZN(n14250) );
  NAND2_X1 U17814 ( .A1(n20771), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14249) );
  AND2_X1 U17815 ( .A1(n14250), .A2(n14249), .ZN(n20805) );
  NOR2_X1 U17816 ( .A1(n14296), .A2(n20805), .ZN(n14290) );
  AOI21_X1 U17817 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n21497), .A(n14290), 
        .ZN(n14251) );
  OAI21_X1 U17818 ( .B1(n14252), .B2(n21499), .A(n14251), .ZN(P1_U2956) );
  INV_X1 U17819 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14256) );
  NAND2_X1 U17820 ( .A1(n20769), .A2(DATAI_5_), .ZN(n14254) );
  NAND2_X1 U17821 ( .A1(n20771), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14253) );
  AND2_X1 U17822 ( .A1(n14254), .A2(n14253), .ZN(n20809) );
  NOR2_X1 U17823 ( .A1(n14296), .A2(n20809), .ZN(n14272) );
  AOI21_X1 U17824 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n21497), .A(n14272), 
        .ZN(n14255) );
  OAI21_X1 U17825 ( .B1(n14256), .B2(n21499), .A(n14255), .ZN(P1_U2957) );
  NAND2_X1 U17826 ( .A1(n20769), .A2(DATAI_7_), .ZN(n14258) );
  NAND2_X1 U17827 ( .A1(n20771), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14257) );
  AND2_X1 U17828 ( .A1(n14258), .A2(n14257), .ZN(n20821) );
  NOR2_X1 U17829 ( .A1(n14296), .A2(n20821), .ZN(n14265) );
  AOI21_X1 U17830 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n21497), .A(n14265), 
        .ZN(n14259) );
  OAI21_X1 U17831 ( .B1(n14260), .B2(n21499), .A(n14259), .ZN(P1_U2959) );
  INV_X1 U17832 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20670) );
  INV_X1 U17833 ( .A(DATAI_8_), .ZN(n14261) );
  MUX2_X1 U17834 ( .A(n14261), .B(n21711), .S(n20771), .Z(n15484) );
  NOR2_X1 U17835 ( .A1(n14296), .A2(n15484), .ZN(n14263) );
  AOI21_X1 U17836 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21497), .A(n14263), 
        .ZN(n14262) );
  OAI21_X1 U17837 ( .B1(n20670), .B2(n21499), .A(n14262), .ZN(P1_U2960) );
  AOI21_X1 U17838 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n21497), .A(n14263), 
        .ZN(n14264) );
  OAI21_X1 U17839 ( .B1(n14718), .B2(n21499), .A(n14264), .ZN(P1_U2945) );
  AOI21_X1 U17840 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n21497), .A(n14265), 
        .ZN(n14266) );
  OAI21_X1 U17841 ( .B1(n14054), .B2(n21499), .A(n14266), .ZN(P1_U2944) );
  NAND2_X1 U17842 ( .A1(n20769), .A2(DATAI_6_), .ZN(n14268) );
  NAND2_X1 U17843 ( .A1(n20771), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14267) );
  AND2_X1 U17844 ( .A1(n14268), .A2(n14267), .ZN(n20813) );
  NOR2_X1 U17845 ( .A1(n14296), .A2(n20813), .ZN(n14270) );
  AOI21_X1 U17846 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n21497), .A(n14270), 
        .ZN(n14269) );
  OAI21_X1 U17847 ( .B1(n15488), .B2(n21499), .A(n14269), .ZN(P1_U2958) );
  AOI21_X1 U17848 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n21497), .A(n14270), 
        .ZN(n14271) );
  OAI21_X1 U17849 ( .B1(n15435), .B2(n21499), .A(n14271), .ZN(P1_U2943) );
  AOI21_X1 U17850 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n21497), .A(n14272), 
        .ZN(n14273) );
  OAI21_X1 U17851 ( .B1(n15439), .B2(n21499), .A(n14273), .ZN(P1_U2942) );
  INV_X1 U17852 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n14277) );
  NAND2_X1 U17853 ( .A1(n20769), .A2(DATAI_3_), .ZN(n14275) );
  NAND2_X1 U17854 ( .A1(n20771), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14274) );
  AND2_X1 U17855 ( .A1(n14275), .A2(n14274), .ZN(n20801) );
  NOR2_X1 U17856 ( .A1(n14296), .A2(n20801), .ZN(n14288) );
  AOI21_X1 U17857 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n21497), .A(n14288), 
        .ZN(n14276) );
  OAI21_X1 U17858 ( .B1(n14277), .B2(n21499), .A(n14276), .ZN(P1_U2955) );
  NOR2_X1 U17859 ( .A1(n14296), .A2(n20797), .ZN(n14286) );
  AOI21_X1 U17860 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n21497), .A(n14286), 
        .ZN(n14278) );
  OAI21_X1 U17861 ( .B1(n20679), .B2(n21499), .A(n14278), .ZN(P1_U2954) );
  INV_X1 U17862 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n14280) );
  NOR2_X1 U17863 ( .A1(n14296), .A2(n20793), .ZN(n14284) );
  AOI21_X1 U17864 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n21497), .A(n14284), 
        .ZN(n14279) );
  OAI21_X1 U17865 ( .B1(n14280), .B2(n21499), .A(n14279), .ZN(P1_U2953) );
  NOR2_X1 U17866 ( .A1(n14296), .A2(n20783), .ZN(n14282) );
  AOI21_X1 U17867 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n21497), .A(n14282), 
        .ZN(n14281) );
  OAI21_X1 U17868 ( .B1(n20684), .B2(n21499), .A(n14281), .ZN(P1_U2952) );
  AOI21_X1 U17869 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n21497), .A(n14282), 
        .ZN(n14283) );
  OAI21_X1 U17870 ( .B1(n15459), .B2(n21499), .A(n14283), .ZN(P1_U2937) );
  AOI21_X1 U17871 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n21497), .A(n14284), 
        .ZN(n14285) );
  OAI21_X1 U17872 ( .B1(n14046), .B2(n21499), .A(n14285), .ZN(P1_U2938) );
  AOI21_X1 U17873 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n21497), .A(n14286), 
        .ZN(n14287) );
  OAI21_X1 U17874 ( .B1(n15451), .B2(n21499), .A(n14287), .ZN(P1_U2939) );
  AOI21_X1 U17875 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n21497), .A(n14288), 
        .ZN(n14289) );
  OAI21_X1 U17876 ( .B1(n14049), .B2(n21499), .A(n14289), .ZN(P1_U2940) );
  AOI21_X1 U17877 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n21497), .A(n14290), 
        .ZN(n14291) );
  OAI21_X1 U17878 ( .B1(n15443), .B2(n21499), .A(n14291), .ZN(P1_U2941) );
  INV_X1 U17879 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14292) );
  NOR2_X1 U17880 ( .A1(n20769), .A2(n14292), .ZN(n14293) );
  AOI21_X1 U17881 ( .B1(DATAI_15_), .B2(n20769), .A(n14293), .ZN(n15466) );
  INV_X1 U17882 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14295) );
  OAI222_X1 U17883 ( .A1(n21499), .A2(n20661), .B1(n14296), .B2(n15466), .C1(
        n14295), .C2(n14294), .ZN(P1_U2967) );
  INV_X1 U17884 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19041) );
  INV_X1 U17885 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18482) );
  NOR2_X1 U17886 ( .A1(n18482), .A2(n18403), .ZN(n14298) );
  AOI21_X1 U17887 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18415), .A(n18419), .ZN(
        n14297) );
  NOR2_X1 U17888 ( .A1(n14298), .A2(n14297), .ZN(n14299) );
  AOI21_X1 U17889 ( .B1(n14300), .B2(n18399), .A(n14299), .ZN(n14301) );
  OAI21_X1 U17890 ( .B1(n18424), .B2(n19041), .A(n14301), .ZN(P3_U2733) );
  INV_X1 U17891 ( .A(n14302), .ZN(n14304) );
  NAND2_X1 U17892 ( .A1(n14304), .A2(n14303), .ZN(n14553) );
  OAI211_X1 U17893 ( .C1(n14304), .C2(n14303), .A(n14553), .B(n16357), .ZN(
        n14306) );
  NAND2_X1 U17894 ( .A1(n16142), .A2(n16350), .ZN(n14305) );
  OAI211_X1 U17895 ( .C1(n16350), .C2(n16132), .A(n14306), .B(n14305), .ZN(
        P2_U2877) );
  INV_X1 U17896 ( .A(n14307), .ZN(n14552) );
  XNOR2_X1 U17897 ( .A(n14553), .B(n14552), .ZN(n14313) );
  AND2_X1 U17898 ( .A1(n14309), .A2(n14308), .ZN(n14310) );
  OR2_X1 U17899 ( .A1(n14310), .A2(n14550), .ZN(n16858) );
  MUX2_X1 U17900 ( .A(n16858), .B(n14311), .S(n16360), .Z(n14312) );
  OAI21_X1 U17901 ( .B1(n14313), .B2(n16353), .A(n14312), .ZN(P2_U2876) );
  NOR2_X1 U17902 ( .A1(n14429), .A2(n14314), .ZN(n14540) );
  XNOR2_X1 U17903 ( .A(n14540), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14320) );
  AND2_X1 U17904 ( .A1(n14316), .A2(n14315), .ZN(n14653) );
  OR2_X1 U17905 ( .A1(n14434), .A2(n14435), .ZN(n14432) );
  AND2_X1 U17906 ( .A1(n14432), .A2(n14317), .ZN(n14318) );
  OR2_X1 U17907 ( .A1(n14653), .A2(n14318), .ZN(n16899) );
  MUX2_X1 U17908 ( .A(n16899), .B(n10593), .S(n16360), .Z(n14319) );
  OAI21_X1 U17909 ( .B1(n14320), .B2(n16353), .A(n14319), .ZN(P2_U2880) );
  AND2_X1 U17910 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17919) );
  INV_X1 U17911 ( .A(n19509), .ZN(n19518) );
  NOR2_X1 U17912 ( .A1(n19626), .A2(n19518), .ZN(n14321) );
  NAND2_X1 U17913 ( .A1(n19065), .A2(n18279), .ZN(n18273) );
  INV_X1 U17914 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17597) );
  INV_X1 U17915 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17997) );
  NAND2_X1 U17916 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n18246) );
  NAND2_X1 U17917 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .ZN(n18093) );
  NAND4_X1 U17918 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n14325)
         );
  INV_X1 U17919 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21756) );
  NAND3_X1 U17920 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18259) );
  INV_X1 U17921 ( .A(n18259), .ZN(n14323) );
  NAND3_X1 U17922 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n14323), .ZN(n18254) );
  OR4_X1 U17923 ( .A1(n17678), .A2(n21756), .A3(n21783), .A4(n18254), .ZN(
        n14324) );
  NOR4_X1 U17924 ( .A1(n18246), .A2(n18093), .A3(n14325), .A4(n14324), .ZN(
        n18031) );
  NAND2_X1 U17925 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18031), .ZN(n18051) );
  NOR3_X1 U17926 ( .A1(n18050), .A2(n18264), .A3(n18051), .ZN(n18035) );
  NAND2_X1 U17927 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18035), .ZN(n17999) );
  NAND2_X1 U17928 ( .A1(n19065), .A2(n18015), .ZN(n17996) );
  NAND2_X1 U17929 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17980), .ZN(n17963) );
  NAND3_X1 U17930 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17939), .ZN(n17925) );
  NAND2_X1 U17931 ( .A1(n18271), .A2(n17925), .ZN(n17929) );
  OAI21_X1 U17932 ( .B1(n17919), .B2(n18273), .A(n17929), .ZN(n17920) );
  INV_X1 U17933 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14327) );
  AOI22_X1 U17934 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18152), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14326) );
  OAI21_X1 U17935 ( .B1(n14388), .B2(n14327), .A(n14326), .ZN(n14328) );
  AOI21_X1 U17936 ( .B1(n18180), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n14328), .ZN(n14331) );
  AOI22_X1 U17937 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U17938 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14329) );
  NAND3_X1 U17939 ( .A1(n14331), .A2(n14330), .A3(n14329), .ZN(n14337) );
  AOI22_X1 U17940 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14335) );
  AOI22_X1 U17941 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U17942 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U17943 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14332) );
  NAND4_X1 U17944 ( .A1(n14335), .A2(n14334), .A3(n14333), .A4(n14332), .ZN(
        n14336) );
  NOR2_X1 U17945 ( .A1(n14337), .A2(n14336), .ZN(n14423) );
  AOI22_X1 U17946 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18194), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17947 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U17948 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U17949 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14338) );
  NAND4_X1 U17950 ( .A1(n14341), .A2(n14340), .A3(n14339), .A4(n14338), .ZN(
        n14351) );
  INV_X1 U17951 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14344) );
  AOI22_X1 U17952 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U17953 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14342) );
  OAI211_X1 U17954 ( .C1(n14344), .C2(n18141), .A(n14343), .B(n14342), .ZN(
        n14349) );
  INV_X1 U17955 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18156) );
  OAI22_X1 U17956 ( .A1(n11711), .A2(n14345), .B1(n13142), .B2(n18156), .ZN(
        n14348) );
  INV_X1 U17957 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18003) );
  INV_X1 U17958 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14346) );
  OAI22_X1 U17959 ( .A1(n18085), .A2(n18003), .B1(n18186), .B2(n14346), .ZN(
        n14347) );
  OR3_X1 U17960 ( .A1(n14349), .A2(n14348), .A3(n14347), .ZN(n14350) );
  NOR2_X1 U17961 ( .A1(n14351), .A2(n14350), .ZN(n17927) );
  AOI22_X1 U17962 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U17963 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14354) );
  AOI22_X1 U17964 ( .A1(n14395), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U17965 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14352) );
  NAND4_X1 U17966 ( .A1(n14355), .A2(n14354), .A3(n14353), .A4(n14352), .ZN(
        n14365) );
  INV_X1 U17967 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U17968 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18152), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U17969 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14356) );
  OAI211_X1 U17970 ( .C1(n18199), .C2(n18141), .A(n14357), .B(n14356), .ZN(
        n14363) );
  OAI22_X1 U17971 ( .A1(n11711), .A2(n18038), .B1(n13041), .B2(n18202), .ZN(
        n14362) );
  INV_X1 U17972 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14360) );
  INV_X1 U17973 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14358) );
  OAI22_X1 U17974 ( .A1(n18186), .A2(n14360), .B1(n14359), .B2(n14358), .ZN(
        n14361) );
  OR3_X1 U17975 ( .A1(n14363), .A2(n14362), .A3(n14361), .ZN(n14364) );
  NOR2_X1 U17976 ( .A1(n14365), .A2(n14364), .ZN(n17936) );
  AOI22_X1 U17977 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14369) );
  INV_X1 U17978 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n21580) );
  AOI22_X1 U17979 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U17980 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17981 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14366) );
  NAND4_X1 U17982 ( .A1(n14369), .A2(n14368), .A3(n14367), .A4(n14366), .ZN(
        n14380) );
  INV_X1 U17983 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17984 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U17985 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14370) );
  OAI211_X1 U17986 ( .C1(n14372), .C2(n18141), .A(n14371), .B(n14370), .ZN(
        n14379) );
  INV_X1 U17987 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14374) );
  OAI22_X1 U17988 ( .A1(n18186), .A2(n14374), .B1(n14388), .B2(n14373), .ZN(
        n14378) );
  INV_X1 U17989 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14376) );
  OAI22_X1 U17990 ( .A1(n14359), .A2(n14376), .B1(n13041), .B2(n14375), .ZN(
        n14377) );
  OR4_X1 U17991 ( .A1(n14380), .A2(n14379), .A3(n14378), .A4(n14377), .ZN(
        n17942) );
  AOI22_X1 U17992 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18229), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U17993 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U17994 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U17995 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14381) );
  NAND4_X1 U17996 ( .A1(n14384), .A2(n14383), .A3(n14382), .A4(n14381), .ZN(
        n14394) );
  INV_X1 U17997 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U17998 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U17999 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14385) );
  OAI211_X1 U18000 ( .C1(n18080), .C2(n14387), .A(n14386), .B(n14385), .ZN(
        n14393) );
  INV_X1 U18001 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14389) );
  INV_X1 U18002 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18082) );
  OAI22_X1 U18003 ( .A1(n18186), .A2(n14389), .B1(n14388), .B2(n18082), .ZN(
        n14392) );
  INV_X1 U18004 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14390) );
  OAI22_X1 U18005 ( .A1(n14359), .A2(n14390), .B1(n13041), .B2(n18081), .ZN(
        n14391) );
  OR4_X1 U18006 ( .A1(n14394), .A2(n14393), .A3(n14392), .A4(n14391), .ZN(
        n17943) );
  NAND2_X1 U18007 ( .A1(n17942), .A2(n17943), .ZN(n17941) );
  NOR2_X1 U18008 ( .A1(n17936), .A2(n17941), .ZN(n17935) );
  AOI22_X1 U18009 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U18010 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U18011 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U18012 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14396) );
  NAND4_X1 U18013 ( .A1(n14399), .A2(n14398), .A3(n14397), .A4(n14396), .ZN(
        n14407) );
  INV_X1 U18014 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U18015 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U18016 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14400) );
  OAI211_X1 U18017 ( .C1(n14402), .C2(n18141), .A(n14401), .B(n14400), .ZN(
        n14406) );
  INV_X1 U18018 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21751) );
  INV_X1 U18019 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18187) );
  OAI22_X1 U18020 ( .A1(n18186), .A2(n21751), .B1(n14388), .B2(n18187), .ZN(
        n14405) );
  INV_X1 U18021 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18185) );
  OAI22_X1 U18022 ( .A1(n14359), .A2(n18185), .B1(n13041), .B2(n14403), .ZN(
        n14404) );
  NAND2_X1 U18023 ( .A1(n17935), .A2(n17932), .ZN(n17931) );
  NOR2_X1 U18024 ( .A1(n17927), .A2(n17931), .ZN(n17926) );
  AOI22_X1 U18025 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U18026 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U18027 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U18028 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14408) );
  NAND4_X1 U18029 ( .A1(n14411), .A2(n14410), .A3(n14409), .A4(n14408), .ZN(
        n14422) );
  INV_X1 U18030 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U18031 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U18032 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14412) );
  OAI211_X1 U18033 ( .C1(n14414), .C2(n18141), .A(n14413), .B(n14412), .ZN(
        n14421) );
  INV_X1 U18034 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14416) );
  INV_X1 U18035 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14415) );
  OAI22_X1 U18036 ( .A1(n18186), .A2(n14416), .B1(n14388), .B2(n14415), .ZN(
        n14420) );
  INV_X1 U18037 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14418) );
  OAI22_X1 U18038 ( .A1(n14359), .A2(n14418), .B1(n13041), .B2(n14417), .ZN(
        n14419) );
  OR4_X1 U18039 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n14419), .ZN(
        n17923) );
  NAND2_X1 U18040 ( .A1(n17926), .A2(n17923), .ZN(n17922) );
  NOR2_X1 U18041 ( .A1(n14423), .A2(n17922), .ZN(n17917) );
  AOI21_X1 U18042 ( .B1(n14423), .B2(n17922), .A(n17917), .ZN(n18296) );
  AOI22_X1 U18043 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17920), .B1(n18296), 
        .B2(n18276), .ZN(n14427) );
  INV_X1 U18044 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14425) );
  INV_X1 U18045 ( .A(n17925), .ZN(n14424) );
  NAND3_X1 U18046 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14425), .A3(n14424), 
        .ZN(n14426) );
  NAND2_X1 U18047 ( .A1(n14427), .A2(n14426), .ZN(P3_U2675) );
  INV_X1 U18048 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14428) );
  NOR2_X1 U18049 ( .A1(n14429), .A2(n14428), .ZN(n14431) );
  INV_X1 U18050 ( .A(n14540), .ZN(n14430) );
  OAI211_X1 U18051 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14431), .A(
        n14430), .B(n16357), .ZN(n14437) );
  INV_X1 U18052 ( .A(n14432), .ZN(n14433) );
  AOI21_X1 U18053 ( .B1(n14435), .B2(n14434), .A(n14433), .ZN(n16197) );
  NAND2_X1 U18054 ( .A1(n16197), .A2(n16350), .ZN(n14436) );
  OAI211_X1 U18055 ( .C1(n16350), .C2(n10574), .A(n14437), .B(n14436), .ZN(
        P2_U2881) );
  INV_X1 U18056 ( .A(n15491), .ZN(n14438) );
  OAI21_X1 U18057 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n20609) );
  INV_X1 U18058 ( .A(n14170), .ZN(n14443) );
  INV_X1 U18059 ( .A(n17355), .ZN(n14441) );
  AOI21_X1 U18060 ( .B1(n14443), .B2(n14442), .A(n14441), .ZN(n20728) );
  AOI22_X1 U18061 ( .A1(n20648), .A2(n20728), .B1(n15404), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14444) );
  OAI21_X1 U18062 ( .B1(n20609), .B2(n15399), .A(n14444), .ZN(P1_U2869) );
  INV_X1 U18063 ( .A(n14445), .ZN(n14446) );
  NAND2_X1 U18064 ( .A1(n11051), .A2(n15048), .ZN(n14513) );
  NAND2_X1 U18065 ( .A1(n14448), .A2(n14447), .ZN(n14482) );
  INV_X1 U18066 ( .A(n10445), .ZN(n14450) );
  NAND2_X1 U18067 ( .A1(n14450), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14451) );
  NAND2_X1 U18068 ( .A1(n12853), .A2(n14451), .ZN(n14452) );
  NAND2_X1 U18069 ( .A1(n14482), .A2(n14452), .ZN(n14457) );
  NAND2_X1 U18070 ( .A1(n14490), .A2(n14491), .ZN(n14479) );
  INV_X1 U18071 ( .A(n14452), .ZN(n14453) );
  NAND2_X1 U18072 ( .A1(n14479), .A2(n14453), .ZN(n14456) );
  NAND2_X1 U18073 ( .A1(n14476), .A2(n14454), .ZN(n14455) );
  NAND3_X1 U18074 ( .A1(n14457), .A2(n14456), .A3(n14455), .ZN(n14458) );
  AOI21_X1 U18075 ( .B1(n10785), .B2(n14473), .A(n14458), .ZN(n17012) );
  NAND2_X1 U18076 ( .A1(n16966), .A2(n14473), .ZN(n14466) );
  INV_X1 U18077 ( .A(n14467), .ZN(n14460) );
  NAND2_X1 U18078 ( .A1(n14460), .A2(n14459), .ZN(n14464) );
  NOR2_X1 U18079 ( .A1(n14461), .A2(n10445), .ZN(n14463) );
  AOI22_X1 U18080 ( .A1(n14464), .A2(n14463), .B1(n14476), .B2(n14462), .ZN(
        n14465) );
  NAND2_X1 U18081 ( .A1(n14466), .A2(n14465), .ZN(n17006) );
  NAND2_X1 U18082 ( .A1(n17006), .A2(n20252), .ZN(n14470) );
  MUX2_X1 U18083 ( .A(n14467), .B(n14476), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14468) );
  AOI21_X1 U18084 ( .B1(n19788), .B2(n14473), .A(n14468), .ZN(n16994) );
  NAND3_X1 U18085 ( .A1(n11449), .A2(n16991), .A3(n11127), .ZN(n14469) );
  NAND4_X1 U18086 ( .A1(n14470), .A2(n16994), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A4(n14469), .ZN(n14471) );
  OAI211_X1 U18087 ( .C1(n20252), .C2(n17006), .A(n14471), .B(n14496), .ZN(
        n14472) );
  AOI21_X1 U18088 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17012), .A(
        n14472), .ZN(n14488) );
  INV_X1 U18089 ( .A(n14473), .ZN(n14485) );
  MUX2_X1 U18090 ( .A(n14474), .B(n10715), .S(n10445), .Z(n14478) );
  XNOR2_X1 U18091 ( .A(n14475), .B(n10715), .ZN(n14477) );
  AOI22_X1 U18092 ( .A1(n14479), .A2(n14478), .B1(n14477), .B2(n14476), .ZN(
        n14484) );
  OAI21_X1 U18093 ( .B1(n14480), .B2(n10715), .A(n10404), .ZN(n14481) );
  NAND2_X1 U18094 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  OAI211_X1 U18095 ( .C1(n10100), .C2(n14485), .A(n14484), .B(n14483), .ZN(
        n17017) );
  MUX2_X1 U18096 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17017), .S(
        n14496), .Z(n14508) );
  MUX2_X1 U18097 ( .A(n10317), .B(n17012), .S(n14496), .Z(n14489) );
  NOR2_X1 U18098 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n14489), .ZN(
        n14486) );
  OR3_X1 U18099 ( .A1(n14488), .A2(n14508), .A3(n14486), .ZN(n14487) );
  AOI22_X1 U18100 ( .A1(n14488), .A2(n14508), .B1(n21570), .B2(n14487), .ZN(
        n14510) );
  INV_X1 U18101 ( .A(n14489), .ZN(n14507) );
  MUX2_X1 U18102 ( .A(n14491), .B(n14490), .S(n14605), .Z(n14495) );
  NAND2_X1 U18103 ( .A1(n14493), .A2(n14492), .ZN(n14494) );
  NAND2_X1 U18104 ( .A1(n14495), .A2(n14494), .ZN(n20504) );
  NOR2_X1 U18105 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n14505) );
  INV_X1 U18106 ( .A(n14496), .ZN(n14497) );
  NAND2_X1 U18107 ( .A1(n14497), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14503) );
  AOI22_X1 U18108 ( .A1(n14501), .A2(n14500), .B1(n14499), .B2(n14498), .ZN(
        n14502) );
  OAI211_X1 U18109 ( .C1(n14505), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        n14506) );
  AOI211_X1 U18110 ( .C1(n14508), .C2(n14507), .A(n20504), .B(n14506), .ZN(
        n14509) );
  OAI21_X1 U18111 ( .B1(n14510), .B2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n14509), .ZN(n14614) );
  OAI21_X1 U18112 ( .B1(n14614), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14512) );
  INV_X1 U18113 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20508) );
  NOR2_X1 U18114 ( .A1(n14511), .A2(n20508), .ZN(n20519) );
  OAI211_X1 U18115 ( .C1(n14514), .C2(n14513), .A(n14512), .B(n20519), .ZN(
        n17045) );
  OAI21_X1 U18116 ( .B1(n17045), .B2(n12673), .A(n14515), .ZN(P2_U3593) );
  OAI222_X1 U18117 ( .A1(n15501), .A2(n20609), .B1(n15499), .B2(n20801), .C1(
        n15497), .C2(n14277), .ZN(P1_U2901) );
  AND2_X1 U18118 ( .A1(n14517), .A2(n14518), .ZN(n14519) );
  NOR2_X1 U18119 ( .A1(n14516), .A2(n14519), .ZN(n16890) );
  INV_X1 U18120 ( .A(n16890), .ZN(n16170) );
  OAI21_X4 U18121 ( .B1(n14521), .B2(n14520), .A(n17047), .ZN(n16451) );
  INV_X1 U18122 ( .A(n11126), .ZN(n14522) );
  NAND2_X1 U18123 ( .A1(n14524), .A2(n14523), .ZN(n14525) );
  INV_X1 U18124 ( .A(n19713), .ZN(n16472) );
  AOI22_X1 U18125 ( .A1(n16472), .A2(n16401), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n16451), .ZN(n14526) );
  OAI21_X1 U18126 ( .B1(n16170), .B2(n16475), .A(n14526), .ZN(P2_U2911) );
  NAND2_X1 U18127 ( .A1(n14583), .A2(n14582), .ZN(n14581) );
  INV_X1 U18128 ( .A(n14528), .ZN(n14529) );
  NAND2_X1 U18129 ( .A1(n14581), .A2(n14529), .ZN(n14530) );
  NAND2_X1 U18130 ( .A1(n14596), .A2(n14530), .ZN(n16815) );
  AOI22_X1 U18131 ( .A1(n16472), .A2(n14926), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n16451), .ZN(n14531) );
  OAI21_X1 U18132 ( .B1(n16815), .B2(n16475), .A(n14531), .ZN(P2_U2905) );
  INV_X1 U18133 ( .A(n14532), .ZN(n16144) );
  AOI22_X1 U18134 ( .A1(n16472), .A2(n16385), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n16451), .ZN(n14533) );
  OAI21_X1 U18135 ( .B1(n16144), .B2(n16475), .A(n14533), .ZN(P2_U2909) );
  INV_X1 U18136 ( .A(n19814), .ZN(n14539) );
  OR2_X1 U18137 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  AND2_X1 U18138 ( .A1(n11145), .A2(n14536), .ZN(n17390) );
  AOI22_X1 U18139 ( .A1(n19705), .A2(n17390), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n16451), .ZN(n14538) );
  NAND2_X1 U18140 ( .A1(n19858), .A2(n17390), .ZN(n19707) );
  OAI211_X1 U18141 ( .C1(n19858), .C2(n17390), .A(n19707), .B(n19709), .ZN(
        n14537) );
  OAI211_X1 U18142 ( .C1(n19713), .C2(n14539), .A(n14538), .B(n14537), .ZN(
        P2_U2919) );
  NAND2_X1 U18143 ( .A1(n14540), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14656) );
  INV_X1 U18144 ( .A(n14541), .ZN(n14657) );
  NOR2_X1 U18145 ( .A1(n14656), .A2(n14657), .ZN(n14655) );
  OAI211_X1 U18146 ( .C1(n14655), .C2(n14542), .A(n16357), .B(n14302), .ZN(
        n14547) );
  INV_X1 U18147 ( .A(n11504), .ZN(n14544) );
  AOI21_X1 U18148 ( .B1(n14545), .B2(n14543), .A(n14544), .ZN(n16871) );
  NAND2_X1 U18149 ( .A1(n16871), .A2(n16350), .ZN(n14546) );
  OAI211_X1 U18150 ( .C1(n16350), .C2(n10213), .A(n14547), .B(n14546), .ZN(
        P2_U2878) );
  NOR2_X1 U18151 ( .A1(n14550), .A2(n14549), .ZN(n14551) );
  OR2_X1 U18152 ( .A1(n14548), .A2(n14551), .ZN(n16844) );
  NOR2_X1 U18153 ( .A1(n14553), .A2(n14552), .ZN(n14555) );
  NAND2_X1 U18154 ( .A1(n14555), .A2(n14554), .ZN(n14643) );
  OAI211_X1 U18155 ( .C1(n14555), .C2(n14554), .A(n14643), .B(n16357), .ZN(
        n14557) );
  NAND2_X1 U18156 ( .A1(n16360), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14556) );
  OAI211_X1 U18157 ( .C1(n16360), .C2(n16844), .A(n14557), .B(n14556), .ZN(
        P2_U2875) );
  INV_X1 U18158 ( .A(n17037), .ZN(n14572) );
  OR2_X1 U18159 ( .A1(n14559), .A2(n14558), .ZN(n14560) );
  NAND2_X1 U18160 ( .A1(n14561), .A2(n14560), .ZN(n20490) );
  XOR2_X1 U18161 ( .A(n20490), .B(n20491), .Z(n14568) );
  OAI21_X1 U18162 ( .B1(n14564), .B2(n14563), .A(n14562), .ZN(n19704) );
  NOR2_X1 U18163 ( .A1(n20479), .A2(n19704), .ZN(n14565) );
  AOI21_X1 U18164 ( .B1(n20479), .B2(n19704), .A(n14565), .ZN(n19708) );
  NAND2_X1 U18165 ( .A1(n19708), .A2(n19707), .ZN(n19706) );
  INV_X1 U18166 ( .A(n14565), .ZN(n14566) );
  NAND2_X1 U18167 ( .A1(n19706), .A2(n14566), .ZN(n14567) );
  NAND2_X1 U18168 ( .A1(n14568), .A2(n14567), .ZN(n16469) );
  OAI21_X1 U18169 ( .B1(n14568), .B2(n14567), .A(n16469), .ZN(n14569) );
  NAND2_X1 U18170 ( .A1(n14569), .A2(n19709), .ZN(n14571) );
  AOI22_X1 U18171 ( .A1(n19705), .A2(n20490), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n16451), .ZN(n14570) );
  OAI211_X1 U18172 ( .C1(n14572), .C2(n19713), .A(n14571), .B(n14570), .ZN(
        P2_U2917) );
  XNOR2_X1 U18173 ( .A(n14573), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14576) );
  INV_X1 U18174 ( .A(n14574), .ZN(n14575) );
  NOR2_X1 U18175 ( .A1(n14576), .A2(n14575), .ZN(n20704) );
  AOI21_X1 U18176 ( .B1(n14576), .B2(n14575), .A(n20704), .ZN(n20730) );
  NAND2_X1 U18177 ( .A1(n20730), .A2(n20710), .ZN(n14580) );
  NAND2_X1 U18178 ( .A1(n20718), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20726) );
  OAI21_X1 U18179 ( .B1(n15577), .B2(n14577), .A(n20726), .ZN(n14578) );
  AOI21_X1 U18180 ( .B1(n20607), .B2(n15586), .A(n14578), .ZN(n14579) );
  OAI211_X1 U18181 ( .C1(n20770), .C2(n20609), .A(n14580), .B(n14579), .ZN(
        P1_U2996) );
  OAI21_X1 U18182 ( .B1(n14583), .B2(n14582), .A(n14581), .ZN(n16834) );
  INV_X1 U18183 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19720) );
  INV_X1 U18184 ( .A(n16363), .ZN(n14584) );
  OAI222_X1 U18185 ( .A1(n16834), .A2(n16475), .B1(n14604), .B2(n19720), .C1(
        n19713), .C2(n14584), .ZN(P2_U2906) );
  XNOR2_X1 U18186 ( .A(n14587), .B(n14585), .ZN(n16848) );
  INV_X1 U18187 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19722) );
  INV_X1 U18188 ( .A(n16370), .ZN(n14586) );
  OAI222_X1 U18189 ( .A1(n16848), .A2(n16475), .B1(n14604), .B2(n19722), .C1(
        n14586), .C2(n19713), .ZN(P2_U2907) );
  INV_X1 U18190 ( .A(n14587), .ZN(n14588) );
  AOI21_X1 U18191 ( .B1(n14590), .B2(n14589), .A(n14588), .ZN(n16860) );
  INV_X1 U18192 ( .A(n16860), .ZN(n14592) );
  INV_X1 U18193 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19724) );
  INV_X1 U18194 ( .A(n16378), .ZN(n14591) );
  OAI222_X1 U18195 ( .A1(n14592), .A2(n16475), .B1(n14604), .B2(n19724), .C1(
        n19713), .C2(n14591), .ZN(P2_U2908) );
  XNOR2_X1 U18196 ( .A(n14593), .B(n14594), .ZN(n16199) );
  INV_X1 U18197 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19733) );
  INV_X1 U18198 ( .A(n19840), .ZN(n14595) );
  OAI222_X1 U18199 ( .A1(n16199), .A2(n16475), .B1(n19733), .B2(n14604), .C1(
        n19713), .C2(n14595), .ZN(P2_U2913) );
  NOR2_X1 U18200 ( .A1(n14596), .A2(n14597), .ZN(n16063) );
  AOI21_X1 U18201 ( .B1(n14597), .B2(n14596), .A(n16063), .ZN(n16805) );
  INV_X1 U18202 ( .A(n16805), .ZN(n16084) );
  OAI222_X1 U18203 ( .A1(n16084), .A2(n16475), .B1(n14604), .B2(n13937), .C1(
        n14598), .C2(n19713), .ZN(P2_U2904) );
  OAI21_X1 U18204 ( .B1(n14516), .B2(n14599), .A(n11517), .ZN(n16875) );
  INV_X1 U18205 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19728) );
  INV_X1 U18206 ( .A(n16393), .ZN(n14600) );
  OAI222_X1 U18207 ( .A1(n16875), .A2(n16475), .B1(n14604), .B2(n19728), .C1(
        n19713), .C2(n14600), .ZN(P2_U2910) );
  OAI21_X1 U18208 ( .B1(n14602), .B2(n14601), .A(n14517), .ZN(n16895) );
  INV_X1 U18209 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n21790) );
  INV_X1 U18210 ( .A(n19849), .ZN(n14603) );
  OAI222_X1 U18211 ( .A1(n16895), .A2(n16475), .B1(n21790), .B2(n14604), .C1(
        n19713), .C2(n14603), .ZN(P2_U2912) );
  NOR2_X1 U18212 ( .A1(n17045), .A2(n20520), .ZN(n17042) );
  NAND2_X1 U18213 ( .A1(n17044), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14607) );
  NAND2_X1 U18214 ( .A1(n14608), .A2(n14607), .ZN(n20517) );
  AOI21_X1 U18215 ( .B1(n17019), .B2(n17044), .A(n20517), .ZN(n14616) );
  INV_X1 U18216 ( .A(n17041), .ZN(n14610) );
  NAND2_X1 U18217 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20508), .ZN(n19859) );
  NOR2_X1 U18218 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19859), .ZN(n14609) );
  NAND2_X1 U18219 ( .A1(n14609), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15040) );
  OAI211_X1 U18220 ( .C1(n20501), .C2(n14611), .A(n14610), .B(n15040), .ZN(
        n14613) );
  NOR2_X1 U18221 ( .A1(n17045), .A2(n17044), .ZN(n14612) );
  AOI211_X1 U18222 ( .C1(n17047), .C2(n14614), .A(n14613), .B(n14612), .ZN(
        n14615) );
  OAI21_X1 U18223 ( .B1(n17042), .B2(n14616), .A(n14615), .ZN(P2_U3176) );
  INV_X1 U18224 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14626) );
  OR2_X1 U18225 ( .A1(n9738), .A2(n14635), .ZN(n14637) );
  AOI21_X1 U18226 ( .B1(n14618), .B2(n14637), .A(n14617), .ZN(n16801) );
  NAND2_X1 U18227 ( .A1(n16801), .A2(n16350), .ZN(n14625) );
  INV_X1 U18228 ( .A(n14639), .ZN(n14623) );
  INV_X1 U18229 ( .A(n14622), .ZN(n14620) );
  NOR2_X1 U18230 ( .A1(n14639), .A2(n14620), .ZN(n14662) );
  INV_X1 U18231 ( .A(n14662), .ZN(n14621) );
  OAI211_X1 U18232 ( .C1(n14623), .C2(n14622), .A(n14621), .B(n16357), .ZN(
        n14624) );
  OAI211_X1 U18233 ( .C1(n16350), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        P2_U2872) );
  INV_X1 U18234 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20627) );
  NOR2_X1 U18235 ( .A1(n20576), .A2(n20627), .ZN(n20740) );
  NOR2_X1 U18236 ( .A1(n15577), .A2(n14627), .ZN(n14628) );
  AOI211_X1 U18237 ( .C1(n15586), .C2(n20624), .A(n20740), .B(n14628), .ZN(
        n14633) );
  OR2_X1 U18238 ( .A1(n14630), .A2(n14629), .ZN(n20739) );
  NAND3_X1 U18239 ( .A1(n20739), .A2(n14631), .A3(n20710), .ZN(n14632) );
  OAI211_X1 U18240 ( .C1(n14634), .C2(n20770), .A(n14633), .B(n14632), .ZN(
        P1_U2997) );
  NAND2_X1 U18241 ( .A1(n9738), .A2(n14635), .ZN(n14636) );
  NAND2_X1 U18242 ( .A1(n14637), .A2(n14636), .ZN(n16821) );
  NOR2_X1 U18243 ( .A1(n14643), .A2(n14638), .ZN(n14644) );
  OAI211_X1 U18244 ( .C1(n14644), .C2(n14640), .A(n16357), .B(n14639), .ZN(
        n14642) );
  NAND2_X1 U18245 ( .A1(n16360), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14641) );
  OAI211_X1 U18246 ( .C1(n16360), .C2(n16821), .A(n14642), .B(n14641), .ZN(
        P2_U2873) );
  INV_X1 U18247 ( .A(n14643), .ZN(n14647) );
  INV_X1 U18248 ( .A(n14644), .ZN(n14645) );
  OAI211_X1 U18249 ( .C1(n14647), .C2(n14646), .A(n14645), .B(n16357), .ZN(
        n14651) );
  OR2_X1 U18250 ( .A1(n14548), .A2(n14648), .ZN(n14649) );
  NAND2_X1 U18251 ( .A1(n16832), .A2(n16350), .ZN(n14650) );
  OAI211_X1 U18252 ( .C1(n16350), .C2(n16101), .A(n14651), .B(n14650), .ZN(
        P2_U2874) );
  OR2_X1 U18253 ( .A1(n14653), .A2(n14652), .ZN(n14654) );
  NAND2_X1 U18254 ( .A1(n14543), .A2(n14654), .ZN(n16883) );
  NOR2_X1 U18255 ( .A1(n16883), .A2(n16360), .ZN(n14659) );
  AOI211_X1 U18256 ( .C1(n14657), .C2(n14656), .A(n16353), .B(n14655), .ZN(
        n14658) );
  AOI211_X1 U18257 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n16360), .A(n14659), .B(
        n14658), .ZN(n14660) );
  INV_X1 U18258 ( .A(n14660), .ZN(P2_U2879) );
  NAND2_X1 U18259 ( .A1(n14662), .A2(n14661), .ZN(n16355) );
  OAI21_X1 U18260 ( .B1(n14662), .B2(n14661), .A(n16355), .ZN(n16463) );
  NOR2_X1 U18261 ( .A1(n14617), .A2(n14664), .ZN(n14665) );
  OR2_X1 U18262 ( .A1(n14663), .A2(n14665), .ZN(n16788) );
  MUX2_X1 U18263 ( .A(n16788), .B(n14666), .S(n16360), .Z(n14667) );
  OAI21_X1 U18264 ( .B1(n16353), .B2(n16463), .A(n14667), .ZN(P2_U2871) );
  XNOR2_X1 U18265 ( .A(n14669), .B(n14668), .ZN(n14670) );
  NOR2_X1 U18266 ( .A1(n14670), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20755) );
  INV_X1 U18267 ( .A(n14670), .ZN(n14671) );
  NOR2_X1 U18268 ( .A1(n14671), .A2(n20767), .ZN(n20754) );
  NOR3_X1 U18269 ( .A1(n20755), .A2(n20754), .A3(n20537), .ZN(n14673) );
  AND2_X1 U18270 ( .A1(n20718), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20763) );
  MUX2_X1 U18271 ( .A(n15586), .B(n20703), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14672) );
  NOR3_X1 U18272 ( .A1(n14673), .A2(n20763), .A3(n14672), .ZN(n14674) );
  OAI21_X1 U18273 ( .B1(n20770), .B2(n15360), .A(n14674), .ZN(P1_U2998) );
  OR2_X1 U18274 ( .A1(n14675), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14679) );
  NAND2_X1 U18275 ( .A1(n14676), .A2(n14679), .ZN(n19474) );
  NOR2_X1 U18276 ( .A1(n17869), .A2(n19474), .ZN(n14678) );
  MUX2_X1 U18277 ( .A(n14678), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n14677), .Z(P3_U3284) );
  OR2_X1 U18278 ( .A1(n14679), .A2(n18207), .ZN(n19022) );
  NOR2_X1 U18279 ( .A1(n19022), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(n14681) );
  NAND2_X1 U18280 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U18281 ( .B1(n14681), .B2(n19606), .A(n19312), .ZN(n19027) );
  INV_X1 U18282 ( .A(n19027), .ZN(n14682) );
  NAND2_X1 U18283 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18691) );
  NAND2_X1 U18284 ( .A1(n19608), .A2(n19020), .ZN(n19620) );
  NOR2_X1 U18285 ( .A1(n18647), .A2(n19620), .ZN(n17258) );
  AOI21_X1 U18286 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17258), .ZN(n17259) );
  NOR2_X1 U18287 ( .A1(n14682), .A2(n17259), .ZN(n14684) );
  NOR2_X1 U18288 ( .A1(n19608), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19069) );
  OR2_X1 U18289 ( .A1(n19069), .A2(n14682), .ZN(n17257) );
  OR2_X1 U18290 ( .A1(n19090), .A2(n17257), .ZN(n14683) );
  MUX2_X1 U18291 ( .A(n14684), .B(n14683), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND3_X1 U18292 ( .A1(n14686), .A2(n13524), .A3(n14685), .ZN(n14691) );
  NOR2_X1 U18293 ( .A1(n14688), .A2(n14687), .ZN(n19470) );
  NAND2_X1 U18294 ( .A1(n19470), .A2(n19464), .ZN(n14689) );
  NAND2_X1 U18295 ( .A1(n14691), .A2(n18760), .ZN(n14707) );
  NOR2_X1 U18296 ( .A1(n18792), .A2(n18725), .ZN(n18623) );
  OAI22_X1 U18297 ( .A1(n17211), .A2(n18701), .B1(n17210), .B2(n18700), .ZN(
        n17120) );
  NOR2_X1 U18298 ( .A1(n14698), .A2(n17120), .ZN(n14693) );
  NAND2_X1 U18299 ( .A1(n18694), .A2(n18772), .ZN(n18615) );
  OAI21_X1 U18300 ( .B1(n14694), .B2(n18648), .A(n18772), .ZN(n14695) );
  AOI21_X1 U18301 ( .B1(n18647), .B2(n11577), .A(n14695), .ZN(n17117) );
  OAI21_X1 U18302 ( .B1(n18615), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17117), .ZN(n17103) );
  NOR2_X1 U18303 ( .A1(n18830), .A2(n9962), .ZN(n18798) );
  OR2_X1 U18304 ( .A1(n13537), .A2(n18701), .ZN(n14696) );
  NAND2_X1 U18305 ( .A1(n18551), .A2(n14697), .ZN(n17104) );
  NOR3_X1 U18306 ( .A1(n17104), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n14698), .ZN(n14705) );
  AND2_X1 U18307 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18620), .ZN(
        n14699) );
  OR2_X1 U18308 ( .A1(n19409), .A2(n14699), .ZN(n18650) );
  NOR2_X1 U18309 ( .A1(n11577), .A2(n18593), .ZN(n17107) );
  OAI211_X1 U18310 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17107), .B(n14700), .ZN(n14702) );
  NAND2_X1 U18311 ( .A1(n9696), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n14701) );
  OAI211_X1 U18312 ( .C1(n18696), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14704) );
  AOI211_X1 U18313 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17103), .A(
        n14705), .B(n14704), .ZN(n14706) );
  OAI211_X1 U18314 ( .C1(n14708), .C2(n14707), .A(n9751), .B(n14706), .ZN(
        P3_U2802) );
  NAND2_X1 U18315 ( .A1(n15154), .A2(n15144), .ZN(n15143) );
  NOR2_X2 U18316 ( .A1(n15143), .A2(n14833), .ZN(n14832) );
  INV_X1 U18317 ( .A(n14709), .ZN(n14710) );
  NOR2_X1 U18318 ( .A1(n14832), .A2(n14710), .ZN(n14712) );
  NAND2_X1 U18319 ( .A1(n14713), .A2(n20710), .ZN(n14717) );
  NOR2_X1 U18320 ( .A1(n20714), .A2(n14730), .ZN(n14714) );
  AOI211_X1 U18321 ( .C1(n20703), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14715), .B(n14714), .ZN(n14716) );
  OAI211_X1 U18322 ( .C1(n20770), .C2(n14753), .A(n14717), .B(n14716), .ZN(
        P1_U2975) );
  NAND2_X1 U18323 ( .A1(n14720), .A2(n20771), .ZN(n14960) );
  OAI22_X1 U18324 ( .A1(n15460), .A2(n15484), .B1(n15497), .B2(n14718), .ZN(
        n14719) );
  AOI21_X1 U18325 ( .B1(n15462), .B2(BUF1_REG_24__SCAN_IN), .A(n14719), .ZN(
        n14722) );
  NAND2_X1 U18326 ( .A1(n15463), .A2(DATAI_24_), .ZN(n14721) );
  OAI211_X1 U18327 ( .C1(n14753), .C2(n15501), .A(n14722), .B(n14721), .ZN(
        P1_U2880) );
  OAI222_X1 U18328 ( .A1(n14753), .A2(n15399), .B1(n14745), .B2(n20653), .C1(
        n15395), .C2(n14726), .ZN(P1_U2848) );
  INV_X1 U18329 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15509) );
  NAND2_X1 U18330 ( .A1(n14802), .A2(n14725), .ZN(n14737) );
  INV_X1 U18331 ( .A(n14726), .ZN(n14751) );
  NAND2_X1 U18332 ( .A1(n20792), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14740) );
  AND2_X1 U18333 ( .A1(n21487), .A2(n20830), .ZN(n17289) );
  NOR2_X1 U18334 ( .A1(n14740), .A2(n17289), .ZN(n14728) );
  INV_X1 U18335 ( .A(n14737), .ZN(n14729) );
  AND2_X2 U18336 ( .A1(n15056), .A2(n14729), .ZN(n20623) );
  INV_X2 U18337 ( .A(n20623), .ZN(n20620) );
  NOR2_X1 U18338 ( .A1(n20620), .A2(n14730), .ZN(n14750) );
  NOR2_X1 U18339 ( .A1(n14731), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14742) );
  INV_X1 U18340 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21419) );
  INV_X1 U18341 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21393) );
  NAND3_X1 U18342 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20597) );
  NOR2_X1 U18343 ( .A1(n21393), .A2(n20597), .ZN(n20596) );
  INV_X1 U18344 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21399) );
  INV_X1 U18345 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21398) );
  NAND2_X1 U18346 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20562) );
  NOR3_X1 U18347 ( .A1(n21399), .A2(n21398), .A3(n20562), .ZN(n15173) );
  NAND2_X1 U18348 ( .A1(n20596), .A2(n15173), .ZN(n15193) );
  AND2_X1 U18349 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15290) );
  AND2_X1 U18350 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n14732) );
  NAND2_X1 U18351 ( .A1(n15290), .A2(n14732), .ZN(n15242) );
  NAND2_X1 U18352 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14733) );
  NOR2_X1 U18353 ( .A1(n15242), .A2(n14733), .ZN(n15212) );
  NAND2_X1 U18354 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15231) );
  INV_X1 U18355 ( .A(n15231), .ZN(n14734) );
  AND2_X1 U18356 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14734), .ZN(n14735) );
  AND2_X1 U18357 ( .A1(n15212), .A2(n14735), .ZN(n15190) );
  NAND3_X1 U18358 ( .A1(n15190), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n15174) );
  NOR3_X1 U18359 ( .A1(n21419), .A2(n15193), .A3(n15174), .ZN(n15163) );
  INV_X1 U18360 ( .A(n15163), .ZN(n15135) );
  INV_X1 U18361 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21422) );
  NOR2_X1 U18362 ( .A1(n15135), .A2(n21422), .ZN(n14736) );
  NAND3_X1 U18363 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(n14736), .ZN(n15121) );
  NOR3_X1 U18364 ( .A1(n21369), .A2(n21660), .A3(n17368), .ZN(n17261) );
  NAND2_X1 U18365 ( .A1(n20576), .A2(n14737), .ZN(n14738) );
  OR2_X1 U18366 ( .A1(n17261), .A2(n14738), .ZN(n14739) );
  INV_X1 U18367 ( .A(n20561), .ZN(n20610) );
  AOI21_X1 U18368 ( .B1(n20612), .B2(n15121), .A(n20610), .ZN(n15137) );
  INV_X1 U18369 ( .A(n14740), .ZN(n14741) );
  NOR2_X1 U18370 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  AND2_X2 U18371 ( .A1(n14744), .A2(n14743), .ZN(n20622) );
  INV_X1 U18372 ( .A(n20622), .ZN(n15356) );
  NOR2_X1 U18373 ( .A1(n15356), .A2(n14745), .ZN(n14747) );
  NOR3_X1 U18374 ( .A1(n20595), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n15121), 
        .ZN(n14746) );
  AOI211_X1 U18375 ( .C1(n20625), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14747), .B(n14746), .ZN(n14748) );
  OAI21_X1 U18376 ( .B1(n15137), .B2(n21426), .A(n14748), .ZN(n14749) );
  AOI211_X1 U18377 ( .C1(n14751), .C2(n20608), .A(n14750), .B(n14749), .ZN(
        n14752) );
  OAI21_X1 U18378 ( .B1(n14753), .B2(n15350), .A(n14752), .ZN(P1_U2816) );
  NAND2_X1 U18379 ( .A1(n14755), .A2(n14754), .ZN(n14759) );
  INV_X1 U18380 ( .A(n16574), .ZN(n14757) );
  INV_X1 U18381 ( .A(n14845), .ZN(n14851) );
  NAND2_X1 U18382 ( .A1(n14850), .A2(n10038), .ZN(n14770) );
  OAI21_X1 U18383 ( .B1(n14663), .B2(n14762), .A(n14761), .ZN(n16361) );
  INV_X1 U18384 ( .A(n16361), .ZN(n14767) );
  INV_X1 U18385 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14765) );
  AOI21_X1 U18386 ( .B1(n15012), .B2(n14765), .A(n14763), .ZN(n16054) );
  NAND2_X1 U18387 ( .A1(n19771), .A2(n16054), .ZN(n14764) );
  NAND2_X1 U18388 ( .A1(n19748), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n14844) );
  OAI211_X1 U18389 ( .C1(n17388), .C2(n14765), .A(n14764), .B(n14844), .ZN(
        n14766) );
  AOI21_X1 U18390 ( .B1(n14767), .B2(n19787), .A(n14766), .ZN(n14768) );
  INV_X1 U18391 ( .A(n14768), .ZN(n14769) );
  OAI21_X1 U18392 ( .B1(n14857), .B2(n19785), .A(n14771), .ZN(P2_U2997) );
  INV_X1 U18393 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14813) );
  OAI22_X1 U18394 ( .A1(n14772), .A2(n15395), .B1(n20653), .B2(n14813), .ZN(
        P1_U2841) );
  XNOR2_X1 U18395 ( .A(n14773), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15507) );
  AOI22_X1 U18396 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14781) );
  AOI22_X1 U18397 ( .A1(n14774), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14780) );
  AOI22_X1 U18398 ( .A1(n14776), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14775), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14779) );
  AOI22_X1 U18399 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11912), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14778) );
  NAND4_X1 U18400 ( .A1(n14781), .A2(n14780), .A3(n14779), .A4(n14778), .ZN(
        n14790) );
  AOI22_X1 U18401 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14782), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14788) );
  AOI22_X1 U18402 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11812), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14787) );
  AOI22_X1 U18403 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12596), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U18404 ( .A1(n14784), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14783), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14785) );
  NAND4_X1 U18405 ( .A1(n14788), .A2(n14787), .A3(n14786), .A4(n14785), .ZN(
        n14789) );
  NOR2_X1 U18406 ( .A1(n14790), .A2(n14789), .ZN(n14794) );
  NOR2_X1 U18407 ( .A1(n14792), .A2(n14791), .ZN(n14793) );
  XNOR2_X1 U18408 ( .A(n14794), .B(n14793), .ZN(n14800) );
  NAND2_X1 U18409 ( .A1(n21306), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14795) );
  OAI211_X1 U18410 ( .C1(n14797), .C2(n14236), .A(n14796), .B(n14795), .ZN(
        n14798) );
  AOI21_X1 U18411 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n14801) );
  AOI21_X1 U18412 ( .B1(n15507), .B2(n14802), .A(n14801), .ZN(n14952) );
  NAND2_X1 U18413 ( .A1(n14951), .A2(n14952), .ZN(n14806) );
  AOI22_X1 U18414 ( .A1(n12320), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14803), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14804) );
  INV_X1 U18415 ( .A(n14804), .ZN(n14805) );
  XNOR2_X2 U18416 ( .A(n14806), .B(n14805), .ZN(n15058) );
  NAND2_X1 U18417 ( .A1(n15058), .A2(n20582), .ZN(n14818) );
  INV_X1 U18418 ( .A(n15361), .ZN(n14811) );
  NAND2_X1 U18419 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14814) );
  INV_X1 U18420 ( .A(n14814), .ZN(n14810) );
  NAND2_X1 U18421 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14807) );
  NOR2_X1 U18422 ( .A1(n15121), .A2(n14807), .ZN(n15113) );
  NAND2_X1 U18423 ( .A1(n15113), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15097) );
  INV_X1 U18424 ( .A(n15097), .ZN(n14808) );
  NAND2_X1 U18425 ( .A1(n20561), .A2(n14808), .ZN(n15114) );
  NAND2_X1 U18426 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14809) );
  OAI21_X1 U18427 ( .B1(n15114), .B2(n14809), .A(n15361), .ZN(n15073) );
  OAI21_X1 U18428 ( .B1(n14811), .B2(n14810), .A(n15073), .ZN(n15065) );
  OAI22_X1 U18429 ( .A1(n15356), .A2(n14813), .B1(n14812), .B2(n20588), .ZN(
        n14816) );
  INV_X1 U18430 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21431) );
  NOR3_X1 U18431 ( .A1(n20595), .A2(n21431), .A3(n15097), .ZN(n15088) );
  NAND2_X1 U18432 ( .A1(n15088), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15075) );
  NOR3_X1 U18433 ( .A1(n15075), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14814), 
        .ZN(n14815) );
  AOI211_X1 U18434 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n15065), .A(n14816), 
        .B(n14815), .ZN(n14817) );
  OAI211_X1 U18435 ( .C1(n14772), .C2(n20638), .A(n14818), .B(n14817), .ZN(
        P1_U2809) );
  XNOR2_X1 U18436 ( .A(n15641), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14819) );
  XNOR2_X1 U18437 ( .A(n15514), .B(n14819), .ZN(n14839) );
  INV_X1 U18438 ( .A(n14820), .ZN(n14825) );
  INV_X1 U18439 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14821) );
  NOR2_X1 U18440 ( .A1(n20576), .A2(n14821), .ZN(n14834) );
  NOR2_X1 U18441 ( .A1(n14822), .A2(n14824), .ZN(n14823) );
  AOI211_X1 U18442 ( .C1(n14825), .C2(n14824), .A(n14834), .B(n14823), .ZN(
        n14831) );
  INV_X1 U18443 ( .A(n15161), .ZN(n15150) );
  OAI21_X1 U18444 ( .B1(n15150), .B2(n15149), .A(n14826), .ZN(n14828) );
  INV_X1 U18445 ( .A(n15130), .ZN(n14827) );
  NAND2_X1 U18446 ( .A1(n14828), .A2(n14827), .ZN(n15378) );
  INV_X1 U18447 ( .A(n15378), .ZN(n14829) );
  NAND2_X1 U18448 ( .A1(n14829), .A2(n20742), .ZN(n14830) );
  OAI211_X1 U18449 ( .C1(n14839), .C2(n20753), .A(n14831), .B(n14830), .ZN(
        P1_U3008) );
  AOI21_X1 U18450 ( .B1(n14833), .B2(n15143), .A(n14832), .ZN(n15377) );
  INV_X1 U18451 ( .A(n15140), .ZN(n14836) );
  AOI21_X1 U18452 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14834), .ZN(n14835) );
  OAI21_X1 U18453 ( .B1(n20714), .B2(n14836), .A(n14835), .ZN(n14837) );
  OAI21_X1 U18454 ( .B1(n14839), .B2(n20537), .A(n14838), .ZN(P1_U2976) );
  AND2_X1 U18455 ( .A1(n14527), .A2(n14841), .ZN(n16065) );
  OR2_X1 U18456 ( .A1(n16065), .A2(n14842), .ZN(n14843) );
  OAI21_X1 U18457 ( .B1(n16361), .B2(n19803), .A(n14844), .ZN(n14847) );
  NOR2_X1 U18458 ( .A1(n16868), .A2(n14845), .ZN(n16796) );
  INV_X1 U18459 ( .A(n16796), .ZN(n14846) );
  INV_X1 U18460 ( .A(n19801), .ZN(n14848) );
  NOR2_X1 U18461 ( .A1(n17406), .A2(n14851), .ZN(n14852) );
  NOR2_X1 U18462 ( .A1(n16872), .A2(n14852), .ZN(n16800) );
  AND2_X1 U18463 ( .A1(n16800), .A2(n10387), .ZN(n14853) );
  NOR2_X1 U18464 ( .A1(n17406), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14854) );
  OAI21_X1 U18465 ( .B1(n16792), .B2(n14854), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14855) );
  OAI211_X1 U18466 ( .C1(n14857), .C2(n17400), .A(n14856), .B(n14855), .ZN(
        P2_U3029) );
  NAND2_X1 U18467 ( .A1(n14859), .A2(n14858), .ZN(n14860) );
  XNOR2_X1 U18468 ( .A(n14860), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14875) );
  XOR2_X1 U18469 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n14861), .Z(
        n16668) );
  XOR2_X1 U18470 ( .A(n16667), .B(n16668), .Z(n14873) );
  NAND2_X1 U18471 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19748), .ZN(n14862) );
  OAI21_X1 U18472 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14863), .A(
        n14862), .ZN(n14864) );
  AOI21_X1 U18473 ( .B1(n16197), .B2(n16967), .A(n14864), .ZN(n14866) );
  NAND2_X1 U18474 ( .A1(n16902), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14865) );
  OAI211_X1 U18475 ( .C1(n16958), .C2(n16199), .A(n14866), .B(n14865), .ZN(
        n14867) );
  AOI21_X1 U18476 ( .B1(n14873), .B2(n11071), .A(n14867), .ZN(n14868) );
  OAI21_X1 U18477 ( .B1(n14875), .B2(n16942), .A(n14868), .ZN(P2_U3040) );
  INV_X1 U18478 ( .A(n16197), .ZN(n14871) );
  OAI21_X1 U18479 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9712), .A(
        n14996), .ZN(n16184) );
  OAI22_X1 U18480 ( .A1(n20420), .A2(n11468), .B1(n19758), .B2(n16184), .ZN(
        n14869) );
  AOI21_X1 U18481 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14869), .ZN(n14870) );
  OAI21_X1 U18482 ( .B1(n14871), .B2(n19774), .A(n14870), .ZN(n14872) );
  AOI21_X1 U18483 ( .B1(n14873), .B2(n19763), .A(n14872), .ZN(n14874) );
  OAI21_X1 U18484 ( .B1(n14875), .B2(n16690), .A(n14874), .ZN(P2_U3008) );
  AOI21_X1 U18485 ( .B1(n15086), .B2(n14876), .A(n15062), .ZN(n15371) );
  INV_X1 U18486 ( .A(n14877), .ZN(n14882) );
  INV_X1 U18487 ( .A(n14878), .ZN(n14880) );
  NAND3_X1 U18488 ( .A1(n15714), .A2(n15706), .A3(n14881), .ZN(n14879) );
  OAI211_X1 U18489 ( .C1(n14882), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14883) );
  AOI21_X1 U18490 ( .B1(n15371), .B2(n20742), .A(n14883), .ZN(n14884) );
  OAI21_X1 U18491 ( .B1(n14885), .B2(n20753), .A(n14884), .ZN(P1_U3002) );
  NOR2_X1 U18492 ( .A1(n14889), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14890) );
  MUX2_X1 U18493 ( .A(n14891), .B(n14890), .S(n9699), .Z(n15047) );
  NAND2_X1 U18494 ( .A1(n15047), .A2(n11177), .ZN(n14892) );
  XNOR2_X1 U18495 ( .A(n14892), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14893) );
  XNOR2_X1 U18496 ( .A(n14894), .B(n14893), .ZN(n14977) );
  INV_X1 U18497 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n21704) );
  AOI22_X1 U18498 ( .A1(n14895), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14896) );
  AOI21_X1 U18499 ( .B1(n14898), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14897), .ZN(n14899) );
  INV_X1 U18500 ( .A(n15053), .ZN(n16280) );
  INV_X1 U18501 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14901) );
  NOR2_X1 U18502 ( .A1(n11468), .A2(n21704), .ZN(n14970) );
  AOI21_X1 U18503 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14970), .ZN(n14902) );
  OAI21_X1 U18504 ( .B1(n19758), .B2(n14986), .A(n14902), .ZN(n14903) );
  AOI21_X1 U18505 ( .B1(n16280), .B2(n19787), .A(n14903), .ZN(n14906) );
  NAND2_X1 U18506 ( .A1(n16485), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14904) );
  NAND2_X1 U18507 ( .A1(n14974), .A2(n19781), .ZN(n14905) );
  OAI211_X1 U18508 ( .C1(n14977), .C2(n19785), .A(n14906), .B(n14905), .ZN(
        P2_U2983) );
  NAND2_X1 U18509 ( .A1(n14907), .A2(n19781), .ZN(n14914) );
  XNOR2_X1 U18510 ( .A(n14908), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15909) );
  AOI21_X1 U18511 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14909), .ZN(n14910) );
  OAI21_X1 U18512 ( .B1(n19758), .B2(n15909), .A(n14910), .ZN(n14911) );
  AOI21_X1 U18513 ( .B1(n14912), .B2(n19787), .A(n14911), .ZN(n14913) );
  OAI211_X1 U18514 ( .C1(n14915), .C2(n19785), .A(n14914), .B(n14913), .ZN(
        P2_U2984) );
  AOI21_X1 U18515 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14916), .ZN(n14919) );
  NOR2_X1 U18516 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n14991), .ZN(
        n14917) );
  NOR2_X1 U18517 ( .A1(n15015), .A2(n14917), .ZN(n16019) );
  NAND2_X1 U18518 ( .A1(n19771), .A2(n16019), .ZN(n14918) );
  OAI211_X1 U18519 ( .C1(n16333), .C2(n19774), .A(n14919), .B(n14918), .ZN(
        n14920) );
  AOI21_X1 U18520 ( .B1(n9755), .B2(n19781), .A(n14920), .ZN(n14921) );
  OAI21_X1 U18521 ( .B1(n14922), .B2(n19785), .A(n14921), .ZN(P2_U2993) );
  INV_X1 U18522 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14929) );
  INV_X1 U18523 ( .A(n14924), .ZN(n14923) );
  NAND2_X1 U18524 ( .A1(n14923), .A2(n17029), .ZN(n16418) );
  NAND2_X1 U18525 ( .A1(n16415), .A2(BUF2_REG_30__SCAN_IN), .ZN(n14928) );
  AOI22_X1 U18526 ( .A1(n16459), .A2(n14926), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n16451), .ZN(n14927) );
  OAI211_X1 U18527 ( .C1(n14929), .C2(n16418), .A(n14928), .B(n14927), .ZN(
        n14930) );
  AOI21_X1 U18528 ( .B1(n15908), .B2(n19705), .A(n14930), .ZN(n14931) );
  OAI21_X1 U18529 ( .B1(n14932), .B2(n16462), .A(n14931), .ZN(P2_U2889) );
  INV_X1 U18530 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14933) );
  NAND2_X1 U18531 ( .A1(n9725), .A2(n14933), .ZN(n14934) );
  NAND2_X1 U18532 ( .A1(n9789), .A2(n14934), .ZN(n16034) );
  NAND2_X1 U18533 ( .A1(n16038), .A2(n19787), .ZN(n14937) );
  AOI21_X1 U18534 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14935), .ZN(n14936) );
  OAI211_X1 U18535 ( .C1(n19758), .C2(n16034), .A(n14937), .B(n14936), .ZN(
        n14938) );
  OAI21_X1 U18536 ( .B1(n14940), .B2(n19785), .A(n14939), .ZN(P2_U2995) );
  NOR2_X1 U18537 ( .A1(n14941), .A2(n9866), .ZN(n17263) );
  NOR3_X1 U18538 ( .A1(n14942), .A2(n17370), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14943) );
  AOI21_X1 U18539 ( .B1(n14944), .B2(n17263), .A(n14943), .ZN(n14950) );
  INV_X1 U18540 ( .A(n20893), .ZN(n14946) );
  OAI22_X1 U18541 ( .A1(n14946), .A2(n14945), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11945), .ZN(n17262) );
  AOI22_X1 U18542 ( .A1(n14948), .A2(n9866), .B1(n14947), .B2(n17262), .ZN(
        n14949) );
  OAI211_X1 U18543 ( .C1(n9866), .C2(n21457), .A(n14950), .B(n14949), .ZN(
        P1_U3474) );
  XOR2_X1 U18544 ( .A(n14952), .B(n14951), .Z(n15511) );
  INV_X1 U18545 ( .A(n15511), .ZN(n15370) );
  OAI22_X1 U18546 ( .A1(n15460), .A2(n15469), .B1(n15497), .B2(n14236), .ZN(
        n14953) );
  AOI21_X1 U18547 ( .B1(n15462), .B2(BUF1_REG_30__SCAN_IN), .A(n14953), .ZN(
        n14955) );
  NAND2_X1 U18548 ( .A1(n15463), .A2(DATAI_30_), .ZN(n14954) );
  OAI211_X1 U18549 ( .C1(n15370), .C2(n15501), .A(n14955), .B(n14954), .ZN(
        P1_U2874) );
  INV_X1 U18550 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n21659) );
  NAND3_X1 U18551 ( .A1(n15058), .A2(n14956), .A3(n15497), .ZN(n14959) );
  AOI22_X1 U18552 ( .A1(n15463), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14957), .ZN(n14958) );
  OAI211_X1 U18553 ( .C1(n14960), .C2(n21659), .A(n14959), .B(n14958), .ZN(
        P1_U2873) );
  AOI222_X1 U18554 ( .A1(n14962), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14961), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11138), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14963) );
  XNOR2_X1 U18555 ( .A(n14964), .B(n14963), .ZN(n15050) );
  NAND2_X1 U18556 ( .A1(n15050), .A2(n19705), .ZN(n14966) );
  AOI22_X1 U18557 ( .A1(n16415), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n16451), .ZN(n14965) );
  OAI211_X1 U18558 ( .C1(n16418), .C2(n21659), .A(n14966), .B(n14965), .ZN(
        P2_U2888) );
  OAI21_X1 U18559 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17406), .A(
        n14967), .ZN(n14971) );
  NOR4_X1 U18560 ( .A1(n16693), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11114), .A4(n14968), .ZN(n14969) );
  AOI211_X1 U18561 ( .C1(n14971), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14970), .B(n14969), .ZN(n14972) );
  OAI21_X1 U18562 ( .B1(n15053), .B2(n19803), .A(n14972), .ZN(n14973) );
  AOI21_X1 U18563 ( .B1(n19792), .B2(n15050), .A(n14973), .ZN(n14976) );
  NAND2_X1 U18564 ( .A1(n14974), .A2(n19796), .ZN(n14975) );
  OAI211_X1 U18565 ( .C1(n14977), .C2(n17400), .A(n14976), .B(n14975), .ZN(
        P2_U3015) );
  NAND2_X1 U18566 ( .A1(n20520), .A2(n20512), .ZN(n14981) );
  INV_X1 U18567 ( .A(n14981), .ZN(n14978) );
  NAND2_X1 U18568 ( .A1(n14979), .A2(n14978), .ZN(n14980) );
  NAND2_X1 U18569 ( .A1(n14981), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14982) );
  NOR2_X1 U18570 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  INV_X1 U18571 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14985) );
  NOR2_X1 U18572 ( .A1(n14989), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14987) );
  OR2_X1 U18573 ( .A1(n14908), .A2(n14987), .ZN(n16482) );
  NOR2_X1 U18574 ( .A1(n15024), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14988) );
  OR2_X1 U18575 ( .A1(n14989), .A2(n14988), .ZN(n16492) );
  INV_X1 U18576 ( .A(n16492), .ZN(n15028) );
  INV_X1 U18577 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14990) );
  NAND2_X1 U18578 ( .A1(n9789), .A2(n14990), .ZN(n14993) );
  AND2_X1 U18579 ( .A1(n14993), .A2(n14992), .ZN(n19670) );
  NOR2_X1 U18580 ( .A1(n19670), .A2(n16019), .ZN(n15014) );
  AOI21_X1 U18581 ( .B1(n15010), .B2(n16590), .A(n15013), .ZN(n16588) );
  NOR2_X1 U18582 ( .A1(n14994), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14995) );
  OR2_X1 U18583 ( .A1(n15006), .A2(n14995), .ZN(n16637) );
  INV_X1 U18584 ( .A(n16637), .ZN(n16119) );
  AND2_X1 U18585 ( .A1(n14996), .A2(n16684), .ZN(n14997) );
  NOR2_X1 U18586 ( .A1(n15001), .A2(n14997), .ZN(n16686) );
  AOI21_X1 U18587 ( .B1(n16201), .B2(n14999), .A(n9712), .ZN(n17374) );
  AOI21_X1 U18588 ( .B1(n17389), .B2(n14998), .A(n15000), .ZN(n17380) );
  MUX2_X1 U18589 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16995) );
  MUX2_X1 U18590 ( .A(n16264), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n16259) );
  OAI21_X1 U18591 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n14998), .ZN(n19769) );
  OAI21_X1 U18592 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n15000), .A(
        n14999), .ZN(n19757) );
  NOR2_X1 U18593 ( .A1(n17374), .A2(n16204), .ZN(n16182) );
  OR2_X1 U18594 ( .A1(n15001), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15002) );
  NAND2_X1 U18595 ( .A1(n15004), .A2(n15002), .ZN(n16672) );
  INV_X1 U18596 ( .A(n16672), .ZN(n16164) );
  NAND2_X1 U18597 ( .A1(n15004), .A2(n15003), .ZN(n15005) );
  NAND2_X1 U18598 ( .A1(n9733), .A2(n15005), .ZN(n16652) );
  INV_X1 U18599 ( .A(n16652), .ZN(n16147) );
  NAND2_X1 U18600 ( .A1(n16129), .A2(n16130), .ZN(n16117) );
  OR2_X1 U18601 ( .A1(n15006), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15007) );
  NAND2_X1 U18602 ( .A1(n9778), .A2(n15007), .ZN(n16627) );
  NAND2_X1 U18603 ( .A1(n16108), .A2(n16627), .ZN(n16096) );
  AND2_X1 U18604 ( .A1(n9778), .A2(n15008), .ZN(n15009) );
  OR2_X1 U18605 ( .A1(n15011), .A2(n15009), .ZN(n16613) );
  INV_X1 U18606 ( .A(n16613), .ZN(n16098) );
  OAI21_X1 U18607 ( .B1(n15011), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15010), .ZN(n16601) );
  OAI21_X1 U18608 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15013), .A(
        n15012), .ZN(n16070) );
  INV_X1 U18609 ( .A(n15015), .ZN(n15016) );
  NAND2_X1 U18610 ( .A1(n15016), .A2(n10277), .ZN(n15017) );
  AND2_X1 U18611 ( .A1(n15017), .A2(n15018), .ZN(n16011) );
  AND2_X1 U18612 ( .A1(n15018), .A2(n16530), .ZN(n15019) );
  NOR2_X1 U18613 ( .A1(n9793), .A2(n15019), .ZN(n16528) );
  OR2_X1 U18614 ( .A1(n15992), .A2(n16528), .ZN(n15981) );
  OR2_X1 U18615 ( .A1(n9793), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15020) );
  AND2_X1 U18616 ( .A1(n15021), .A2(n15020), .ZN(n16519) );
  NAND2_X1 U18617 ( .A1(n15021), .A2(n15970), .ZN(n15022) );
  NAND2_X1 U18618 ( .A1(n15023), .A2(n15022), .ZN(n16511) );
  INV_X1 U18619 ( .A(n15024), .ZN(n15027) );
  NAND2_X1 U18620 ( .A1(n15025), .A2(n15944), .ZN(n15026) );
  NAND2_X1 U18621 ( .A1(n15027), .A2(n15026), .ZN(n16502) );
  AOI21_X1 U18622 ( .B1(n15946), .B2(n16502), .A(n17002), .ZN(n15928) );
  OAI211_X1 U18623 ( .C1(n17002), .C2(n16482), .A(n15920), .B(n15909), .ZN(
        n15911) );
  INV_X1 U18624 ( .A(n15029), .ZN(n15031) );
  NOR2_X1 U18625 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15030) );
  NOR2_X1 U18626 ( .A1(n15911), .A2(n16219), .ZN(n15046) );
  INV_X1 U18627 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15044) );
  INV_X1 U18628 ( .A(n15032), .ZN(n15035) );
  OAI21_X1 U18629 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20509), .A(n15044), 
        .ZN(n15033) );
  INV_X1 U18630 ( .A(n15033), .ZN(n15034) );
  NAND2_X1 U18631 ( .A1(n15035), .A2(n15034), .ZN(n15036) );
  NAND2_X1 U18632 ( .A1(n15037), .A2(n15036), .ZN(n15039) );
  INV_X1 U18633 ( .A(n15048), .ZN(n15038) );
  AND3_X1 U18634 ( .A1(n11468), .A2(n17049), .A3(n15040), .ZN(n15041) );
  AND2_X2 U18635 ( .A1(n19664), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19671) );
  AOI22_X1 U18636 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        n16249), .B2(P2_REIP_REG_31__SCAN_IN), .ZN(n15043) );
  OAI21_X1 U18637 ( .B1(n15044), .B2(n19667), .A(n15043), .ZN(n15045) );
  AOI211_X1 U18638 ( .C1(n15047), .C2(n19676), .A(n15046), .B(n15045), .ZN(
        n15052) );
  NAND2_X1 U18639 ( .A1(n15050), .A2(n19674), .ZN(n15051) );
  OAI211_X1 U18640 ( .C1(n15053), .C2(n16254), .A(n15052), .B(n15051), .ZN(
        P2_U2824) );
  AOI21_X1 U18641 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15054), .ZN(n15055) );
  OAI21_X1 U18642 ( .B1(n15056), .B2(n20714), .A(n15055), .ZN(n15057) );
  OAI22_X1 U18643 ( .A1(n15062), .A2(n13375), .B1(n15061), .B2(n15086), .ZN(
        n15064) );
  XNOR2_X1 U18644 ( .A(n15064), .B(n15063), .ZN(n15702) );
  INV_X1 U18645 ( .A(n15507), .ZN(n15069) );
  NOR2_X1 U18646 ( .A1(n15075), .A2(n21434), .ZN(n15066) );
  OAI21_X1 U18647 ( .B1(n15066), .B2(P1_REIP_REG_30__SCAN_IN), .A(n15065), 
        .ZN(n15068) );
  AOI22_X1 U18648 ( .A1(n20622), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20625), .ZN(n15067) );
  OAI211_X1 U18649 ( .C1(n20620), .C2(n15069), .A(n15068), .B(n15067), .ZN(
        n15070) );
  AOI21_X1 U18650 ( .B1(n15702), .B2(n20608), .A(n15070), .ZN(n15071) );
  OAI21_X1 U18651 ( .B1(n15370), .B2(n15350), .A(n15071), .ZN(P1_U2810) );
  INV_X1 U18652 ( .A(n15072), .ZN(n15412) );
  INV_X1 U18653 ( .A(n15073), .ZN(n15087) );
  AOI22_X1 U18654 ( .A1(n20622), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20625), .ZN(n15074) );
  OAI21_X1 U18655 ( .B1(n15075), .B2(P1_REIP_REG_29__SCAN_IN), .A(n15074), 
        .ZN(n15076) );
  AOI21_X1 U18656 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n15087), .A(n15076), 
        .ZN(n15077) );
  OAI21_X1 U18657 ( .B1(n15078), .B2(n20620), .A(n15077), .ZN(n15079) );
  AOI21_X1 U18658 ( .B1(n15371), .B2(n20608), .A(n15079), .ZN(n15080) );
  OAI21_X1 U18659 ( .B1(n15412), .B2(n15350), .A(n15080), .ZN(P1_U2811) );
  OR2_X1 U18660 ( .A1(n9716), .A2(n15084), .ZN(n15085) );
  AND2_X1 U18661 ( .A1(n15086), .A2(n15085), .ZN(n15710) );
  INV_X1 U18662 ( .A(n15521), .ZN(n15091) );
  AOI22_X1 U18663 ( .A1(n20622), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20625), .ZN(n15090) );
  OAI21_X1 U18664 ( .B1(n15088), .B2(P1_REIP_REG_28__SCAN_IN), .A(n15087), 
        .ZN(n15089) );
  OAI211_X1 U18665 ( .C1(n20620), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        n15092) );
  AOI21_X1 U18666 ( .B1(n15710), .B2(n20608), .A(n15092), .ZN(n15093) );
  OAI21_X1 U18667 ( .B1(n15524), .B2(n15350), .A(n15093), .ZN(P1_U2812) );
  NAND2_X1 U18668 ( .A1(n15154), .A2(n15094), .ZN(n15106) );
  AOI21_X1 U18669 ( .B1(n15096), .B2(n15106), .A(n15095), .ZN(n15536) );
  INV_X1 U18670 ( .A(n15536), .ZN(n15420) );
  INV_X1 U18671 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15101) );
  NAND3_X1 U18672 ( .A1(n15361), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15114), 
        .ZN(n15100) );
  NOR2_X1 U18673 ( .A1(n15097), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15098) );
  AOI22_X1 U18674 ( .A1(n20612), .A2(n15098), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20625), .ZN(n15099) );
  OAI211_X1 U18675 ( .C1(n15101), .C2(n15356), .A(n15100), .B(n15099), .ZN(
        n15102) );
  AOI21_X1 U18676 ( .B1(n20623), .B2(n15532), .A(n15102), .ZN(n15105) );
  AOI21_X1 U18677 ( .B1(n15103), .B2(n15111), .A(n9716), .ZN(n15720) );
  NAND2_X1 U18678 ( .A1(n15720), .A2(n20608), .ZN(n15104) );
  OAI211_X1 U18679 ( .C1(n15420), .C2(n15350), .A(n15105), .B(n15104), .ZN(
        P1_U2813) );
  INV_X1 U18680 ( .A(n15106), .ZN(n15107) );
  AOI21_X1 U18681 ( .B1(n15109), .B2(n15108), .A(n15107), .ZN(n15544) );
  INV_X1 U18682 ( .A(n15544), .ZN(n15424) );
  AOI21_X1 U18683 ( .B1(n15112), .B2(n15110), .A(n10225), .ZN(n15728) );
  AOI22_X1 U18684 ( .A1(n20622), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20625), .ZN(n15117) );
  AND2_X1 U18685 ( .A1(n20612), .A2(n15113), .ZN(n15115) );
  OAI211_X1 U18686 ( .C1(n15115), .C2(P1_REIP_REG_26__SCAN_IN), .A(n15361), 
        .B(n15114), .ZN(n15116) );
  OAI211_X1 U18687 ( .C1(n20620), .C2(n15542), .A(n15117), .B(n15116), .ZN(
        n15118) );
  AOI21_X1 U18688 ( .B1(n15728), .B2(n20608), .A(n15118), .ZN(n15119) );
  OAI21_X1 U18689 ( .B1(n15424), .B2(n15350), .A(n15119), .ZN(P1_U2814) );
  INV_X1 U18690 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U18691 ( .A1(n20622), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20625), .ZN(n15124) );
  OAI21_X1 U18692 ( .B1(n15121), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n15122) );
  OAI211_X1 U18693 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n20612), .B(n15122), .ZN(n15123) );
  OAI211_X1 U18694 ( .C1(n15137), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        n15126) );
  AOI21_X1 U18695 ( .B1(n20623), .B2(n15127), .A(n15126), .ZN(n15134) );
  INV_X1 U18696 ( .A(n15110), .ZN(n15132) );
  AOI21_X1 U18697 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(n15131) );
  NOR2_X1 U18698 ( .A1(n15132), .A2(n15131), .ZN(n15736) );
  NAND2_X1 U18699 ( .A1(n15736), .A2(n20608), .ZN(n15133) );
  OAI211_X1 U18700 ( .C1(n15120), .C2(n15350), .A(n15134), .B(n15133), .ZN(
        P1_U2815) );
  NAND2_X1 U18701 ( .A1(n15377), .A2(n20582), .ZN(n15142) );
  INV_X1 U18702 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15559) );
  NOR3_X1 U18703 ( .A1(n20595), .A2(n15559), .A3(n15135), .ZN(n15145) );
  AOI21_X1 U18704 ( .B1(n15145), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U18705 ( .A1(n20622), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20625), .ZN(n15136) );
  OAI21_X1 U18706 ( .B1(n15138), .B2(n15137), .A(n15136), .ZN(n15139) );
  AOI21_X1 U18707 ( .B1(n15140), .B2(n20623), .A(n15139), .ZN(n15141) );
  OAI211_X1 U18708 ( .C1(n15378), .C2(n20638), .A(n15142), .B(n15141), .ZN(
        P1_U2817) );
  OAI21_X1 U18709 ( .B1(n15154), .B2(n15144), .A(n15143), .ZN(n15554) );
  OAI21_X1 U18710 ( .B1(n20595), .B2(n15163), .A(n20561), .ZN(n15175) );
  AOI21_X1 U18711 ( .B1(n20612), .B2(n15559), .A(n15175), .ZN(n15148) );
  AOI22_X1 U18712 ( .A1(n20622), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20625), .ZN(n15147) );
  NAND2_X1 U18713 ( .A1(n15145), .A2(n21422), .ZN(n15146) );
  OAI211_X1 U18714 ( .C1(n15148), .C2(n21422), .A(n15147), .B(n15146), .ZN(
        n15152) );
  XNOR2_X1 U18715 ( .A(n15150), .B(n15149), .ZN(n15749) );
  NOR2_X1 U18716 ( .A1(n15749), .A2(n20638), .ZN(n15151) );
  AOI211_X1 U18717 ( .C1(n20623), .C2(n15551), .A(n15152), .B(n15151), .ZN(
        n15153) );
  OAI21_X1 U18718 ( .B1(n15554), .B2(n15350), .A(n15153), .ZN(P1_U2818) );
  INV_X1 U18719 ( .A(n15154), .ZN(n15158) );
  OR2_X1 U18720 ( .A1(n15156), .A2(n15155), .ZN(n15157) );
  INV_X1 U18721 ( .A(n15188), .ZN(n15160) );
  AOI21_X1 U18722 ( .B1(n15160), .B2(n15172), .A(n15159), .ZN(n15162) );
  OR2_X1 U18723 ( .A1(n15162), .A2(n15161), .ZN(n15381) );
  INV_X1 U18724 ( .A(n15381), .ZN(n15755) );
  INV_X1 U18725 ( .A(n15564), .ZN(n15168) );
  INV_X1 U18726 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15560) );
  NAND3_X1 U18727 ( .A1(n20612), .A2(n15163), .A3(n15559), .ZN(n15165) );
  NAND2_X1 U18728 ( .A1(n20622), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n15164) );
  OAI211_X1 U18729 ( .C1(n20588), .C2(n15560), .A(n15165), .B(n15164), .ZN(
        n15166) );
  AOI21_X1 U18730 ( .B1(n15175), .B2(P1_REIP_REG_21__SCAN_IN), .A(n15166), 
        .ZN(n15167) );
  OAI21_X1 U18731 ( .B1(n20620), .B2(n15168), .A(n15167), .ZN(n15169) );
  AOI21_X1 U18732 ( .B1(n15755), .B2(n20608), .A(n15169), .ZN(n15170) );
  OAI21_X1 U18733 ( .B1(n15561), .B2(n15350), .A(n15170), .ZN(P1_U2819) );
  XOR2_X1 U18734 ( .A(n15171), .B(n9737), .Z(n15572) );
  INV_X1 U18735 ( .A(n15572), .ZN(n15447) );
  XNOR2_X1 U18736 ( .A(n15188), .B(n15172), .ZN(n15764) );
  AOI22_X1 U18737 ( .A1(n20622), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20625), .ZN(n15178) );
  NAND2_X1 U18738 ( .A1(n20586), .A2(n15173), .ZN(n20560) );
  NOR2_X1 U18739 ( .A1(n20560), .A2(n15174), .ZN(n15176) );
  OAI21_X1 U18740 ( .B1(n15176), .B2(P1_REIP_REG_20__SCAN_IN), .A(n15175), 
        .ZN(n15177) );
  OAI211_X1 U18741 ( .C1(n20620), .C2(n15570), .A(n15178), .B(n15177), .ZN(
        n15179) );
  AOI21_X1 U18742 ( .B1(n15764), .B2(n20608), .A(n15179), .ZN(n15180) );
  OAI21_X1 U18743 ( .B1(n15447), .B2(n15350), .A(n15180), .ZN(P1_U2820) );
  NAND2_X1 U18744 ( .A1(n15181), .A2(n15182), .ZN(n15183) );
  NAND2_X1 U18745 ( .A1(n9737), .A2(n15183), .ZN(n15578) );
  INV_X1 U18746 ( .A(n15185), .ZN(n15203) );
  INV_X1 U18747 ( .A(n15186), .ZN(n15187) );
  OAI21_X1 U18748 ( .B1(n15184), .B2(n15203), .A(n15187), .ZN(n15189) );
  AND2_X1 U18749 ( .A1(n15189), .A2(n15188), .ZN(n15772) );
  INV_X1 U18750 ( .A(n15581), .ZN(n15199) );
  OAI21_X1 U18751 ( .B1(n20588), .B2(n15576), .A(n20576), .ZN(n15192) );
  INV_X1 U18752 ( .A(n15190), .ZN(n15195) );
  INV_X1 U18753 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21417) );
  NOR4_X1 U18754 ( .A1(n20560), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15195), 
        .A4(n21417), .ZN(n15191) );
  AOI211_X1 U18755 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n20622), .A(n15192), .B(
        n15191), .ZN(n15198) );
  NOR3_X1 U18756 ( .A1(n20560), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n15195), 
        .ZN(n15205) );
  INV_X1 U18757 ( .A(n15193), .ZN(n15194) );
  NAND2_X1 U18758 ( .A1(n20561), .A2(n15194), .ZN(n15232) );
  NAND2_X1 U18759 ( .A1(n15361), .A2(n15232), .ZN(n20553) );
  NAND2_X1 U18760 ( .A1(n15361), .A2(n15195), .ZN(n15196) );
  NAND2_X1 U18761 ( .A1(n20553), .A2(n15196), .ZN(n15211) );
  OAI21_X1 U18762 ( .B1(n15205), .B2(n15211), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15197) );
  OAI211_X1 U18763 ( .C1(n20620), .C2(n15199), .A(n15198), .B(n15197), .ZN(
        n15200) );
  AOI21_X1 U18764 ( .B1(n20608), .B2(n15772), .A(n15200), .ZN(n15201) );
  OAI21_X1 U18765 ( .B1(n15578), .B2(n15350), .A(n15201), .ZN(P1_U2821) );
  OAI21_X1 U18766 ( .B1(n15213), .B2(n15202), .A(n15181), .ZN(n15589) );
  XNOR2_X1 U18767 ( .A(n15184), .B(n15203), .ZN(n15792) );
  OAI21_X1 U18768 ( .B1(n20588), .B2(n15204), .A(n20576), .ZN(n15206) );
  AOI211_X1 U18769 ( .C1(n20622), .C2(P1_EBX_REG_18__SCAN_IN), .A(n15206), .B(
        n15205), .ZN(n15208) );
  AOI22_X1 U18770 ( .A1(n20623), .A2(n15585), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n15211), .ZN(n15207) );
  OAI211_X1 U18771 ( .C1(n15792), .C2(n20638), .A(n15208), .B(n15207), .ZN(
        n15209) );
  INV_X1 U18772 ( .A(n15209), .ZN(n15210) );
  OAI21_X1 U18773 ( .B1(n15589), .B2(n15350), .A(n15210), .ZN(P1_U2822) );
  INV_X1 U18774 ( .A(n15211), .ZN(n15225) );
  INV_X1 U18775 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21402) );
  AOI21_X1 U18776 ( .B1(n15274), .B2(n15212), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n15224) );
  AOI21_X1 U18777 ( .B1(n15214), .B2(n15228), .A(n15213), .ZN(n15604) );
  NAND2_X1 U18778 ( .A1(n15604), .A2(n20582), .ZN(n15223) );
  OR2_X1 U18779 ( .A1(n15237), .A2(n15215), .ZN(n15216) );
  NAND2_X1 U18780 ( .A1(n15184), .A2(n15216), .ZN(n15795) );
  INV_X1 U18781 ( .A(n15602), .ZN(n15219) );
  NAND2_X1 U18782 ( .A1(n20622), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n15217) );
  OAI211_X1 U18783 ( .C1(n20588), .C2(n21646), .A(n15217), .B(n20576), .ZN(
        n15218) );
  AOI21_X1 U18784 ( .B1(n20623), .B2(n15219), .A(n15218), .ZN(n15220) );
  OAI21_X1 U18785 ( .B1(n15795), .B2(n20638), .A(n15220), .ZN(n15221) );
  INV_X1 U18786 ( .A(n15221), .ZN(n15222) );
  OAI211_X1 U18787 ( .C1(n15225), .C2(n15224), .A(n15223), .B(n15222), .ZN(
        P1_U2823) );
  INV_X1 U18788 ( .A(n15226), .ZN(n15229) );
  OAI21_X1 U18789 ( .B1(n15229), .B2(n12479), .A(n15228), .ZN(n15612) );
  INV_X1 U18790 ( .A(n15612), .ZN(n15248) );
  NOR2_X1 U18791 ( .A1(n15242), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15230) );
  NAND2_X1 U18792 ( .A1(n15274), .A2(n15230), .ZN(n15259) );
  NOR2_X1 U18793 ( .A1(n15232), .A2(n15231), .ZN(n15291) );
  INV_X1 U18794 ( .A(n15291), .ZN(n15233) );
  NAND2_X1 U18795 ( .A1(n15361), .A2(n15233), .ZN(n15337) );
  NAND2_X1 U18796 ( .A1(n15361), .A2(n15242), .ZN(n15234) );
  AND2_X1 U18797 ( .A1(n15337), .A2(n15234), .ZN(n15253) );
  INV_X1 U18798 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21413) );
  AOI21_X1 U18799 ( .B1(n15259), .B2(n15253), .A(n21413), .ZN(n15247) );
  NOR2_X1 U18800 ( .A1(n15255), .A2(n15235), .ZN(n15236) );
  OR2_X1 U18801 ( .A1(n15237), .A2(n15236), .ZN(n15811) );
  INV_X1 U18802 ( .A(n15608), .ZN(n15241) );
  NAND2_X1 U18803 ( .A1(n20622), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15238) );
  OAI211_X1 U18804 ( .C1(n20588), .C2(n15239), .A(n15238), .B(n20576), .ZN(
        n15240) );
  AOI21_X1 U18805 ( .B1(n20623), .B2(n15241), .A(n15240), .ZN(n15245) );
  INV_X1 U18806 ( .A(n15242), .ZN(n15243) );
  NAND4_X1 U18807 ( .A1(n15274), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n15243), 
        .A4(n21413), .ZN(n15244) );
  OAI211_X1 U18808 ( .C1(n15811), .C2(n20638), .A(n15245), .B(n15244), .ZN(
        n15246) );
  AOI211_X1 U18809 ( .C1(n15248), .C2(n20582), .A(n15247), .B(n15246), .ZN(
        n15249) );
  INV_X1 U18810 ( .A(n15249), .ZN(P1_U2824) );
  NAND2_X1 U18811 ( .A1(n15250), .A2(n15251), .ZN(n15252) );
  AND2_X1 U18812 ( .A1(n15226), .A2(n15252), .ZN(n15623) );
  INV_X1 U18813 ( .A(n15621), .ZN(n15254) );
  INV_X1 U18814 ( .A(n15253), .ZN(n15275) );
  AOI22_X1 U18815 ( .A1(n20623), .A2(n15254), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15275), .ZN(n15263) );
  AOI21_X1 U18816 ( .B1(n15256), .B2(n15267), .A(n15255), .ZN(n15817) );
  NAND2_X1 U18817 ( .A1(n20622), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15257) );
  OAI211_X1 U18818 ( .C1(n20588), .C2(n15258), .A(n15257), .B(n20576), .ZN(
        n15261) );
  INV_X1 U18819 ( .A(n15259), .ZN(n15260) );
  AOI211_X1 U18820 ( .C1(n15817), .C2(n20608), .A(n15261), .B(n15260), .ZN(
        n15262) );
  OAI211_X1 U18821 ( .C1(n15467), .C2(n15350), .A(n15263), .B(n15262), .ZN(
        P1_U2825) );
  OR2_X1 U18822 ( .A1(n15264), .A2(n15265), .ZN(n15266) );
  INV_X1 U18823 ( .A(n15267), .ZN(n15268) );
  AOI21_X1 U18824 ( .B1(n15269), .B2(n15289), .A(n15268), .ZN(n15824) );
  NAND2_X1 U18825 ( .A1(n20622), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n15270) );
  OAI211_X1 U18826 ( .C1(n20588), .C2(n15271), .A(n15270), .B(n20576), .ZN(
        n15273) );
  NOR2_X1 U18827 ( .A1(n20620), .A2(n15629), .ZN(n15272) );
  AOI211_X1 U18828 ( .C1(n15824), .C2(n20608), .A(n15273), .B(n15272), .ZN(
        n15278) );
  NAND2_X1 U18829 ( .A1(n15274), .A2(n15290), .ZN(n15296) );
  INV_X1 U18830 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21408) );
  NOR2_X1 U18831 ( .A1(n15296), .A2(n21408), .ZN(n15276) );
  OAI21_X1 U18832 ( .B1(n15276), .B2(P1_REIP_REG_14__SCAN_IN), .A(n15275), 
        .ZN(n15277) );
  OAI211_X1 U18833 ( .C1(n15470), .C2(n15350), .A(n15278), .B(n15277), .ZN(
        P1_U2826) );
  INV_X1 U18834 ( .A(n15329), .ZN(n15283) );
  INV_X1 U18835 ( .A(n15281), .ZN(n15316) );
  AOI21_X1 U18836 ( .B1(n15283), .B2(n15282), .A(n9742), .ZN(n15303) );
  INV_X1 U18837 ( .A(n15284), .ZN(n15302) );
  NOR2_X1 U18838 ( .A1(n15303), .A2(n15302), .ZN(n15301) );
  INV_X1 U18839 ( .A(n15264), .ZN(n15285) );
  OAI21_X1 U18840 ( .B1(n15301), .B2(n15286), .A(n15285), .ZN(n15648) );
  INV_X1 U18841 ( .A(n15633), .ZN(n15299) );
  NAND2_X1 U18842 ( .A1(n15306), .A2(n15287), .ZN(n15288) );
  NAND2_X1 U18843 ( .A1(n15289), .A2(n15288), .ZN(n15836) );
  NAND2_X1 U18844 ( .A1(n15291), .A2(n15290), .ZN(n15312) );
  NAND3_X1 U18845 ( .A1(n15361), .A2(P1_REIP_REG_13__SCAN_IN), .A3(n15312), 
        .ZN(n15295) );
  NAND2_X1 U18846 ( .A1(n20625), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15292) );
  NAND2_X1 U18847 ( .A1(n15292), .A2(n20576), .ZN(n15293) );
  AOI21_X1 U18848 ( .B1(n20622), .B2(P1_EBX_REG_13__SCAN_IN), .A(n15293), .ZN(
        n15294) );
  OAI211_X1 U18849 ( .C1(n15836), .C2(n20638), .A(n15295), .B(n15294), .ZN(
        n15298) );
  NOR2_X1 U18850 ( .A1(n15296), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15297) );
  AOI211_X1 U18851 ( .C1(n20623), .C2(n15299), .A(n15298), .B(n15297), .ZN(
        n15300) );
  OAI21_X1 U18852 ( .B1(n15648), .B2(n15350), .A(n15300), .ZN(P1_U2827) );
  AOI21_X1 U18853 ( .B1(n15303), .B2(n15302), .A(n15301), .ZN(n15655) );
  INV_X1 U18854 ( .A(n15655), .ZN(n15474) );
  INV_X1 U18855 ( .A(n15653), .ZN(n15311) );
  OR2_X1 U18856 ( .A1(n10397), .A2(n15304), .ZN(n15305) );
  NAND2_X1 U18857 ( .A1(n15306), .A2(n15305), .ZN(n15846) );
  OAI21_X1 U18858 ( .B1(n20588), .B2(n15307), .A(n20576), .ZN(n15308) );
  AOI21_X1 U18859 ( .B1(n20622), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15308), .ZN(
        n15309) );
  OAI21_X1 U18860 ( .B1(n20638), .B2(n15846), .A(n15309), .ZN(n15310) );
  AOI21_X1 U18861 ( .B1(n20623), .B2(n15311), .A(n15310), .ZN(n15315) );
  INV_X1 U18862 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21406) );
  NOR2_X1 U18863 ( .A1(n15328), .A2(n21406), .ZN(n15313) );
  OAI211_X1 U18864 ( .C1(n15313), .C2(P1_REIP_REG_12__SCAN_IN), .A(n15361), 
        .B(n15312), .ZN(n15314) );
  OAI211_X1 U18865 ( .C1(n15474), .C2(n15350), .A(n15315), .B(n15314), .ZN(
        P1_U2828) );
  AOI21_X1 U18866 ( .B1(n15317), .B2(n15316), .A(n9742), .ZN(n15664) );
  NAND2_X1 U18867 ( .A1(n15664), .A2(n20582), .ZN(n15327) );
  INV_X1 U18868 ( .A(n15662), .ZN(n15325) );
  NAND2_X1 U18869 ( .A1(n20625), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15318) );
  NAND2_X1 U18870 ( .A1(n15318), .A2(n20576), .ZN(n15319) );
  AOI21_X1 U18871 ( .B1(n20622), .B2(P1_EBX_REG_11__SCAN_IN), .A(n15319), .ZN(
        n15323) );
  AND2_X1 U18872 ( .A1(n9794), .A2(n15320), .ZN(n15321) );
  OR2_X1 U18873 ( .A1(n10397), .A2(n15321), .ZN(n15392) );
  INV_X1 U18874 ( .A(n15392), .ZN(n15860) );
  NAND2_X1 U18875 ( .A1(n15860), .A2(n20608), .ZN(n15322) );
  OAI211_X1 U18876 ( .C1(n15337), .C2(n21406), .A(n15323), .B(n15322), .ZN(
        n15324) );
  AOI21_X1 U18877 ( .B1(n20623), .B2(n15325), .A(n15324), .ZN(n15326) );
  OAI211_X1 U18878 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15328), .A(n15327), 
        .B(n15326), .ZN(P1_U2829) );
  OAI21_X1 U18879 ( .B1(n15482), .B2(n15330), .A(n15329), .ZN(n15677) );
  NOR2_X1 U18880 ( .A1(n21402), .A2(n20560), .ZN(n15336) );
  NAND2_X1 U18881 ( .A1(n15331), .A2(n15332), .ZN(n15333) );
  NAND2_X1 U18882 ( .A1(n9794), .A2(n15333), .ZN(n15872) );
  AOI22_X1 U18883 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20625), .B1(
        P1_EBX_REG_10__SCAN_IN), .B2(n20622), .ZN(n15334) );
  OAI211_X1 U18884 ( .C1(n15872), .C2(n20638), .A(n15334), .B(n20576), .ZN(
        n15335) );
  AOI21_X1 U18885 ( .B1(n15336), .B2(n21403), .A(n15335), .ZN(n15341) );
  INV_X1 U18886 ( .A(n15673), .ZN(n15339) );
  NOR2_X1 U18887 ( .A1(n15337), .A2(n21403), .ZN(n15338) );
  AOI21_X1 U18888 ( .B1(n20623), .B2(n15339), .A(n15338), .ZN(n15340) );
  OAI211_X1 U18889 ( .C1(n15677), .C2(n15350), .A(n15341), .B(n15340), .ZN(
        P1_U2830) );
  INV_X1 U18890 ( .A(n15480), .ZN(n15342) );
  OAI21_X1 U18891 ( .B1(n15280), .B2(n15343), .A(n15342), .ZN(n15695) );
  NOR2_X1 U18892 ( .A1(n21399), .A2(n20553), .ZN(n15348) );
  XOR2_X1 U18893 ( .A(n15879), .B(n9792), .Z(n17325) );
  AOI22_X1 U18894 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(n20622), .B1(n20608), .B2(
        n17325), .ZN(n15344) );
  OAI211_X1 U18895 ( .C1(n20588), .C2(n12360), .A(n15344), .B(n20576), .ZN(
        n15347) );
  INV_X1 U18896 ( .A(n20562), .ZN(n20563) );
  NAND4_X1 U18897 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20563), .A3(n20586), 
        .A4(n21399), .ZN(n15345) );
  OAI21_X1 U18898 ( .B1(n15691), .B2(n20620), .A(n15345), .ZN(n15346) );
  NOR3_X1 U18899 ( .A1(n15348), .A2(n15347), .A3(n15346), .ZN(n15349) );
  OAI21_X1 U18900 ( .B1(n15695), .B2(n15350), .A(n15349), .ZN(P1_U2832) );
  OAI21_X1 U18901 ( .B1(n15351), .B2(n15353), .A(n15350), .ZN(n20633) );
  INV_X1 U18902 ( .A(n20633), .ZN(n15368) );
  NOR2_X1 U18903 ( .A1(n15353), .A2(n15352), .ZN(n20626) );
  AOI22_X1 U18904 ( .A1(n20626), .A2(n21256), .B1(n20610), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n15354) );
  OAI21_X1 U18905 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15357) );
  NOR2_X1 U18906 ( .A1(n20595), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20611) );
  AOI211_X1 U18907 ( .C1(n20608), .C2(n20758), .A(n15357), .B(n20611), .ZN(
        n15359) );
  MUX2_X1 U18908 ( .A(n20620), .B(n20588), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15358) );
  OAI211_X1 U18909 ( .C1(n15368), .C2(n15360), .A(n15359), .B(n15358), .ZN(
        P1_U2839) );
  NAND2_X1 U18910 ( .A1(n20620), .A2(n20588), .ZN(n15365) );
  AOI22_X1 U18911 ( .A1(n20622), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n20893), .B2(
        n20626), .ZN(n15363) );
  NAND2_X1 U18912 ( .A1(n15361), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15362) );
  OAI211_X1 U18913 ( .C1(n20638), .C2(n15891), .A(n15363), .B(n15362), .ZN(
        n15364) );
  AOI21_X1 U18914 ( .B1(n15365), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n15364), .ZN(n15366) );
  OAI21_X1 U18915 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(P1_U2840) );
  AOI22_X1 U18916 ( .A1(n15702), .A2(n20648), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15404), .ZN(n15369) );
  OAI21_X1 U18917 ( .B1(n15370), .B2(n15399), .A(n15369), .ZN(P1_U2842) );
  AOI22_X1 U18918 ( .A1(n15371), .A2(n20648), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n15404), .ZN(n15372) );
  OAI21_X1 U18919 ( .B1(n15412), .B2(n15399), .A(n15372), .ZN(P1_U2843) );
  AOI22_X1 U18920 ( .A1(n15710), .A2(n20648), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15404), .ZN(n15373) );
  OAI21_X1 U18921 ( .B1(n15524), .B2(n15399), .A(n15373), .ZN(P1_U2844) );
  AOI22_X1 U18922 ( .A1(n15720), .A2(n20648), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n15404), .ZN(n15374) );
  OAI21_X1 U18923 ( .B1(n15420), .B2(n15399), .A(n15374), .ZN(P1_U2845) );
  AOI22_X1 U18924 ( .A1(n15728), .A2(n20648), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n15404), .ZN(n15375) );
  OAI21_X1 U18925 ( .B1(n15424), .B2(n15399), .A(n15375), .ZN(P1_U2846) );
  AOI22_X1 U18926 ( .A1(n15736), .A2(n20648), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n15404), .ZN(n15376) );
  OAI21_X1 U18927 ( .B1(n15120), .B2(n15399), .A(n15376), .ZN(P1_U2847) );
  INV_X1 U18928 ( .A(n15377), .ZN(n15434) );
  INV_X1 U18929 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15379) );
  OAI222_X1 U18930 ( .A1(n15434), .A2(n15399), .B1(n15379), .B2(n20653), .C1(
        n15378), .C2(n15395), .ZN(P1_U2849) );
  INV_X1 U18931 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15380) );
  OAI222_X1 U18932 ( .A1(n15554), .A2(n15399), .B1(n15380), .B2(n20653), .C1(
        n15395), .C2(n15749), .ZN(P1_U2850) );
  INV_X1 U18933 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15382) );
  OAI222_X1 U18934 ( .A1(n15561), .A2(n15399), .B1(n15382), .B2(n20653), .C1(
        n15381), .C2(n15395), .ZN(P1_U2851) );
  AOI22_X1 U18935 ( .A1(n15764), .A2(n20648), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n15404), .ZN(n15383) );
  OAI21_X1 U18936 ( .B1(n15447), .B2(n15399), .A(n15383), .ZN(P1_U2852) );
  INV_X1 U18937 ( .A(n15772), .ZN(n15384) );
  OAI222_X1 U18938 ( .A1(n15578), .A2(n15399), .B1(n21676), .B2(n20653), .C1(
        n15384), .C2(n15395), .ZN(P1_U2853) );
  OAI222_X1 U18939 ( .A1(n15589), .A2(n15399), .B1(n15385), .B2(n20653), .C1(
        n15395), .C2(n15792), .ZN(P1_U2854) );
  INV_X1 U18940 ( .A(n15604), .ZN(n15458) );
  INV_X1 U18941 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15386) );
  OAI222_X1 U18942 ( .A1(n15399), .A2(n15458), .B1(n15386), .B2(n20653), .C1(
        n15795), .C2(n15395), .ZN(P1_U2855) );
  OAI222_X1 U18943 ( .A1(n15612), .A2(n15399), .B1(n15387), .B2(n20653), .C1(
        n15811), .C2(n15395), .ZN(P1_U2856) );
  AOI22_X1 U18944 ( .A1(n15817), .A2(n20648), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15404), .ZN(n15388) );
  OAI21_X1 U18945 ( .B1(n15467), .B2(n15399), .A(n15388), .ZN(P1_U2857) );
  AOI22_X1 U18946 ( .A1(n15824), .A2(n20648), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15404), .ZN(n15389) );
  OAI21_X1 U18947 ( .B1(n15470), .B2(n15399), .A(n15389), .ZN(P1_U2858) );
  INV_X1 U18948 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15390) );
  OAI222_X1 U18949 ( .A1(n15648), .A2(n15399), .B1(n15390), .B2(n20653), .C1(
        n15836), .C2(n15395), .ZN(P1_U2859) );
  INV_X1 U18950 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15391) );
  OAI222_X1 U18951 ( .A1(n15474), .A2(n15399), .B1(n15391), .B2(n20653), .C1(
        n15846), .C2(n15395), .ZN(P1_U2860) );
  INV_X1 U18952 ( .A(n15664), .ZN(n15477) );
  INV_X1 U18953 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15393) );
  OAI222_X1 U18954 ( .A1(n15477), .A2(n15399), .B1(n15393), .B2(n20653), .C1(
        n15392), .C2(n15395), .ZN(P1_U2861) );
  OAI22_X1 U18955 ( .A1(n15872), .A2(n15395), .B1(n15394), .B2(n20653), .ZN(
        n15396) );
  INV_X1 U18956 ( .A(n15396), .ZN(n15397) );
  OAI21_X1 U18957 ( .B1(n15677), .B2(n15399), .A(n15397), .ZN(P1_U2862) );
  AOI22_X1 U18958 ( .A1(n17325), .A2(n20648), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n15404), .ZN(n15398) );
  OAI21_X1 U18959 ( .B1(n15695), .B2(n15399), .A(n15398), .ZN(P1_U2864) );
  XOR2_X1 U18960 ( .A(n15496), .B(n15400), .Z(n20583) );
  INV_X1 U18961 ( .A(n20583), .ZN(n15489) );
  AND2_X1 U18962 ( .A1(n17356), .A2(n15401), .ZN(n15402) );
  NOR2_X1 U18963 ( .A1(n17340), .A2(n15402), .ZN(n20578) );
  AOI22_X1 U18964 ( .A1(n20578), .A2(n20648), .B1(n15404), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n15403) );
  OAI21_X1 U18965 ( .B1(n15489), .B2(n15399), .A(n15403), .ZN(P1_U2866) );
  XOR2_X1 U18966 ( .A(n15490), .B(n15491), .Z(n20708) );
  INV_X1 U18967 ( .A(n20708), .ZN(n15500) );
  XOR2_X1 U18968 ( .A(n17354), .B(n17355), .Z(n20719) );
  AOI22_X1 U18969 ( .A1(n20648), .A2(n20719), .B1(n15404), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n15405) );
  OAI21_X1 U18970 ( .B1(n15500), .B2(n15399), .A(n15405), .ZN(P1_U2868) );
  NAND2_X1 U18971 ( .A1(n20769), .A2(DATAI_13_), .ZN(n15407) );
  NAND2_X1 U18972 ( .A1(n20771), .A2(BUF1_REG_13__SCAN_IN), .ZN(n15406) );
  AND2_X1 U18973 ( .A1(n15407), .A2(n15406), .ZN(n20688) );
  OAI22_X1 U18974 ( .A1(n15460), .A2(n20688), .B1(n15497), .B2(n15408), .ZN(
        n15409) );
  AOI21_X1 U18975 ( .B1(n15462), .B2(BUF1_REG_29__SCAN_IN), .A(n15409), .ZN(
        n15411) );
  NAND2_X1 U18976 ( .A1(n15463), .A2(DATAI_29_), .ZN(n15410) );
  OAI211_X1 U18977 ( .C1(n15412), .C2(n15501), .A(n15411), .B(n15410), .ZN(
        P1_U2875) );
  OAI22_X1 U18978 ( .A1(n15460), .A2(n15473), .B1(n15497), .B2(n15413), .ZN(
        n15414) );
  AOI21_X1 U18979 ( .B1(n15462), .B2(BUF1_REG_28__SCAN_IN), .A(n15414), .ZN(
        n15416) );
  NAND2_X1 U18980 ( .A1(n15463), .A2(DATAI_28_), .ZN(n15415) );
  OAI211_X1 U18981 ( .C1(n15524), .C2(n15501), .A(n15416), .B(n15415), .ZN(
        P1_U2876) );
  OAI22_X1 U18982 ( .A1(n15460), .A2(n15476), .B1(n15497), .B2(n14241), .ZN(
        n15417) );
  AOI21_X1 U18983 ( .B1(n15462), .B2(BUF1_REG_27__SCAN_IN), .A(n15417), .ZN(
        n15419) );
  NAND2_X1 U18984 ( .A1(n15463), .A2(DATAI_27_), .ZN(n15418) );
  OAI211_X1 U18985 ( .C1(n15420), .C2(n15501), .A(n15419), .B(n15418), .ZN(
        P1_U2877) );
  OAI22_X1 U18986 ( .A1(n15460), .A2(n15478), .B1(n15497), .B2(n14041), .ZN(
        n15421) );
  AOI21_X1 U18987 ( .B1(n15462), .B2(BUF1_REG_26__SCAN_IN), .A(n15421), .ZN(
        n15423) );
  NAND2_X1 U18988 ( .A1(n15463), .A2(DATAI_26_), .ZN(n15422) );
  OAI211_X1 U18989 ( .C1(n15424), .C2(n15501), .A(n15423), .B(n15422), .ZN(
        P1_U2878) );
  NAND2_X1 U18990 ( .A1(n20769), .A2(DATAI_9_), .ZN(n15426) );
  NAND2_X1 U18991 ( .A1(n20771), .A2(BUF1_REG_9__SCAN_IN), .ZN(n15425) );
  AND2_X1 U18992 ( .A1(n15426), .A2(n15425), .ZN(n20685) );
  OAI22_X1 U18993 ( .A1(n15460), .A2(n20685), .B1(n15497), .B2(n15427), .ZN(
        n15428) );
  AOI21_X1 U18994 ( .B1(n15462), .B2(BUF1_REG_25__SCAN_IN), .A(n15428), .ZN(
        n15430) );
  NAND2_X1 U18995 ( .A1(n15463), .A2(DATAI_25_), .ZN(n15429) );
  OAI211_X1 U18996 ( .C1(n15120), .C2(n15501), .A(n15430), .B(n15429), .ZN(
        P1_U2879) );
  OAI22_X1 U18997 ( .A1(n15460), .A2(n20821), .B1(n15497), .B2(n14054), .ZN(
        n15431) );
  AOI21_X1 U18998 ( .B1(n15462), .B2(BUF1_REG_23__SCAN_IN), .A(n15431), .ZN(
        n15433) );
  NAND2_X1 U18999 ( .A1(n15463), .A2(DATAI_23_), .ZN(n15432) );
  OAI211_X1 U19000 ( .C1(n15434), .C2(n15501), .A(n15433), .B(n15432), .ZN(
        P1_U2881) );
  OAI22_X1 U19001 ( .A1(n15460), .A2(n20813), .B1(n15497), .B2(n15435), .ZN(
        n15436) );
  AOI21_X1 U19002 ( .B1(n15462), .B2(BUF1_REG_22__SCAN_IN), .A(n15436), .ZN(
        n15438) );
  NAND2_X1 U19003 ( .A1(n15463), .A2(DATAI_22_), .ZN(n15437) );
  OAI211_X1 U19004 ( .C1(n15554), .C2(n15501), .A(n15438), .B(n15437), .ZN(
        P1_U2882) );
  OAI22_X1 U19005 ( .A1(n15460), .A2(n20809), .B1(n15497), .B2(n15439), .ZN(
        n15440) );
  AOI21_X1 U19006 ( .B1(n15462), .B2(BUF1_REG_21__SCAN_IN), .A(n15440), .ZN(
        n15442) );
  NAND2_X1 U19007 ( .A1(n15463), .A2(DATAI_21_), .ZN(n15441) );
  OAI211_X1 U19008 ( .C1(n15561), .C2(n15501), .A(n15442), .B(n15441), .ZN(
        P1_U2883) );
  OAI22_X1 U19009 ( .A1(n15460), .A2(n20805), .B1(n15497), .B2(n15443), .ZN(
        n15444) );
  AOI21_X1 U19010 ( .B1(n15462), .B2(BUF1_REG_20__SCAN_IN), .A(n15444), .ZN(
        n15446) );
  NAND2_X1 U19011 ( .A1(n15463), .A2(DATAI_20_), .ZN(n15445) );
  OAI211_X1 U19012 ( .C1(n15447), .C2(n15501), .A(n15446), .B(n15445), .ZN(
        P1_U2884) );
  OAI22_X1 U19013 ( .A1(n15460), .A2(n20801), .B1(n15497), .B2(n14049), .ZN(
        n15448) );
  AOI21_X1 U19014 ( .B1(n15462), .B2(BUF1_REG_19__SCAN_IN), .A(n15448), .ZN(
        n15450) );
  NAND2_X1 U19015 ( .A1(n15463), .A2(DATAI_19_), .ZN(n15449) );
  OAI211_X1 U19016 ( .C1(n15578), .C2(n15501), .A(n15450), .B(n15449), .ZN(
        P1_U2885) );
  OAI22_X1 U19017 ( .A1(n15460), .A2(n20797), .B1(n15497), .B2(n15451), .ZN(
        n15452) );
  AOI21_X1 U19018 ( .B1(n15462), .B2(BUF1_REG_18__SCAN_IN), .A(n15452), .ZN(
        n15454) );
  NAND2_X1 U19019 ( .A1(n15463), .A2(DATAI_18_), .ZN(n15453) );
  OAI211_X1 U19020 ( .C1(n15589), .C2(n15501), .A(n15454), .B(n15453), .ZN(
        P1_U2886) );
  OAI22_X1 U19021 ( .A1(n15460), .A2(n20793), .B1(n15497), .B2(n14046), .ZN(
        n15455) );
  AOI21_X1 U19022 ( .B1(n15462), .B2(BUF1_REG_17__SCAN_IN), .A(n15455), .ZN(
        n15457) );
  NAND2_X1 U19023 ( .A1(n15463), .A2(DATAI_17_), .ZN(n15456) );
  OAI211_X1 U19024 ( .C1(n15458), .C2(n15501), .A(n15457), .B(n15456), .ZN(
        P1_U2887) );
  OAI22_X1 U19025 ( .A1(n15460), .A2(n20783), .B1(n15497), .B2(n15459), .ZN(
        n15461) );
  AOI21_X1 U19026 ( .B1(n15462), .B2(BUF1_REG_16__SCAN_IN), .A(n15461), .ZN(
        n15465) );
  NAND2_X1 U19027 ( .A1(n15463), .A2(DATAI_16_), .ZN(n15464) );
  OAI211_X1 U19028 ( .C1(n15612), .C2(n15501), .A(n15465), .B(n15464), .ZN(
        P1_U2888) );
  OAI222_X1 U19029 ( .A1(n15501), .A2(n15467), .B1(n15499), .B2(n15466), .C1(
        n20661), .C2(n15497), .ZN(P1_U2889) );
  INV_X1 U19030 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15468) );
  OAI222_X1 U19031 ( .A1(n15470), .A2(n15501), .B1(n15469), .B2(n15499), .C1(
        n15468), .C2(n15497), .ZN(P1_U2890) );
  INV_X1 U19032 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15471) );
  OAI222_X1 U19033 ( .A1(n15648), .A2(n15501), .B1(n20688), .B2(n15499), .C1(
        n15471), .C2(n15497), .ZN(P1_U2891) );
  INV_X1 U19034 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15472) );
  OAI222_X1 U19035 ( .A1(n15474), .A2(n15501), .B1(n15473), .B2(n15499), .C1(
        n15472), .C2(n15497), .ZN(P1_U2892) );
  INV_X1 U19036 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15475) );
  OAI222_X1 U19037 ( .A1(n15477), .A2(n15501), .B1(n15476), .B2(n15499), .C1(
        n15475), .C2(n15497), .ZN(P1_U2893) );
  OAI222_X1 U19038 ( .A1(n15677), .A2(n15501), .B1(n15497), .B2(n14248), .C1(
        n15478), .C2(n15499), .ZN(P1_U2894) );
  NOR2_X1 U19039 ( .A1(n15480), .A2(n15479), .ZN(n15481) );
  INV_X1 U19040 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15483) );
  OAI222_X1 U19041 ( .A1(n15684), .A2(n15501), .B1(n20685), .B2(n15499), .C1(
        n15483), .C2(n15497), .ZN(P1_U2895) );
  OAI222_X1 U19042 ( .A1(n15695), .A2(n15501), .B1(n15484), .B2(n15499), .C1(
        n20670), .C2(n15497), .ZN(P1_U2896) );
  AOI21_X1 U19043 ( .B1(n15486), .B2(n15485), .A(n15280), .ZN(n20644) );
  INV_X1 U19044 ( .A(n20644), .ZN(n15487) );
  OAI222_X1 U19045 ( .A1(n15501), .A2(n15487), .B1(n20821), .B2(n15499), .C1(
        n15497), .C2(n14260), .ZN(P1_U2897) );
  OAI222_X1 U19046 ( .A1(n15501), .A2(n15489), .B1(n15488), .B2(n15497), .C1(
        n20813), .C2(n15499), .ZN(P1_U2898) );
  NAND2_X1 U19047 ( .A1(n15491), .A2(n15490), .ZN(n15494) );
  INV_X1 U19048 ( .A(n15492), .ZN(n15493) );
  NAND2_X1 U19049 ( .A1(n15494), .A2(n15493), .ZN(n15495) );
  AND2_X1 U19050 ( .A1(n15496), .A2(n15495), .ZN(n20650) );
  INV_X1 U19051 ( .A(n20650), .ZN(n15498) );
  OAI222_X1 U19052 ( .A1(n15501), .A2(n15498), .B1(n15499), .B2(n20809), .C1(
        n15497), .C2(n14256), .ZN(P1_U2899) );
  OAI222_X1 U19053 ( .A1(n15501), .A2(n15500), .B1(n15497), .B2(n14252), .C1(
        n20805), .C2(n15499), .ZN(P1_U2900) );
  NOR2_X1 U19054 ( .A1(n15503), .A2(n15502), .ZN(n15504) );
  NAND2_X1 U19055 ( .A1(n15507), .A2(n15586), .ZN(n15508) );
  NAND2_X1 U19056 ( .A1(n20718), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15696) );
  OAI211_X1 U19057 ( .C1(n15577), .C2(n15509), .A(n15508), .B(n15696), .ZN(
        n15510) );
  AOI21_X1 U19058 ( .B1(n15511), .B2(n20709), .A(n15510), .ZN(n15512) );
  OAI21_X1 U19059 ( .B1(n15704), .B2(n20537), .A(n15512), .ZN(P1_U2969) );
  NAND2_X1 U19060 ( .A1(n15657), .A2(n15513), .ZN(n15539) );
  NAND2_X1 U19061 ( .A1(n15514), .A2(n15539), .ZN(n15518) );
  OAI21_X1 U19062 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15515), .A(
        n15518), .ZN(n15517) );
  INV_X1 U19063 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15717) );
  MUX2_X1 U19064 ( .A(n15717), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15657), .Z(n15516) );
  OAI211_X1 U19065 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15518), .A(
        n15517), .B(n15516), .ZN(n15520) );
  XNOR2_X1 U19066 ( .A(n15520), .B(n15519), .ZN(n15713) );
  INV_X1 U19067 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21433) );
  NOR2_X1 U19068 ( .A1(n20576), .A2(n21433), .ZN(n15709) );
  AOI21_X1 U19069 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15709), .ZN(n15523) );
  NAND2_X1 U19070 ( .A1(n15521), .A2(n15586), .ZN(n15522) );
  OAI211_X1 U19071 ( .C1(n15524), .C2(n20770), .A(n15523), .B(n15522), .ZN(
        n15525) );
  INV_X1 U19072 ( .A(n15525), .ZN(n15526) );
  OAI21_X1 U19073 ( .B1(n20537), .B2(n15713), .A(n15526), .ZN(P1_U2971) );
  NAND2_X1 U19074 ( .A1(n15528), .A2(n12192), .ZN(n15529) );
  NAND2_X1 U19075 ( .A1(n15530), .A2(n15529), .ZN(n15531) );
  NAND2_X1 U19076 ( .A1(n15532), .A2(n15586), .ZN(n15533) );
  NAND2_X1 U19077 ( .A1(n20718), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15716) );
  OAI211_X1 U19078 ( .C1(n15577), .C2(n15534), .A(n15533), .B(n15716), .ZN(
        n15535) );
  AOI21_X1 U19079 ( .B1(n15536), .B2(n20709), .A(n15535), .ZN(n15537) );
  OAI21_X1 U19080 ( .B1(n15722), .B2(n20537), .A(n15537), .ZN(P1_U2972) );
  OAI211_X1 U19081 ( .C1(n12192), .C2(n15514), .A(n15538), .B(n15539), .ZN(
        n15540) );
  XNOR2_X1 U19082 ( .A(n15540), .B(n21717), .ZN(n15730) );
  INV_X1 U19083 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21429) );
  NOR2_X1 U19084 ( .A1(n20576), .A2(n21429), .ZN(n15724) );
  AOI21_X1 U19085 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15724), .ZN(n15541) );
  OAI21_X1 U19086 ( .B1(n15542), .B2(n20714), .A(n15541), .ZN(n15543) );
  AOI21_X1 U19087 ( .B1(n15544), .B2(n20709), .A(n15543), .ZN(n15545) );
  OAI21_X1 U19088 ( .B1(n20537), .B2(n15730), .A(n15545), .ZN(P1_U2973) );
  NAND2_X1 U19089 ( .A1(n15546), .A2(n15547), .ZN(n15548) );
  XNOR2_X1 U19090 ( .A(n15548), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15739) );
  NAND2_X1 U19091 ( .A1(n15739), .A2(n20710), .ZN(n15553) );
  NOR2_X1 U19092 ( .A1(n20576), .A2(n21422), .ZN(n15745) );
  NOR2_X1 U19093 ( .A1(n15577), .A2(n15549), .ZN(n15550) );
  AOI211_X1 U19094 ( .C1(n15586), .C2(n15551), .A(n15745), .B(n15550), .ZN(
        n15552) );
  OAI211_X1 U19095 ( .C1(n20770), .C2(n15554), .A(n15553), .B(n15552), .ZN(
        P1_U2977) );
  INV_X1 U19096 ( .A(n15758), .ZN(n15741) );
  NOR2_X1 U19097 ( .A1(n15555), .A2(n15741), .ZN(n15557) );
  MUX2_X1 U19098 ( .A(n15557), .B(n15556), .S(n12192), .Z(n15558) );
  XNOR2_X1 U19099 ( .A(n15558), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15757) );
  OR2_X1 U19100 ( .A1(n20576), .A2(n15559), .ZN(n15750) );
  OAI21_X1 U19101 ( .B1(n15577), .B2(n15560), .A(n15750), .ZN(n15563) );
  NOR2_X1 U19102 ( .A1(n15561), .A2(n20770), .ZN(n15562) );
  AOI211_X1 U19103 ( .C1(n15586), .C2(n15564), .A(n15563), .B(n15562), .ZN(
        n15565) );
  OAI21_X1 U19104 ( .B1(n20537), .B2(n15757), .A(n15565), .ZN(P1_U2978) );
  INV_X1 U19105 ( .A(n15555), .ZN(n15775) );
  NAND2_X1 U19106 ( .A1(n15775), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15567) );
  MUX2_X1 U19107 ( .A(n15566), .B(n15567), .S(n15657), .Z(n15568) );
  XOR2_X1 U19108 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n15568), .Z(
        n15766) );
  NOR2_X1 U19109 ( .A1(n20576), .A2(n21419), .ZN(n15763) );
  AOI21_X1 U19110 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15763), .ZN(n15569) );
  OAI21_X1 U19111 ( .B1(n20714), .B2(n15570), .A(n15569), .ZN(n15571) );
  AOI21_X1 U19112 ( .B1(n15572), .B2(n20709), .A(n15571), .ZN(n15573) );
  OAI21_X1 U19113 ( .B1(n15766), .B2(n20537), .A(n15573), .ZN(P1_U2979) );
  NOR2_X1 U19114 ( .A1(n15641), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15574) );
  MUX2_X1 U19115 ( .A(n15657), .B(n15574), .S(n15555), .Z(n15575) );
  XNOR2_X1 U19116 ( .A(n15575), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15774) );
  NAND2_X1 U19117 ( .A1(n20718), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15768) );
  OAI21_X1 U19118 ( .B1(n15577), .B2(n15576), .A(n15768), .ZN(n15580) );
  NOR2_X1 U19119 ( .A1(n15578), .A2(n20770), .ZN(n15579) );
  AOI211_X1 U19120 ( .C1(n15586), .C2(n15581), .A(n15580), .B(n15579), .ZN(
        n15582) );
  OAI21_X1 U19121 ( .B1(n20537), .B2(n15774), .A(n15582), .ZN(P1_U2980) );
  NOR2_X1 U19122 ( .A1(n15583), .A2(n15584), .ZN(n15776) );
  NOR3_X1 U19123 ( .A1(n15776), .A2(n15775), .A3(n20537), .ZN(n15591) );
  NOR2_X1 U19124 ( .A1(n20576), .A2(n21417), .ZN(n15789) );
  AOI21_X1 U19125 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15789), .ZN(n15588) );
  NAND2_X1 U19126 ( .A1(n15586), .A2(n15585), .ZN(n15587) );
  OAI211_X1 U19127 ( .C1(n15589), .C2(n20770), .A(n15588), .B(n15587), .ZN(
        n15590) );
  OR2_X1 U19128 ( .A1(n15591), .A2(n15590), .ZN(P1_U2981) );
  NAND2_X1 U19129 ( .A1(n15657), .A2(n15592), .ZN(n15678) );
  INV_X1 U19130 ( .A(n15593), .ZN(n15595) );
  NAND2_X1 U19131 ( .A1(n15641), .A2(n15806), .ZN(n15616) );
  OAI21_X1 U19132 ( .B1(n15615), .B2(n15597), .A(n15616), .ZN(n15606) );
  XNOR2_X1 U19133 ( .A(n15641), .B(n15805), .ZN(n15607) );
  NOR2_X1 U19134 ( .A1(n15606), .A2(n15607), .ZN(n15599) );
  NOR2_X1 U19135 ( .A1(n15599), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15598) );
  MUX2_X1 U19136 ( .A(n15599), .B(n15598), .S(n12192), .Z(n15600) );
  XNOR2_X1 U19137 ( .A(n15600), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15801) );
  INV_X1 U19138 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21415) );
  NOR2_X1 U19139 ( .A1(n20576), .A2(n21415), .ZN(n15797) );
  AOI21_X1 U19140 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15797), .ZN(n15601) );
  OAI21_X1 U19141 ( .B1(n20714), .B2(n15602), .A(n15601), .ZN(n15603) );
  AOI21_X1 U19142 ( .B1(n15604), .B2(n20709), .A(n15603), .ZN(n15605) );
  OAI21_X1 U19143 ( .B1(n15801), .B2(n20537), .A(n15605), .ZN(P1_U2982) );
  XOR2_X1 U19144 ( .A(n15607), .B(n15606), .Z(n15802) );
  NAND2_X1 U19145 ( .A1(n15802), .A2(n20710), .ZN(n15611) );
  NOR2_X1 U19146 ( .A1(n20576), .A2(n21413), .ZN(n15808) );
  NOR2_X1 U19147 ( .A1(n20714), .A2(n15608), .ZN(n15609) );
  AOI211_X1 U19148 ( .C1(n20703), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15808), .B(n15609), .ZN(n15610) );
  OAI211_X1 U19149 ( .C1(n20770), .C2(n15612), .A(n15611), .B(n15610), .ZN(
        P1_U2983) );
  INV_X1 U19150 ( .A(n15613), .ZN(n15614) );
  NOR2_X1 U19151 ( .A1(n15615), .A2(n15614), .ZN(n15619) );
  NAND2_X1 U19152 ( .A1(n15617), .A2(n15616), .ZN(n15618) );
  XNOR2_X1 U19153 ( .A(n15619), .B(n15618), .ZN(n15819) );
  INV_X1 U19154 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21766) );
  NOR2_X1 U19155 ( .A1(n20576), .A2(n21766), .ZN(n15812) );
  AOI21_X1 U19156 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15812), .ZN(n15620) );
  OAI21_X1 U19157 ( .B1(n20714), .B2(n15621), .A(n15620), .ZN(n15622) );
  AOI21_X1 U19158 ( .B1(n15623), .B2(n20709), .A(n15622), .ZN(n15624) );
  OAI21_X1 U19159 ( .B1(n15819), .B2(n20537), .A(n15624), .ZN(P1_U2984) );
  AOI21_X1 U19160 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n12192), .A(
        n15625), .ZN(n15627) );
  XNOR2_X1 U19161 ( .A(n15641), .B(n15820), .ZN(n15626) );
  XNOR2_X1 U19162 ( .A(n15627), .B(n15626), .ZN(n15827) );
  INV_X1 U19163 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21409) );
  NOR2_X1 U19164 ( .A1(n20576), .A2(n21409), .ZN(n15822) );
  AOI21_X1 U19165 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15822), .ZN(n15628) );
  OAI21_X1 U19166 ( .B1(n20714), .B2(n15629), .A(n15628), .ZN(n15630) );
  AOI21_X1 U19167 ( .B1(n15631), .B2(n20709), .A(n15630), .ZN(n15632) );
  OAI21_X1 U19168 ( .B1(n15827), .B2(n20537), .A(n15632), .ZN(P1_U2985) );
  NOR2_X1 U19169 ( .A1(n20576), .A2(n21408), .ZN(n15831) );
  NOR2_X1 U19170 ( .A1(n20714), .A2(n15633), .ZN(n15634) );
  AOI211_X1 U19171 ( .C1(n20703), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15831), .B(n15634), .ZN(n15647) );
  OR2_X1 U19172 ( .A1(n15667), .A2(n15635), .ZN(n15639) );
  INV_X1 U19173 ( .A(n15636), .ZN(n15637) );
  OR2_X1 U19174 ( .A1(n15657), .A2(n15637), .ZN(n15638) );
  NAND2_X1 U19175 ( .A1(n15639), .A2(n15638), .ZN(n15651) );
  NOR2_X1 U19176 ( .A1(n15641), .A2(n15852), .ZN(n15642) );
  OR2_X1 U19177 ( .A1(n15643), .A2(n15642), .ZN(n15650) );
  NOR2_X1 U19178 ( .A1(n15651), .A2(n15650), .ZN(n15649) );
  NOR2_X1 U19179 ( .A1(n15649), .A2(n15643), .ZN(n15645) );
  XNOR2_X1 U19180 ( .A(n15645), .B(n15644), .ZN(n15828) );
  NAND2_X1 U19181 ( .A1(n15828), .A2(n20710), .ZN(n15646) );
  OAI211_X1 U19182 ( .C1(n15648), .C2(n20770), .A(n15647), .B(n15646), .ZN(
        P1_U2986) );
  AOI21_X1 U19183 ( .B1(n15651), .B2(n15650), .A(n15649), .ZN(n15856) );
  INV_X1 U19184 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21407) );
  NOR2_X1 U19185 ( .A1(n20576), .A2(n21407), .ZN(n15848) );
  AOI21_X1 U19186 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15848), .ZN(n15652) );
  OAI21_X1 U19187 ( .B1(n20714), .B2(n15653), .A(n15652), .ZN(n15654) );
  AOI21_X1 U19188 ( .B1(n15655), .B2(n20709), .A(n15654), .ZN(n15656) );
  OAI21_X1 U19189 ( .B1(n15856), .B2(n20537), .A(n15656), .ZN(P1_U2987) );
  NAND2_X1 U19190 ( .A1(n15657), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15659) );
  INV_X1 U19191 ( .A(n15668), .ZN(n15658) );
  NAND3_X1 U19192 ( .A1(n15658), .A2(n12192), .A3(n15666), .ZN(n15671) );
  OAI21_X1 U19193 ( .B1(n15667), .B2(n15659), .A(n15671), .ZN(n15660) );
  XNOR2_X1 U19194 ( .A(n15660), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15865) );
  NOR2_X1 U19195 ( .A1(n20576), .A2(n21406), .ZN(n15859) );
  AOI21_X1 U19196 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15859), .ZN(n15661) );
  OAI21_X1 U19197 ( .B1(n20714), .B2(n15662), .A(n15661), .ZN(n15663) );
  AOI21_X1 U19198 ( .B1(n15664), .B2(n20709), .A(n15663), .ZN(n15665) );
  OAI21_X1 U19199 ( .B1(n15865), .B2(n20537), .A(n15665), .ZN(P1_U2988) );
  XNOR2_X1 U19200 ( .A(n15667), .B(n15666), .ZN(n15670) );
  NAND2_X1 U19201 ( .A1(n15668), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15669) );
  MUX2_X1 U19202 ( .A(n15670), .B(n15669), .S(n12192), .Z(n15672) );
  NAND2_X1 U19203 ( .A1(n15672), .A2(n15671), .ZN(n15866) );
  NAND2_X1 U19204 ( .A1(n15866), .A2(n20710), .ZN(n15676) );
  NOR2_X1 U19205 ( .A1(n20576), .A2(n21403), .ZN(n15874) );
  NOR2_X1 U19206 ( .A1(n20714), .A2(n15673), .ZN(n15674) );
  AOI211_X1 U19207 ( .C1(n20703), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15874), .B(n15674), .ZN(n15675) );
  OAI211_X1 U19208 ( .C1(n20770), .C2(n15677), .A(n15676), .B(n15675), .ZN(
        P1_U2989) );
  NAND2_X1 U19209 ( .A1(n15679), .A2(n15678), .ZN(n15683) );
  NAND2_X1 U19210 ( .A1(n15680), .A2(n15681), .ZN(n15682) );
  XOR2_X1 U19211 ( .A(n15683), .B(n15682), .Z(n15889) );
  NAND2_X1 U19212 ( .A1(n20718), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15882) );
  NAND2_X1 U19213 ( .A1(n20703), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15685) );
  OAI211_X1 U19214 ( .C1(n20714), .C2(n20557), .A(n15882), .B(n15685), .ZN(
        n15686) );
  AOI21_X1 U19215 ( .B1(n20640), .B2(n20709), .A(n15686), .ZN(n15687) );
  OAI21_X1 U19216 ( .B1(n15889), .B2(n20537), .A(n15687), .ZN(P1_U2990) );
  XNOR2_X1 U19217 ( .A(n15689), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15690) );
  XNOR2_X1 U19218 ( .A(n15688), .B(n15690), .ZN(n17335) );
  NAND2_X1 U19219 ( .A1(n17335), .A2(n20710), .ZN(n15694) );
  AND2_X1 U19220 ( .A1(n20718), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n17324) );
  NOR2_X1 U19221 ( .A1(n20714), .A2(n15691), .ZN(n15692) );
  AOI211_X1 U19222 ( .C1(n20703), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17324), .B(n15692), .ZN(n15693) );
  OAI211_X1 U19223 ( .C1(n20770), .C2(n15695), .A(n15694), .B(n15693), .ZN(
        P1_U2991) );
  INV_X1 U19224 ( .A(n15696), .ZN(n15701) );
  AOI21_X1 U19225 ( .B1(n15699), .B2(n15698), .A(n15697), .ZN(n15700) );
  AOI211_X1 U19226 ( .C1(n15702), .C2(n20742), .A(n15701), .B(n15700), .ZN(
        n15703) );
  OAI21_X1 U19227 ( .B1(n15704), .B2(n20753), .A(n15703), .ZN(P1_U3001) );
  INV_X1 U19228 ( .A(n15714), .ZN(n15707) );
  NOR3_X1 U19229 ( .A1(n15707), .A2(n15706), .A3(n15705), .ZN(n15708) );
  AOI211_X1 U19230 ( .C1(n10186), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15709), .B(n15708), .ZN(n15712) );
  NAND2_X1 U19231 ( .A1(n15710), .A2(n20742), .ZN(n15711) );
  OAI211_X1 U19232 ( .C1(n15713), .C2(n20753), .A(n15712), .B(n15711), .ZN(
        P1_U3003) );
  NAND2_X1 U19233 ( .A1(n15714), .A2(n15717), .ZN(n15715) );
  OAI211_X1 U19234 ( .C1(n15718), .C2(n15717), .A(n15716), .B(n15715), .ZN(
        n15719) );
  AOI21_X1 U19235 ( .B1(n15720), .B2(n20742), .A(n15719), .ZN(n15721) );
  OAI21_X1 U19236 ( .B1(n15722), .B2(n20753), .A(n15721), .ZN(P1_U3004) );
  INV_X1 U19237 ( .A(n15723), .ZN(n15734) );
  XNOR2_X1 U19238 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15726) );
  AOI21_X1 U19239 ( .B1(n15731), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15724), .ZN(n15725) );
  OAI21_X1 U19240 ( .B1(n15734), .B2(n15726), .A(n15725), .ZN(n15727) );
  AOI21_X1 U19241 ( .B1(n15728), .B2(n20742), .A(n15727), .ZN(n15729) );
  OAI21_X1 U19242 ( .B1(n15730), .B2(n20753), .A(n15729), .ZN(P1_U3005) );
  NAND2_X1 U19243 ( .A1(n15731), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15733) );
  OAI211_X1 U19244 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15734), .A(
        n15733), .B(n15732), .ZN(n15735) );
  AOI21_X1 U19245 ( .B1(n15736), .B2(n20742), .A(n15735), .ZN(n15737) );
  OAI21_X1 U19246 ( .B1(n15738), .B2(n20753), .A(n15737), .ZN(P1_U3006) );
  NAND2_X1 U19247 ( .A1(n15739), .A2(n20738), .ZN(n15748) );
  NAND2_X1 U19248 ( .A1(n15758), .A2(n15752), .ZN(n15740) );
  OR2_X1 U19249 ( .A1(n15770), .A2(n15740), .ZN(n15751) );
  AND2_X1 U19250 ( .A1(n20757), .A2(n15741), .ZN(n15742) );
  NOR2_X1 U19251 ( .A1(n15767), .A2(n15742), .ZN(n15753) );
  NAND2_X1 U19252 ( .A1(n15751), .A2(n15753), .ZN(n15746) );
  NOR3_X1 U19253 ( .A1(n15770), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15743), .ZN(n15744) );
  AOI211_X1 U19254 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15746), .A(
        n15745), .B(n15744), .ZN(n15747) );
  OAI211_X1 U19255 ( .C1(n15749), .C2(n20760), .A(n15748), .B(n15747), .ZN(
        P1_U3009) );
  OAI211_X1 U19256 ( .C1(n15753), .C2(n15752), .A(n15751), .B(n15750), .ZN(
        n15754) );
  AOI21_X1 U19257 ( .B1(n15755), .B2(n20742), .A(n15754), .ZN(n15756) );
  OAI21_X1 U19258 ( .B1(n15757), .B2(n20753), .A(n15756), .ZN(P1_U3010) );
  INV_X1 U19259 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15761) );
  AOI21_X1 U19260 ( .B1(n15785), .B2(n15779), .A(n15758), .ZN(n15759) );
  OAI22_X1 U19261 ( .A1(n15759), .A2(n15767), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15760) );
  AOI21_X1 U19262 ( .B1(n15761), .B2(n15770), .A(n15760), .ZN(n15762) );
  AOI211_X1 U19263 ( .C1(n15764), .C2(n20742), .A(n15763), .B(n15762), .ZN(
        n15765) );
  OAI21_X1 U19264 ( .B1(n15766), .B2(n20753), .A(n15765), .ZN(P1_U3011) );
  NAND2_X1 U19265 ( .A1(n15767), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15769) );
  OAI211_X1 U19266 ( .C1(n15770), .C2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15769), .B(n15768), .ZN(n15771) );
  AOI21_X1 U19267 ( .B1(n15772), .B2(n20742), .A(n15771), .ZN(n15773) );
  OAI21_X1 U19268 ( .B1(n15774), .B2(n20753), .A(n15773), .ZN(P1_U3012) );
  OR3_X1 U19269 ( .A1(n15776), .A2(n15775), .A3(n20753), .ZN(n15791) );
  NOR2_X1 U19270 ( .A1(n15777), .A2(n15833), .ZN(n15778) );
  OR2_X1 U19271 ( .A1(n15779), .A2(n15778), .ZN(n15783) );
  OR2_X1 U19272 ( .A1(n15781), .A2(n15780), .ZN(n15782) );
  AND4_X1 U19273 ( .A1(n15784), .A2(n15895), .A3(n15783), .A4(n15782), .ZN(
        n15829) );
  OAI21_X1 U19274 ( .B1(n15785), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15829), .ZN(n15823) );
  AOI21_X1 U19275 ( .B1(n15820), .B2(n20757), .A(n15823), .ZN(n15803) );
  OAI21_X1 U19276 ( .B1(n15786), .B2(n17334), .A(n15803), .ZN(n15799) );
  INV_X1 U19277 ( .A(n15786), .ZN(n15787) );
  NOR3_X1 U19278 ( .A1(n15815), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15787), .ZN(n15788) );
  AOI211_X1 U19279 ( .C1(n15799), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15789), .B(n15788), .ZN(n15790) );
  OAI211_X1 U19280 ( .C1(n15792), .C2(n20760), .A(n15791), .B(n15790), .ZN(
        P1_U3013) );
  INV_X1 U19281 ( .A(n15804), .ZN(n15794) );
  OAI21_X1 U19282 ( .B1(n15815), .B2(n15794), .A(n15793), .ZN(n15798) );
  NOR2_X1 U19283 ( .A1(n15795), .A2(n20760), .ZN(n15796) );
  AOI211_X1 U19284 ( .C1(n15799), .C2(n15798), .A(n15797), .B(n15796), .ZN(
        n15800) );
  OAI21_X1 U19285 ( .B1(n15801), .B2(n20753), .A(n15800), .ZN(P1_U3014) );
  NAND2_X1 U19286 ( .A1(n15802), .A2(n20738), .ZN(n15810) );
  INV_X1 U19287 ( .A(n15803), .ZN(n15813) );
  AOI211_X1 U19288 ( .C1(n15806), .C2(n15805), .A(n15804), .B(n15815), .ZN(
        n15807) );
  AOI211_X1 U19289 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15813), .A(
        n15808), .B(n15807), .ZN(n15809) );
  OAI211_X1 U19290 ( .C1(n20760), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        P1_U3015) );
  AOI21_X1 U19291 ( .B1(n15813), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15812), .ZN(n15814) );
  OAI21_X1 U19292 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15815), .A(
        n15814), .ZN(n15816) );
  AOI21_X1 U19293 ( .B1(n20742), .B2(n15817), .A(n15816), .ZN(n15818) );
  OAI21_X1 U19294 ( .B1(n15819), .B2(n20753), .A(n15818), .ZN(P1_U3016) );
  AND3_X1 U19295 ( .A1(n15832), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15820), .ZN(n15821) );
  AOI211_X1 U19296 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15823), .A(
        n15822), .B(n15821), .ZN(n15826) );
  NAND2_X1 U19297 ( .A1(n15824), .A2(n20742), .ZN(n15825) );
  OAI211_X1 U19298 ( .C1(n15827), .C2(n20753), .A(n15826), .B(n15825), .ZN(
        P1_U3017) );
  NAND2_X1 U19299 ( .A1(n15828), .A2(n20738), .ZN(n15835) );
  NOR2_X1 U19300 ( .A1(n15829), .A2(n15833), .ZN(n15830) );
  AOI211_X1 U19301 ( .C1(n15833), .C2(n15832), .A(n15831), .B(n15830), .ZN(
        n15834) );
  OAI211_X1 U19302 ( .C1(n20760), .C2(n15836), .A(n15835), .B(n15834), .ZN(
        P1_U3018) );
  INV_X1 U19303 ( .A(n20735), .ZN(n15841) );
  NOR2_X1 U19304 ( .A1(n15841), .A2(n15837), .ZN(n15869) );
  INV_X1 U19305 ( .A(n15838), .ZN(n15862) );
  INV_X1 U19306 ( .A(n15839), .ZN(n15853) );
  OAI22_X1 U19307 ( .A1(n15841), .A2(n15862), .B1(n15840), .B2(n15853), .ZN(
        n15845) );
  INV_X1 U19308 ( .A(n15842), .ZN(n15843) );
  NAND2_X1 U19309 ( .A1(n20736), .A2(n15843), .ZN(n15844) );
  NAND2_X1 U19310 ( .A1(n20750), .A2(n15844), .ZN(n17331) );
  NOR3_X1 U19311 ( .A1(n15869), .A2(n15845), .A3(n17331), .ZN(n15857) );
  OAI21_X1 U19312 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n20743), .A(
        n15857), .ZN(n15849) );
  NOR2_X1 U19313 ( .A1(n15846), .A2(n20760), .ZN(n15847) );
  AOI211_X1 U19314 ( .C1(n15849), .C2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15848), .B(n15847), .ZN(n15855) );
  INV_X1 U19315 ( .A(n20720), .ZN(n15850) );
  NAND3_X1 U19316 ( .A1(n17348), .A2(n15853), .A3(n15852), .ZN(n15854) );
  OAI211_X1 U19317 ( .C1(n15856), .C2(n20753), .A(n15855), .B(n15854), .ZN(
        P1_U3019) );
  NOR2_X1 U19318 ( .A1(n15857), .A2(n15861), .ZN(n15858) );
  AOI211_X1 U19319 ( .C1(n20742), .C2(n15860), .A(n15859), .B(n15858), .ZN(
        n15864) );
  NAND3_X1 U19320 ( .A1(n17348), .A2(n15862), .A3(n15861), .ZN(n15863) );
  OAI211_X1 U19321 ( .C1(n15865), .C2(n20753), .A(n15864), .B(n15863), .ZN(
        P1_U3020) );
  XNOR2_X1 U19322 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15877) );
  NAND2_X1 U19323 ( .A1(n17348), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17347) );
  OR2_X1 U19324 ( .A1(n17347), .A2(n17323), .ZN(n15884) );
  NAND2_X1 U19325 ( .A1(n15866), .A2(n20738), .ZN(n15876) );
  INV_X1 U19326 ( .A(n15867), .ZN(n15868) );
  OAI21_X1 U19327 ( .B1(n15869), .B2(n15868), .A(n20757), .ZN(n15871) );
  INV_X1 U19328 ( .A(n17331), .ZN(n15870) );
  NAND2_X1 U19329 ( .A1(n15871), .A2(n15870), .ZN(n15887) );
  NOR2_X1 U19330 ( .A1(n15872), .A2(n20760), .ZN(n15873) );
  AOI211_X1 U19331 ( .C1(n15887), .C2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15874), .B(n15873), .ZN(n15875) );
  OAI211_X1 U19332 ( .C1(n15877), .C2(n15884), .A(n15876), .B(n15875), .ZN(
        P1_U3021) );
  INV_X1 U19333 ( .A(n15331), .ZN(n15881) );
  AOI21_X1 U19334 ( .B1(n9792), .B2(n15879), .A(n15878), .ZN(n15880) );
  NOR2_X1 U19335 ( .A1(n15881), .A2(n15880), .ZN(n20639) );
  INV_X1 U19336 ( .A(n20639), .ZN(n15883) );
  OAI21_X1 U19337 ( .B1(n15883), .B2(n20760), .A(n15882), .ZN(n15886) );
  NOR2_X1 U19338 ( .A1(n15884), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15885) );
  AOI211_X1 U19339 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15887), .A(
        n15886), .B(n15885), .ZN(n15888) );
  OAI21_X1 U19340 ( .B1(n15889), .B2(n20753), .A(n15888), .ZN(P1_U3022) );
  NAND2_X1 U19341 ( .A1(n15890), .A2(n20738), .ZN(n15899) );
  INV_X1 U19342 ( .A(n15891), .ZN(n15893) );
  AOI21_X1 U19343 ( .B1(n20742), .B2(n15893), .A(n15892), .ZN(n15898) );
  OAI21_X1 U19344 ( .B1(n15894), .B2(n20736), .A(n20734), .ZN(n20766) );
  INV_X1 U19345 ( .A(n15895), .ZN(n20752) );
  OAI21_X1 U19346 ( .B1(n20752), .B2(n15896), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15897) );
  NAND4_X1 U19347 ( .A1(n15899), .A2(n15898), .A3(n20766), .A4(n15897), .ZN(
        P1_U3031) );
  INV_X1 U19348 ( .A(n15900), .ZN(n15901) );
  NAND2_X1 U19349 ( .A1(n15901), .A2(n17366), .ZN(n17297) );
  AOI22_X1 U19350 ( .A1(n20774), .A2(n9694), .B1(n20893), .B2(n15902), .ZN(
        n15903) );
  NAND2_X1 U19351 ( .A1(n17297), .A2(n15903), .ZN(n15904) );
  MUX2_X1 U19352 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15904), .S(
        n21475), .Z(P1_U3478) );
  AND2_X1 U19353 ( .A1(n9694), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20969) );
  NAND2_X1 U19354 ( .A1(n20971), .A2(n20969), .ZN(n21312) );
  MUX2_X1 U19355 ( .A(n21312), .B(n20898), .S(n21065), .Z(n15906) );
  OAI21_X1 U19356 ( .B1(n21465), .B2(n13843), .A(n15906), .ZN(n15907) );
  MUX2_X1 U19357 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15907), .S(
        n21475), .Z(P1_U3476) );
  NAND2_X1 U19358 ( .A1(n15908), .A2(n19674), .ZN(n15916) );
  INV_X1 U19359 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15914) );
  AOI21_X1 U19360 ( .B1(n15920), .B2(n16482), .A(n15909), .ZN(n15910) );
  NOR2_X1 U19361 ( .A1(n15910), .A2(n17049), .ZN(n15912) );
  AOI22_X1 U19362 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        n16249), .B2(P2_REIP_REG_30__SCAN_IN), .ZN(n15913) );
  OAI21_X1 U19363 ( .B1(n15919), .B2(n15918), .A(n11444), .ZN(n16697) );
  AOI22_X1 U19364 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n16249), .B2(P2_REIP_REG_29__SCAN_IN), .ZN(n15922) );
  NAND2_X1 U19365 ( .A1(n16272), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15921) );
  NAND2_X1 U19366 ( .A1(n11539), .A2(n15924), .ZN(n15925) );
  NAND2_X1 U19367 ( .A1(n16699), .A2(n19674), .ZN(n15927) );
  XNOR2_X1 U19368 ( .A(n15928), .B(n16492), .ZN(n15929) );
  NAND2_X1 U19369 ( .A1(n15929), .A2(n19681), .ZN(n15931) );
  AOI22_X1 U19370 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n16249), .B2(P2_REIP_REG_28__SCAN_IN), .ZN(n15930) );
  OAI211_X1 U19371 ( .C1(n19667), .C2(n15932), .A(n15931), .B(n15930), .ZN(
        n15935) );
  NOR2_X1 U19372 ( .A1(n15933), .A2(n16254), .ZN(n15934) );
  AOI211_X1 U19373 ( .C1(n19676), .C2(n15936), .A(n15935), .B(n15934), .ZN(
        n15937) );
  OAI21_X1 U19374 ( .B1(n16373), .B2(n16267), .A(n15937), .ZN(P2_U2827) );
  NOR2_X1 U19375 ( .A1(n13555), .A2(n15938), .ZN(n15939) );
  OR2_X1 U19376 ( .A1(n11540), .A2(n15939), .ZN(n16704) );
  AND2_X1 U19377 ( .A1(n15941), .A2(n15940), .ZN(n15942) );
  OR2_X1 U19378 ( .A1(n15942), .A2(n11545), .ZN(n16711) );
  INV_X1 U19379 ( .A(n16711), .ZN(n15953) );
  NOR2_X1 U19380 ( .A1(n15943), .A2(n16270), .ZN(n15952) );
  AOI21_X1 U19381 ( .B1(n15946), .B2(n19681), .A(n19669), .ZN(n15950) );
  OAI22_X1 U19382 ( .A1(n16202), .A2(n15944), .B1(n20455), .B2(n19664), .ZN(
        n15948) );
  INV_X1 U19383 ( .A(n16502), .ZN(n15945) );
  NOR3_X1 U19384 ( .A1(n15946), .A2(n15945), .A3(n16219), .ZN(n15947) );
  AOI211_X1 U19385 ( .C1(n16272), .C2(P2_EBX_REG_27__SCAN_IN), .A(n15948), .B(
        n15947), .ZN(n15949) );
  OAI21_X1 U19386 ( .B1(n15950), .B2(n16502), .A(n15949), .ZN(n15951) );
  AOI211_X1 U19387 ( .C1(n15953), .C2(n19678), .A(n15952), .B(n15951), .ZN(
        n15954) );
  OAI21_X1 U19388 ( .B1(n16704), .B2(n16267), .A(n15954), .ZN(P2_U2828) );
  XNOR2_X1 U19389 ( .A(n15955), .B(n10421), .ZN(n15959) );
  OAI22_X1 U19390 ( .A1(n16202), .A2(n15956), .B1(n20452), .B2(n19664), .ZN(
        n15957) );
  AOI21_X1 U19391 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16272), .A(n15957), .ZN(
        n15958) );
  OAI21_X1 U19392 ( .B1(n17049), .B2(n15959), .A(n15958), .ZN(n15960) );
  AOI21_X1 U19393 ( .B1(n15961), .B2(n19676), .A(n15960), .ZN(n15963) );
  NAND2_X1 U19394 ( .A1(n16390), .A2(n19674), .ZN(n15962) );
  OAI211_X1 U19395 ( .C1(n16304), .C2(n16254), .A(n15963), .B(n15962), .ZN(
        P2_U2829) );
  OAI21_X1 U19396 ( .B1(n13025), .B2(n15964), .A(n13560), .ZN(n16722) );
  INV_X1 U19397 ( .A(n13556), .ZN(n15965) );
  AOI21_X1 U19398 ( .B1(n15966), .B2(n13032), .A(n15965), .ZN(n16724) );
  NAND2_X1 U19399 ( .A1(n16724), .A2(n19674), .ZN(n15977) );
  XNOR2_X1 U19400 ( .A(n15967), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n15975) );
  NOR2_X1 U19401 ( .A1(n17002), .A2(n15968), .ZN(n15969) );
  XOR2_X1 U19402 ( .A(n16511), .B(n15969), .Z(n15973) );
  OAI22_X1 U19403 ( .A1(n16202), .A2(n15970), .B1(n20451), .B2(n19664), .ZN(
        n15971) );
  AOI21_X1 U19404 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16272), .A(n15971), .ZN(
        n15972) );
  OAI21_X1 U19405 ( .B1(n17049), .B2(n15973), .A(n15972), .ZN(n15974) );
  AOI21_X1 U19406 ( .B1(n15975), .B2(n19676), .A(n15974), .ZN(n15976) );
  OAI211_X1 U19407 ( .C1(n16722), .C2(n16254), .A(n15977), .B(n15976), .ZN(
        P2_U2830) );
  INV_X1 U19408 ( .A(n16521), .ZN(n15978) );
  NAND2_X1 U19409 ( .A1(n15978), .A2(n19678), .ZN(n15989) );
  OAI22_X1 U19410 ( .A1(n16202), .A2(n10278), .B1(n15979), .B2(n19667), .ZN(
        n15987) );
  INV_X1 U19411 ( .A(n16519), .ZN(n15980) );
  NAND3_X1 U19412 ( .A1(n16273), .A2(n15980), .A3(n15981), .ZN(n15984) );
  NOR2_X1 U19413 ( .A1(n15981), .A2(n17049), .ZN(n15982) );
  OAI21_X1 U19414 ( .B1(n19669), .B2(n15982), .A(n16519), .ZN(n15983) );
  OAI211_X1 U19415 ( .C1(n19664), .C2(n15985), .A(n15984), .B(n15983), .ZN(
        n15986) );
  OAI211_X1 U19416 ( .C1(n16267), .C2(n16403), .A(n15989), .B(n15988), .ZN(
        P2_U2831) );
  AOI21_X1 U19417 ( .B1(n15991), .B2(n15990), .A(n13026), .ZN(n16535) );
  INV_X1 U19418 ( .A(n16535), .ZN(n16736) );
  NAND2_X1 U19419 ( .A1(n16146), .A2(n15992), .ZN(n15993) );
  XOR2_X1 U19420 ( .A(n16528), .B(n15993), .Z(n15996) );
  OAI22_X1 U19421 ( .A1(n16202), .A2(n16530), .B1(n20448), .B2(n19664), .ZN(
        n15994) );
  AOI21_X1 U19422 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16272), .A(n15994), .ZN(
        n15995) );
  OAI21_X1 U19423 ( .B1(n17049), .B2(n15996), .A(n15995), .ZN(n15997) );
  AOI21_X1 U19424 ( .B1(n15998), .B2(n19676), .A(n15997), .ZN(n16003) );
  AOI21_X1 U19425 ( .B1(n16001), .B2(n15999), .A(n16000), .ZN(n16741) );
  NAND2_X1 U19426 ( .A1(n16741), .A2(n19674), .ZN(n16002) );
  OAI211_X1 U19427 ( .C1(n16736), .C2(n16254), .A(n16003), .B(n16002), .ZN(
        P2_U2832) );
  AOI21_X1 U19428 ( .B1(n16004), .B2(n11566), .A(n10301), .ZN(n16752) );
  INV_X1 U19429 ( .A(n16752), .ZN(n16422) );
  INV_X1 U19430 ( .A(n15990), .ZN(n16005) );
  AOI21_X1 U19431 ( .B1(n16006), .B2(n9754), .A(n16005), .ZN(n16556) );
  AOI22_X1 U19432 ( .A1(n16272), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19671), .ZN(n16013) );
  OAI21_X1 U19433 ( .B1(n17049), .B2(n16007), .A(n16216), .ZN(n16010) );
  INV_X1 U19434 ( .A(n16011), .ZN(n16554) );
  NAND3_X1 U19435 ( .A1(n16273), .A2(n16554), .A3(n16007), .ZN(n16008) );
  OAI21_X1 U19436 ( .B1(n19664), .B2(n20446), .A(n16008), .ZN(n16009) );
  AOI21_X1 U19437 ( .B1(n16011), .B2(n16010), .A(n16009), .ZN(n16012) );
  OAI211_X1 U19438 ( .C1(n16014), .C2(n16270), .A(n16013), .B(n16012), .ZN(
        n16015) );
  AOI21_X1 U19439 ( .B1(n16556), .B2(n19678), .A(n16015), .ZN(n16016) );
  OAI21_X1 U19440 ( .B1(n16422), .B2(n16267), .A(n16016), .ZN(P2_U2833) );
  NOR2_X1 U19441 ( .A1(n16017), .A2(n16270), .ZN(n16024) );
  INV_X1 U19442 ( .A(n19670), .ZN(n19683) );
  NAND2_X1 U19443 ( .A1(n19683), .A2(n19684), .ZN(n16018) );
  NAND2_X1 U19444 ( .A1(n16146), .A2(n16018), .ZN(n19680) );
  XOR2_X1 U19445 ( .A(n16019), .B(n19680), .Z(n16022) );
  AOI22_X1 U19446 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16249), .B2(P2_REIP_REG_21__SCAN_IN), .ZN(n16021) );
  NAND2_X1 U19447 ( .A1(n16272), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16020) );
  OAI211_X1 U19448 ( .C1(n16022), .C2(n17049), .A(n16021), .B(n16020), .ZN(
        n16023) );
  AOI211_X1 U19449 ( .C1(n16025), .C2(n19678), .A(n16024), .B(n16023), .ZN(
        n16026) );
  OAI21_X1 U19450 ( .B1(n16429), .B2(n16267), .A(n16026), .ZN(P2_U2834) );
  INV_X1 U19451 ( .A(n16027), .ZN(n16444) );
  NOR2_X1 U19452 ( .A1(n16028), .A2(n16270), .ZN(n16037) );
  AOI21_X1 U19453 ( .B1(n19681), .B2(n16029), .A(n19669), .ZN(n16035) );
  INV_X1 U19454 ( .A(n16034), .ZN(n16030) );
  NOR3_X1 U19455 ( .A1(n16219), .A2(n16030), .A3(n16029), .ZN(n16031) );
  AOI211_X1 U19456 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16031), .ZN(n16033) );
  AOI22_X1 U19457 ( .A1(n16272), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19671), .ZN(n16032) );
  OAI211_X1 U19458 ( .C1(n16035), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        n16036) );
  AOI211_X1 U19459 ( .C1(n16038), .C2(n19678), .A(n16037), .B(n16036), .ZN(
        n16039) );
  OAI21_X1 U19460 ( .B1(n16444), .B2(n16267), .A(n16039), .ZN(P2_U2836) );
  OAI21_X1 U19461 ( .B1(n11343), .B2(n10412), .A(n16040), .ZN(n16781) );
  NAND2_X1 U19462 ( .A1(n16779), .A2(n19678), .ZN(n16050) );
  AOI21_X1 U19463 ( .B1(n19681), .B2(n16051), .A(n19669), .ZN(n16046) );
  INV_X1 U19464 ( .A(n16045), .ZN(n16041) );
  NOR3_X1 U19465 ( .A1(n16219), .A2(n16041), .A3(n16051), .ZN(n16042) );
  AOI211_X1 U19466 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16042), .ZN(n16044) );
  AOI22_X1 U19467 ( .A1(n16272), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19671), .ZN(n16043) );
  OAI211_X1 U19468 ( .C1(n16046), .C2(n16045), .A(n16044), .B(n16043), .ZN(
        n16047) );
  AOI21_X1 U19469 ( .B1(n16048), .B2(n19676), .A(n16047), .ZN(n16049) );
  OAI211_X1 U19470 ( .C1(n16267), .C2(n16781), .A(n16050), .B(n16049), .ZN(
        P2_U2837) );
  INV_X1 U19471 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n16057) );
  AOI211_X1 U19472 ( .C1(n16054), .C2(n16052), .A(n16051), .B(n16219), .ZN(
        n16053) );
  AOI211_X1 U19473 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16053), .ZN(n16056) );
  AOI22_X1 U19474 ( .A1(n16054), .A2(n19669), .B1(n19671), .B2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16055) );
  OAI211_X1 U19475 ( .C1(n16057), .C2(n19667), .A(n16056), .B(n16055), .ZN(
        n16058) );
  AOI21_X1 U19476 ( .B1(n16059), .B2(n19676), .A(n16058), .ZN(n16061) );
  NAND2_X1 U19477 ( .A1(n16450), .A2(n19674), .ZN(n16060) );
  OAI211_X1 U19478 ( .C1(n16361), .C2(n16254), .A(n16061), .B(n16060), .ZN(
        P2_U2838) );
  NOR2_X1 U19479 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  AOI21_X1 U19480 ( .B1(n19681), .B2(n16075), .A(n19669), .ZN(n16069) );
  INV_X1 U19481 ( .A(n16070), .ZN(n16577) );
  NOR3_X1 U19482 ( .A1(n16219), .A2(n16075), .A3(n16577), .ZN(n16066) );
  AOI211_X1 U19483 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16066), .ZN(n16068) );
  AOI22_X1 U19484 ( .A1(n16272), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19671), .ZN(n16067) );
  OAI211_X1 U19485 ( .C1(n16070), .C2(n16069), .A(n16068), .B(n16067), .ZN(
        n16072) );
  NOR2_X1 U19486 ( .A1(n16788), .A2(n16254), .ZN(n16071) );
  AOI211_X1 U19487 ( .C1(n19676), .C2(n16073), .A(n16072), .B(n16071), .ZN(
        n16074) );
  OAI21_X1 U19488 ( .B1(n16786), .B2(n16267), .A(n16074), .ZN(P2_U2839) );
  AOI22_X1 U19489 ( .A1(n16272), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19671), .ZN(n16080) );
  OAI21_X1 U19490 ( .B1(n19664), .B2(n20435), .A(n11468), .ZN(n16078) );
  AOI211_X1 U19491 ( .C1(n16076), .C2(n16588), .A(n16075), .B(n16219), .ZN(
        n16077) );
  AOI211_X1 U19492 ( .C1(n19669), .C2(n16588), .A(n16078), .B(n16077), .ZN(
        n16079) );
  OAI211_X1 U19493 ( .C1(n16081), .C2(n16270), .A(n16080), .B(n16079), .ZN(
        n16082) );
  AOI21_X1 U19494 ( .B1(n16801), .B2(n19678), .A(n16082), .ZN(n16083) );
  OAI21_X1 U19495 ( .B1(n16084), .B2(n16267), .A(n16083), .ZN(P2_U2840) );
  NOR2_X1 U19496 ( .A1(n16085), .A2(n17002), .ZN(n16094) );
  XOR2_X1 U19497 ( .A(n16601), .B(n16094), .Z(n16089) );
  NAND2_X1 U19498 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16086) );
  OAI211_X1 U19499 ( .C1(n20433), .C2(n19664), .A(n16086), .B(n11468), .ZN(
        n16087) );
  AOI21_X1 U19500 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n16272), .A(n16087), .ZN(
        n16088) );
  OAI21_X1 U19501 ( .B1(n16089), .B2(n17049), .A(n16088), .ZN(n16091) );
  NOR2_X1 U19502 ( .A1(n16821), .A2(n16254), .ZN(n16090) );
  AOI211_X1 U19503 ( .C1(n19676), .C2(n16092), .A(n16091), .B(n16090), .ZN(
        n16093) );
  OAI21_X1 U19504 ( .B1(n16815), .B2(n16267), .A(n16093), .ZN(P2_U2841) );
  NAND2_X1 U19505 ( .A1(n16832), .A2(n19678), .ZN(n16105) );
  INV_X1 U19506 ( .A(n16094), .ZN(n16095) );
  AOI211_X1 U19507 ( .C1(n16098), .C2(n16096), .A(n17049), .B(n16095), .ZN(
        n16097) );
  AOI211_X1 U19508 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16097), .ZN(n16100) );
  AOI22_X1 U19509 ( .A1(n16098), .A2(n19669), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19671), .ZN(n16099) );
  OAI211_X1 U19510 ( .C1(n16101), .C2(n19667), .A(n16100), .B(n16099), .ZN(
        n16102) );
  AOI21_X1 U19511 ( .B1(n19676), .B2(n16103), .A(n16102), .ZN(n16104) );
  OAI211_X1 U19512 ( .C1(n16267), .C2(n16834), .A(n16105), .B(n16104), .ZN(
        P2_U2842) );
  INV_X1 U19513 ( .A(n16844), .ZN(n16115) );
  NOR2_X1 U19514 ( .A1(n16106), .A2(n16270), .ZN(n16114) );
  AOI21_X1 U19515 ( .B1(n16108), .B2(n19681), .A(n19669), .ZN(n16112) );
  INV_X1 U19516 ( .A(n16627), .ZN(n16107) );
  NOR3_X1 U19517 ( .A1(n16108), .A2(n16219), .A3(n16107), .ZN(n16109) );
  AOI211_X1 U19518 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16109), .ZN(n16111) );
  AOI22_X1 U19519 ( .A1(n16272), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19671), .ZN(n16110) );
  OAI211_X1 U19520 ( .C1(n16112), .C2(n16627), .A(n16111), .B(n16110), .ZN(
        n16113) );
  AOI211_X1 U19521 ( .C1(n16115), .C2(n19678), .A(n16114), .B(n16113), .ZN(
        n16116) );
  OAI21_X1 U19522 ( .B1(n16848), .B2(n16267), .A(n16116), .ZN(P2_U2843) );
  INV_X1 U19523 ( .A(n16117), .ZN(n16118) );
  AOI21_X1 U19524 ( .B1(n19681), .B2(n16118), .A(n19669), .ZN(n16123) );
  NOR3_X1 U19525 ( .A1(n16219), .A2(n16119), .A3(n16118), .ZN(n16120) );
  AOI211_X1 U19526 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n16249), .A(n19748), 
        .B(n16120), .ZN(n16122) );
  AOI22_X1 U19527 ( .A1(n16272), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19671), .ZN(n16121) );
  OAI211_X1 U19528 ( .C1(n16123), .C2(n16637), .A(n16122), .B(n16121), .ZN(
        n16124) );
  AOI21_X1 U19529 ( .B1(n16125), .B2(n19676), .A(n16124), .ZN(n16127) );
  NAND2_X1 U19530 ( .A1(n16860), .A2(n19674), .ZN(n16126) );
  OAI211_X1 U19531 ( .C1(n16858), .C2(n16254), .A(n16127), .B(n16126), .ZN(
        P2_U2844) );
  NAND2_X1 U19532 ( .A1(n16129), .A2(n19681), .ZN(n16128) );
  AOI21_X1 U19533 ( .B1(n16216), .B2(n16128), .A(n16130), .ZN(n16141) );
  INV_X1 U19534 ( .A(n16129), .ZN(n16131) );
  NAND2_X1 U19535 ( .A1(n16131), .A2(n16130), .ZN(n16139) );
  OAI22_X1 U19536 ( .A1(n16133), .A2(n16270), .B1(n16132), .B2(n19667), .ZN(
        n16134) );
  INV_X1 U19537 ( .A(n16134), .ZN(n16135) );
  OAI211_X1 U19538 ( .C1(n20426), .C2(n19664), .A(n16135), .B(n11468), .ZN(
        n16136) );
  INV_X1 U19539 ( .A(n16136), .ZN(n16138) );
  NAND2_X1 U19540 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16137) );
  OAI211_X1 U19541 ( .C1(n16219), .C2(n16139), .A(n16138), .B(n16137), .ZN(
        n16140) );
  AOI211_X1 U19542 ( .C1(n16142), .C2(n19678), .A(n16141), .B(n16140), .ZN(
        n16143) );
  OAI21_X1 U19543 ( .B1(n16144), .B2(n16267), .A(n16143), .ZN(P2_U2845) );
  NAND2_X1 U19544 ( .A1(n16146), .A2(n16145), .ZN(n16148) );
  XNOR2_X1 U19545 ( .A(n16148), .B(n16147), .ZN(n16152) );
  OAI21_X1 U19546 ( .B1(n19664), .B2(n20424), .A(n11468), .ZN(n16149) );
  AOI21_X1 U19547 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19671), .A(
        n16149), .ZN(n16150) );
  OAI21_X1 U19548 ( .B1(n10213), .B2(n19667), .A(n16150), .ZN(n16151) );
  AOI21_X1 U19549 ( .B1(n19681), .B2(n16152), .A(n16151), .ZN(n16153) );
  OAI21_X1 U19550 ( .B1(n16154), .B2(n16270), .A(n16153), .ZN(n16155) );
  AOI21_X1 U19551 ( .B1(n16871), .B2(n19678), .A(n16155), .ZN(n16156) );
  OAI21_X1 U19552 ( .B1(n16875), .B2(n16267), .A(n16156), .ZN(P2_U2846) );
  INV_X1 U19553 ( .A(n16883), .ZN(n16168) );
  OAI21_X1 U19554 ( .B1(n17049), .B2(n16159), .A(n16216), .ZN(n16163) );
  OAI22_X1 U19555 ( .A1(n16202), .A2(n16158), .B1(n16157), .B2(n19667), .ZN(
        n16162) );
  INV_X1 U19556 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n16671) );
  NAND3_X1 U19557 ( .A1(n16273), .A2(n16672), .A3(n16159), .ZN(n16160) );
  OAI211_X1 U19558 ( .C1(n16671), .C2(n19664), .A(n16160), .B(n11468), .ZN(
        n16161) );
  AOI211_X1 U19559 ( .C1(n16164), .C2(n16163), .A(n16162), .B(n16161), .ZN(
        n16165) );
  OAI21_X1 U19560 ( .B1(n16166), .B2(n16270), .A(n16165), .ZN(n16167) );
  AOI21_X1 U19561 ( .B1(n16168), .B2(n19678), .A(n16167), .ZN(n16169) );
  OAI21_X1 U19562 ( .B1(n16170), .B2(n16267), .A(n16169), .ZN(P2_U2847) );
  INV_X1 U19563 ( .A(n16899), .ZN(n16180) );
  OAI21_X1 U19564 ( .B1(n16172), .B2(n17049), .A(n16216), .ZN(n16176) );
  OAI22_X1 U19565 ( .A1(n16202), .A2(n16684), .B1(n10593), .B2(n19667), .ZN(
        n16175) );
  INV_X1 U19566 ( .A(n16686), .ZN(n16171) );
  NAND3_X1 U19567 ( .A1(n16273), .A2(n16172), .A3(n16171), .ZN(n16173) );
  OAI211_X1 U19568 ( .C1(n21760), .C2(n19664), .A(n16173), .B(n11468), .ZN(
        n16174) );
  AOI211_X1 U19569 ( .C1(n16686), .C2(n16176), .A(n16175), .B(n16174), .ZN(
        n16177) );
  OAI21_X1 U19570 ( .B1(n16178), .B2(n16270), .A(n16177), .ZN(n16179) );
  AOI21_X1 U19571 ( .B1(n16180), .B2(n19678), .A(n16179), .ZN(n16181) );
  OAI21_X1 U19572 ( .B1(n16895), .B2(n16267), .A(n16181), .ZN(P2_U2848) );
  INV_X1 U19573 ( .A(n16182), .ZN(n16183) );
  NAND2_X1 U19574 ( .A1(n16184), .A2(n16183), .ZN(n16190) );
  NOR2_X1 U19575 ( .A1(n17049), .A2(n16183), .ZN(n16186) );
  INV_X1 U19576 ( .A(n16184), .ZN(n16185) );
  OAI21_X1 U19577 ( .B1(n19669), .B2(n16186), .A(n16185), .ZN(n16189) );
  OAI21_X1 U19578 ( .B1(n20420), .B2(n19664), .A(n11468), .ZN(n16187) );
  INV_X1 U19579 ( .A(n16187), .ZN(n16188) );
  OAI211_X1 U19580 ( .C1(n16219), .C2(n16190), .A(n16189), .B(n16188), .ZN(
        n16193) );
  NAND2_X1 U19581 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16191) );
  OAI21_X1 U19582 ( .B1(n19667), .B2(n10574), .A(n16191), .ZN(n16192) );
  NOR2_X1 U19583 ( .A1(n16193), .A2(n16192), .ZN(n16194) );
  OAI21_X1 U19584 ( .B1(n16195), .B2(n16270), .A(n16194), .ZN(n16196) );
  AOI21_X1 U19585 ( .B1(n16197), .B2(n19678), .A(n16196), .ZN(n16198) );
  OAI21_X1 U19586 ( .B1(n16267), .B2(n16199), .A(n16198), .ZN(P2_U2849) );
  XNOR2_X1 U19587 ( .A(n16200), .B(n10418), .ZN(n16918) );
  INV_X1 U19588 ( .A(n16918), .ZN(n16476) );
  OAI21_X1 U19589 ( .B1(n16204), .B2(n17049), .A(n16216), .ZN(n16209) );
  OAI22_X1 U19590 ( .A1(n16202), .A2(n16201), .B1(n11371), .B2(n19667), .ZN(
        n16208) );
  INV_X1 U19591 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16206) );
  INV_X1 U19592 ( .A(n17374), .ZN(n16203) );
  NAND3_X1 U19593 ( .A1(n16273), .A2(n16204), .A3(n16203), .ZN(n16205) );
  OAI211_X1 U19594 ( .C1(n16206), .C2(n19664), .A(n16205), .B(n11468), .ZN(
        n16207) );
  AOI211_X1 U19595 ( .C1(n17374), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        n16210) );
  OAI21_X1 U19596 ( .B1(n16211), .B2(n16270), .A(n16210), .ZN(n16212) );
  AOI21_X1 U19597 ( .B1(n17376), .B2(n19678), .A(n16212), .ZN(n16213) );
  OAI21_X1 U19598 ( .B1(n16476), .B2(n16267), .A(n16213), .ZN(P2_U2850) );
  INV_X1 U19599 ( .A(n19753), .ZN(n16228) );
  OR2_X1 U19600 ( .A1(n16231), .A2(n16230), .ZN(n16233) );
  NAND2_X1 U19601 ( .A1(n16233), .A2(n16214), .ZN(n16215) );
  NAND2_X1 U19602 ( .A1(n16200), .A2(n16215), .ZN(n19689) );
  NOR2_X1 U19603 ( .A1(n19689), .A2(n16267), .ZN(n16227) );
  INV_X1 U19604 ( .A(n19757), .ZN(n16223) );
  INV_X1 U19605 ( .A(n16218), .ZN(n16217) );
  OAI21_X1 U19606 ( .B1(n17049), .B2(n16217), .A(n16216), .ZN(n16222) );
  INV_X1 U19607 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20417) );
  OAI21_X1 U19608 ( .B1(n19664), .B2(n20417), .A(n11468), .ZN(n16221) );
  NOR3_X1 U19609 ( .A1(n16219), .A2(n16218), .A3(n16223), .ZN(n16220) );
  AOI211_X1 U19610 ( .C1(n16223), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        n16225) );
  AOI22_X1 U19611 ( .A1(n16272), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19671), .ZN(n16224) );
  OAI211_X1 U19612 ( .C1(n16932), .C2(n16270), .A(n16225), .B(n16224), .ZN(
        n16226) );
  AOI211_X1 U19613 ( .C1(n16228), .C2(n19678), .A(n16227), .B(n16226), .ZN(
        n16229) );
  OAI21_X1 U19614 ( .B1(n19691), .B2(n16279), .A(n16229), .ZN(P2_U2851) );
  NAND2_X1 U19615 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  NAND2_X1 U19616 ( .A1(n16233), .A2(n16232), .ZN(n16957) );
  INV_X1 U19617 ( .A(n16234), .ZN(n16243) );
  NAND2_X1 U19618 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16235) );
  OAI21_X1 U19619 ( .B1(n19667), .B2(n10491), .A(n16235), .ZN(n16242) );
  INV_X1 U19620 ( .A(n17380), .ZN(n16236) );
  NAND3_X1 U19621 ( .A1(n16273), .A2(n16237), .A3(n16236), .ZN(n16240) );
  NOR2_X1 U19622 ( .A1(n16237), .A2(n17049), .ZN(n16238) );
  OAI21_X1 U19623 ( .B1(n19669), .B2(n16238), .A(n17380), .ZN(n16239) );
  OAI211_X1 U19624 ( .C1(n10772), .C2(n19664), .A(n16240), .B(n16239), .ZN(
        n16241) );
  AOI211_X1 U19625 ( .C1(n16243), .C2(n19676), .A(n16242), .B(n16241), .ZN(
        n16244) );
  OAI21_X1 U19626 ( .B1(n16957), .B2(n16267), .A(n16244), .ZN(n16245) );
  AOI21_X1 U19627 ( .B1(n16246), .B2(n19678), .A(n16245), .ZN(n16247) );
  OAI21_X1 U19628 ( .B1(n20124), .B2(n16279), .A(n16247), .ZN(P2_U2852) );
  NOR2_X1 U19629 ( .A1(n17002), .A2(n16248), .ZN(n16261) );
  XOR2_X1 U19630 ( .A(n19769), .B(n16261), .Z(n16253) );
  AOI22_X1 U19631 ( .A1(n19671), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16249), .B2(P2_REIP_REG_2__SCAN_IN), .ZN(n16252) );
  AOI22_X1 U19632 ( .A1(n16272), .A2(P2_EBX_REG_2__SCAN_IN), .B1(n16250), .B2(
        n19676), .ZN(n16251) );
  OAI211_X1 U19633 ( .C1(n16253), .C2(n17049), .A(n16252), .B(n16251), .ZN(
        n16256) );
  NOR2_X1 U19634 ( .A1(n19802), .A2(n16254), .ZN(n16255) );
  AOI211_X1 U19635 ( .C1(n19674), .C2(n20490), .A(n16256), .B(n16255), .ZN(
        n16257) );
  OAI21_X1 U19636 ( .B1(n17015), .B2(n16279), .A(n16257), .ZN(P2_U2853) );
  INV_X1 U19637 ( .A(n19704), .ZN(n16989) );
  OAI22_X1 U19638 ( .A1(n16270), .A2(n16258), .B1(n20412), .B2(n19664), .ZN(
        n16263) );
  NAND2_X1 U19639 ( .A1(n16995), .A2(n16259), .ZN(n16260) );
  NAND2_X1 U19640 ( .A1(n16261), .A2(n16260), .ZN(n17004) );
  NOR2_X1 U19641 ( .A1(n17004), .A2(n17049), .ZN(n16262) );
  AOI211_X1 U19642 ( .C1(n16264), .C2(n19669), .A(n16263), .B(n16262), .ZN(
        n16266) );
  AOI22_X1 U19643 ( .A1(n16272), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n19671), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16265) );
  OAI211_X1 U19644 ( .C1(n16989), .C2(n16267), .A(n16266), .B(n16265), .ZN(
        n16268) );
  AOI21_X1 U19645 ( .B1(n19678), .B2(n16966), .A(n16268), .ZN(n16269) );
  OAI21_X1 U19646 ( .B1(n19957), .B2(n16279), .A(n16269), .ZN(P2_U2854) );
  OAI22_X1 U19647 ( .A1(n16270), .A2(n17392), .B1(n10758), .B2(n19664), .ZN(
        n16271) );
  AOI21_X1 U19648 ( .B1(n19674), .B2(n17390), .A(n16271), .ZN(n16276) );
  AOI22_X1 U19649 ( .A1(n16273), .A2(n16995), .B1(n16272), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n16275) );
  OAI21_X1 U19650 ( .B1(n19669), .B2(n19671), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16274) );
  NAND3_X1 U19651 ( .A1(n16276), .A2(n16275), .A3(n16274), .ZN(n16277) );
  AOI21_X1 U19652 ( .B1(n19788), .B2(n19678), .A(n16277), .ZN(n16278) );
  OAI21_X1 U19653 ( .B1(n20090), .B2(n16279), .A(n16278), .ZN(P2_U2855) );
  MUX2_X1 U19654 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16280), .S(n16350), .Z(
        P2_U2856) );
  OR2_X1 U19655 ( .A1(n16282), .A2(n16281), .ZN(n16362) );
  NAND3_X1 U19656 ( .A1(n16362), .A2(n16283), .A3(n16357), .ZN(n16285) );
  NAND2_X1 U19657 ( .A1(n16360), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16284) );
  OAI211_X1 U19658 ( .C1(n16360), .C2(n16697), .A(n16285), .B(n16284), .ZN(
        P2_U2858) );
  NOR2_X1 U19659 ( .A1(n16287), .A2(n16286), .ZN(n16289) );
  XNOR2_X1 U19660 ( .A(n16289), .B(n16288), .ZN(n16377) );
  NOR2_X1 U19661 ( .A1(n15933), .A2(n16360), .ZN(n16290) );
  AOI21_X1 U19662 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16360), .A(n16290), .ZN(
        n16291) );
  OAI21_X1 U19663 ( .B1(n16377), .B2(n16353), .A(n16291), .ZN(P2_U2859) );
  OAI21_X1 U19664 ( .B1(n16294), .B2(n16293), .A(n16292), .ZN(n16384) );
  NOR2_X1 U19665 ( .A1(n16711), .A2(n16360), .ZN(n16295) );
  AOI21_X1 U19666 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16360), .A(n16295), .ZN(
        n16296) );
  OAI21_X1 U19667 ( .B1(n16353), .B2(n16384), .A(n16296), .ZN(P2_U2860) );
  NOR2_X1 U19668 ( .A1(n16297), .A2(n16308), .ZN(n16307) );
  NOR2_X1 U19669 ( .A1(n16307), .A2(n16298), .ZN(n16303) );
  NOR2_X1 U19670 ( .A1(n11127), .A2(n16299), .ZN(n16300) );
  XNOR2_X1 U19671 ( .A(n16301), .B(n16300), .ZN(n16302) );
  XNOR2_X1 U19672 ( .A(n16303), .B(n16302), .ZN(n16392) );
  NOR2_X1 U19673 ( .A1(n16304), .A2(n16360), .ZN(n16305) );
  AOI21_X1 U19674 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16360), .A(n16305), .ZN(
        n16306) );
  OAI21_X1 U19675 ( .B1(n16392), .B2(n16353), .A(n16306), .ZN(P2_U2861) );
  AOI21_X1 U19676 ( .B1(n16297), .B2(n16308), .A(n16307), .ZN(n16398) );
  NAND2_X1 U19677 ( .A1(n16398), .A2(n16357), .ZN(n16310) );
  NAND2_X1 U19678 ( .A1(n16360), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16309) );
  OAI211_X1 U19679 ( .C1(n16722), .C2(n16360), .A(n16310), .B(n16309), .ZN(
        P2_U2862) );
  INV_X1 U19680 ( .A(n16311), .ZN(n16314) );
  XOR2_X1 U19681 ( .A(n16313), .B(n16311), .Z(n16323) );
  NAND2_X1 U19682 ( .A1(n11051), .A2(n16312), .ZN(n16322) );
  NOR2_X1 U19683 ( .A1(n16323), .A2(n16322), .ZN(n16321) );
  AOI21_X1 U19684 ( .B1(n16314), .B2(n16313), .A(n16321), .ZN(n16318) );
  XNOR2_X1 U19685 ( .A(n16316), .B(n16315), .ZN(n16317) );
  XNOR2_X1 U19686 ( .A(n16318), .B(n16317), .ZN(n16407) );
  NOR2_X1 U19687 ( .A1(n16521), .A2(n16360), .ZN(n16319) );
  AOI21_X1 U19688 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16360), .A(n16319), .ZN(
        n16320) );
  OAI21_X1 U19689 ( .B1(n16407), .B2(n16353), .A(n16320), .ZN(P2_U2863) );
  AOI21_X1 U19690 ( .B1(n16323), .B2(n16322), .A(n16321), .ZN(n16412) );
  NAND2_X1 U19691 ( .A1(n16412), .A2(n16357), .ZN(n16325) );
  NAND2_X1 U19692 ( .A1(n16360), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16324) );
  OAI211_X1 U19693 ( .C1(n16736), .C2(n16360), .A(n16325), .B(n16324), .ZN(
        P2_U2864) );
  INV_X1 U19694 ( .A(n16556), .ZN(n16750) );
  NAND2_X1 U19695 ( .A1(n16338), .A2(n16330), .ZN(n16329) );
  NAND2_X1 U19696 ( .A1(n16329), .A2(n16326), .ZN(n16327) );
  AND2_X1 U19697 ( .A1(n16311), .A2(n16327), .ZN(n16420) );
  AOI22_X1 U19698 ( .A1(n16420), .A2(n16357), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16360), .ZN(n16328) );
  OAI21_X1 U19699 ( .B1(n16750), .B2(n16360), .A(n16328), .ZN(P2_U2865) );
  OAI21_X1 U19700 ( .B1(n16338), .B2(n16330), .A(n16329), .ZN(n16331) );
  INV_X1 U19701 ( .A(n16331), .ZN(n16427) );
  AOI22_X1 U19702 ( .A1(n16427), .A2(n16357), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16360), .ZN(n16332) );
  OAI21_X1 U19703 ( .B1(n16333), .B2(n16360), .A(n16332), .ZN(P2_U2866) );
  OAI21_X1 U19704 ( .B1(n16335), .B2(n16334), .A(n11568), .ZN(n19672) );
  INV_X1 U19705 ( .A(n16336), .ZN(n16340) );
  INV_X1 U19706 ( .A(n16337), .ZN(n16339) );
  AOI21_X1 U19707 ( .B1(n16340), .B2(n16339), .A(n16338), .ZN(n16436) );
  AOI22_X1 U19708 ( .A1(n16436), .A2(n16357), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n16360), .ZN(n16341) );
  OAI21_X1 U19709 ( .B1(n19672), .B2(n16360), .A(n16341), .ZN(P2_U2867) );
  INV_X1 U19710 ( .A(n16342), .ZN(n16344) );
  INV_X1 U19711 ( .A(n16343), .ZN(n16348) );
  AOI21_X1 U19712 ( .B1(n16344), .B2(n16348), .A(n16337), .ZN(n16442) );
  AOI22_X1 U19713 ( .A1(n16442), .A2(n16357), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16360), .ZN(n16345) );
  OAI21_X1 U19714 ( .B1(n16346), .B2(n16360), .A(n16345), .ZN(P2_U2868) );
  INV_X1 U19715 ( .A(n16347), .ZN(n16356) );
  NOR2_X1 U19716 ( .A1(n16355), .A2(n16356), .ZN(n16354) );
  OAI21_X1 U19717 ( .B1(n16354), .B2(n16349), .A(n16348), .ZN(n16446) );
  NAND2_X1 U19718 ( .A1(n16779), .A2(n16350), .ZN(n16352) );
  NAND2_X1 U19719 ( .A1(n16360), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16351) );
  OAI211_X1 U19720 ( .C1(n16446), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        P2_U2869) );
  AOI21_X1 U19721 ( .B1(n16356), .B2(n16355), .A(n16354), .ZN(n16456) );
  NAND2_X1 U19722 ( .A1(n16456), .A2(n16357), .ZN(n16359) );
  NAND2_X1 U19723 ( .A1(n16360), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16358) );
  OAI211_X1 U19724 ( .C1(n16361), .C2(n16360), .A(n16359), .B(n16358), .ZN(
        P2_U2870) );
  NAND3_X1 U19725 ( .A1(n16362), .A2(n16283), .A3(n19709), .ZN(n16369) );
  INV_X1 U19726 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16366) );
  AOI22_X1 U19727 ( .A1(n16459), .A2(n16363), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n16451), .ZN(n16365) );
  NAND2_X1 U19728 ( .A1(n16415), .A2(BUF2_REG_29__SCAN_IN), .ZN(n16364) );
  OAI211_X1 U19729 ( .C1(n16366), .C2(n16418), .A(n16365), .B(n16364), .ZN(
        n16367) );
  AOI21_X1 U19730 ( .B1(n16699), .B2(n19705), .A(n16367), .ZN(n16368) );
  NAND2_X1 U19731 ( .A1(n16369), .A2(n16368), .ZN(P2_U2890) );
  INV_X1 U19732 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16372) );
  AOI22_X1 U19733 ( .A1(n16459), .A2(n16370), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n16451), .ZN(n16371) );
  OAI21_X1 U19734 ( .B1(n16418), .B2(n16372), .A(n16371), .ZN(n16375) );
  NOR2_X1 U19735 ( .A1(n16373), .A2(n16468), .ZN(n16374) );
  OAI21_X1 U19736 ( .B1(n16377), .B2(n16462), .A(n16376), .ZN(P2_U2891) );
  INV_X1 U19737 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16380) );
  AOI22_X1 U19738 ( .A1(n16459), .A2(n16378), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n16451), .ZN(n16379) );
  OAI21_X1 U19739 ( .B1(n16418), .B2(n16380), .A(n16379), .ZN(n16382) );
  NOR2_X1 U19740 ( .A1(n16704), .A2(n16468), .ZN(n16381) );
  AOI211_X1 U19741 ( .C1(n16415), .C2(BUF2_REG_27__SCAN_IN), .A(n16382), .B(
        n16381), .ZN(n16383) );
  OAI21_X1 U19742 ( .B1(n16462), .B2(n16384), .A(n16383), .ZN(P2_U2892) );
  INV_X1 U19743 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16388) );
  AOI22_X1 U19744 ( .A1(n16459), .A2(n16385), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n16451), .ZN(n16387) );
  NAND2_X1 U19745 ( .A1(n16415), .A2(BUF2_REG_26__SCAN_IN), .ZN(n16386) );
  OAI211_X1 U19746 ( .C1(n16388), .C2(n16418), .A(n16387), .B(n16386), .ZN(
        n16389) );
  AOI21_X1 U19747 ( .B1(n16390), .B2(n19705), .A(n16389), .ZN(n16391) );
  OAI21_X1 U19748 ( .B1(n16392), .B2(n16462), .A(n16391), .ZN(P2_U2893) );
  INV_X1 U19749 ( .A(n16724), .ZN(n16400) );
  INV_X1 U19750 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U19751 ( .A1(n16459), .A2(n16393), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n16451), .ZN(n16395) );
  NAND2_X1 U19752 ( .A1(n16466), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16394) );
  OAI211_X1 U19753 ( .C1(n16461), .C2(n16396), .A(n16395), .B(n16394), .ZN(
        n16397) );
  AOI21_X1 U19754 ( .B1(n16398), .B2(n19709), .A(n16397), .ZN(n16399) );
  OAI21_X1 U19755 ( .B1(n16400), .B2(n16468), .A(n16399), .ZN(P2_U2894) );
  INV_X1 U19756 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n21666) );
  AOI22_X1 U19757 ( .A1(n16459), .A2(n16401), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n16451), .ZN(n16402) );
  OAI21_X1 U19758 ( .B1(n16418), .B2(n21666), .A(n16402), .ZN(n16405) );
  NOR2_X1 U19759 ( .A1(n16403), .A2(n16468), .ZN(n16404) );
  AOI211_X1 U19760 ( .C1(n16415), .C2(BUF2_REG_24__SCAN_IN), .A(n16405), .B(
        n16404), .ZN(n16406) );
  OAI21_X1 U19761 ( .B1(n16407), .B2(n16462), .A(n16406), .ZN(P2_U2895) );
  INV_X1 U19762 ( .A(n16741), .ZN(n16414) );
  INV_X1 U19763 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16410) );
  AOI22_X1 U19764 ( .A1(n16459), .A2(n19849), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n16451), .ZN(n16409) );
  NAND2_X1 U19765 ( .A1(n16466), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16408) );
  OAI211_X1 U19766 ( .C1(n16461), .C2(n16410), .A(n16409), .B(n16408), .ZN(
        n16411) );
  AOI21_X1 U19767 ( .B1(n16412), .B2(n19709), .A(n16411), .ZN(n16413) );
  OAI21_X1 U19768 ( .B1(n16414), .B2(n16468), .A(n16413), .ZN(P2_U2896) );
  INV_X1 U19769 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n17419) );
  NAND2_X1 U19770 ( .A1(n16415), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U19771 ( .A1(n16459), .A2(n19840), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n16451), .ZN(n16416) );
  OAI211_X1 U19772 ( .C1(n17419), .C2(n16418), .A(n16417), .B(n16416), .ZN(
        n16419) );
  AOI21_X1 U19773 ( .B1(n16420), .B2(n19709), .A(n16419), .ZN(n16421) );
  OAI21_X1 U19774 ( .B1(n16422), .B2(n16468), .A(n16421), .ZN(P2_U2897) );
  INV_X1 U19775 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16425) );
  AOI22_X1 U19776 ( .A1(n16459), .A2(n19835), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n16451), .ZN(n16424) );
  NAND2_X1 U19777 ( .A1(n16466), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16423) );
  OAI211_X1 U19778 ( .C1(n16461), .C2(n16425), .A(n16424), .B(n16423), .ZN(
        n16426) );
  AOI21_X1 U19779 ( .B1(n16427), .B2(n19709), .A(n16426), .ZN(n16428) );
  OAI21_X1 U19780 ( .B1(n16429), .B2(n16468), .A(n16428), .ZN(P2_U2898) );
  OAI21_X1 U19781 ( .B1(n16431), .B2(n16430), .A(n11565), .ZN(n19673) );
  INV_X1 U19782 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19783 ( .A1(n16459), .A2(n19830), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n16451), .ZN(n16433) );
  NAND2_X1 U19784 ( .A1(n16466), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16432) );
  OAI211_X1 U19785 ( .C1(n16461), .C2(n16434), .A(n16433), .B(n16432), .ZN(
        n16435) );
  AOI21_X1 U19786 ( .B1(n16436), .B2(n19709), .A(n16435), .ZN(n16437) );
  OAI21_X1 U19787 ( .B1(n19673), .B2(n16468), .A(n16437), .ZN(P2_U2899) );
  INV_X1 U19788 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16440) );
  AOI22_X1 U19789 ( .A1(n16459), .A2(n19825), .B1(P2_EAX_REG_19__SCAN_IN), 
        .B2(n16451), .ZN(n16439) );
  NAND2_X1 U19790 ( .A1(n16466), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16438) );
  OAI211_X1 U19791 ( .C1(n16461), .C2(n16440), .A(n16439), .B(n16438), .ZN(
        n16441) );
  AOI21_X1 U19792 ( .B1(n16442), .B2(n19709), .A(n16441), .ZN(n16443) );
  OAI21_X1 U19793 ( .B1(n16444), .B2(n16468), .A(n16443), .ZN(P2_U2900) );
  AOI22_X1 U19794 ( .A1(n16459), .A2(n17037), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n16451), .ZN(n16445) );
  OAI21_X1 U19795 ( .B1(n16461), .B2(n19040), .A(n16445), .ZN(n16448) );
  NOR2_X1 U19796 ( .A1(n16446), .A2(n16462), .ZN(n16447) );
  AOI211_X1 U19797 ( .C1(BUF1_REG_18__SCAN_IN), .C2(n16466), .A(n16448), .B(
        n16447), .ZN(n16449) );
  OAI21_X1 U19798 ( .B1(n16781), .B2(n16468), .A(n16449), .ZN(P2_U2901) );
  INV_X1 U19799 ( .A(n16450), .ZN(n16458) );
  INV_X1 U19800 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U19801 ( .A1(n16459), .A2(n19820), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n16451), .ZN(n16453) );
  NAND2_X1 U19802 ( .A1(n16466), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16452) );
  OAI211_X1 U19803 ( .C1(n16461), .C2(n16454), .A(n16453), .B(n16452), .ZN(
        n16455) );
  AOI21_X1 U19804 ( .B1(n16456), .B2(n19709), .A(n16455), .ZN(n16457) );
  OAI21_X1 U19805 ( .B1(n16458), .B2(n16468), .A(n16457), .ZN(P2_U2902) );
  AOI22_X1 U19806 ( .A1(n16459), .A2(n19814), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n16451), .ZN(n16460) );
  OAI21_X1 U19807 ( .B1(n16461), .B2(n19815), .A(n16460), .ZN(n16465) );
  NOR2_X1 U19808 ( .A1(n16463), .A2(n16462), .ZN(n16464) );
  AOI211_X1 U19809 ( .C1(BUF1_REG_16__SCAN_IN), .C2(n16466), .A(n16465), .B(
        n16464), .ZN(n16467) );
  OAI21_X1 U19810 ( .B1(n16786), .B2(n16468), .A(n16467), .ZN(P2_U2903) );
  INV_X1 U19811 ( .A(n16957), .ZN(n20485) );
  OAI21_X1 U19812 ( .B1(n20491), .B2(n20490), .A(n16469), .ZN(n19698) );
  XNOR2_X1 U19813 ( .A(n20486), .B(n16957), .ZN(n19699) );
  NAND2_X1 U19814 ( .A1(n19698), .A2(n19699), .ZN(n19697) );
  OAI21_X1 U19815 ( .B1(n20485), .B2(n20486), .A(n19697), .ZN(n16470) );
  NAND2_X1 U19816 ( .A1(n16470), .A2(n19689), .ZN(n19692) );
  INV_X1 U19817 ( .A(n19691), .ZN(n16471) );
  NAND3_X1 U19818 ( .A1(n19692), .A2(n16471), .A3(n19709), .ZN(n16474) );
  AOI22_X1 U19819 ( .A1(n16472), .A2(n19835), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n16451), .ZN(n16473) );
  OAI211_X1 U19820 ( .C1(n16476), .C2(n16475), .A(n16474), .B(n16473), .ZN(
        P2_U2914) );
  NAND2_X1 U19821 ( .A1(n16478), .A2(n16477), .ZN(n16480) );
  XOR2_X1 U19822 ( .A(n16480), .B(n16479), .Z(n16703) );
  INV_X1 U19823 ( .A(n16697), .ZN(n16484) );
  NAND2_X1 U19824 ( .A1(n19748), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16691) );
  NAND2_X1 U19825 ( .A1(n19779), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16481) );
  OAI211_X1 U19826 ( .C1(n19758), .C2(n16482), .A(n16691), .B(n16481), .ZN(
        n16483) );
  AOI21_X1 U19827 ( .B1(n16484), .B2(n19787), .A(n16483), .ZN(n16489) );
  NOR2_X2 U19828 ( .A1(n16487), .A2(n16486), .ZN(n16700) );
  NAND2_X1 U19829 ( .A1(n16700), .A2(n19781), .ZN(n16488) );
  OAI211_X1 U19830 ( .C1(n16703), .C2(n19785), .A(n16489), .B(n16488), .ZN(
        P2_U2985) );
  NAND2_X1 U19831 ( .A1(n19779), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16490) );
  OAI211_X1 U19832 ( .C1(n19758), .C2(n16492), .A(n16491), .B(n16490), .ZN(
        n16494) );
  NOR2_X1 U19833 ( .A1(n15933), .A2(n19774), .ZN(n16493) );
  AOI211_X1 U19834 ( .C1(n16495), .C2(n19781), .A(n16494), .B(n16493), .ZN(
        n16496) );
  OAI21_X1 U19835 ( .B1(n16497), .B2(n19785), .A(n16496), .ZN(P2_U2986) );
  XNOR2_X1 U19836 ( .A(n16498), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16716) );
  OR2_X1 U19837 ( .A1(n11468), .A2(n20455), .ZN(n16706) );
  NAND2_X1 U19838 ( .A1(n19779), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16501) );
  OAI211_X1 U19839 ( .C1(n19758), .C2(n16502), .A(n16706), .B(n16501), .ZN(
        n16504) );
  NOR2_X1 U19840 ( .A1(n16711), .A2(n19774), .ZN(n16503) );
  AOI211_X1 U19841 ( .C1(n16714), .C2(n19781), .A(n16504), .B(n16503), .ZN(
        n16505) );
  OAI21_X1 U19842 ( .B1(n16716), .B2(n19785), .A(n16505), .ZN(P2_U2987) );
  INV_X1 U19843 ( .A(n16506), .ZN(n16507) );
  NOR2_X1 U19844 ( .A1(n16508), .A2(n16507), .ZN(n16509) );
  XNOR2_X1 U19845 ( .A(n9739), .B(n16509), .ZN(n16728) );
  INV_X1 U19846 ( .A(n16722), .ZN(n16513) );
  NAND2_X1 U19847 ( .A1(n19748), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U19848 ( .A1(n19779), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16510) );
  OAI211_X1 U19849 ( .C1(n19758), .C2(n16511), .A(n16721), .B(n16510), .ZN(
        n16512) );
  AOI21_X1 U19850 ( .B1(n16513), .B2(n19787), .A(n16512), .ZN(n16516) );
  NAND2_X1 U19851 ( .A1(n16514), .A2(n16717), .ZN(n16725) );
  NAND3_X1 U19852 ( .A1(n9743), .A2(n19781), .A3(n16725), .ZN(n16515) );
  OAI211_X1 U19853 ( .C1(n19785), .C2(n16728), .A(n16516), .B(n16515), .ZN(
        P2_U2989) );
  OAI21_X1 U19854 ( .B1(n17388), .B2(n10278), .A(n16517), .ZN(n16518) );
  AOI21_X1 U19855 ( .B1(n19771), .B2(n16519), .A(n16518), .ZN(n16520) );
  OAI21_X1 U19856 ( .B1(n16521), .B2(n19774), .A(n16520), .ZN(n16522) );
  AOI21_X1 U19857 ( .B1(n16523), .B2(n19763), .A(n16522), .ZN(n16524) );
  OAI21_X1 U19858 ( .B1(n16690), .B2(n16525), .A(n16524), .ZN(P2_U2990) );
  INV_X1 U19859 ( .A(n16526), .ZN(n16527) );
  OAI21_X1 U19860 ( .B1(n16557), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16527), .ZN(n16743) );
  NAND2_X1 U19861 ( .A1(n19771), .A2(n16528), .ZN(n16529) );
  NAND2_X1 U19862 ( .A1(n19748), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16729) );
  OAI211_X1 U19863 ( .C1(n17388), .C2(n16530), .A(n16529), .B(n16729), .ZN(
        n16534) );
  AND2_X1 U19864 ( .A1(n16532), .A2(n16531), .ZN(n16737) );
  NOR3_X1 U19865 ( .A1(n16738), .A2(n16737), .A3(n19785), .ZN(n16533) );
  AOI211_X1 U19866 ( .C1(n19787), .C2(n16535), .A(n16534), .B(n16533), .ZN(
        n16536) );
  OAI21_X1 U19867 ( .B1(n16690), .B2(n16743), .A(n16536), .ZN(P2_U2991) );
  NOR2_X1 U19868 ( .A1(n16538), .A2(n16537), .ZN(n16552) );
  AOI21_X1 U19869 ( .B1(n16539), .B2(n16620), .A(n16540), .ZN(n16550) );
  INV_X1 U19870 ( .A(n16541), .ZN(n16547) );
  NAND2_X1 U19871 ( .A1(n16543), .A2(n16607), .ZN(n16546) );
  OR4_X1 U19872 ( .A1(n16547), .A2(n16546), .A3(n16545), .A4(n16544), .ZN(
        n16548) );
  NOR4_X1 U19873 ( .A1(n16550), .A2(n16549), .A3(n11560), .A4(n16548), .ZN(
        n16551) );
  XOR2_X1 U19874 ( .A(n16552), .B(n16551), .Z(n16757) );
  NOR2_X1 U19875 ( .A1(n11468), .A2(n20446), .ZN(n16744) );
  AOI21_X1 U19876 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16744), .ZN(n16553) );
  OAI21_X1 U19877 ( .B1(n19758), .B2(n16554), .A(n16553), .ZN(n16555) );
  AOI21_X1 U19878 ( .B1(n16556), .B2(n19787), .A(n16555), .ZN(n16559) );
  INV_X1 U19879 ( .A(n16557), .ZN(n16754) );
  NAND3_X1 U19880 ( .A1(n16754), .A2(n19781), .A3(n16753), .ZN(n16558) );
  OAI211_X1 U19881 ( .C1(n16757), .C2(n19785), .A(n16559), .B(n16558), .ZN(
        P2_U2992) );
  INV_X1 U19882 ( .A(n16560), .ZN(n16564) );
  OAI21_X1 U19883 ( .B1(n11560), .B2(n16562), .A(n16561), .ZN(n16563) );
  OAI21_X1 U19884 ( .B1(n16564), .B2(n11560), .A(n16563), .ZN(n16769) );
  INV_X1 U19885 ( .A(n16565), .ZN(n16567) );
  NOR2_X1 U19886 ( .A1(n11468), .A2(n19665), .ZN(n16763) );
  AOI21_X1 U19887 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16763), .ZN(n16569) );
  NAND2_X1 U19888 ( .A1(n19771), .A2(n19670), .ZN(n16568) );
  OAI211_X1 U19889 ( .C1(n19672), .C2(n19774), .A(n16569), .B(n16568), .ZN(
        n16570) );
  AOI21_X1 U19890 ( .B1(n16767), .B2(n19781), .A(n16570), .ZN(n16571) );
  OAI21_X1 U19891 ( .B1(n16769), .B2(n19785), .A(n16571), .ZN(P2_U2994) );
  XNOR2_X1 U19892 ( .A(n16592), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16581) );
  NOR2_X1 U19893 ( .A1(n16574), .A2(n16573), .ZN(n16791) );
  INV_X1 U19894 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16575) );
  OR2_X1 U19895 ( .A1(n11468), .A2(n20437), .ZN(n16787) );
  OAI21_X1 U19896 ( .B1(n17388), .B2(n16575), .A(n16787), .ZN(n16576) );
  AOI21_X1 U19897 ( .B1(n19771), .B2(n16577), .A(n16576), .ZN(n16578) );
  OAI21_X1 U19898 ( .B1(n16788), .B2(n19774), .A(n16578), .ZN(n16579) );
  AOI21_X1 U19899 ( .B1(n16791), .B2(n19763), .A(n16579), .ZN(n16580) );
  OAI21_X1 U19900 ( .B1(n16690), .B2(n16581), .A(n16580), .ZN(P2_U2998) );
  INV_X1 U19901 ( .A(n16597), .ZN(n16583) );
  AOI21_X1 U19902 ( .B1(n16600), .B2(n16598), .A(n16583), .ZN(n16587) );
  NAND2_X1 U19903 ( .A1(n16585), .A2(n16584), .ZN(n16586) );
  XNOR2_X1 U19904 ( .A(n16587), .B(n16586), .ZN(n16809) );
  NAND2_X1 U19905 ( .A1(n16588), .A2(n19771), .ZN(n16589) );
  NAND2_X1 U19906 ( .A1(n19748), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16798) );
  OAI211_X1 U19907 ( .C1(n17388), .C2(n16590), .A(n16589), .B(n16798), .ZN(
        n16591) );
  AOI21_X1 U19908 ( .B1(n16801), .B2(n19787), .A(n16591), .ZN(n16594) );
  AOI21_X1 U19909 ( .B1(n16799), .B2(n16596), .A(n16592), .ZN(n16806) );
  NAND2_X1 U19910 ( .A1(n16806), .A2(n19781), .ZN(n16593) );
  OAI211_X1 U19911 ( .C1(n16809), .C2(n19785), .A(n16594), .B(n16593), .ZN(
        P2_U2999) );
  INV_X1 U19912 ( .A(n16818), .ZN(n16595) );
  OAI21_X1 U19913 ( .B1(n16610), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16596), .ZN(n16827) );
  NAND2_X1 U19914 ( .A1(n16598), .A2(n16597), .ZN(n16599) );
  XNOR2_X1 U19915 ( .A(n16600), .B(n16599), .ZN(n16810) );
  NOR2_X1 U19916 ( .A1(n11468), .A2(n20433), .ZN(n16816) );
  NOR2_X1 U19917 ( .A1(n19758), .A2(n16601), .ZN(n16602) );
  AOI211_X1 U19918 ( .C1(n19779), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16816), .B(n16602), .ZN(n16603) );
  OAI21_X1 U19919 ( .B1(n16821), .B2(n19774), .A(n16603), .ZN(n16604) );
  AOI21_X1 U19920 ( .B1(n16810), .B2(n19763), .A(n16604), .ZN(n16605) );
  OAI21_X1 U19921 ( .B1(n16827), .B2(n16690), .A(n16605), .ZN(P2_U3000) );
  NAND2_X1 U19922 ( .A1(n16607), .A2(n16606), .ZN(n16608) );
  XNOR2_X1 U19923 ( .A(n16609), .B(n16608), .ZN(n16840) );
  NOR2_X1 U19924 ( .A1(n16611), .A2(n16610), .ZN(n16828) );
  NAND2_X1 U19925 ( .A1(n16828), .A2(n19781), .ZN(n16616) );
  NOR2_X1 U19926 ( .A1(n11468), .A2(n21718), .ZN(n16831) );
  AOI21_X1 U19927 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16831), .ZN(n16612) );
  OAI21_X1 U19928 ( .B1(n19758), .B2(n16613), .A(n16612), .ZN(n16614) );
  AOI21_X1 U19929 ( .B1(n16832), .B2(n19787), .A(n16614), .ZN(n16615) );
  OAI211_X1 U19930 ( .C1(n19785), .C2(n16840), .A(n16616), .B(n16615), .ZN(
        P2_U3001) );
  XNOR2_X1 U19931 ( .A(n16632), .B(n10204), .ZN(n16852) );
  INV_X1 U19932 ( .A(n16617), .ZN(n16619) );
  NOR2_X1 U19933 ( .A1(n16619), .A2(n16618), .ZN(n16626) );
  AND2_X1 U19934 ( .A1(n16621), .A2(n16620), .ZN(n16624) );
  OR2_X1 U19935 ( .A1(n16539), .A2(n16622), .ZN(n16623) );
  OAI22_X1 U19936 ( .A1(n16626), .A2(n16625), .B1(n16624), .B2(n16623), .ZN(
        n16850) );
  NOR2_X1 U19937 ( .A1(n11468), .A2(n20430), .ZN(n16841) );
  NOR2_X1 U19938 ( .A1(n19758), .A2(n16627), .ZN(n16628) );
  AOI211_X1 U19939 ( .C1(n19779), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16841), .B(n16628), .ZN(n16629) );
  OAI21_X1 U19940 ( .B1(n16844), .B2(n19774), .A(n16629), .ZN(n16630) );
  AOI21_X1 U19941 ( .B1(n16850), .B2(n19763), .A(n16630), .ZN(n16631) );
  OAI21_X1 U19942 ( .B1(n16852), .B2(n16690), .A(n16631), .ZN(P2_U3002) );
  OAI21_X1 U19943 ( .B1(n16633), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16632), .ZN(n16867) );
  NAND2_X1 U19944 ( .A1(n16635), .A2(n16634), .ZN(n16636) );
  XOR2_X1 U19945 ( .A(n16636), .B(n11553), .Z(n16865) );
  NOR2_X1 U19946 ( .A1(n11468), .A2(n20428), .ZN(n16853) );
  NOR2_X1 U19947 ( .A1(n19758), .A2(n16637), .ZN(n16638) );
  AOI211_X1 U19948 ( .C1(n19779), .C2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16853), .B(n16638), .ZN(n16639) );
  OAI21_X1 U19949 ( .B1(n16858), .B2(n19774), .A(n16639), .ZN(n16640) );
  AOI21_X1 U19950 ( .B1(n16865), .B2(n19763), .A(n16640), .ZN(n16641) );
  OAI21_X1 U19951 ( .B1(n16867), .B2(n16690), .A(n16641), .ZN(P2_U3003) );
  OAI21_X1 U19952 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16643), .A(
        n16642), .ZN(n16879) );
  INV_X1 U19953 ( .A(n16644), .ZN(n16649) );
  NAND2_X1 U19954 ( .A1(n16648), .A2(n16645), .ZN(n16646) );
  AOI22_X1 U19955 ( .A1(n16649), .A2(n16648), .B1(n16647), .B2(n16646), .ZN(
        n16877) );
  NAND2_X1 U19956 ( .A1(n16871), .A2(n19787), .ZN(n16651) );
  NOR2_X1 U19957 ( .A1(n11468), .A2(n20424), .ZN(n16870) );
  AOI21_X1 U19958 ( .B1(n19779), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16870), .ZN(n16650) );
  OAI211_X1 U19959 ( .C1(n19758), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        n16653) );
  AOI21_X1 U19960 ( .B1(n16877), .B2(n19763), .A(n16653), .ZN(n16654) );
  OAI21_X1 U19961 ( .B1(n16879), .B2(n16690), .A(n16654), .ZN(P2_U3005) );
  AND2_X1 U19962 ( .A1(n16656), .A2(n16655), .ZN(n16659) );
  XNOR2_X1 U19963 ( .A(n16659), .B(n16657), .ZN(n16677) );
  AOI22_X1 U19964 ( .A1(n16677), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16659), .B2(n16658), .ZN(n16662) );
  XNOR2_X1 U19965 ( .A(n16660), .B(n16886), .ZN(n16661) );
  XNOR2_X1 U19966 ( .A(n16662), .B(n16661), .ZN(n16894) );
  NAND2_X1 U19967 ( .A1(n16664), .A2(n16663), .ZN(n16670) );
  INV_X1 U19968 ( .A(n16665), .ZN(n16666) );
  AOI21_X1 U19969 ( .B1(n16668), .B2(n16667), .A(n16666), .ZN(n16681) );
  NAND2_X1 U19970 ( .A1(n16681), .A2(n16678), .ZN(n16683) );
  NAND2_X1 U19971 ( .A1(n16683), .A2(n16679), .ZN(n16669) );
  XOR2_X1 U19972 ( .A(n16670), .B(n16669), .Z(n16891) );
  NOR2_X1 U19973 ( .A1(n11468), .A2(n16671), .ZN(n16880) );
  NOR2_X1 U19974 ( .A1(n19758), .A2(n16672), .ZN(n16673) );
  AOI211_X1 U19975 ( .C1(n19779), .C2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16880), .B(n16673), .ZN(n16674) );
  OAI21_X1 U19976 ( .B1(n16883), .B2(n19774), .A(n16674), .ZN(n16675) );
  AOI21_X1 U19977 ( .B1(n16891), .B2(n19763), .A(n16675), .ZN(n16676) );
  OAI21_X1 U19978 ( .B1(n16894), .B2(n16690), .A(n16676), .ZN(P2_U3006) );
  XNOR2_X1 U19979 ( .A(n16677), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16906) );
  INV_X1 U19980 ( .A(n16679), .ZN(n16682) );
  AND2_X1 U19981 ( .A1(n16679), .A2(n16678), .ZN(n16680) );
  OAI22_X1 U19982 ( .A1(n16683), .A2(n16682), .B1(n16681), .B2(n16680), .ZN(
        n16903) );
  NOR2_X1 U19983 ( .A1(n11468), .A2(n21760), .ZN(n16896) );
  NOR2_X1 U19984 ( .A1(n17388), .A2(n16684), .ZN(n16685) );
  AOI211_X1 U19985 ( .C1(n16686), .C2(n19771), .A(n16896), .B(n16685), .ZN(
        n16687) );
  OAI21_X1 U19986 ( .B1(n16899), .B2(n19774), .A(n16687), .ZN(n16688) );
  AOI21_X1 U19987 ( .B1(n16903), .B2(n19763), .A(n16688), .ZN(n16689) );
  OAI21_X1 U19988 ( .B1(n16906), .B2(n16690), .A(n16689), .ZN(P2_U3007) );
  XNOR2_X1 U19989 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16692) );
  OAI21_X1 U19990 ( .B1(n16693), .B2(n16692), .A(n16691), .ZN(n16694) );
  AOI21_X1 U19991 ( .B1(n16695), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16694), .ZN(n16696) );
  OAI21_X1 U19992 ( .B1(n16697), .B2(n19803), .A(n16696), .ZN(n16698) );
  AOI21_X1 U19993 ( .B1(n19792), .B2(n16699), .A(n16698), .ZN(n16702) );
  NAND2_X1 U19994 ( .A1(n16700), .A2(n19796), .ZN(n16701) );
  OAI211_X1 U19995 ( .C1(n16703), .C2(n17400), .A(n16702), .B(n16701), .ZN(
        P2_U3017) );
  NOR2_X1 U19996 ( .A1(n16704), .A2(n16958), .ZN(n16713) );
  OR3_X1 U19997 ( .A1(n16718), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16705), .ZN(n16707) );
  NAND2_X1 U19998 ( .A1(n16707), .A2(n16706), .ZN(n16708) );
  AOI21_X1 U19999 ( .B1(n16709), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16708), .ZN(n16710) );
  OAI21_X1 U20000 ( .B1(n16711), .B2(n19803), .A(n16710), .ZN(n16712) );
  OAI21_X1 U20001 ( .B1(n16716), .B2(n17400), .A(n16715), .ZN(P2_U3019) );
  MUX2_X1 U20002 ( .A(n16719), .B(n16718), .S(n16717), .Z(n16720) );
  OAI211_X1 U20003 ( .C1(n16722), .C2(n19803), .A(n16721), .B(n16720), .ZN(
        n16723) );
  AOI21_X1 U20004 ( .B1(n19792), .B2(n16724), .A(n16723), .ZN(n16727) );
  NAND3_X1 U20005 ( .A1(n9743), .A2(n19796), .A3(n16725), .ZN(n16726) );
  OAI211_X1 U20006 ( .C1(n16728), .C2(n17400), .A(n16727), .B(n16726), .ZN(
        P2_U3021) );
  INV_X1 U20007 ( .A(n16729), .ZN(n16734) );
  INV_X1 U20008 ( .A(n16730), .ZN(n16731) );
  AOI211_X1 U20009 ( .C1(n16732), .C2(n21707), .A(n16731), .B(n16747), .ZN(
        n16733) );
  AOI211_X1 U20010 ( .C1(n16745), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16734), .B(n16733), .ZN(n16735) );
  OAI21_X1 U20011 ( .B1(n16736), .B2(n19803), .A(n16735), .ZN(n16740) );
  NOR3_X1 U20012 ( .A1(n16738), .A2(n16737), .A3(n17400), .ZN(n16739) );
  AOI211_X1 U20013 ( .C1(n19792), .C2(n16741), .A(n16740), .B(n16739), .ZN(
        n16742) );
  OAI21_X1 U20014 ( .B1(n16942), .B2(n16743), .A(n16742), .ZN(P2_U3023) );
  INV_X1 U20015 ( .A(n16744), .ZN(n16749) );
  INV_X1 U20016 ( .A(n16745), .ZN(n16746) );
  MUX2_X1 U20017 ( .A(n16747), .B(n16746), .S(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n16748) );
  OAI211_X1 U20018 ( .C1(n16750), .C2(n19803), .A(n16749), .B(n16748), .ZN(
        n16751) );
  AOI21_X1 U20019 ( .B1(n19792), .B2(n16752), .A(n16751), .ZN(n16756) );
  NAND3_X1 U20020 ( .A1(n16754), .A2(n19796), .A3(n16753), .ZN(n16755) );
  NOR2_X1 U20021 ( .A1(n19672), .A2(n19803), .ZN(n16764) );
  AOI21_X1 U20022 ( .B1(n16777), .B2(n16759), .A(n16758), .ZN(n16762) );
  NOR3_X1 U20023 ( .A1(n16760), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16868), .ZN(n16761) );
  NOR4_X1 U20024 ( .A1(n16764), .A2(n16763), .A3(n16762), .A4(n16761), .ZN(
        n16765) );
  OAI21_X1 U20025 ( .B1(n16958), .B2(n19673), .A(n16765), .ZN(n16766) );
  OAI21_X1 U20026 ( .B1(n16769), .B2(n17400), .A(n16768), .ZN(P2_U3026) );
  INV_X1 U20027 ( .A(n16770), .ZN(n16783) );
  INV_X1 U20028 ( .A(n16771), .ZN(n16775) );
  NAND3_X1 U20029 ( .A1(n16773), .A2(n16772), .A3(n16776), .ZN(n16774) );
  OAI211_X1 U20030 ( .C1(n16777), .C2(n16776), .A(n16775), .B(n16774), .ZN(
        n16778) );
  AOI21_X1 U20031 ( .B1(n16779), .B2(n16967), .A(n16778), .ZN(n16780) );
  OAI21_X1 U20032 ( .B1(n16958), .B2(n16781), .A(n16780), .ZN(n16782) );
  AOI21_X1 U20033 ( .B1(n16783), .B2(n19796), .A(n16782), .ZN(n16784) );
  NOR2_X1 U20034 ( .A1(n16786), .A2(n16958), .ZN(n16790) );
  OAI21_X1 U20035 ( .B1(n16788), .B2(n19803), .A(n16787), .ZN(n16789) );
  AOI211_X1 U20036 ( .C1(n16791), .C2(n11071), .A(n16790), .B(n16789), .ZN(
        n16794) );
  NAND2_X1 U20037 ( .A1(n16792), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16793) );
  OAI211_X1 U20038 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16795), .A(
        n16794), .B(n16793), .ZN(P2_U3030) );
  NAND2_X1 U20039 ( .A1(n16796), .A2(n16799), .ZN(n16797) );
  OAI211_X1 U20040 ( .C1(n16800), .C2(n16799), .A(n16798), .B(n16797), .ZN(
        n16804) );
  INV_X1 U20041 ( .A(n16801), .ZN(n16802) );
  NOR2_X1 U20042 ( .A1(n16802), .A2(n19803), .ZN(n16803) );
  AOI211_X1 U20043 ( .C1(n16805), .C2(n19792), .A(n16804), .B(n16803), .ZN(
        n16808) );
  NAND2_X1 U20044 ( .A1(n16806), .A2(n19796), .ZN(n16807) );
  OAI211_X1 U20045 ( .C1(n16809), .C2(n17400), .A(n16808), .B(n16807), .ZN(
        P2_U3031) );
  AND2_X1 U20046 ( .A1(n16810), .A2(n11071), .ZN(n16825) );
  INV_X1 U20047 ( .A(n16813), .ZN(n16854) );
  NAND2_X1 U20048 ( .A1(n16811), .A2(n16854), .ZN(n16812) );
  NAND2_X1 U20049 ( .A1(n16862), .A2(n16812), .ZN(n16846) );
  INV_X1 U20050 ( .A(n16842), .ZN(n16830) );
  NOR2_X1 U20051 ( .A1(n16830), .A2(n16818), .ZN(n16814) );
  OR2_X1 U20052 ( .A1(n16846), .A2(n16814), .ZN(n16837) );
  AND2_X1 U20053 ( .A1(n16837), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16824) );
  NOR2_X1 U20054 ( .A1(n16815), .A2(n16958), .ZN(n16823) );
  INV_X1 U20055 ( .A(n16816), .ZN(n16820) );
  NAND3_X1 U20056 ( .A1(n16842), .A2(n16818), .A3(n16817), .ZN(n16819) );
  OAI211_X1 U20057 ( .C1(n16821), .C2(n19803), .A(n16820), .B(n16819), .ZN(
        n16822) );
  NOR4_X1 U20058 ( .A1(n16825), .A2(n16824), .A3(n16823), .A4(n16822), .ZN(
        n16826) );
  OAI21_X1 U20059 ( .B1(n16942), .B2(n16827), .A(n16826), .ZN(P2_U3032) );
  NAND2_X1 U20060 ( .A1(n16828), .A2(n19796), .ZN(n16839) );
  OAI21_X1 U20061 ( .B1(n16830), .B2(n10204), .A(n16829), .ZN(n16836) );
  AOI21_X1 U20062 ( .B1(n16832), .B2(n16967), .A(n16831), .ZN(n16833) );
  OAI21_X1 U20063 ( .B1(n16958), .B2(n16834), .A(n16833), .ZN(n16835) );
  AOI21_X1 U20064 ( .B1(n16837), .B2(n16836), .A(n16835), .ZN(n16838) );
  AOI21_X1 U20065 ( .B1(n16842), .B2(n10204), .A(n16841), .ZN(n16843) );
  OAI21_X1 U20066 ( .B1(n16844), .B2(n19803), .A(n16843), .ZN(n16845) );
  AOI21_X1 U20067 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16846), .A(
        n16845), .ZN(n16847) );
  OAI21_X1 U20068 ( .B1(n16848), .B2(n16958), .A(n16847), .ZN(n16849) );
  AOI21_X1 U20069 ( .B1(n16850), .B2(n11071), .A(n16849), .ZN(n16851) );
  OAI21_X1 U20070 ( .B1(n16852), .B2(n16942), .A(n16851), .ZN(P2_U3034) );
  INV_X1 U20071 ( .A(n16853), .ZN(n16857) );
  OAI211_X1 U20072 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16855), .B(n16854), .ZN(
        n16856) );
  OAI211_X1 U20073 ( .C1(n16858), .C2(n19803), .A(n16857), .B(n16856), .ZN(
        n16859) );
  AOI21_X1 U20074 ( .B1(n19792), .B2(n16860), .A(n16859), .ZN(n16861) );
  OAI21_X1 U20075 ( .B1(n16863), .B2(n16862), .A(n16861), .ZN(n16864) );
  AOI21_X1 U20076 ( .B1(n16865), .B2(n11071), .A(n16864), .ZN(n16866) );
  OAI21_X1 U20077 ( .B1(n16867), .B2(n16942), .A(n16866), .ZN(P2_U3035) );
  NOR2_X1 U20078 ( .A1(n16868), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16869) );
  AOI211_X1 U20079 ( .C1(n16871), .C2(n16967), .A(n16870), .B(n16869), .ZN(
        n16874) );
  NAND2_X1 U20080 ( .A1(n16872), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16873) );
  OAI211_X1 U20081 ( .C1(n16958), .C2(n16875), .A(n16874), .B(n16873), .ZN(
        n16876) );
  AOI21_X1 U20082 ( .B1(n16877), .B2(n11071), .A(n16876), .ZN(n16878) );
  OAI21_X1 U20083 ( .B1(n16879), .B2(n16942), .A(n16878), .ZN(P2_U3037) );
  INV_X1 U20084 ( .A(n16880), .ZN(n16882) );
  NAND4_X1 U20085 ( .A1(n16886), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n16884), .ZN(n16881) );
  OAI211_X1 U20086 ( .C1(n16883), .C2(n19803), .A(n16882), .B(n16881), .ZN(
        n16889) );
  INV_X1 U20087 ( .A(n16902), .ZN(n16887) );
  NAND3_X1 U20088 ( .A1(n16885), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16884), .ZN(n16898) );
  AOI21_X1 U20089 ( .B1(n16887), .B2(n16898), .A(n16886), .ZN(n16888) );
  AOI211_X1 U20090 ( .C1(n19792), .C2(n16890), .A(n16889), .B(n16888), .ZN(
        n16893) );
  NAND2_X1 U20091 ( .A1(n16891), .A2(n11071), .ZN(n16892) );
  OAI211_X1 U20092 ( .C1(n16894), .C2(n16942), .A(n16893), .B(n16892), .ZN(
        P2_U3038) );
  NOR2_X1 U20093 ( .A1(n16895), .A2(n16958), .ZN(n16901) );
  INV_X1 U20094 ( .A(n16896), .ZN(n16897) );
  OAI211_X1 U20095 ( .C1(n16899), .C2(n19803), .A(n16898), .B(n16897), .ZN(
        n16900) );
  AOI211_X1 U20096 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16902), .A(
        n16901), .B(n16900), .ZN(n16905) );
  NAND2_X1 U20097 ( .A1(n16903), .A2(n11071), .ZN(n16904) );
  OAI211_X1 U20098 ( .C1(n16906), .C2(n16942), .A(n16905), .B(n16904), .ZN(
        P2_U3039) );
  OAI21_X1 U20099 ( .B1(n9765), .B2(n16908), .A(n16907), .ZN(n16909) );
  OAI21_X1 U20100 ( .B1(n16910), .B2(n9765), .A(n16909), .ZN(n16911) );
  INV_X1 U20101 ( .A(n16911), .ZN(n17375) );
  NAND2_X1 U20102 ( .A1(n17375), .A2(n19796), .ZN(n16925) );
  INV_X1 U20103 ( .A(n16936), .ZN(n16917) );
  NOR2_X1 U20104 ( .A1(n16206), .A2(n11468), .ZN(n16916) );
  INV_X1 U20105 ( .A(n16912), .ZN(n16938) );
  AOI211_X1 U20106 ( .C1(n16914), .C2(n16937), .A(n16913), .B(n16938), .ZN(
        n16915) );
  AOI211_X1 U20107 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n16917), .A(
        n16916), .B(n16915), .ZN(n16924) );
  AOI22_X1 U20108 ( .A1(n17376), .A2(n16967), .B1(n19792), .B2(n16918), .ZN(
        n16923) );
  INV_X1 U20109 ( .A(n16919), .ZN(n16920) );
  XNOR2_X1 U20110 ( .A(n16921), .B(n16920), .ZN(n17377) );
  NAND2_X1 U20111 ( .A1(n17377), .A2(n11071), .ZN(n16922) );
  NAND4_X1 U20112 ( .A1(n16925), .A2(n16924), .A3(n16923), .A4(n16922), .ZN(
        P2_U3041) );
  XNOR2_X1 U20113 ( .A(n16926), .B(n16937), .ZN(n19749) );
  INV_X1 U20114 ( .A(n19749), .ZN(n16943) );
  INV_X1 U20115 ( .A(n16927), .ZN(n16929) );
  NAND2_X1 U20116 ( .A1(n16929), .A2(n16928), .ZN(n16945) );
  NAND2_X1 U20117 ( .A1(n16927), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16944) );
  NAND2_X1 U20118 ( .A1(n16944), .A2(n16930), .ZN(n16931) );
  NAND2_X1 U20119 ( .A1(n16945), .A2(n16931), .ZN(n16934) );
  XNOR2_X1 U20120 ( .A(n16932), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16933) );
  XNOR2_X1 U20121 ( .A(n16934), .B(n16933), .ZN(n19750) );
  NAND2_X1 U20122 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19748), .ZN(n16935) );
  OAI221_X1 U20123 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16938), .C1(
        n16937), .C2(n16936), .A(n16935), .ZN(n16940) );
  OAI22_X1 U20124 ( .A1(n16958), .A2(n19689), .B1(n19753), .B2(n19803), .ZN(
        n16939) );
  AOI211_X1 U20125 ( .C1(n19750), .C2(n11071), .A(n16940), .B(n16939), .ZN(
        n16941) );
  OAI21_X1 U20126 ( .B1(n16943), .B2(n16942), .A(n16941), .ZN(P2_U3042) );
  NAND2_X1 U20127 ( .A1(n16945), .A2(n16944), .ZN(n16947) );
  XNOR2_X1 U20128 ( .A(n16947), .B(n16946), .ZN(n17385) );
  AND3_X1 U20129 ( .A1(n17382), .A2(n19796), .A3(n17381), .ZN(n16960) );
  INV_X1 U20130 ( .A(n16950), .ZN(n16951) );
  NAND2_X1 U20131 ( .A1(n16970), .A2(n16951), .ZN(n16953) );
  MUX2_X1 U20132 ( .A(n16953), .B(n16952), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n16956) );
  OAI22_X1 U20133 ( .A1(n19803), .A2(n10100), .B1(n10772), .B2(n11468), .ZN(
        n16954) );
  INV_X1 U20134 ( .A(n16954), .ZN(n16955) );
  OAI211_X1 U20135 ( .C1(n16958), .C2(n16957), .A(n16956), .B(n16955), .ZN(
        n16959) );
  AOI211_X1 U20136 ( .C1(n17385), .C2(n11071), .A(n16960), .B(n16959), .ZN(
        n16961) );
  INV_X1 U20137 ( .A(n16961), .ZN(P2_U3043) );
  OAI22_X1 U20138 ( .A1(n19806), .A2(n16963), .B1(n17400), .B2(n16962), .ZN(
        n16964) );
  AOI211_X1 U20139 ( .C1(n16967), .C2(n16966), .A(n16965), .B(n16964), .ZN(
        n16973) );
  AOI22_X1 U20140 ( .A1(n19796), .A2(n16968), .B1(n19792), .B2(n19704), .ZN(
        n16972) );
  OAI211_X1 U20141 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16970), .B(n16969), .ZN(n16971) );
  NAND3_X1 U20142 ( .A1(n16973), .A2(n16972), .A3(n16971), .ZN(P2_U3045) );
  INV_X1 U20143 ( .A(n16986), .ZN(n16977) );
  INV_X1 U20144 ( .A(n16974), .ZN(n20259) );
  AOI21_X1 U20145 ( .B1(n16975), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n20259), 
        .ZN(n16976) );
  OAI21_X1 U20146 ( .B1(n20090), .B2(n16977), .A(n16976), .ZN(n16983) );
  OAI21_X1 U20147 ( .B1(n20501), .B2(P2_FLUSH_REG_SCAN_IN), .A(n16980), .ZN(
        n16981) );
  INV_X1 U20148 ( .A(n16981), .ZN(n16982) );
  MUX2_X1 U20149 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16983), .S(
        n20495), .Z(P2_U3605) );
  INV_X1 U20150 ( .A(n20476), .ZN(n16987) );
  INV_X1 U20151 ( .A(n16984), .ZN(n16985) );
  NAND2_X1 U20152 ( .A1(n16986), .A2(n16985), .ZN(n20480) );
  MUX2_X1 U20153 ( .A(n16987), .B(n20480), .S(n20479), .Z(n16988) );
  OAI21_X1 U20154 ( .B1(n16989), .B2(n12673), .A(n16988), .ZN(n16990) );
  MUX2_X1 U20155 ( .A(n16990), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n20498), .Z(P2_U3604) );
  NAND3_X1 U20156 ( .A1(n11449), .A2(n11138), .A3(n16991), .ZN(n16992) );
  OAI211_X1 U20157 ( .C1(n16994), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n16993), 
        .B(n16992), .ZN(n16999) );
  MUX2_X1 U20158 ( .A(n16995), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(
        n17002), .Z(n16996) );
  NAND2_X1 U20159 ( .A1(n16996), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17010) );
  INV_X1 U20160 ( .A(n17019), .ZN(n16997) );
  AOI22_X1 U20161 ( .A1(n16999), .A2(n17010), .B1(n16998), .B2(n16997), .ZN(
        n17001) );
  NAND2_X1 U20162 ( .A1(n17020), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17000) );
  OAI21_X1 U20163 ( .B1(n17001), .B2(n17020), .A(n17000), .ZN(P2_U3601) );
  INV_X1 U20164 ( .A(n17010), .ZN(n17005) );
  NAND2_X1 U20165 ( .A1(n17002), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17003) );
  AND2_X1 U20166 ( .A1(n17004), .A2(n17003), .ZN(n17011) );
  AOI22_X1 U20167 ( .A1(n17006), .A2(n17009), .B1(n17005), .B2(n17011), .ZN(
        n17007) );
  OAI21_X1 U20168 ( .B1(n19957), .B2(n17019), .A(n17007), .ZN(n17008) );
  MUX2_X1 U20169 ( .A(n17008), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n17020), .Z(P2_U3600) );
  INV_X1 U20170 ( .A(n17009), .ZN(n17043) );
  OAI22_X1 U20171 ( .A1(n17012), .A2(n17043), .B1(n17011), .B2(n17010), .ZN(
        n17013) );
  INV_X1 U20172 ( .A(n17013), .ZN(n17014) );
  OAI21_X1 U20173 ( .B1(n17015), .B2(n17019), .A(n17014), .ZN(n17016) );
  MUX2_X1 U20174 ( .A(n17016), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17020), .Z(P2_U3599) );
  INV_X1 U20175 ( .A(n17017), .ZN(n17018) );
  OAI22_X1 U20176 ( .A1(n20124), .A2(n17019), .B1(n17018), .B2(n17043), .ZN(
        n17021) );
  MUX2_X1 U20177 ( .A(n17021), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17020), .Z(P2_U3596) );
  NAND2_X1 U20178 ( .A1(n21570), .A2(n20497), .ZN(n19919) );
  INV_X1 U20179 ( .A(n19848), .ZN(n17030) );
  OAI21_X1 U20180 ( .B1(n17033), .B2(n20508), .A(n12673), .ZN(n17026) );
  INV_X1 U20181 ( .A(n20484), .ZN(n20478) );
  NOR3_X1 U20182 ( .A1(n20389), .A2(n19880), .A3(n20478), .ZN(n17022) );
  AND2_X1 U20183 ( .A1(n20484), .A2(n20512), .ZN(n20091) );
  NOR2_X1 U20184 ( .A1(n17022), .A2(n20091), .ZN(n17036) );
  AND2_X1 U20185 ( .A1(n17030), .A2(n20328), .ZN(n17035) );
  INV_X1 U20186 ( .A(n17035), .ZN(n17023) );
  NOR2_X1 U20187 ( .A1(n17036), .A2(n17023), .ZN(n17024) );
  INV_X1 U20188 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17040) );
  INV_X1 U20189 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21597) );
  OAI22_X2 U20190 ( .A1(n21597), .A2(n19851), .B1(n19040), .B2(n19850), .ZN(
        n20354) );
  INV_X1 U20191 ( .A(n20389), .ZN(n17031) );
  OR2_X1 U20192 ( .A1(n19847), .A2(n10734), .ZN(n19871) );
  OAI22_X1 U20193 ( .A1(n17031), .A2(n20308), .B1(n17030), .B2(n19871), .ZN(
        n17032) );
  AOI21_X1 U20194 ( .B1(n19880), .B2(n20354), .A(n17032), .ZN(n17039) );
  OAI21_X1 U20195 ( .B1(n17033), .B2(n19848), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17034) );
  NAND2_X1 U20196 ( .A1(n19853), .A2(n20352), .ZN(n17038) );
  OAI211_X1 U20197 ( .C1(n19857), .C2(n17040), .A(n17039), .B(n17038), .ZN(
        P2_U3050) );
  OAI21_X1 U20198 ( .B1(n17042), .B2(n17041), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n17050) );
  NOR3_X1 U20199 ( .A1(n20509), .A2(n17044), .A3(n17043), .ZN(n17046) );
  OAI21_X1 U20200 ( .B1(n17047), .B2(n17046), .A(n17045), .ZN(n17048) );
  NAND3_X1 U20201 ( .A1(n17050), .A2(n17049), .A3(n17048), .ZN(P2_U3177) );
  OAI21_X1 U20202 ( .B1(n17052), .B2(n17063), .A(n17051), .ZN(n17069) );
  INV_X1 U20203 ( .A(n17089), .ZN(n17054) );
  NOR2_X1 U20204 ( .A1(n17054), .A2(n18648), .ZN(n17056) );
  INV_X1 U20205 ( .A(n18772), .ZN(n17055) );
  AOI211_X1 U20206 ( .C1(n19409), .C2(n17053), .A(n17056), .B(n17055), .ZN(
        n17092) );
  INV_X1 U20207 ( .A(n17092), .ZN(n17057) );
  AOI21_X1 U20208 ( .B1(n18620), .B2(n10088), .A(n17057), .ZN(n17077) );
  INV_X1 U20209 ( .A(n17053), .ZN(n17058) );
  NAND2_X1 U20210 ( .A1(n18650), .A2(n17058), .ZN(n17075) );
  XOR2_X1 U20211 ( .A(n17067), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17060) );
  OAI21_X1 U20212 ( .B1(n17075), .B2(n17060), .A(n17059), .ZN(n17061) );
  AOI21_X1 U20213 ( .B1(n18714), .B2(n11593), .A(n17061), .ZN(n17066) );
  OAI21_X1 U20214 ( .B1(n17096), .B2(n17063), .A(n17062), .ZN(n17064) );
  NAND2_X1 U20215 ( .A1(n17064), .A2(n18725), .ZN(n17065) );
  OAI211_X1 U20216 ( .C1(n17077), .C2(n17067), .A(n17066), .B(n17065), .ZN(
        n17068) );
  AOI21_X1 U20217 ( .B1(n17069), .B2(n18792), .A(n17068), .ZN(n17070) );
  OAI21_X1 U20218 ( .B1(n17071), .B2(n18748), .A(n17070), .ZN(P3_U2799) );
  AND2_X1 U20219 ( .A1(n17187), .A2(n18792), .ZN(n17088) );
  INV_X1 U20220 ( .A(n17088), .ZN(n17074) );
  NAND2_X1 U20221 ( .A1(n17189), .A2(n18725), .ZN(n17097) );
  NAND2_X1 U20222 ( .A1(n17074), .A2(n17097), .ZN(n17099) );
  NOR3_X1 U20223 ( .A1(n17104), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n10165), .ZN(n17082) );
  INV_X1 U20224 ( .A(n17075), .ZN(n17076) );
  NAND2_X1 U20225 ( .A1(n17076), .A2(n17505), .ZN(n17080) );
  NOR2_X1 U20226 ( .A1(n10420), .A2(n21720), .ZN(n17194) );
  NOR2_X1 U20227 ( .A1(n10415), .A2(n17194), .ZN(n17079) );
  OR2_X1 U20228 ( .A1(n17077), .A2(n17505), .ZN(n17078) );
  NAND3_X1 U20229 ( .A1(n17080), .A2(n17079), .A3(n17078), .ZN(n17081) );
  AOI21_X1 U20230 ( .B1(n17099), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17083), .ZN(n17084) );
  OAI21_X1 U20231 ( .B1(n17197), .B2(n18748), .A(n17084), .ZN(P3_U2800) );
  OAI21_X1 U20232 ( .B1(n17086), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17085), .ZN(n17208) );
  NAND2_X1 U20233 ( .A1(n17088), .A2(n17087), .ZN(n17095) );
  AOI21_X1 U20234 ( .B1(n9821), .B2(n19409), .A(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17091) );
  OR3_X1 U20235 ( .A1(n17089), .A2(n18615), .A3(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17090) );
  NAND2_X1 U20236 ( .A1(n9696), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17203) );
  OAI211_X1 U20237 ( .C1(n17092), .C2(n17091), .A(n17090), .B(n17203), .ZN(
        n17093) );
  AOI21_X1 U20238 ( .B1(n18714), .B2(n17515), .A(n17093), .ZN(n17094) );
  OAI211_X1 U20239 ( .C1(n17097), .C2(n17096), .A(n17095), .B(n17094), .ZN(
        n17098) );
  AOI21_X1 U20240 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17099), .A(
        n17098), .ZN(n17100) );
  OAI21_X1 U20241 ( .B1(n18748), .B2(n17208), .A(n17100), .ZN(P3_U2801) );
  NAND2_X1 U20242 ( .A1(n17101), .A2(n13524), .ZN(n17102) );
  XNOR2_X1 U20243 ( .A(n17102), .B(n18703), .ZN(n17225) );
  INV_X1 U20244 ( .A(n17538), .ZN(n17109) );
  NAND2_X1 U20245 ( .A1(n17103), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17108) );
  NAND2_X1 U20246 ( .A1(n9696), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17209) );
  OAI21_X1 U20247 ( .B1(n17104), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17209), .ZN(n17105) );
  XOR2_X1 U20248 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n17110), .Z(
        n18799) );
  INV_X1 U20249 ( .A(n17111), .ZN(n17112) );
  NOR3_X1 U20250 ( .A1(n17113), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n17112), .ZN(n17119) );
  AOI21_X1 U20251 ( .B1(n17114), .B2(n19409), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17116) );
  OAI21_X1 U20252 ( .B1(n18714), .B2(n18620), .A(n17550), .ZN(n17115) );
  NAND2_X1 U20253 ( .A1(n9696), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18801) );
  OAI211_X1 U20254 ( .C1(n17117), .C2(n17116), .A(n17115), .B(n18801), .ZN(
        n17118) );
  AOI211_X1 U20255 ( .C1(n17120), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17119), .B(n17118), .ZN(n17121) );
  OAI21_X1 U20256 ( .B1(n18748), .B2(n18799), .A(n17121), .ZN(P3_U2804) );
  OAI21_X1 U20257 ( .B1(n18587), .B2(n18734), .A(n18636), .ZN(n17122) );
  XOR2_X1 U20258 ( .A(n17122), .B(n18637), .Z(n17236) );
  INV_X1 U20259 ( .A(n17236), .ZN(n17128) );
  INV_X1 U20260 ( .A(n18601), .ZN(n18659) );
  AOI22_X1 U20261 ( .A1(n18792), .A2(n17226), .B1(n18725), .B2(n18899), .ZN(
        n18658) );
  OAI21_X1 U20262 ( .B1(n17229), .B2(n18659), .A(n18658), .ZN(n17130) );
  INV_X1 U20263 ( .A(n17229), .ZN(n18588) );
  NOR2_X1 U20264 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18588), .ZN(
        n17234) );
  AOI22_X1 U20265 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17130), .B1(
        n18601), .B2(n17234), .ZN(n17127) );
  NOR2_X1 U20266 ( .A1(n18593), .A2(n17123), .ZN(n18630) );
  INV_X1 U20267 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17649) );
  AOI21_X1 U20268 ( .B1(n18647), .B2(n17123), .A(n17055), .ZN(n17134) );
  OAI21_X1 U20269 ( .B1(n17131), .B2(n18648), .A(n17134), .ZN(n18634) );
  INV_X1 U20270 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19569) );
  NOR2_X1 U20271 ( .A1(n17649), .A2(n17124), .ZN(n17628) );
  INV_X1 U20272 ( .A(n17628), .ZN(n17629) );
  OAI21_X1 U20273 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17131), .A(
        n17629), .ZN(n17643) );
  OAI22_X1 U20274 ( .A1(n10420), .A2(n19569), .B1(n18696), .B2(n17643), .ZN(
        n17125) );
  AOI221_X1 U20275 ( .B1(n18630), .B2(n17649), .C1(n18634), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17125), .ZN(n17126) );
  OAI211_X1 U20276 ( .C1(n18748), .C2(n17128), .A(n17127), .B(n17126), .ZN(
        P3_U2812) );
  XNOR2_X1 U20277 ( .A(n17129), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17245) );
  INV_X1 U20278 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18894) );
  NOR2_X1 U20279 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18894), .ZN(
        n17242) );
  AOI22_X1 U20280 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17130), .B1(
        n18601), .B2(n17242), .ZN(n17138) );
  AOI21_X1 U20281 ( .B1(n17132), .B2(n17650), .A(n17131), .ZN(n17653) );
  AOI21_X1 U20282 ( .B1(n17133), .B2(n19409), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17135) );
  NAND2_X1 U20283 ( .A1(n9696), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17243) );
  OAI21_X1 U20284 ( .B1(n17135), .B2(n17134), .A(n17243), .ZN(n17136) );
  AOI21_X1 U20285 ( .B1(n17653), .B2(n18790), .A(n17136), .ZN(n17137) );
  OAI211_X1 U20286 ( .C1(n18748), .C2(n17245), .A(n17138), .B(n17137), .ZN(
        P3_U2813) );
  NAND2_X1 U20287 ( .A1(n17139), .A2(n18956), .ZN(n17142) );
  XNOR2_X1 U20288 ( .A(n17142), .B(n18734), .ZN(n19001) );
  INV_X1 U20289 ( .A(n19001), .ZN(n17149) );
  AOI21_X1 U20290 ( .B1(n17141), .B2(n18993), .A(n17140), .ZN(n18997) );
  INV_X1 U20291 ( .A(n17142), .ZN(n18995) );
  AOI22_X1 U20292 ( .A1(n18997), .A2(n18792), .B1(n18725), .B2(n18995), .ZN(
        n17148) );
  INV_X1 U20293 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17760) );
  INV_X1 U20294 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17768) );
  NOR2_X1 U20295 ( .A1(n17143), .A2(n17768), .ZN(n17144) );
  NAND2_X1 U20296 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17144), .ZN(
        n17150) );
  NOR2_X1 U20297 ( .A1(n17760), .A2(n17150), .ZN(n17742) );
  AOI21_X1 U20298 ( .B1(n17760), .B2(n17150), .A(n17742), .ZN(n17753) );
  AOI21_X1 U20299 ( .B1(n18647), .B2(n17143), .A(n17055), .ZN(n18690) );
  NAND2_X1 U20300 ( .A1(n9696), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n19004) );
  OAI211_X1 U20301 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17144), .A(
        n19409), .B(n17743), .ZN(n17145) );
  OAI211_X1 U20302 ( .C1(n18690), .C2(n17760), .A(n19004), .B(n17145), .ZN(
        n17146) );
  AOI21_X1 U20303 ( .B1(n17753), .B2(n18790), .A(n17146), .ZN(n17147) );
  OAI211_X1 U20304 ( .C1(n17149), .C2(n18748), .A(n17148), .B(n17147), .ZN(
        P3_U2822) );
  NAND2_X1 U20305 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17151), .ZN(
        n17792) );
  NOR2_X1 U20306 ( .A1(n21610), .A2(n17792), .ZN(n17782) );
  OAI21_X1 U20307 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17782), .A(
        n17150), .ZN(n17771) );
  NAND2_X1 U20308 ( .A1(n19409), .A2(n17151), .ZN(n18765) );
  NOR2_X1 U20309 ( .A1(n21610), .A2(n18765), .ZN(n18753) );
  INV_X1 U20310 ( .A(n18690), .ZN(n17153) );
  AOI221_X1 U20311 ( .B1(n18753), .B2(n17768), .C1(n17153), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17152), .ZN(n17157) );
  INV_X1 U20312 ( .A(n18786), .ZN(n17181) );
  AOI22_X1 U20313 ( .A1(n17155), .A2(n18792), .B1(n17181), .B2(n17154), .ZN(
        n17156) );
  OAI211_X1 U20314 ( .C1(n18776), .C2(n17771), .A(n17157), .B(n17156), .ZN(
        P3_U2823) );
  OAI21_X1 U20315 ( .B1(n18786), .B2(n17159), .A(n17158), .ZN(n17164) );
  NOR2_X1 U20316 ( .A1(n17860), .A2(n17169), .ZN(n17160) );
  INV_X1 U20317 ( .A(n17161), .ZN(n17808) );
  NAND2_X1 U20318 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17808), .ZN(
        n17806) );
  OAI21_X1 U20319 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17160), .A(
        n17806), .ZN(n17821) );
  AOI21_X1 U20320 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18772), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17162) );
  AOI21_X1 U20321 ( .B1(n18647), .B2(n17161), .A(n17055), .ZN(n18795) );
  OAI22_X1 U20322 ( .A1(n18776), .A2(n17821), .B1(n17162), .B2(n18795), .ZN(
        n17163) );
  AOI211_X1 U20323 ( .C1(n18792), .C2(n17165), .A(n17164), .B(n17163), .ZN(
        n17166) );
  INV_X1 U20324 ( .A(n17166), .ZN(P3_U2827) );
  NAND2_X1 U20325 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17055), .ZN(
        n17168) );
  OAI211_X1 U20326 ( .C1(n19313), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17168), .B(n17167), .ZN(n17172) );
  AOI22_X1 U20327 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17169), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17860), .ZN(n17841) );
  OAI22_X1 U20328 ( .A1(n18776), .A2(n17841), .B1(n18701), .B2(n17170), .ZN(
        n17171) );
  AOI211_X1 U20329 ( .C1(n17181), .C2(n17173), .A(n17172), .B(n17171), .ZN(
        n17174) );
  INV_X1 U20330 ( .A(n17174), .ZN(P3_U2828) );
  XNOR2_X1 U20331 ( .A(n17176), .B(n17175), .ZN(n17247) );
  XOR2_X1 U20332 ( .A(n17177), .B(n17176), .Z(n17251) );
  NAND2_X1 U20333 ( .A1(n17181), .A2(n17251), .ZN(n17178) );
  NAND2_X1 U20334 ( .A1(n9696), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17246) );
  OAI211_X1 U20335 ( .C1(n17247), .C2(n18701), .A(n17178), .B(n17246), .ZN(
        n17179) );
  AOI21_X1 U20336 ( .B1(n18764), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n17179), .ZN(n17180) );
  OAI21_X1 U20337 ( .B1(n18776), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n17180), .ZN(P3_U2829) );
  NAND2_X1 U20338 ( .A1(n17181), .A2(n17186), .ZN(n17185) );
  NAND3_X1 U20339 ( .A1(n18425), .A2(n18648), .A3(n18772), .ZN(n17183) );
  AOI21_X1 U20340 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17183), .A(
        n17182), .ZN(n17184) );
  OAI211_X1 U20341 ( .C1(n17186), .C2(n18701), .A(n17185), .B(n17184), .ZN(
        P3_U2830) );
  INV_X1 U20342 ( .A(n17187), .ZN(n17188) );
  NOR2_X1 U20343 ( .A1(n17188), .A2(n17248), .ZN(n17190) );
  OAI21_X1 U20344 ( .B1(n17190), .B2(n18926), .A(n17189), .ZN(n17201) );
  NAND2_X1 U20345 ( .A1(n17201), .A2(n17191), .ZN(n17195) );
  INV_X1 U20346 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17192) );
  NOR3_X1 U20347 ( .A1(n17204), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17192), .ZN(n17193) );
  AOI211_X1 U20348 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17195), .A(
        n17194), .B(n17193), .ZN(n17196) );
  OAI21_X1 U20349 ( .B1(n17197), .B2(n18976), .A(n17196), .ZN(P3_U2832) );
  NAND3_X1 U20350 ( .A1(n17198), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17216), .ZN(n17199) );
  AOI21_X1 U20351 ( .B1(n19010), .B2(n17199), .A(n19008), .ZN(n17200) );
  OAI211_X1 U20352 ( .C1(n17202), .C2(n19006), .A(n17201), .B(n17200), .ZN(
        n17206) );
  OAI21_X1 U20353 ( .B1(n17204), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17203), .ZN(n17205) );
  AOI21_X1 U20354 ( .B1(n17206), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17205), .ZN(n17207) );
  OAI21_X1 U20355 ( .B1(n18976), .B2(n17208), .A(n17207), .ZN(P3_U2833) );
  INV_X1 U20356 ( .A(n17209), .ZN(n17223) );
  INV_X1 U20357 ( .A(n18822), .ZN(n17213) );
  OAI22_X1 U20358 ( .A1(n17211), .A2(n18933), .B1(n17210), .B2(n18931), .ZN(
        n17212) );
  AOI21_X1 U20359 ( .B1(n17214), .B2(n17213), .A(n17212), .ZN(n17219) );
  NOR2_X1 U20360 ( .A1(n17228), .A2(n17215), .ZN(n18821) );
  AOI21_X1 U20361 ( .B1(n18810), .B2(n18821), .A(n18822), .ZN(n18806) );
  INV_X1 U20362 ( .A(n17216), .ZN(n17217) );
  NOR2_X1 U20363 ( .A1(n18806), .A2(n17217), .ZN(n17218) );
  INV_X1 U20364 ( .A(n18797), .ZN(n18835) );
  AOI21_X1 U20365 ( .B1(n18835), .B2(n17220), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17221) );
  AOI211_X1 U20366 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18804), .A(
        n19006), .B(n17221), .ZN(n17222) );
  OAI21_X1 U20367 ( .B1(n17225), .B2(n18976), .A(n17224), .ZN(P3_U2835) );
  AOI22_X1 U20368 ( .A1(n19465), .A2(n17226), .B1(n18996), .B2(n18899), .ZN(
        n18854) );
  NAND2_X1 U20369 ( .A1(n18951), .A2(n18854), .ZN(n18893) );
  NOR2_X1 U20370 ( .A1(n17228), .A2(n17227), .ZN(n17230) );
  NOR2_X1 U20371 ( .A1(n19465), .A2(n18996), .ZN(n18957) );
  OAI22_X1 U20372 ( .A1(n18822), .A2(n17230), .B1(n17229), .B2(n18957), .ZN(
        n17231) );
  AOI211_X2 U20373 ( .C1(n10299), .C2(n17232), .A(n18893), .B(n17231), .ZN(
        n17240) );
  AOI221_X1 U20374 ( .B1(n18822), .B2(n17240), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17240), .A(n9696), .ZN(
        n17235) );
  NOR2_X1 U20375 ( .A1(n18980), .A2(n17233), .ZN(n18994) );
  NOR2_X1 U20376 ( .A1(n18644), .A2(n18992), .ZN(n18895) );
  AOI22_X1 U20377 ( .A1(n17236), .A2(n19002), .B1(n9696), .B2(
        P3_REIP_REG_18__SCAN_IN), .ZN(n17237) );
  NAND2_X1 U20378 ( .A1(n17238), .A2(n17237), .ZN(P3_U2844) );
  NOR3_X1 U20379 ( .A1(n9696), .A2(n17240), .A3(n17239), .ZN(n17241) );
  AOI21_X1 U20380 ( .B1(n18895), .B2(n17242), .A(n17241), .ZN(n17244) );
  OAI211_X1 U20381 ( .C1(n18976), .C2(n17245), .A(n17244), .B(n17243), .ZN(
        P3_U2845) );
  INV_X1 U20382 ( .A(n17246), .ZN(n17250) );
  NOR2_X1 U20383 ( .A1(n17248), .A2(n17247), .ZN(n17249) );
  AOI211_X1 U20384 ( .C1(n17252), .C2(n17251), .A(n17250), .B(n17249), .ZN(
        n17256) );
  OAI211_X1 U20385 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18981), .A(
        n19010), .B(n13253), .ZN(n17255) );
  OAI21_X1 U20386 ( .B1(n17253), .B2(n19008), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17254) );
  NAND3_X1 U20387 ( .A1(n17256), .A2(n17255), .A3(n17254), .ZN(P3_U2861) );
  NAND2_X1 U20388 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19175) );
  AOI221_X1 U20389 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19175), .C1(n17258), 
        .C2(n19175), .A(n17257), .ZN(n19026) );
  NOR2_X1 U20390 ( .A1(n17259), .A2(n19478), .ZN(n17260) );
  OAI21_X1 U20391 ( .B1(n17260), .B2(n19090), .A(n19027), .ZN(n19024) );
  AOI22_X1 U20392 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19026), .B1(
        n19024), .B2(n19028), .ZN(P3_U2865) );
  INV_X1 U20393 ( .A(n17261), .ZN(n17304) );
  NOR3_X1 U20394 ( .A1(n17263), .A2(n21677), .A3(n17262), .ZN(n17268) );
  AOI21_X1 U20395 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17268), .A(
        n17264), .ZN(n17266) );
  NAND2_X1 U20396 ( .A1(n17266), .A2(n17265), .ZN(n17267) );
  OAI21_X1 U20397 ( .B1(n17268), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17267), .ZN(n17270) );
  INV_X1 U20398 ( .A(n17270), .ZN(n17269) );
  NOR2_X1 U20399 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17269), .ZN(
        n17271) );
  OAI22_X1 U20400 ( .A1(n17272), .A2(n17271), .B1(n17270), .B2(n21066), .ZN(
        n17274) );
  AOI21_X1 U20401 ( .B1(n17274), .B2(n17273), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17276) );
  NOR2_X1 U20402 ( .A1(n17274), .A2(n17273), .ZN(n17275) );
  INV_X1 U20403 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20768) );
  OAI21_X1 U20404 ( .B1(n17276), .B2(n17275), .A(n20768), .ZN(n17286) );
  INV_X1 U20405 ( .A(n17277), .ZN(n17281) );
  OAI21_X1 U20406 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17278), .ZN(n17279) );
  AND4_X1 U20407 ( .A1(n17282), .A2(n17281), .A3(n17280), .A4(n17279), .ZN(
        n17283) );
  AND2_X1 U20408 ( .A1(n17284), .A2(n17283), .ZN(n17285) );
  INV_X1 U20409 ( .A(n17298), .ZN(n17294) );
  OAI21_X1 U20410 ( .B1(n17287), .B2(n21487), .A(n21370), .ZN(n17293) );
  INV_X1 U20411 ( .A(n17288), .ZN(n17291) );
  NAND3_X1 U20412 ( .A1(n17291), .A2(n17290), .A3(n17289), .ZN(n17292) );
  NAND2_X1 U20413 ( .A1(n17293), .A2(n17292), .ZN(n17365) );
  NOR3_X1 U20414 ( .A1(n17295), .A2(n21660), .A3(n17368), .ZN(n17296) );
  NOR2_X1 U20415 ( .A1(n17371), .A2(n17296), .ZN(n17302) );
  OAI21_X1 U20416 ( .B1(n17298), .B2(n21370), .A(n17297), .ZN(n17299) );
  AOI21_X1 U20417 ( .B1(n21378), .B2(n21306), .A(n17299), .ZN(n17300) );
  NAND2_X1 U20418 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17300), .ZN(n17301) );
  OAI22_X1 U20419 ( .A1(n17302), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n17371), 
        .B2(n17301), .ZN(n17303) );
  NAND2_X1 U20420 ( .A1(n17304), .A2(n17303), .ZN(P1_U3161) );
  INV_X1 U20421 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20529) );
  INV_X1 U20422 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21380) );
  INV_X1 U20423 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21383) );
  NOR2_X1 U20424 ( .A1(n21380), .A2(n21383), .ZN(n21376) );
  INV_X1 U20425 ( .A(HOLD), .ZN(n21372) );
  NOR2_X1 U20426 ( .A1(n20529), .A2(n21372), .ZN(n21374) );
  OAI22_X1 U20427 ( .A1(n21376), .A2(n21374), .B1(n21388), .B2(n21372), .ZN(
        n17305) );
  OAI211_X1 U20428 ( .C1(n21487), .C2(n20529), .A(n17306), .B(n17305), .ZN(
        P1_U3195) );
  INV_X1 U20429 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17477) );
  NOR2_X1 U20430 ( .A1(n20675), .A2(n17477), .ZN(P1_U2905) );
  AND2_X1 U20431 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20498), .ZN(
        P2_U3047) );
  AOI22_X1 U20432 ( .A1(n20703), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20718), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17312) );
  NAND2_X1 U20433 ( .A1(n17309), .A2(n17308), .ZN(n17310) );
  XNOR2_X1 U20434 ( .A(n17307), .B(n17310), .ZN(n17344) );
  AOI22_X1 U20435 ( .A1(n20709), .A2(n20644), .B1(n17344), .B2(n20710), .ZN(
        n17311) );
  OAI211_X1 U20436 ( .C1(n20714), .C2(n20565), .A(n17312), .B(n17311), .ZN(
        P1_U2992) );
  AOI22_X1 U20437 ( .A1(n20703), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20718), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17316) );
  XNOR2_X1 U20438 ( .A(n12153), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17314) );
  XNOR2_X1 U20439 ( .A(n17313), .B(n17314), .ZN(n17349) );
  AOI22_X1 U20440 ( .A1(n17349), .A2(n20710), .B1(n20583), .B2(n20709), .ZN(
        n17315) );
  OAI211_X1 U20441 ( .C1(n20714), .C2(n20580), .A(n17316), .B(n17315), .ZN(
        P1_U2993) );
  AOI22_X1 U20442 ( .A1(n20703), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20718), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17322) );
  OR2_X1 U20443 ( .A1(n17318), .A2(n17317), .ZN(n17319) );
  AND2_X1 U20444 ( .A1(n17320), .A2(n17319), .ZN(n17359) );
  AOI22_X1 U20445 ( .A1(n17359), .A2(n20710), .B1(n20709), .B2(n20650), .ZN(
        n17321) );
  OAI211_X1 U20446 ( .C1(n20714), .C2(n20587), .A(n17322), .B(n17321), .ZN(
        P1_U2994) );
  OAI21_X1 U20447 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17323), .ZN(n17338) );
  AOI21_X1 U20448 ( .B1(n17325), .B2(n20742), .A(n17324), .ZN(n17337) );
  NAND2_X1 U20449 ( .A1(n17326), .A2(n20715), .ZN(n17362) );
  INV_X1 U20450 ( .A(n17362), .ZN(n17332) );
  INV_X1 U20451 ( .A(n20715), .ZN(n17327) );
  NAND2_X1 U20452 ( .A1(n20735), .A2(n17327), .ZN(n17329) );
  NAND2_X1 U20453 ( .A1(n20735), .A2(n17328), .ZN(n20721) );
  NAND2_X1 U20454 ( .A1(n17329), .A2(n20721), .ZN(n17330) );
  OR2_X1 U20455 ( .A1(n17331), .A2(n17330), .ZN(n17358) );
  AOI21_X1 U20456 ( .B1(n17333), .B2(n17332), .A(n17358), .ZN(n17351) );
  OAI21_X1 U20457 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17334), .A(
        n17351), .ZN(n17343) );
  AOI22_X1 U20458 ( .A1(n17335), .A2(n20738), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17343), .ZN(n17336) );
  OAI211_X1 U20459 ( .C1(n17347), .C2(n17338), .A(n17337), .B(n17336), .ZN(
        P1_U3023) );
  INV_X1 U20460 ( .A(n17339), .ZN(n17342) );
  INV_X1 U20461 ( .A(n17340), .ZN(n17341) );
  AOI21_X1 U20462 ( .B1(n17342), .B2(n17341), .A(n9792), .ZN(n20643) );
  AOI22_X1 U20463 ( .A1(n20643), .A2(n20742), .B1(n20718), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20464 ( .A1(n17344), .A2(n20738), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17343), .ZN(n17345) );
  OAI211_X1 U20465 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17347), .A(
        n17346), .B(n17345), .ZN(P1_U3024) );
  INV_X1 U20466 ( .A(n17348), .ZN(n17352) );
  AOI222_X1 U20467 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20718), .B1(n20742), 
        .B2(n20578), .C1(n20738), .C2(n17349), .ZN(n17350) );
  OAI221_X1 U20468 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17352), .C1(
        n12150), .C2(n17351), .A(n17350), .ZN(P1_U3025) );
  OAI21_X1 U20469 ( .B1(n17355), .B2(n17354), .A(n17353), .ZN(n17357) );
  AND2_X1 U20470 ( .A1(n17357), .A2(n17356), .ZN(n20647) );
  AOI22_X1 U20471 ( .A1(n20742), .A2(n20647), .B1(n20718), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U20472 ( .A1(n17359), .A2(n20738), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17358), .ZN(n17360) );
  OAI211_X1 U20473 ( .C1(n20733), .C2(n17362), .A(n17361), .B(n17360), .ZN(
        P1_U3026) );
  NAND4_X1 U20474 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n21306), .A4(n21487), .ZN(n17363) );
  NAND2_X1 U20475 ( .A1(n17364), .A2(n17363), .ZN(n21368) );
  OAI21_X1 U20476 ( .B1(n17366), .B2(n21368), .A(n17365), .ZN(n17367) );
  OAI221_X1 U20477 ( .B1(n17368), .B2(n21660), .C1(n17368), .C2(n21487), .A(
        n17367), .ZN(n17369) );
  AOI221_X1 U20478 ( .B1(n17371), .B2(n17370), .C1(n21369), .C2(n17370), .A(
        n17369), .ZN(P1_U3162) );
  NOR2_X1 U20479 ( .A1(n17371), .A2(n21369), .ZN(n17373) );
  OAI21_X1 U20480 ( .B1(n17373), .B2(n21660), .A(n17372), .ZN(P1_U3466) );
  AOI22_X1 U20481 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19748), .B1(n19771), 
        .B2(n17374), .ZN(n17379) );
  AOI222_X1 U20482 ( .A1(n17377), .A2(n19763), .B1(n19787), .B2(n17376), .C1(
        n19781), .C2(n17375), .ZN(n17378) );
  OAI211_X1 U20483 ( .C1(n17388), .C2(n16201), .A(n17379), .B(n17378), .ZN(
        P2_U3009) );
  AOI22_X1 U20484 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19748), .B1(n19771), 
        .B2(n17380), .ZN(n17387) );
  NAND3_X1 U20485 ( .A1(n17382), .A2(n17381), .A3(n19781), .ZN(n17383) );
  OAI21_X1 U20486 ( .B1(n19774), .B2(n10100), .A(n17383), .ZN(n17384) );
  AOI21_X1 U20487 ( .B1(n17385), .B2(n19763), .A(n17384), .ZN(n17386) );
  OAI211_X1 U20488 ( .C1(n17389), .C2(n17388), .A(n17387), .B(n17386), .ZN(
        P2_U3011) );
  INV_X1 U20489 ( .A(n19806), .ZN(n17391) );
  AOI22_X1 U20490 ( .A1(n17391), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19792), .B2(n17390), .ZN(n17405) );
  NAND2_X1 U20491 ( .A1(n17392), .A2(n17395), .ZN(n17393) );
  NAND2_X1 U20492 ( .A1(n17394), .A2(n17393), .ZN(n19784) );
  NAND2_X1 U20493 ( .A1(n17396), .A2(n17395), .ZN(n17397) );
  AND2_X1 U20494 ( .A1(n17398), .A2(n17397), .ZN(n19780) );
  NAND2_X1 U20495 ( .A1(n19796), .A2(n19780), .ZN(n17399) );
  OAI21_X1 U20496 ( .B1(n17400), .B2(n19784), .A(n17399), .ZN(n17403) );
  OR2_X1 U20497 ( .A1(n11468), .A2(n10758), .ZN(n19782) );
  OAI21_X1 U20498 ( .B1(n19803), .B2(n17401), .A(n19782), .ZN(n17402) );
  NOR2_X1 U20499 ( .A1(n17403), .A2(n17402), .ZN(n17404) );
  OAI211_X1 U20500 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17406), .A(
        n17405), .B(n17404), .ZN(P2_U3046) );
  NOR3_X1 U20501 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17408) );
  NOR4_X1 U20502 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17407) );
  NAND4_X1 U20503 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17408), .A3(n17407), .A4(
        U215), .ZN(U213) );
  INV_X1 U20504 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19715) );
  INV_X2 U20505 ( .A(U214), .ZN(n17445) );
  OAI222_X1 U20506 ( .A1(U212), .A2(n19715), .B1(n17442), .B2(n21659), .C1(
        U214), .C2(n17477), .ZN(U216) );
  AOI22_X1 U20507 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17443), .ZN(n17410) );
  OAI21_X1 U20508 ( .B1(n14929), .B2(n17442), .A(n17410), .ZN(U217) );
  AOI222_X1 U20509 ( .A1(n17443), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n17444), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n17445), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n17411) );
  INV_X1 U20510 ( .A(n17411), .ZN(U218) );
  AOI22_X1 U20511 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17443), .ZN(n17412) );
  OAI21_X1 U20512 ( .B1(n16372), .B2(n17442), .A(n17412), .ZN(U219) );
  AOI22_X1 U20513 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17443), .ZN(n17413) );
  OAI21_X1 U20514 ( .B1(n16380), .B2(n17442), .A(n17413), .ZN(U220) );
  AOI22_X1 U20515 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17443), .ZN(n17414) );
  OAI21_X1 U20516 ( .B1(n16388), .B2(n17442), .A(n17414), .ZN(U221) );
  INV_X1 U20517 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n21594) );
  INV_X1 U20518 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17415) );
  INV_X1 U20519 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n21587) );
  OAI222_X1 U20520 ( .A1(U214), .A2(n21594), .B1(n17442), .B2(n17415), .C1(
        U212), .C2(n21587), .ZN(U222) );
  AOI22_X1 U20521 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17443), .ZN(n17416) );
  OAI21_X1 U20522 ( .B1(n21666), .B2(n17442), .A(n17416), .ZN(U223) );
  INV_X1 U20523 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U20524 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17443), .ZN(n17417) );
  OAI21_X1 U20525 ( .B1(n19852), .B2(n17442), .A(n17417), .ZN(U224) );
  AOI22_X1 U20526 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17443), .ZN(n17418) );
  OAI21_X1 U20527 ( .B1(n17419), .B2(n17442), .A(n17418), .ZN(U225) );
  INV_X1 U20528 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19836) );
  AOI22_X1 U20529 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17443), .ZN(n17420) );
  OAI21_X1 U20530 ( .B1(n19836), .B2(n17442), .A(n17420), .ZN(U226) );
  INV_X1 U20531 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U20532 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17443), .ZN(n17421) );
  OAI21_X1 U20533 ( .B1(n19831), .B2(n17442), .A(n17421), .ZN(U227) );
  INV_X1 U20534 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U20535 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17443), .ZN(n17422) );
  OAI21_X1 U20536 ( .B1(n19826), .B2(n17442), .A(n17422), .ZN(U228) );
  INV_X1 U20537 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n17463) );
  INV_X1 U20538 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n21744) );
  OAI222_X1 U20539 ( .A1(U212), .A2(n17463), .B1(n17442), .B2(n21597), .C1(
        U214), .C2(n21744), .ZN(U229) );
  INV_X1 U20540 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U20541 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17443), .ZN(n17423) );
  OAI21_X1 U20542 ( .B1(n19821), .B2(n17442), .A(n17423), .ZN(U230) );
  INV_X1 U20543 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n19816) );
  AOI22_X1 U20544 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17443), .ZN(n17424) );
  OAI21_X1 U20545 ( .B1(n19816), .B2(n17433), .A(n17424), .ZN(U231) );
  AOI22_X1 U20546 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17443), .ZN(n17425) );
  OAI21_X1 U20547 ( .B1(n14292), .B2(n17433), .A(n17425), .ZN(U232) );
  AOI22_X1 U20548 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17443), .ZN(n17426) );
  OAI21_X1 U20549 ( .B1(n13963), .B2(n17442), .A(n17426), .ZN(U233) );
  AOI22_X1 U20550 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17443), .ZN(n17427) );
  OAI21_X1 U20551 ( .B1(n13982), .B2(n17442), .A(n17427), .ZN(U234) );
  AOI22_X1 U20552 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17443), .ZN(n17428) );
  OAI21_X1 U20553 ( .B1(n13976), .B2(n17433), .A(n17428), .ZN(U235) );
  AOI22_X1 U20554 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17443), .ZN(n17429) );
  OAI21_X1 U20555 ( .B1(n13988), .B2(n17442), .A(n17429), .ZN(U236) );
  INV_X1 U20556 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17455) );
  INV_X1 U20557 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n21586) );
  OAI222_X1 U20558 ( .A1(U212), .A2(n17455), .B1(n17442), .B2(n17430), .C1(
        U214), .C2(n21586), .ZN(U237) );
  AOI22_X1 U20559 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17443), .ZN(n17431) );
  OAI21_X1 U20560 ( .B1(n13959), .B2(n17442), .A(n17431), .ZN(U238) );
  AOI22_X1 U20561 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17443), .ZN(n17432) );
  OAI21_X1 U20562 ( .B1(n21711), .B2(n17433), .A(n17432), .ZN(U239) );
  INV_X1 U20563 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n21577) );
  AOI22_X1 U20564 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17444), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17445), .ZN(n17434) );
  OAI21_X1 U20565 ( .B1(n21577), .B2(U212), .A(n17434), .ZN(U240) );
  INV_X1 U20566 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20567 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n17444), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17445), .ZN(n17435) );
  OAI21_X1 U20568 ( .B1(n17452), .B2(U212), .A(n17435), .ZN(U241) );
  INV_X1 U20569 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n21754) );
  AOI22_X1 U20570 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17444), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17443), .ZN(n17436) );
  OAI21_X1 U20571 ( .B1(n21754), .B2(U214), .A(n17436), .ZN(U242) );
  AOI22_X1 U20572 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17443), .ZN(n17437) );
  OAI21_X1 U20573 ( .B1(n13944), .B2(n17442), .A(n17437), .ZN(U243) );
  INV_X1 U20574 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U20575 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17444), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17445), .ZN(n17438) );
  OAI21_X1 U20576 ( .B1(n17449), .B2(U212), .A(n17438), .ZN(U244) );
  AOI22_X1 U20577 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17443), .ZN(n17439) );
  OAI21_X1 U20578 ( .B1(n17440), .B2(n17442), .A(n17439), .ZN(U245) );
  INV_X1 U20579 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n21663) );
  AOI22_X1 U20580 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17445), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17443), .ZN(n17441) );
  OAI21_X1 U20581 ( .B1(n21663), .B2(n17442), .A(n17441), .ZN(U246) );
  AOI222_X1 U20582 ( .A1(n17445), .A2(P1_DATAO_REG_0__SCAN_IN), .B1(n17444), 
        .B2(BUF1_REG_0__SCAN_IN), .C1(n17443), .C2(P2_DATAO_REG_0__SCAN_IN), 
        .ZN(n17446) );
  INV_X1 U20583 ( .A(n17446), .ZN(U247) );
  INV_X1 U20584 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n21641) );
  AOI22_X1 U20585 ( .A1(n17471), .A2(n21641), .B1(n19029), .B2(U215), .ZN(U251) );
  OAI22_X1 U20586 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17471), .ZN(n17447) );
  INV_X1 U20587 ( .A(n17447), .ZN(U252) );
  INV_X1 U20588 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20589 ( .A1(n17471), .A2(n17448), .B1(n19041), .B2(U215), .ZN(U253) );
  INV_X1 U20590 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19045) );
  AOI22_X1 U20591 ( .A1(n17471), .A2(n17449), .B1(n19045), .B2(U215), .ZN(U254) );
  INV_X1 U20592 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17450) );
  INV_X1 U20593 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19050) );
  AOI22_X1 U20594 ( .A1(n17471), .A2(n17450), .B1(n19050), .B2(U215), .ZN(U255) );
  INV_X1 U20595 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17451) );
  INV_X1 U20596 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19054) );
  AOI22_X1 U20597 ( .A1(n17471), .A2(n17451), .B1(n19054), .B2(U215), .ZN(U256) );
  INV_X1 U20598 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21656) );
  AOI22_X1 U20599 ( .A1(n17471), .A2(n17452), .B1(n21656), .B2(U215), .ZN(U257) );
  AOI22_X1 U20600 ( .A1(n17471), .A2(n21577), .B1(n19062), .B2(U215), .ZN(U258) );
  INV_X1 U20601 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17453) );
  INV_X1 U20602 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U20603 ( .A1(n17471), .A2(n17453), .B1(n18517), .B2(U215), .ZN(U259) );
  INV_X1 U20604 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17454) );
  INV_X1 U20605 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18519) );
  AOI22_X1 U20606 ( .A1(n17471), .A2(n17454), .B1(n18519), .B2(U215), .ZN(U260) );
  INV_X1 U20607 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18521) );
  AOI22_X1 U20608 ( .A1(n17471), .A2(n17455), .B1(n18521), .B2(U215), .ZN(U261) );
  OAI22_X1 U20609 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17471), .ZN(n17456) );
  INV_X1 U20610 ( .A(n17456), .ZN(U262) );
  INV_X1 U20611 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17457) );
  INV_X1 U20612 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18525) );
  AOI22_X1 U20613 ( .A1(n17471), .A2(n17457), .B1(n18525), .B2(U215), .ZN(U263) );
  INV_X1 U20614 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17458) );
  INV_X1 U20615 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18529) );
  AOI22_X1 U20616 ( .A1(n17471), .A2(n17458), .B1(n18529), .B2(U215), .ZN(U264) );
  OAI22_X1 U20617 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17471), .ZN(n17459) );
  INV_X1 U20618 ( .A(n17459), .ZN(U265) );
  OAI22_X1 U20619 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17471), .ZN(n17460) );
  INV_X1 U20620 ( .A(n17460), .ZN(U266) );
  INV_X1 U20621 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n17461) );
  INV_X1 U20622 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U20623 ( .A1(n17471), .A2(n17461), .B1(n19815), .B2(U215), .ZN(U267) );
  INV_X1 U20624 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20625 ( .A1(n17471), .A2(n17462), .B1(n16454), .B2(U215), .ZN(U268) );
  AOI22_X1 U20626 ( .A1(n17471), .A2(n17463), .B1(n19040), .B2(U215), .ZN(U269) );
  INV_X1 U20627 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U20628 ( .A1(n17471), .A2(n17464), .B1(n16440), .B2(U215), .ZN(U270) );
  INV_X1 U20629 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n17465) );
  AOI22_X1 U20630 ( .A1(n17471), .A2(n17465), .B1(n16434), .B2(U215), .ZN(U271) );
  INV_X1 U20631 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U20632 ( .A1(n17471), .A2(n17466), .B1(n16425), .B2(U215), .ZN(U272) );
  OAI22_X1 U20633 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17471), .ZN(n17467) );
  INV_X1 U20634 ( .A(n17467), .ZN(U273) );
  INV_X1 U20635 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20636 ( .A1(n17471), .A2(n17468), .B1(n16410), .B2(U215), .ZN(U274) );
  OAI22_X1 U20637 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17471), .ZN(n17469) );
  INV_X1 U20638 ( .A(n17469), .ZN(U275) );
  OAI22_X1 U20639 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17471), .ZN(n17470) );
  INV_X1 U20640 ( .A(n17470), .ZN(U276) );
  OAI22_X1 U20641 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17471), .ZN(n17472) );
  INV_X1 U20642 ( .A(n17472), .ZN(U277) );
  INV_X1 U20643 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n17473) );
  INV_X1 U20644 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21578) );
  AOI22_X1 U20645 ( .A1(n17471), .A2(n17473), .B1(n21578), .B2(U215), .ZN(U278) );
  INV_X1 U20646 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17474) );
  AOI22_X1 U20647 ( .A1(n17471), .A2(n17474), .B1(n19049), .B2(U215), .ZN(U279) );
  OAI22_X1 U20648 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17471), .ZN(n17475) );
  INV_X1 U20649 ( .A(n17475), .ZN(U280) );
  INV_X1 U20650 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17476) );
  INV_X1 U20651 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n21630) );
  AOI22_X1 U20652 ( .A1(n17471), .A2(n17476), .B1(n21630), .B2(U215), .ZN(U281) );
  INV_X1 U20653 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19061) );
  AOI22_X1 U20654 ( .A1(n17471), .A2(n19715), .B1(n19061), .B2(U215), .ZN(U282) );
  AOI222_X1 U20655 ( .A1(n17477), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19715), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n18427), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17478) );
  INV_X2 U20656 ( .A(n17480), .ZN(n17479) );
  INV_X1 U20657 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19554) );
  INV_X1 U20658 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20427) );
  AOI22_X1 U20659 ( .A1(n17479), .A2(n19554), .B1(n20427), .B2(n17480), .ZN(
        U347) );
  INV_X1 U20660 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19552) );
  INV_X1 U20661 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20425) );
  AOI22_X1 U20662 ( .A1(n17478), .A2(n19552), .B1(n20425), .B2(n17480), .ZN(
        U348) );
  INV_X1 U20663 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19550) );
  INV_X1 U20664 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20423) );
  AOI22_X1 U20665 ( .A1(n17479), .A2(n19550), .B1(n20423), .B2(n17480), .ZN(
        U349) );
  INV_X1 U20666 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19549) );
  INV_X1 U20667 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20422) );
  AOI22_X1 U20668 ( .A1(n17479), .A2(n19549), .B1(n20422), .B2(n17480), .ZN(
        U350) );
  INV_X1 U20669 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19547) );
  INV_X1 U20670 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U20671 ( .A1(n17479), .A2(n19547), .B1(n20421), .B2(n17480), .ZN(
        U351) );
  INV_X1 U20672 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19545) );
  INV_X1 U20673 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20419) );
  AOI22_X1 U20674 ( .A1(n17479), .A2(n19545), .B1(n20419), .B2(n17480), .ZN(
        U352) );
  INV_X1 U20675 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19544) );
  INV_X1 U20676 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U20677 ( .A1(n17479), .A2(n19544), .B1(n20418), .B2(n17480), .ZN(
        U353) );
  INV_X1 U20678 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19542) );
  INV_X1 U20679 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20416) );
  AOI22_X1 U20680 ( .A1(n17479), .A2(n19542), .B1(n20416), .B2(n17480), .ZN(
        U354) );
  INV_X1 U20681 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19592) );
  INV_X1 U20682 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20463) );
  AOI22_X1 U20683 ( .A1(n17479), .A2(n19592), .B1(n20463), .B2(n17480), .ZN(
        U355) );
  INV_X1 U20684 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19589) );
  INV_X1 U20685 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20460) );
  AOI22_X1 U20686 ( .A1(n17479), .A2(n19589), .B1(n20460), .B2(n17480), .ZN(
        U356) );
  INV_X1 U20687 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19586) );
  INV_X1 U20688 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20457) );
  AOI22_X1 U20689 ( .A1(n17479), .A2(n19586), .B1(n20457), .B2(n17480), .ZN(
        U357) );
  INV_X1 U20690 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n21710) );
  INV_X1 U20691 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20454) );
  AOI22_X1 U20692 ( .A1(n17479), .A2(n21710), .B1(n20454), .B2(n17480), .ZN(
        U358) );
  INV_X1 U20693 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19584) );
  INV_X1 U20694 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20453) );
  AOI22_X1 U20695 ( .A1(n17479), .A2(n19584), .B1(n20453), .B2(n17480), .ZN(
        U359) );
  INV_X1 U20696 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19582) );
  INV_X1 U20697 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21738) );
  AOI22_X1 U20698 ( .A1(n17479), .A2(n19582), .B1(n21738), .B2(n17480), .ZN(
        U360) );
  INV_X1 U20699 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19581) );
  INV_X1 U20700 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20450) );
  AOI22_X1 U20701 ( .A1(n17479), .A2(n19581), .B1(n20450), .B2(n17480), .ZN(
        U361) );
  INV_X1 U20702 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19578) );
  INV_X1 U20703 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20449) );
  AOI22_X1 U20704 ( .A1(n17479), .A2(n19578), .B1(n20449), .B2(n17480), .ZN(
        U362) );
  INV_X1 U20705 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19577) );
  INV_X1 U20706 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20447) );
  AOI22_X1 U20707 ( .A1(n17479), .A2(n19577), .B1(n20447), .B2(n17480), .ZN(
        U363) );
  INV_X1 U20708 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19574) );
  INV_X1 U20709 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20445) );
  AOI22_X1 U20710 ( .A1(n17479), .A2(n19574), .B1(n20445), .B2(n17480), .ZN(
        U364) );
  INV_X1 U20711 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19540) );
  INV_X1 U20712 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20415) );
  AOI22_X1 U20713 ( .A1(n17479), .A2(n19540), .B1(n20415), .B2(n17480), .ZN(
        U365) );
  INV_X1 U20714 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19573) );
  INV_X1 U20715 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20443) );
  AOI22_X1 U20716 ( .A1(n17479), .A2(n19573), .B1(n20443), .B2(n17480), .ZN(
        U366) );
  INV_X1 U20717 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19572) );
  INV_X1 U20718 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21600) );
  AOI22_X1 U20719 ( .A1(n17479), .A2(n19572), .B1(n21600), .B2(n17480), .ZN(
        U367) );
  INV_X1 U20720 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19570) );
  INV_X1 U20721 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20441) );
  AOI22_X1 U20722 ( .A1(n17479), .A2(n19570), .B1(n20441), .B2(n17480), .ZN(
        U368) );
  INV_X1 U20723 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19568) );
  INV_X1 U20724 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20440) );
  AOI22_X1 U20725 ( .A1(n17479), .A2(n19568), .B1(n20440), .B2(n17480), .ZN(
        U369) );
  INV_X1 U20726 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19565) );
  INV_X1 U20727 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20438) );
  AOI22_X1 U20728 ( .A1(n17479), .A2(n19565), .B1(n20438), .B2(n17480), .ZN(
        U370) );
  INV_X1 U20729 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19564) );
  INV_X1 U20730 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20436) );
  AOI22_X1 U20731 ( .A1(n17478), .A2(n19564), .B1(n20436), .B2(n17480), .ZN(
        U371) );
  INV_X1 U20732 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19561) );
  INV_X1 U20733 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20434) );
  AOI22_X1 U20734 ( .A1(n17478), .A2(n19561), .B1(n20434), .B2(n17480), .ZN(
        U372) );
  INV_X1 U20735 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19560) );
  INV_X1 U20736 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20432) );
  AOI22_X1 U20737 ( .A1(n17479), .A2(n19560), .B1(n20432), .B2(n17480), .ZN(
        U373) );
  INV_X1 U20738 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19557) );
  INV_X1 U20739 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20431) );
  AOI22_X1 U20740 ( .A1(n17479), .A2(n19557), .B1(n20431), .B2(n17480), .ZN(
        U374) );
  INV_X1 U20741 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19556) );
  INV_X1 U20742 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20429) );
  AOI22_X1 U20743 ( .A1(n17478), .A2(n19556), .B1(n20429), .B2(n17480), .ZN(
        U375) );
  INV_X1 U20744 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19538) );
  INV_X1 U20745 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20413) );
  AOI22_X1 U20746 ( .A1(n17479), .A2(n19538), .B1(n20413), .B2(n17480), .ZN(
        U376) );
  INV_X1 U20747 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17482) );
  NAND2_X1 U20748 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19537), .ZN(n19527) );
  NAND2_X1 U20749 ( .A1(n17483), .A2(n17481), .ZN(n19523) );
  INV_X1 U20750 ( .A(n19605), .ZN(n19602) );
  OAI21_X1 U20751 ( .B1(n17483), .B2(n17482), .A(n19602), .ZN(P3_U2633) );
  AND2_X1 U20752 ( .A1(n19509), .A2(n19473), .ZN(n17484) );
  INV_X1 U20753 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n17485) );
  NAND2_X1 U20754 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19639), .ZN(n19517) );
  OAI21_X1 U20755 ( .B1(n17484), .B2(n17485), .A(n19517), .ZN(P3_U2634) );
  AOI22_X1 U20756 ( .A1(n19635), .A2(n17485), .B1(P3_D_C_N_REG_SCAN_IN), .B2(
        n19616), .ZN(n17486) );
  OAI21_X1 U20757 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n19522), .A(n17486), 
        .ZN(P3_U2635) );
  INV_X1 U20758 ( .A(n19522), .ZN(n17487) );
  OAI21_X1 U20759 ( .B1(n17487), .B2(BS16), .A(n19605), .ZN(n19603) );
  OAI21_X1 U20760 ( .B1(n19605), .B2(n19625), .A(n19603), .ZN(P3_U2636) );
  AOI21_X1 U20761 ( .B1(n19473), .B2(n19472), .A(n19518), .ZN(n19618) );
  OAI21_X1 U20762 ( .B1(n19618), .B2(n19021), .A(n17488), .ZN(P3_U2637) );
  NOR4_X1 U20763 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17492) );
  NOR4_X1 U20764 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17491) );
  NOR4_X1 U20765 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17490) );
  NOR4_X1 U20766 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17489) );
  NAND4_X1 U20767 ( .A1(n17492), .A2(n17491), .A3(n17490), .A4(n17489), .ZN(
        n17498) );
  NOR4_X1 U20768 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_31__SCAN_IN), .A3(P3_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n17496) );
  AOI211_X1 U20769 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_15__SCAN_IN), .B(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n17495) );
  NOR4_X1 U20770 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17494) );
  NOR4_X1 U20771 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17493) );
  NAND4_X1 U20772 ( .A1(n17496), .A2(n17495), .A3(n17494), .A4(n17493), .ZN(
        n17497) );
  NOR2_X1 U20773 ( .A1(n17498), .A2(n17497), .ZN(n19615) );
  INV_X1 U20774 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19598) );
  NOR3_X1 U20775 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17500) );
  OAI21_X1 U20776 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17500), .A(n19615), .ZN(
        n17499) );
  OAI21_X1 U20777 ( .B1(n19615), .B2(n19598), .A(n17499), .ZN(P3_U2638) );
  INV_X1 U20778 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19609) );
  INV_X1 U20779 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19604) );
  AOI21_X1 U20780 ( .B1(n19609), .B2(n19604), .A(n17500), .ZN(n17501) );
  INV_X1 U20781 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19595) );
  INV_X1 U20782 ( .A(n19615), .ZN(n19611) );
  AOI22_X1 U20783 ( .A1(n19615), .A2(n17501), .B1(n19595), .B2(n19611), .ZN(
        P3_U2639) );
  NAND2_X1 U20784 ( .A1(n17829), .A2(n17502), .ZN(n17519) );
  OAI22_X1 U20785 ( .A1(n17523), .A2(n21720), .B1(n17505), .B2(n17852), .ZN(
        n17506) );
  INV_X1 U20786 ( .A(n17506), .ZN(n17507) );
  OAI21_X1 U20787 ( .B1(n17804), .B2(n17508), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17509) );
  OAI211_X1 U20788 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17519), .A(n17510), .B(
        n17509), .ZN(P3_U2641) );
  INV_X1 U20789 ( .A(n17512), .ZN(n17513) );
  AOI211_X1 U20790 ( .C1(n17515), .C2(n17514), .A(n17513), .B(n17823), .ZN(
        n17517) );
  OAI22_X1 U20791 ( .A1(n10088), .A2(n17852), .B1(n17865), .B2(n17875), .ZN(
        n17516) );
  AOI211_X1 U20792 ( .C1(n17518), .C2(n19588), .A(n17517), .B(n17516), .ZN(
        n17522) );
  INV_X1 U20793 ( .A(n17519), .ZN(n17520) );
  OAI21_X1 U20794 ( .B1(n17525), .B2(n17875), .A(n17520), .ZN(n17521) );
  OAI211_X1 U20795 ( .C1(n17523), .C2(n19588), .A(n17522), .B(n17521), .ZN(
        P3_U2642) );
  OAI21_X1 U20796 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n17524), .ZN(n17535) );
  AOI22_X1 U20797 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17844), .B1(
        n17804), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17534) );
  AOI211_X1 U20798 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17542), .A(n17525), .B(
        n17864), .ZN(n17532) );
  INV_X1 U20799 ( .A(n17526), .ZN(n17529) );
  INV_X1 U20800 ( .A(n17527), .ZN(n17528) );
  AOI211_X1 U20801 ( .C1(n17530), .C2(n17529), .A(n17528), .B(n17823), .ZN(
        n17531) );
  OAI211_X1 U20802 ( .C1(n17539), .C2(n17535), .A(n17534), .B(n17533), .ZN(
        P3_U2643) );
  INV_X1 U20803 ( .A(n17553), .ZN(n17546) );
  INV_X1 U20804 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19585) );
  AOI211_X1 U20805 ( .C1(n17538), .C2(n17537), .A(n17536), .B(n17823), .ZN(
        n17541) );
  OAI22_X1 U20806 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17539), .B1(n17543), 
        .B2(n17865), .ZN(n17540) );
  AOI211_X1 U20807 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17541), .B(n17540), .ZN(n17545) );
  OAI211_X1 U20808 ( .C1(n17547), .C2(n17543), .A(n17829), .B(n17542), .ZN(
        n17544) );
  OAI211_X1 U20809 ( .C1(n17546), .C2(n19585), .A(n17545), .B(n17544), .ZN(
        P3_U2644) );
  AOI22_X1 U20810 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17844), .B1(
        n17804), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17555) );
  AOI211_X1 U20811 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17563), .A(n17547), .B(
        n17864), .ZN(n17552) );
  AOI211_X1 U20812 ( .C1(n17550), .C2(n17549), .A(n17548), .B(n17823), .ZN(
        n17551) );
  AOI211_X1 U20813 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17553), .A(n17552), 
        .B(n17551), .ZN(n17554) );
  OAI211_X1 U20814 ( .C1(n17557), .C2(n17556), .A(n17555), .B(n17554), .ZN(
        P3_U2645) );
  AOI22_X1 U20815 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17844), .B1(
        n17804), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n17568) );
  INV_X1 U20816 ( .A(n17558), .ZN(n17570) );
  OAI21_X1 U20817 ( .B1(n17570), .B2(n17857), .A(n17868), .ZN(n17579) );
  NOR2_X1 U20818 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17857), .ZN(n17569) );
  AOI211_X1 U20819 ( .C1(n17561), .C2(n17560), .A(n17559), .B(n17823), .ZN(
        n17562) );
  AOI221_X1 U20820 ( .B1(n17579), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n17569), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n17562), .ZN(n17567) );
  OAI211_X1 U20821 ( .C1(n17571), .C2(n17874), .A(n17829), .B(n17563), .ZN(
        n17566) );
  INV_X1 U20822 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21627) );
  NAND3_X1 U20823 ( .A1(n17846), .A2(n17564), .A3(n21627), .ZN(n17565) );
  NAND4_X1 U20824 ( .A1(n17568), .A2(n17567), .A3(n17566), .A4(n17565), .ZN(
        P3_U2646) );
  AOI22_X1 U20825 ( .A1(n17804), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17570), 
        .B2(n17569), .ZN(n17577) );
  AOI211_X1 U20826 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17585), .A(n17571), .B(
        n17864), .ZN(n17575) );
  AOI211_X1 U20827 ( .C1(n18555), .C2(n17573), .A(n17572), .B(n17823), .ZN(
        n17574) );
  AOI211_X1 U20828 ( .C1(n17579), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17575), 
        .B(n17574), .ZN(n17576) );
  OAI211_X1 U20829 ( .C1(n18557), .C2(n17852), .A(n17577), .B(n17576), .ZN(
        P3_U2647) );
  AOI21_X1 U20830 ( .B1(n17846), .B2(n17578), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n17590) );
  INV_X1 U20831 ( .A(n17579), .ZN(n17589) );
  AOI211_X1 U20832 ( .C1(n17582), .C2(n17581), .A(n17580), .B(n17823), .ZN(
        n17584) );
  NOR2_X1 U20833 ( .A1(n17865), .A2(n17586), .ZN(n17583) );
  AOI211_X1 U20834 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17584), .B(n17583), .ZN(n17588) );
  OAI211_X1 U20835 ( .C1(n17593), .C2(n17586), .A(n17829), .B(n17585), .ZN(
        n17587) );
  OAI211_X1 U20836 ( .C1(n17590), .C2(n17589), .A(n17588), .B(n17587), .ZN(
        P3_U2648) );
  INV_X1 U20837 ( .A(n17592), .ZN(n17591) );
  AOI21_X1 U20838 ( .B1(n17846), .B2(n17591), .A(n17851), .ZN(n17624) );
  INV_X1 U20839 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19575) );
  NAND3_X1 U20840 ( .A1(n17846), .A2(n17592), .A3(n19575), .ZN(n17608) );
  AOI211_X1 U20841 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17611), .A(n17593), .B(
        n17864), .ZN(n17602) );
  INV_X1 U20842 ( .A(n17594), .ZN(n17595) );
  AOI211_X1 U20843 ( .C1(n18589), .C2(n17595), .A(n9805), .B(n17823), .ZN(
        n17601) );
  NOR3_X1 U20844 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17857), .A3(n17596), 
        .ZN(n17600) );
  OAI22_X1 U20845 ( .A1(n17598), .A2(n17852), .B1(n17865), .B2(n17597), .ZN(
        n17599) );
  NOR4_X1 U20846 ( .A1(n17602), .A2(n17601), .A3(n17600), .A4(n17599), .ZN(
        n17603) );
  OAI221_X1 U20847 ( .B1(n19576), .B2(n17624), .C1(n19576), .C2(n17608), .A(
        n17603), .ZN(P3_U2649) );
  INV_X1 U20848 ( .A(n17604), .ZN(n17605) );
  AOI211_X1 U20849 ( .C1(n17607), .C2(n17606), .A(n17605), .B(n17823), .ZN(
        n17610) );
  OAI21_X1 U20850 ( .B1(n17979), .B2(n17865), .A(n17608), .ZN(n17609) );
  AOI211_X1 U20851 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17610), .B(n17609), .ZN(n17613) );
  OAI211_X1 U20852 ( .C1(n17617), .C2(n17979), .A(n17829), .B(n17611), .ZN(
        n17612) );
  OAI211_X1 U20853 ( .C1(n17624), .C2(n19575), .A(n17613), .B(n17612), .ZN(
        P3_U2650) );
  INV_X1 U20854 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19567) );
  INV_X1 U20855 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19566) );
  INV_X1 U20856 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19563) );
  NAND2_X1 U20857 ( .A1(n17846), .A2(n17614), .ZN(n17701) );
  INV_X1 U20858 ( .A(n17701), .ZN(n17685) );
  NAND3_X1 U20859 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17685), .ZN(n17682) );
  NOR4_X1 U20860 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n19567), .A3(n17636), 
        .A4(n17660), .ZN(n17622) );
  AOI211_X1 U20861 ( .C1(n18621), .C2(n17616), .A(n17615), .B(n17823), .ZN(
        n17621) );
  AOI211_X1 U20862 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17631), .A(n17617), .B(
        n17864), .ZN(n17620) );
  OAI22_X1 U20863 ( .A1(n17618), .A2(n17852), .B1(n17865), .B2(n17997), .ZN(
        n17619) );
  NOR4_X1 U20864 ( .A1(n17622), .A2(n17621), .A3(n17620), .A4(n17619), .ZN(
        n17623) );
  OAI21_X1 U20865 ( .B1(n21741), .B2(n17624), .A(n17623), .ZN(P3_U2651) );
  OR2_X1 U20866 ( .A1(n17851), .A2(n17625), .ZN(n17684) );
  NAND2_X1 U20867 ( .A1(n17857), .A2(n17868), .ZN(n17866) );
  OAI21_X1 U20868 ( .B1(n17626), .B2(n17684), .A(n17866), .ZN(n17659) );
  INV_X1 U20869 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19571) );
  OAI21_X1 U20870 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17628), .A(
        n17627), .ZN(n18632) );
  OAI21_X1 U20871 ( .B1(n17629), .B2(n17666), .A(n11593), .ZN(n17642) );
  OAI21_X1 U20872 ( .B1(n18632), .B2(n17642), .A(n17837), .ZN(n17630) );
  AOI21_X1 U20873 ( .B1(n18632), .B2(n17642), .A(n17630), .ZN(n17635) );
  OAI211_X1 U20874 ( .C1(n17639), .C2(n17633), .A(n17829), .B(n17631), .ZN(
        n17632) );
  OAI211_X1 U20875 ( .C1(n17865), .C2(n17633), .A(n10420), .B(n17632), .ZN(
        n17634) );
  AOI211_X1 U20876 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17635), .B(n17634), .ZN(n17638) );
  NOR2_X1 U20877 ( .A1(n19567), .A2(n17660), .ZN(n17645) );
  OAI211_X1 U20878 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n17645), .B(n17636), .ZN(n17637) );
  OAI211_X1 U20879 ( .C1(n17659), .C2(n19571), .A(n17638), .B(n17637), .ZN(
        P3_U2652) );
  AOI211_X1 U20880 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17654), .A(n17639), .B(
        n17864), .ZN(n17640) );
  AOI211_X1 U20881 ( .C1(n17804), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9696), .B(
        n17640), .ZN(n17648) );
  INV_X1 U20882 ( .A(n17659), .ZN(n17646) );
  NAND2_X1 U20883 ( .A1(n17837), .A2(n17820), .ZN(n17856) );
  OAI221_X1 U20884 ( .B1(n17643), .B2(n17667), .C1(n17643), .C2(n17649), .A(
        n17837), .ZN(n17641) );
  AOI22_X1 U20885 ( .A1(n17643), .A2(n17642), .B1(n17856), .B2(n17641), .ZN(
        n17644) );
  AOI221_X1 U20886 ( .B1(n17646), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n17645), 
        .C2(n19569), .A(n17644), .ZN(n17647) );
  OAI211_X1 U20887 ( .C1(n17649), .C2(n17852), .A(n17648), .B(n17647), .ZN(
        P3_U2653) );
  OAI21_X1 U20888 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17672), .A(
        n17650), .ZN(n18655) );
  AOI21_X1 U20889 ( .B1(n17667), .B2(n18655), .A(n17820), .ZN(n17652) );
  OAI21_X1 U20890 ( .B1(n17653), .B2(n17652), .A(n17837), .ZN(n17651) );
  AOI21_X1 U20891 ( .B1(n17653), .B2(n17652), .A(n17651), .ZN(n17657) );
  OAI211_X1 U20892 ( .C1(n17661), .C2(n18050), .A(n17829), .B(n17654), .ZN(
        n17655) );
  OAI211_X1 U20893 ( .C1(n17865), .C2(n18050), .A(n10420), .B(n17655), .ZN(
        n17656) );
  AOI211_X1 U20894 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n17657), .B(n17656), .ZN(n17658) );
  OAI221_X1 U20895 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n17660), .C1(n19567), 
        .C2(n17659), .A(n17658), .ZN(P3_U2654) );
  NAND2_X1 U20896 ( .A1(n17866), .A2(n17684), .ZN(n17696) );
  AOI221_X1 U20897 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n19566), .C2(n19563), .A(n17682), .ZN(n17665) );
  AOI211_X1 U20898 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17676), .A(n17661), .B(
        n17864), .ZN(n17664) );
  INV_X1 U20899 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17662) );
  INV_X1 U20900 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n18071) );
  OAI22_X1 U20901 ( .A1(n17662), .A2(n17852), .B1(n17865), .B2(n18071), .ZN(
        n17663) );
  NOR4_X1 U20902 ( .A1(n9696), .A2(n17665), .A3(n17664), .A4(n17663), .ZN(
        n17671) );
  NAND2_X1 U20903 ( .A1(n11593), .A2(n17666), .ZN(n17669) );
  OAI21_X1 U20904 ( .B1(n17667), .B2(n17820), .A(n18655), .ZN(n17668) );
  OAI211_X1 U20905 ( .C1(n18655), .C2(n17669), .A(n17837), .B(n17668), .ZN(
        n17670) );
  OAI211_X1 U20906 ( .C1(n19566), .C2(n17696), .A(n17671), .B(n17670), .ZN(
        P3_U2655) );
  AOI21_X1 U20907 ( .B1(n18664), .B2(n17690), .A(n17672), .ZN(n17673) );
  INV_X1 U20908 ( .A(n17673), .ZN(n18661) );
  OAI21_X1 U20909 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17690), .A(
        n11593), .ZN(n17675) );
  OAI21_X1 U20910 ( .B1(n18661), .B2(n17675), .A(n17837), .ZN(n17674) );
  AOI21_X1 U20911 ( .B1(n18661), .B2(n17675), .A(n17674), .ZN(n17680) );
  OAI211_X1 U20912 ( .C1(n17683), .C2(n17678), .A(n17829), .B(n17676), .ZN(
        n17677) );
  OAI211_X1 U20913 ( .C1(n17865), .C2(n17678), .A(n10420), .B(n17677), .ZN(
        n17679) );
  AOI211_X1 U20914 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17680), .B(n17679), .ZN(n17681) );
  OAI221_X1 U20915 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17682), .C1(n19563), 
        .C2(n17696), .A(n17681), .ZN(P3_U2656) );
  INV_X1 U20916 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19562) );
  AOI211_X1 U20917 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17705), .A(n17683), .B(
        n17864), .ZN(n17688) );
  INV_X1 U20918 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18112) );
  NAND3_X1 U20919 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17685), .A3(n17684), 
        .ZN(n17686) );
  OAI211_X1 U20920 ( .C1(n17865), .C2(n18112), .A(n10420), .B(n17686), .ZN(
        n17687) );
  AOI211_X1 U20921 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17688), .B(n17687), .ZN(n17695) );
  NAND2_X1 U20922 ( .A1(n10099), .A2(n17782), .ZN(n18693) );
  INV_X1 U20923 ( .A(n18693), .ZN(n17698) );
  NAND2_X1 U20924 ( .A1(n18689), .A2(n17698), .ZN(n17697) );
  INV_X1 U20925 ( .A(n17697), .ZN(n17691) );
  OAI21_X1 U20926 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17691), .A(
        n17690), .ZN(n18682) );
  OAI21_X1 U20927 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17697), .A(
        n11593), .ZN(n17693) );
  AOI21_X1 U20928 ( .B1(n18682), .B2(n17693), .A(n17823), .ZN(n17692) );
  OAI21_X1 U20929 ( .B1(n18682), .B2(n17693), .A(n17692), .ZN(n17694) );
  OAI211_X1 U20930 ( .C1(n17696), .C2(n19562), .A(n17695), .B(n17694), .ZN(
        P3_U2657) );
  NOR2_X1 U20931 ( .A1(n18710), .A2(n18693), .ZN(n17710) );
  OAI21_X1 U20932 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17710), .A(
        n17697), .ZN(n18695) );
  NAND2_X1 U20933 ( .A1(n17698), .A2(n17854), .ZN(n17711) );
  OAI21_X1 U20934 ( .B1(n18710), .B2(n17711), .A(n11593), .ZN(n17700) );
  OAI21_X1 U20935 ( .B1(n18695), .B2(n17700), .A(n17837), .ZN(n17699) );
  AOI21_X1 U20936 ( .B1(n18695), .B2(n17700), .A(n17699), .ZN(n17704) );
  AOI21_X1 U20937 ( .B1(n17846), .B2(n17714), .A(n17851), .ZN(n17721) );
  NAND2_X1 U20938 ( .A1(n17846), .A2(n19558), .ZN(n17713) );
  INV_X1 U20939 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19559) );
  AOI21_X1 U20940 ( .B1(n17721), .B2(n17713), .A(n19559), .ZN(n17703) );
  OAI22_X1 U20941 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17701), .B1(n17865), 
        .B2(n18129), .ZN(n17702) );
  NOR4_X1 U20942 ( .A1(n9696), .A2(n17704), .A3(n17703), .A4(n17702), .ZN(
        n17707) );
  OAI211_X1 U20943 ( .C1(n17708), .C2(n18129), .A(n17829), .B(n17705), .ZN(
        n17706) );
  OAI211_X1 U20944 ( .C1(n17852), .C2(n18697), .A(n17707), .B(n17706), .ZN(
        P3_U2658) );
  AOI211_X1 U20945 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17724), .A(n17708), .B(
        n17864), .ZN(n17709) );
  AOI21_X1 U20946 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17804), .A(n17709), .ZN(
        n17718) );
  AOI21_X1 U20947 ( .B1(n18710), .B2(n18693), .A(n17710), .ZN(n18713) );
  NAND2_X1 U20948 ( .A1(n11593), .A2(n17711), .ZN(n17712) );
  XNOR2_X1 U20949 ( .A(n18713), .B(n17712), .ZN(n17716) );
  OAI22_X1 U20950 ( .A1(n18710), .A2(n17852), .B1(n17714), .B2(n17713), .ZN(
        n17715) );
  AOI211_X1 U20951 ( .C1(n17837), .C2(n17716), .A(n9696), .B(n17715), .ZN(
        n17717) );
  OAI211_X1 U20952 ( .C1(n19558), .C2(n17721), .A(n17718), .B(n17717), .ZN(
        P3_U2659) );
  INV_X1 U20953 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21725) );
  INV_X1 U20954 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19553) );
  NOR2_X1 U20955 ( .A1(n21725), .A2(n19553), .ZN(n17735) );
  NOR3_X1 U20956 ( .A1(n17857), .A2(n19551), .A3(n17754), .ZN(n17750) );
  AOI21_X1 U20957 ( .B1(n17735), .B2(n17750), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17722) );
  INV_X1 U20958 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18740) );
  NAND2_X1 U20959 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17742), .ZN(
        n17741) );
  NOR2_X1 U20960 ( .A1(n18740), .A2(n17741), .ZN(n17731) );
  AOI21_X1 U20961 ( .B1(n17731), .B2(n17854), .A(n17820), .ZN(n17719) );
  OAI21_X1 U20962 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17731), .A(
        n18693), .ZN(n18721) );
  XOR2_X1 U20963 ( .A(n17719), .B(n18721), .Z(n17720) );
  OAI22_X1 U20964 ( .A1(n17722), .A2(n17721), .B1(n17823), .B2(n17720), .ZN(
        n17723) );
  AOI211_X1 U20965 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17844), .A(
        n9696), .B(n17723), .ZN(n17726) );
  OAI211_X1 U20966 ( .C1(n17727), .C2(n21783), .A(n17829), .B(n17724), .ZN(
        n17725) );
  OAI211_X1 U20967 ( .C1(n21783), .C2(n17865), .A(n17726), .B(n17725), .ZN(
        P3_U2660) );
  AOI211_X1 U20968 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17728), .A(n17727), .B(
        n17864), .ZN(n17729) );
  AOI211_X1 U20969 ( .C1(n17804), .C2(P3_EBX_REG_10__SCAN_IN), .A(n9696), .B(
        n17729), .ZN(n17739) );
  OAI21_X1 U20970 ( .B1(n17730), .B2(n17857), .A(n17868), .ZN(n17755) );
  AOI21_X1 U20971 ( .B1(n18740), .B2(n17741), .A(n17731), .ZN(n18743) );
  NAND2_X1 U20972 ( .A1(n17782), .A2(n17854), .ZN(n17772) );
  INV_X1 U20973 ( .A(n17772), .ZN(n17784) );
  AOI21_X1 U20974 ( .B1(n18720), .B2(n17784), .A(n17820), .ZN(n17744) );
  INV_X1 U20975 ( .A(n18743), .ZN(n17733) );
  INV_X1 U20976 ( .A(n17744), .ZN(n17732) );
  AOI221_X1 U20977 ( .B1(n18743), .B2(n17744), .C1(n17733), .C2(n17732), .A(
        n17823), .ZN(n17737) );
  INV_X1 U20978 ( .A(n17750), .ZN(n17734) );
  AOI211_X1 U20979 ( .C1(n21725), .C2(n19553), .A(n17735), .B(n17734), .ZN(
        n17736) );
  AOI211_X1 U20980 ( .C1(n17755), .C2(P3_REIP_REG_10__SCAN_IN), .A(n17737), 
        .B(n17736), .ZN(n17738) );
  OAI211_X1 U20981 ( .C1(n18740), .C2(n17852), .A(n17739), .B(n17738), .ZN(
        P3_U2661) );
  NOR2_X1 U20982 ( .A1(n17746), .A2(n17864), .ZN(n17757) );
  AOI22_X1 U20983 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17844), .B1(
        n17757), .B2(n17740), .ZN(n17752) );
  OAI21_X1 U20984 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17742), .A(
        n17741), .ZN(n18755) );
  NOR2_X1 U20985 ( .A1(n17743), .A2(n17772), .ZN(n17745) );
  OAI211_X1 U20986 ( .C1(n17745), .C2(n18755), .A(n17837), .B(n17744), .ZN(
        n17748) );
  OAI221_X1 U20987 ( .B1(n17804), .B2(n17829), .C1(n17804), .C2(n17746), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n17747) );
  OAI211_X1 U20988 ( .C1(n17856), .C2(n18755), .A(n17748), .B(n17747), .ZN(
        n17749) );
  AOI221_X1 U20989 ( .B1(n17755), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n17750), 
        .C2(n21725), .A(n17749), .ZN(n17751) );
  NAND3_X1 U20990 ( .A1(n17752), .A2(n17751), .A3(n10420), .ZN(P3_U2662) );
  AOI21_X1 U20991 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17784), .A(
        n17820), .ZN(n17774) );
  XNOR2_X1 U20992 ( .A(n17774), .B(n17753), .ZN(n17763) );
  NOR2_X1 U20993 ( .A1(n17857), .A2(n17754), .ZN(n17756) );
  OAI21_X1 U20994 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n17756), .A(n17755), .ZN(
        n17759) );
  OAI21_X1 U20995 ( .B1(n17764), .B2(n18238), .A(n17757), .ZN(n17758) );
  OAI211_X1 U20996 ( .C1(n17852), .C2(n17760), .A(n17759), .B(n17758), .ZN(
        n17761) );
  AOI211_X1 U20997 ( .C1(n17804), .C2(P3_EBX_REG_8__SCAN_IN), .A(n9696), .B(
        n17761), .ZN(n17762) );
  OAI21_X1 U20998 ( .B1(n17763), .B2(n17823), .A(n17762), .ZN(P3_U2663) );
  AOI221_X1 U20999 ( .B1(n19546), .B2(n17846), .C1(n17783), .C2(n17846), .A(
        n17851), .ZN(n17778) );
  AOI211_X1 U21000 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17765), .A(n17764), .B(
        n17864), .ZN(n17770) );
  NAND3_X1 U21001 ( .A1(n17846), .A2(n17766), .A3(n19548), .ZN(n17767) );
  OAI211_X1 U21002 ( .C1(n17768), .C2(n17852), .A(n10420), .B(n17767), .ZN(
        n17769) );
  AOI211_X1 U21003 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17804), .A(n17770), .B(
        n17769), .ZN(n17777) );
  INV_X1 U21004 ( .A(n17771), .ZN(n17775) );
  INV_X1 U21005 ( .A(n17856), .ZN(n17815) );
  AOI21_X1 U21006 ( .B1(n17775), .B2(n17772), .A(n17823), .ZN(n17773) );
  OAI22_X1 U21007 ( .A1(n17775), .A2(n17774), .B1(n17815), .B2(n17773), .ZN(
        n17776) );
  OAI211_X1 U21008 ( .C1(n17778), .C2(n19548), .A(n17777), .B(n17776), .ZN(
        P3_U2664) );
  AND2_X1 U21009 ( .A1(n17783), .A2(n17846), .ZN(n17790) );
  NOR2_X1 U21010 ( .A1(n17851), .A2(n17790), .ZN(n17793) );
  AOI211_X1 U21011 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17796), .A(n17779), .B(
        n17864), .ZN(n17781) );
  INV_X1 U21012 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18092) );
  OAI22_X1 U21013 ( .A1(n21610), .A2(n17852), .B1(n17865), .B2(n18092), .ZN(
        n17780) );
  NOR3_X1 U21014 ( .A1(n9696), .A2(n17781), .A3(n17780), .ZN(n17789) );
  AOI21_X1 U21015 ( .B1(n21610), .B2(n17792), .A(n17782), .ZN(n18768) );
  NAND2_X1 U21016 ( .A1(n17837), .A2(n17854), .ZN(n17855) );
  OAI21_X1 U21017 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17855), .A(
        n17856), .ZN(n17787) );
  NOR3_X1 U21018 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17857), .A3(n17783), .ZN(
        n17786) );
  NOR3_X1 U21019 ( .A1(n18768), .A2(n17784), .A3(n17853), .ZN(n17785) );
  AOI211_X1 U21020 ( .C1(n18768), .C2(n17787), .A(n17786), .B(n17785), .ZN(
        n17788) );
  OAI211_X1 U21021 ( .C1(n17793), .C2(n19546), .A(n17789), .B(n17788), .ZN(
        P3_U2665) );
  AOI22_X1 U21022 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17844), .B1(
        n17804), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n17800) );
  AOI21_X1 U21023 ( .B1(n17791), .B2(n17790), .A(n9696), .ZN(n17799) );
  NOR2_X1 U21024 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17860), .ZN(
        n17838) );
  AOI21_X1 U21025 ( .B1(n18773), .B2(n17838), .A(n17820), .ZN(n17810) );
  AND2_X1 U21026 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18773), .ZN(
        n17805) );
  OAI21_X1 U21027 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17805), .A(
        n17792), .ZN(n18775) );
  XNOR2_X1 U21028 ( .A(n17810), .B(n18775), .ZN(n17795) );
  INV_X1 U21029 ( .A(n17793), .ZN(n17794) );
  AOI22_X1 U21030 ( .A1(n17837), .A2(n17795), .B1(P3_REIP_REG_5__SCAN_IN), 
        .B2(n17794), .ZN(n17798) );
  OAI211_X1 U21031 ( .C1(n17801), .C2(n18091), .A(n17829), .B(n17796), .ZN(
        n17797) );
  NAND4_X1 U21032 ( .A1(n17800), .A2(n17799), .A3(n17798), .A4(n17797), .ZN(
        P3_U2666) );
  AOI211_X1 U21033 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17828), .A(n17801), .B(
        n17864), .ZN(n17803) );
  NOR3_X1 U21034 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17857), .A3(n17818), .ZN(
        n17802) );
  AOI211_X1 U21035 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17804), .A(n17803), .B(
        n17802), .ZN(n17817) );
  AOI21_X1 U21036 ( .B1(n21640), .B2(n17806), .A(n17805), .ZN(n18791) );
  INV_X1 U21037 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21648) );
  NAND2_X1 U21038 ( .A1(n19035), .A2(n19642), .ZN(n17872) );
  AOI21_X1 U21039 ( .B1(n21648), .B2(n14359), .A(n17872), .ZN(n17807) );
  OR2_X1 U21040 ( .A1(n17807), .A2(n9696), .ZN(n17814) );
  NAND2_X1 U21041 ( .A1(n17808), .A2(n21640), .ZN(n18785) );
  INV_X1 U21042 ( .A(n18785), .ZN(n17811) );
  INV_X1 U21043 ( .A(n18791), .ZN(n17809) );
  AOI22_X1 U21044 ( .A1(n17838), .A2(n17811), .B1(n17810), .B2(n17809), .ZN(
        n17812) );
  AOI21_X1 U21045 ( .B1(n17846), .B2(n17818), .A(n17851), .ZN(n17824) );
  OAI22_X1 U21046 ( .A1(n17812), .A2(n17823), .B1(n17824), .B2(n19543), .ZN(
        n17813) );
  AOI211_X1 U21047 ( .C1(n18791), .C2(n17815), .A(n17814), .B(n17813), .ZN(
        n17816) );
  OAI211_X1 U21048 ( .C1(n21640), .C2(n17852), .A(n17817), .B(n17816), .ZN(
        P3_U2667) );
  INV_X1 U21049 ( .A(n17872), .ZN(n17850) );
  NAND2_X1 U21050 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17845) );
  NAND2_X1 U21051 ( .A1(n17846), .A2(n17818), .ZN(n17819) );
  OAI22_X1 U21052 ( .A1(n17865), .A2(n18255), .B1(n17845), .B2(n17819), .ZN(
        n17826) );
  INV_X1 U21053 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19541) );
  AOI21_X1 U21054 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17838), .A(
        n17820), .ZN(n17836) );
  XOR2_X1 U21055 ( .A(n17836), .B(n17821), .Z(n17822) );
  OAI22_X1 U21056 ( .A1(n17824), .A2(n19541), .B1(n17823), .B2(n17822), .ZN(
        n17825) );
  AOI211_X1 U21057 ( .C1(n17827), .C2(n17850), .A(n17826), .B(n17825), .ZN(
        n17831) );
  OAI211_X1 U21058 ( .C1(n17833), .C2(n18255), .A(n17829), .B(n17828), .ZN(
        n17830) );
  OAI211_X1 U21059 ( .C1(n17852), .C2(n17832), .A(n17831), .B(n17830), .ZN(
        P3_U2668) );
  INV_X1 U21060 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18263) );
  INV_X1 U21061 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n21726) );
  INV_X1 U21062 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18278) );
  NAND2_X1 U21063 ( .A1(n21726), .A2(n18278), .ZN(n17834) );
  AOI211_X1 U21064 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17834), .A(n17833), .B(
        n17864), .ZN(n17843) );
  AOI22_X1 U21065 ( .A1(n17851), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n17850), 
        .B2(n17835), .ZN(n17840) );
  OAI211_X1 U21066 ( .C1(n17838), .C2(n17841), .A(n17837), .B(n17836), .ZN(
        n17839) );
  OAI211_X1 U21067 ( .C1(n17856), .C2(n17841), .A(n17840), .B(n17839), .ZN(
        n17842) );
  AOI211_X1 U21068 ( .C1(n17844), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17843), .B(n17842), .ZN(n17848) );
  OAI211_X1 U21069 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17846), .B(n17845), .ZN(n17847) );
  OAI211_X1 U21070 ( .C1(n18263), .C2(n17865), .A(n17848), .B(n17847), .ZN(
        P3_U2669) );
  NAND2_X1 U21071 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .ZN(n18265) );
  OAI21_X1 U21072 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n18265), .ZN(n18274) );
  AOI22_X1 U21073 ( .A1(n17851), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17850), 
        .B2(n17849), .ZN(n17863) );
  OAI21_X1 U21074 ( .B1(n17854), .B2(n17853), .A(n17852), .ZN(n17861) );
  NAND2_X1 U21075 ( .A1(n17856), .A2(n17855), .ZN(n17859) );
  OAI22_X1 U21076 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17857), .B1(n17865), 
        .B2(n21726), .ZN(n17858) );
  AOI221_X1 U21077 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17861), .C1(
        n17860), .C2(n17859), .A(n17858), .ZN(n17862) );
  OAI211_X1 U21078 ( .C1(n17864), .C2(n18274), .A(n17863), .B(n17862), .ZN(
        P3_U2670) );
  NAND2_X1 U21079 ( .A1(n17865), .A2(n17864), .ZN(n17867) );
  AOI22_X1 U21080 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17867), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17866), .ZN(n17871) );
  NAND3_X1 U21081 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17869), .A3(
        n17868), .ZN(n17870) );
  OAI211_X1 U21082 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17872), .A(
        n17871), .B(n17870), .ZN(P3_U2671) );
  INV_X1 U21083 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17930) );
  NAND4_X1 U21084 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_20__SCAN_IN), .A4(n18015), .ZN(n17873) );
  NOR4_X1 U21085 ( .A1(n17875), .A2(n17930), .A3(n17874), .A4(n17873), .ZN(
        n17876) );
  NAND4_X1 U21086 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17919), .A4(n17876), .ZN(n17879) );
  NOR2_X1 U21087 ( .A1(n17880), .A2(n17879), .ZN(n17914) );
  NAND2_X1 U21088 ( .A1(n18271), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17878) );
  NAND2_X1 U21089 ( .A1(n17914), .A2(n19065), .ZN(n17877) );
  OAI22_X1 U21090 ( .A1(n17914), .A2(n17878), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17877), .ZN(P3_U2672) );
  NAND2_X1 U21091 ( .A1(n17880), .A2(n17879), .ZN(n17881) );
  NAND2_X1 U21092 ( .A1(n17881), .A2(n18269), .ZN(n17913) );
  INV_X1 U21093 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17884) );
  AOI22_X1 U21094 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17883) );
  NAND2_X1 U21095 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n17882) );
  OAI211_X1 U21096 ( .C1(n18141), .C2(n17884), .A(n17883), .B(n17882), .ZN(
        n17885) );
  INV_X1 U21097 ( .A(n17885), .ZN(n17889) );
  AOI22_X1 U21098 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17888) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18229), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17887) );
  NAND3_X1 U21100 ( .A1(n17889), .A2(n17888), .A3(n17887), .ZN(n17896) );
  AOI22_X1 U21101 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U21102 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18152), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U21103 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17892) );
  AOI22_X1 U21104 ( .A1(n14395), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17891) );
  NAND4_X1 U21105 ( .A1(n17894), .A2(n17893), .A3(n17892), .A4(n17891), .ZN(
        n17895) );
  NOR2_X1 U21106 ( .A1(n17896), .A2(n17895), .ZN(n17912) );
  AOI22_X1 U21107 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17901) );
  AOI22_X1 U21108 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17900) );
  AOI22_X1 U21109 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17899) );
  AOI22_X1 U21110 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17898) );
  NAND4_X1 U21111 ( .A1(n17901), .A2(n17900), .A3(n17899), .A4(n17898), .ZN(
        n17911) );
  INV_X1 U21112 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U21113 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17903) );
  NAND2_X1 U21114 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n17902) );
  OAI211_X1 U21115 ( .C1(n17904), .C2(n18141), .A(n17903), .B(n17902), .ZN(
        n17910) );
  INV_X1 U21116 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17905) );
  OAI22_X1 U21117 ( .A1(n21584), .A2(n18186), .B1(n14388), .B2(n17905), .ZN(
        n17909) );
  INV_X1 U21118 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17907) );
  OAI22_X1 U21119 ( .A1(n14359), .A2(n17907), .B1(n13041), .B2(n17906), .ZN(
        n17908) );
  NAND2_X1 U21120 ( .A1(n17917), .A2(n17916), .ZN(n17915) );
  XNOR2_X1 U21121 ( .A(n17912), .B(n17915), .ZN(n18290) );
  OAI22_X1 U21122 ( .A1(n17914), .A2(n17913), .B1(n18290), .B2(n18269), .ZN(
        P3_U2673) );
  OAI21_X1 U21123 ( .B1(n17917), .B2(n17916), .A(n17915), .ZN(n18295) );
  NOR2_X1 U21124 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17925), .ZN(n17918) );
  AOI22_X1 U21125 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17920), .B1(n17919), 
        .B2(n17918), .ZN(n17921) );
  OAI21_X1 U21126 ( .B1(n18295), .B2(n18269), .A(n17921), .ZN(P3_U2674) );
  OAI21_X1 U21127 ( .B1(n17926), .B2(n17923), .A(n17922), .ZN(n18304) );
  NAND3_X1 U21128 ( .A1(n17925), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18269), 
        .ZN(n17924) );
  OAI221_X1 U21129 ( .B1(n17925), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18269), 
        .C2(n18304), .A(n17924), .ZN(P3_U2676) );
  NAND2_X1 U21130 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17939), .ZN(n17933) );
  AOI21_X1 U21131 ( .B1(n17927), .B2(n17931), .A(n17926), .ZN(n18305) );
  NAND2_X1 U21132 ( .A1(n18305), .A2(n18276), .ZN(n17928) );
  OAI221_X1 U21133 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17933), .C1(n17930), 
        .C2(n17929), .A(n17928), .ZN(P3_U2677) );
  OAI21_X1 U21134 ( .B1(n17935), .B2(n17932), .A(n17931), .ZN(n18313) );
  OAI211_X1 U21135 ( .C1(n17939), .C2(P3_EBX_REG_25__SCAN_IN), .A(n18271), .B(
        n17933), .ZN(n17934) );
  OAI21_X1 U21136 ( .B1(n18269), .B2(n18313), .A(n17934), .ZN(P3_U2678) );
  AOI21_X1 U21137 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18271), .A(n17945), .ZN(
        n17938) );
  AOI21_X1 U21138 ( .B1(n17936), .B2(n17941), .A(n17935), .ZN(n18314) );
  INV_X1 U21139 ( .A(n18314), .ZN(n17937) );
  OAI22_X1 U21140 ( .A1(n17939), .A2(n17938), .B1(n18271), .B2(n17937), .ZN(
        P3_U2679) );
  AOI21_X1 U21141 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18271), .A(n17940), .ZN(
        n17944) );
  OAI21_X1 U21142 ( .B1(n17943), .B2(n17942), .A(n17941), .ZN(n18323) );
  OAI22_X1 U21143 ( .A1(n17945), .A2(n17944), .B1(n18271), .B2(n18323), .ZN(
        P3_U2680) );
  INV_X1 U21144 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17948) );
  NAND2_X1 U21145 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n17947) );
  NAND2_X1 U21146 ( .A1(n18216), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n17946) );
  OAI211_X1 U21147 ( .C1(n17948), .C2(n18141), .A(n17947), .B(n17946), .ZN(
        n17949) );
  INV_X1 U21148 ( .A(n17949), .ZN(n17954) );
  AOI22_X1 U21149 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17953) );
  AOI22_X1 U21150 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17952) );
  INV_X1 U21151 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17950) );
  OR2_X1 U21152 ( .A1(n18224), .A2(n17950), .ZN(n17951) );
  NAND4_X1 U21153 ( .A1(n17954), .A2(n17953), .A3(n17952), .A4(n17951), .ZN(
        n17960) );
  AOI22_X1 U21154 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U21155 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17957) );
  AOI22_X1 U21156 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17956) );
  AOI22_X1 U21157 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17955) );
  NAND4_X1 U21158 ( .A1(n17958), .A2(n17957), .A3(n17956), .A4(n17955), .ZN(
        n17959) );
  OR2_X1 U21159 ( .A1(n17960), .A2(n17959), .ZN(n18324) );
  INV_X1 U21160 ( .A(n18324), .ZN(n17962) );
  NAND3_X1 U21161 ( .A1(n17963), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18269), 
        .ZN(n17961) );
  OAI221_X1 U21162 ( .B1(n17963), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18269), 
        .C2(n17962), .A(n17961), .ZN(P3_U2681) );
  INV_X1 U21163 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17966) );
  AOI22_X1 U21164 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17965) );
  NAND2_X1 U21165 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n17964) );
  OAI211_X1 U21166 ( .C1(n17966), .C2(n9702), .A(n17965), .B(n17964), .ZN(
        n17972) );
  INV_X1 U21167 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18122) );
  INV_X1 U21168 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17967) );
  OAI22_X1 U21169 ( .A1(n18203), .A2(n18122), .B1(n13142), .B2(n17967), .ZN(
        n17971) );
  OAI22_X1 U21170 ( .A1(n18200), .A2(n17969), .B1(n18198), .B2(n17968), .ZN(
        n17970) );
  OR3_X1 U21171 ( .A1(n17972), .A2(n17971), .A3(n17970), .ZN(n17978) );
  AOI22_X1 U21172 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17976) );
  AOI22_X1 U21173 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17975) );
  AOI22_X1 U21174 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U21175 ( .A1(n9707), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17973) );
  NAND4_X1 U21176 ( .A1(n17976), .A2(n17975), .A3(n17974), .A4(n17973), .ZN(
        n17977) );
  NOR2_X1 U21177 ( .A1(n17978), .A2(n17977), .ZN(n18332) );
  AOI21_X1 U21178 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18015), .A(n18276), .ZN(
        n17982) );
  AOI22_X1 U21179 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17982), .B1(n17980), 
        .B2(n17979), .ZN(n17981) );
  OAI21_X1 U21180 ( .B1(n18332), .B2(n18269), .A(n17981), .ZN(P3_U2682) );
  INV_X1 U21181 ( .A(n17982), .ZN(n17998) );
  AOI22_X1 U21182 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U21183 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U21184 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U21185 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17983) );
  NAND4_X1 U21186 ( .A1(n17986), .A2(n17985), .A3(n17984), .A4(n17983), .ZN(
        n17994) );
  INV_X1 U21187 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17989) );
  AOI22_X1 U21188 ( .A1(n17890), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17988) );
  NAND2_X1 U21189 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n17987) );
  OAI211_X1 U21190 ( .C1(n17989), .C2(n18141), .A(n17988), .B(n17987), .ZN(
        n17993) );
  AOI22_X1 U21191 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U21192 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17990) );
  NAND2_X1 U21193 ( .A1(n17991), .A2(n17990), .ZN(n17992) );
  OR3_X1 U21194 ( .A1(n17994), .A2(n17993), .A3(n17992), .ZN(n18335) );
  NAND2_X1 U21195 ( .A1(n18276), .A2(n18335), .ZN(n17995) );
  OAI221_X1 U21196 ( .B1(n17998), .B2(n17997), .C1(n17998), .C2(n17996), .A(
        n17995), .ZN(P3_U2683) );
  INV_X1 U21197 ( .A(n17999), .ZN(n18000) );
  OAI21_X1 U21198 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18000), .A(n18271), .ZN(
        n18014) );
  AOI22_X1 U21199 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18002) );
  NAND2_X1 U21200 ( .A1(n9707), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n18001) );
  OAI211_X1 U21201 ( .C1(n18003), .C2(n18224), .A(n18002), .B(n18001), .ZN(
        n18004) );
  INV_X1 U21202 ( .A(n18004), .ZN(n18007) );
  AOI22_X1 U21203 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18006) );
  AOI22_X1 U21204 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18005) );
  NAND3_X1 U21205 ( .A1(n18007), .A2(n18006), .A3(n18005), .ZN(n18013) );
  AOI22_X1 U21206 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18011) );
  AOI22_X1 U21207 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18010) );
  AOI22_X1 U21208 ( .A1(n13086), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U21209 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18008) );
  NAND4_X1 U21210 ( .A1(n18011), .A2(n18010), .A3(n18009), .A4(n18008), .ZN(
        n18012) );
  NOR2_X1 U21211 ( .A1(n18013), .A2(n18012), .ZN(n18344) );
  OAI22_X1 U21212 ( .A1(n18015), .A2(n18014), .B1(n18344), .B2(n18269), .ZN(
        P3_U2684) );
  NAND2_X1 U21213 ( .A1(n18269), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U21214 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18207), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U21215 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18018) );
  AOI22_X1 U21216 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18017) );
  AOI22_X1 U21217 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18016) );
  NAND4_X1 U21218 ( .A1(n18019), .A2(n18018), .A3(n18017), .A4(n18016), .ZN(
        n18030) );
  INV_X1 U21219 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U21220 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18021) );
  NAND2_X1 U21221 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n18020) );
  OAI211_X1 U21222 ( .C1(n18022), .C2(n18141), .A(n18021), .B(n18020), .ZN(
        n18029) );
  INV_X1 U21223 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18024) );
  INV_X1 U21224 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18023) );
  OAI22_X1 U21225 ( .A1(n18186), .A2(n18024), .B1(n14388), .B2(n18023), .ZN(
        n18028) );
  INV_X1 U21226 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18026) );
  OAI22_X1 U21227 ( .A1(n14359), .A2(n18026), .B1(n13041), .B2(n18025), .ZN(
        n18027) );
  OR4_X1 U21228 ( .A1(n18030), .A2(n18029), .A3(n18028), .A4(n18027), .ZN(
        n18345) );
  INV_X1 U21229 ( .A(n18273), .ZN(n18275) );
  NAND2_X1 U21230 ( .A1(n18031), .A2(n18275), .ZN(n18072) );
  NOR2_X1 U21231 ( .A1(n18071), .A2(n18072), .ZN(n18049) );
  NOR2_X1 U21232 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18050), .ZN(n18032) );
  AOI22_X1 U21233 ( .A1(n18276), .A2(n18345), .B1(n18049), .B2(n18032), .ZN(
        n18033) );
  OAI21_X1 U21234 ( .B1(n18035), .B2(n18034), .A(n18033), .ZN(P3_U2685) );
  AOI22_X1 U21235 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18037) );
  NAND2_X1 U21236 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n18036) );
  OAI211_X1 U21237 ( .C1(n18038), .C2(n13041), .A(n18037), .B(n18036), .ZN(
        n18039) );
  INV_X1 U21238 ( .A(n18039), .ZN(n18042) );
  AOI22_X1 U21239 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18041) );
  AOI22_X1 U21240 ( .A1(n9707), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9701), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18040) );
  NAND3_X1 U21241 ( .A1(n18042), .A2(n18041), .A3(n18040), .ZN(n18048) );
  AOI22_X1 U21242 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18046) );
  AOI22_X1 U21243 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18045) );
  AOI22_X1 U21244 ( .A1(n14395), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18152), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18044) );
  AOI22_X1 U21245 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13929), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18043) );
  NAND4_X1 U21246 ( .A1(n18046), .A2(n18045), .A3(n18044), .A4(n18043), .ZN(
        n18047) );
  NOR2_X1 U21247 ( .A1(n18048), .A2(n18047), .ZN(n18356) );
  NOR2_X1 U21248 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18049), .ZN(n18053) );
  AOI211_X1 U21249 ( .C1(n19065), .C2(n18051), .A(n18050), .B(n18264), .ZN(
        n18052) );
  OAI22_X1 U21250 ( .A1(n18356), .A2(n18269), .B1(n18053), .B2(n18052), .ZN(
        P3_U2686) );
  NAND2_X1 U21251 ( .A1(n18271), .A2(n18072), .ZN(n18095) );
  AOI22_X1 U21252 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18057) );
  AOI22_X1 U21253 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18056) );
  AOI22_X1 U21254 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18055) );
  AOI22_X1 U21255 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18054) );
  NAND4_X1 U21256 ( .A1(n18057), .A2(n18056), .A3(n18055), .A4(n18054), .ZN(
        n18069) );
  AOI22_X1 U21257 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18060) );
  NAND2_X1 U21258 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n18059) );
  OAI211_X1 U21259 ( .C1(n18061), .C2(n18141), .A(n18060), .B(n18059), .ZN(
        n18068) );
  INV_X1 U21260 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18063) );
  OAI22_X1 U21261 ( .A1(n18186), .A2(n18063), .B1(n14388), .B2(n18062), .ZN(
        n18067) );
  INV_X1 U21262 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18065) );
  INV_X1 U21263 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18064) );
  OAI22_X1 U21264 ( .A1(n14359), .A2(n18065), .B1(n13041), .B2(n18064), .ZN(
        n18066) );
  OR4_X1 U21265 ( .A1(n18069), .A2(n18068), .A3(n18067), .A4(n18066), .ZN(
        n18357) );
  NAND2_X1 U21266 ( .A1(n18276), .A2(n18357), .ZN(n18070) );
  OAI221_X1 U21267 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18072), .C1(n18071), 
        .C2(n18095), .A(n18070), .ZN(P3_U2687) );
  AOI22_X1 U21268 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18076) );
  AOI22_X1 U21269 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U21270 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U21271 ( .A1(n9707), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18073) );
  NAND4_X1 U21272 ( .A1(n18076), .A2(n18075), .A3(n18074), .A4(n18073), .ZN(
        n18090) );
  INV_X1 U21273 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18230), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18078) );
  NAND2_X1 U21275 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n18077) );
  OAI211_X1 U21276 ( .C1(n18080), .C2(n18079), .A(n18078), .B(n18077), .ZN(
        n18088) );
  OAI22_X1 U21277 ( .A1(n11711), .A2(n18082), .B1(n13142), .B2(n18081), .ZN(
        n18087) );
  INV_X1 U21278 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18083) );
  OAI22_X1 U21279 ( .A1(n18085), .A2(n18084), .B1(n18186), .B2(n18083), .ZN(
        n18086) );
  OR3_X1 U21280 ( .A1(n18088), .A2(n18087), .A3(n18086), .ZN(n18089) );
  NOR2_X1 U21281 ( .A1(n18090), .A2(n18089), .ZN(n18370) );
  NOR2_X1 U21282 ( .A1(n18112), .A2(n18129), .ZN(n18094) );
  NOR3_X1 U21283 ( .A1(n18091), .A2(n18264), .A3(n18254), .ZN(n18248) );
  INV_X1 U21284 ( .A(n18248), .ZN(n18250) );
  NOR2_X1 U21285 ( .A1(n18092), .A2(n18250), .ZN(n18243) );
  NAND2_X1 U21286 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n18243), .ZN(n18237) );
  NAND3_X1 U21287 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n18173), .ZN(n18169) );
  AOI21_X1 U21288 ( .B1(n18094), .B2(n18131), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n18096) );
  OAI22_X1 U21289 ( .A1(n18370), .A2(n18269), .B1(n18096), .B2(n18095), .ZN(
        P3_U2688) );
  INV_X1 U21290 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18099) );
  NAND2_X1 U21291 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n18098) );
  NAND2_X1 U21292 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n18097) );
  OAI211_X1 U21293 ( .C1(n18099), .C2(n18141), .A(n18098), .B(n18097), .ZN(
        n18100) );
  INV_X1 U21294 ( .A(n18100), .ZN(n18105) );
  AOI22_X1 U21295 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18104) );
  AOI22_X1 U21296 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18103) );
  INV_X1 U21297 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18101) );
  OR2_X1 U21298 ( .A1(n18224), .A2(n18101), .ZN(n18102) );
  NAND4_X1 U21299 ( .A1(n18105), .A2(n18104), .A3(n18103), .A4(n18102), .ZN(
        n18111) );
  AOI22_X1 U21300 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18207), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18109) );
  AOI22_X1 U21301 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18108) );
  AOI22_X1 U21302 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18107) );
  AOI22_X1 U21303 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18106) );
  NAND4_X1 U21304 ( .A1(n18109), .A2(n18108), .A3(n18107), .A4(n18106), .ZN(
        n18110) );
  OR2_X1 U21305 ( .A1(n18111), .A2(n18110), .ZN(n18374) );
  INV_X1 U21306 ( .A(n18374), .ZN(n18115) );
  INV_X1 U21307 ( .A(n18131), .ZN(n18130) );
  OAI211_X1 U21308 ( .C1(n18129), .C2(n18130), .A(P3_EBX_REG_14__SCAN_IN), .B(
        n18269), .ZN(n18114) );
  NAND4_X1 U21309 ( .A1(n19065), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n18131), 
        .A4(n18112), .ZN(n18113) );
  OAI211_X1 U21310 ( .C1(n18115), .C2(n18271), .A(n18114), .B(n18113), .ZN(
        P3_U2689) );
  AOI22_X1 U21311 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U21312 ( .A1(n13086), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U21313 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18117) );
  AOI22_X1 U21314 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18116) );
  NAND4_X1 U21315 ( .A1(n18119), .A2(n18118), .A3(n18117), .A4(n18116), .ZN(
        n18128) );
  AOI22_X1 U21316 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18194), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18121) );
  NAND2_X1 U21317 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n18120) );
  OAI211_X1 U21318 ( .C1(n18122), .C2(n18141), .A(n18121), .B(n18120), .ZN(
        n18123) );
  INV_X1 U21319 ( .A(n18123), .ZN(n18126) );
  AOI22_X1 U21320 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U21321 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18124) );
  NAND3_X1 U21322 ( .A1(n18126), .A2(n18125), .A3(n18124), .ZN(n18127) );
  NOR2_X1 U21323 ( .A1(n18128), .A2(n18127), .ZN(n18378) );
  AOI21_X1 U21324 ( .B1(n18271), .B2(n18130), .A(n18129), .ZN(n18133) );
  AOI21_X1 U21325 ( .B1(n19065), .B2(n18131), .A(P3_EBX_REG_13__SCAN_IN), .ZN(
        n18132) );
  OAI22_X1 U21326 ( .A1(n18378), .A2(n18271), .B1(n18133), .B2(n18132), .ZN(
        P3_U2690) );
  AOI22_X1 U21327 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U21328 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18220), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18137) );
  AOI22_X1 U21329 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18136) );
  AOI22_X1 U21330 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18135) );
  NAND4_X1 U21331 ( .A1(n18138), .A2(n18137), .A3(n18136), .A4(n18135), .ZN(
        n18148) );
  INV_X1 U21332 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U21333 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13086), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18140) );
  NAND2_X1 U21334 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n18139) );
  OAI211_X1 U21335 ( .C1(n18142), .C2(n18141), .A(n18140), .B(n18139), .ZN(
        n18143) );
  INV_X1 U21336 ( .A(n18143), .ZN(n18146) );
  AOI22_X1 U21337 ( .A1(n9701), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18145) );
  AOI22_X1 U21338 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18144) );
  NAND3_X1 U21339 ( .A1(n18146), .A2(n18145), .A3(n18144), .ZN(n18147) );
  NOR2_X1 U21340 ( .A1(n18148), .A2(n18147), .ZN(n18383) );
  INV_X1 U21341 ( .A(n18169), .ZN(n18149) );
  OAI33_X1 U21342 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18364), .A3(n18169), 
        .B1(n21756), .B2(n18276), .B3(n18149), .ZN(n18150) );
  INV_X1 U21343 ( .A(n18150), .ZN(n18151) );
  OAI21_X1 U21344 ( .B1(n18383), .B2(n18269), .A(n18151), .ZN(P3_U2691) );
  NAND2_X1 U21345 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n18155) );
  NAND2_X1 U21346 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n18154) );
  OAI211_X1 U21347 ( .C1(n18156), .C2(n18141), .A(n18155), .B(n18154), .ZN(
        n18157) );
  INV_X1 U21348 ( .A(n18157), .ZN(n18162) );
  AOI22_X1 U21349 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U21350 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18160) );
  INV_X1 U21351 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18260) );
  OR2_X1 U21352 ( .A1(n18224), .A2(n18260), .ZN(n18159) );
  NAND4_X1 U21353 ( .A1(n18162), .A2(n18161), .A3(n18160), .A4(n18159), .ZN(
        n18168) );
  AOI22_X1 U21354 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18166) );
  AOI22_X1 U21355 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13086), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18165) );
  AOI22_X1 U21356 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18164) );
  AOI22_X1 U21357 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18163) );
  NAND4_X1 U21358 ( .A1(n18166), .A2(n18165), .A3(n18164), .A4(n18163), .ZN(
        n18167) );
  OR2_X1 U21359 ( .A1(n18168), .A2(n18167), .ZN(n18386) );
  INV_X1 U21360 ( .A(n18386), .ZN(n18172) );
  AOI21_X1 U21361 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18173), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n18171) );
  NAND2_X1 U21362 ( .A1(n18271), .A2(n18169), .ZN(n18170) );
  OAI22_X1 U21363 ( .A1(n18172), .A2(n18271), .B1(n18171), .B2(n18170), .ZN(
        P3_U2692) );
  NAND2_X1 U21364 ( .A1(n19065), .A2(n18173), .ZN(n18193) );
  NOR2_X1 U21365 ( .A1(n18276), .A2(n18173), .ZN(n18214) );
  AOI22_X1 U21366 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18179) );
  AOI22_X1 U21367 ( .A1(n17886), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18178) );
  AOI22_X1 U21368 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U21369 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18176) );
  NAND4_X1 U21370 ( .A1(n18179), .A2(n18178), .A3(n18177), .A4(n18176), .ZN(
        n18191) );
  INV_X1 U21371 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U21372 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18182) );
  NAND2_X1 U21373 ( .A1(n18180), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n18181) );
  OAI211_X1 U21374 ( .C1(n18183), .C2(n18141), .A(n18182), .B(n18181), .ZN(
        n18190) );
  INV_X1 U21375 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18184) );
  OAI22_X1 U21376 ( .A1(n18186), .A2(n18185), .B1(n14388), .B2(n18184), .ZN(
        n18189) );
  OAI22_X1 U21377 ( .A1(n21564), .A2(n14359), .B1(n13041), .B2(n18187), .ZN(
        n18188) );
  OR4_X1 U21378 ( .A1(n18191), .A2(n18190), .A3(n18189), .A4(n18188), .ZN(
        n18389) );
  AOI22_X1 U21379 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18214), .B1(n18276), 
        .B2(n18389), .ZN(n18192) );
  OAI21_X1 U21380 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18193), .A(n18192), .ZN(
        P3_U2693) );
  INV_X1 U21381 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18272) );
  AOI22_X1 U21382 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18216), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18196) );
  NAND2_X1 U21383 ( .A1(n18194), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n18195) );
  OAI211_X1 U21384 ( .C1(n18272), .C2(n18224), .A(n18196), .B(n18195), .ZN(
        n18206) );
  OAI22_X1 U21385 ( .A1(n18200), .A2(n18199), .B1(n18198), .B2(n18197), .ZN(
        n18205) );
  INV_X1 U21386 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18201) );
  OAI22_X1 U21387 ( .A1(n18203), .A2(n18202), .B1(n9702), .B2(n18201), .ZN(
        n18204) );
  OR3_X1 U21388 ( .A1(n18206), .A2(n18205), .A3(n18204), .ZN(n18213) );
  AOI22_X1 U21389 ( .A1(n11663), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18221), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U21390 ( .A1(n18207), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U21391 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U21392 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18208) );
  NAND4_X1 U21393 ( .A1(n18211), .A2(n18210), .A3(n18209), .A4(n18208), .ZN(
        n18212) );
  NOR2_X1 U21394 ( .A1(n18213), .A2(n18212), .ZN(n18395) );
  NOR2_X1 U21395 ( .A1(n18238), .A2(n18237), .ZN(n18241) );
  OAI21_X1 U21396 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18241), .A(n18214), .ZN(
        n18215) );
  OAI21_X1 U21397 ( .B1(n18395), .B2(n18269), .A(n18215), .ZN(P3_U2694) );
  NAND2_X1 U21398 ( .A1(n18152), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n18218) );
  NAND2_X1 U21399 ( .A1(n18216), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n18217) );
  OAI211_X1 U21400 ( .C1(n21580), .C2(n18141), .A(n18218), .B(n18217), .ZN(
        n18219) );
  INV_X1 U21401 ( .A(n18219), .ZN(n18228) );
  AOI22_X1 U21402 ( .A1(n18221), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9707), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18227) );
  AOI22_X1 U21403 ( .A1(n13929), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18222), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18226) );
  OR2_X1 U21404 ( .A1(n18224), .A2(n18223), .ZN(n18225) );
  NAND4_X1 U21405 ( .A1(n18228), .A2(n18227), .A3(n18226), .A4(n18225), .ZN(
        n18236) );
  AOI22_X1 U21406 ( .A1(n18229), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18234) );
  AOI22_X1 U21407 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14395), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U21408 ( .A1(n18175), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13047), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U21409 ( .A1(n18230), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18231) );
  NAND4_X1 U21410 ( .A1(n18234), .A2(n18233), .A3(n18232), .A4(n18231), .ZN(
        n18235) );
  OR2_X1 U21411 ( .A1(n18236), .A2(n18235), .ZN(n18398) );
  INV_X1 U21412 ( .A(n18398), .ZN(n18242) );
  AOI21_X1 U21413 ( .B1(n18238), .B2(n18237), .A(n18276), .ZN(n18239) );
  INV_X1 U21414 ( .A(n18239), .ZN(n18240) );
  OAI22_X1 U21415 ( .A1(n18242), .A2(n18271), .B1(n18241), .B2(n18240), .ZN(
        P3_U2695) );
  OR3_X1 U21416 ( .A1(n18254), .A2(n18273), .A3(P3_EBX_REG_7__SCAN_IN), .ZN(
        n18245) );
  NOR2_X1 U21417 ( .A1(n18276), .A2(n18243), .ZN(n18247) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18276), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n18247), .ZN(n18244) );
  OAI21_X1 U21419 ( .B1(n18246), .B2(n18245), .A(n18244), .ZN(P3_U2696) );
  OAI21_X1 U21420 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18248), .A(n18247), .ZN(
        n18249) );
  OAI21_X1 U21421 ( .B1(n18269), .B2(n18101), .A(n18249), .ZN(P3_U2697) );
  NOR2_X1 U21422 ( .A1(n18264), .A2(n18254), .ZN(n18251) );
  OAI21_X1 U21423 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18251), .A(n18250), .ZN(
        n18252) );
  AOI22_X1 U21424 ( .A1(n18276), .A2(n18253), .B1(n18252), .B2(n18269), .ZN(
        P3_U2698) );
  NOR2_X1 U21425 ( .A1(n18254), .A2(n18273), .ZN(n18258) );
  NOR3_X1 U21426 ( .A1(n18255), .A2(n18259), .A3(n18273), .ZN(n18262) );
  AOI21_X1 U21427 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18271), .A(n18262), .ZN(
        n18257) );
  INV_X1 U21428 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18256) );
  OAI22_X1 U21429 ( .A1(n18258), .A2(n18257), .B1(n18256), .B2(n18269), .ZN(
        P3_U2699) );
  NOR2_X1 U21430 ( .A1(n18259), .A2(n18273), .ZN(n18266) );
  AOI21_X1 U21431 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18271), .A(n18266), .ZN(
        n18261) );
  OAI22_X1 U21432 ( .A1(n18262), .A2(n18261), .B1(n18260), .B2(n18269), .ZN(
        P3_U2700) );
  OAI221_X1 U21433 ( .B1(n18265), .B2(n18264), .C1(n19065), .C2(n18264), .A(
        n18263), .ZN(n18268) );
  INV_X1 U21434 ( .A(n18266), .ZN(n18267) );
  OAI211_X1 U21435 ( .C1(n18269), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n18268), .B(n18267), .ZN(n18270) );
  INV_X1 U21436 ( .A(n18270), .ZN(P3_U2701) );
  OAI222_X1 U21437 ( .A1(n18274), .A2(n18273), .B1(n21726), .B2(n18279), .C1(
        n18272), .C2(n18271), .ZN(P3_U2702) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18276), .B1(
        n18275), .B2(n18278), .ZN(n18277) );
  OAI21_X1 U21439 ( .B1(n18279), .B2(n18278), .A(n18277), .ZN(P3_U2703) );
  INV_X1 U21440 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18431) );
  INV_X1 U21441 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18434) );
  INV_X1 U21442 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18438) );
  NAND2_X1 U21443 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .ZN(n18404) );
  NAND4_X1 U21444 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n18280) );
  NOR3_X1 U21445 ( .A1(n18281), .A2(n18404), .A3(n18280), .ZN(n18371) );
  NAND2_X1 U21446 ( .A1(n18282), .A2(n18371), .ZN(n18400) );
  NAND2_X1 U21447 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n18381) );
  NAND4_X1 U21448 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n18283)
         );
  OR4_X2 U21449 ( .A1(n18400), .A2(n18470), .A3(n18381), .A4(n18283), .ZN(
        n18365) );
  INV_X1 U21450 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18448) );
  INV_X1 U21451 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18450) );
  NOR2_X1 U21452 ( .A1(n18448), .A2(n18450), .ZN(n18325) );
  NAND4_X1 U21453 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n18325), .ZN(n18330) );
  NOR2_X2 U21454 ( .A1(n18434), .A2(n18306), .ZN(n18300) );
  NAND3_X1 U21455 ( .A1(n18415), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n18287), 
        .ZN(n18285) );
  NOR2_X2 U21456 ( .A1(n19058), .A2(n18415), .ZN(n18358) );
  NAND2_X1 U21457 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18358), .ZN(n18284) );
  OAI211_X1 U21458 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n18287), .A(n18285), .B(
        n18284), .ZN(P3_U2704) );
  AOI22_X1 U21459 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18358), .ZN(n18289) );
  OAI211_X1 U21460 ( .C1(n18290), .C2(n18421), .A(n18289), .B(n18288), .ZN(
        P3_U2705) );
  AOI22_X1 U21461 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18358), .ZN(n18294) );
  AOI211_X1 U21462 ( .C1(n18431), .C2(n18297), .A(n18291), .B(n18346), .ZN(
        n18292) );
  INV_X1 U21463 ( .A(n18292), .ZN(n18293) );
  OAI211_X1 U21464 ( .C1(n18295), .C2(n18421), .A(n18294), .B(n18293), .ZN(
        P3_U2706) );
  INV_X1 U21465 ( .A(n18358), .ZN(n18331) );
  AOI22_X1 U21466 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18351), .B1(n18399), .B2(
        n18296), .ZN(n18299) );
  OAI211_X1 U21467 ( .C1(n18300), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18415), .B(
        n18297), .ZN(n18298) );
  OAI211_X1 U21468 ( .C1(n18331), .C2(n19049), .A(n18299), .B(n18298), .ZN(
        P3_U2707) );
  AOI22_X1 U21469 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18358), .ZN(n18303) );
  AOI211_X1 U21470 ( .C1(n18434), .C2(n18306), .A(n18300), .B(n18346), .ZN(
        n18301) );
  INV_X1 U21471 ( .A(n18301), .ZN(n18302) );
  OAI211_X1 U21472 ( .C1(n18304), .C2(n18421), .A(n18303), .B(n18302), .ZN(
        P3_U2708) );
  AOI22_X1 U21473 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18358), .B1(n18399), .B2(
        n18305), .ZN(n18308) );
  OAI211_X1 U21474 ( .C1(n18309), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18415), .B(
        n18306), .ZN(n18307) );
  OAI211_X1 U21475 ( .C1(n18363), .C2(n18521), .A(n18308), .B(n18307), .ZN(
        P3_U2709) );
  AOI22_X1 U21476 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18358), .ZN(n18312) );
  AOI211_X1 U21477 ( .C1(n18438), .C2(n18315), .A(n18309), .B(n18346), .ZN(
        n18310) );
  INV_X1 U21478 ( .A(n18310), .ZN(n18311) );
  OAI211_X1 U21479 ( .C1(n18313), .C2(n18421), .A(n18312), .B(n18311), .ZN(
        P3_U2710) );
  AOI22_X1 U21480 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18358), .B1(n18399), .B2(
        n18314), .ZN(n18318) );
  OAI211_X1 U21481 ( .C1(n18316), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18415), .B(
        n18315), .ZN(n18317) );
  OAI211_X1 U21482 ( .C1(n18363), .C2(n18517), .A(n18318), .B(n18317), .ZN(
        P3_U2711) );
  AOI22_X1 U21483 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18358), .ZN(n18322) );
  OAI211_X1 U21484 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18320), .A(n18415), .B(
        n18319), .ZN(n18321) );
  OAI211_X1 U21485 ( .C1(n18323), .C2(n18421), .A(n18322), .B(n18321), .ZN(
        P3_U2712) );
  NAND2_X1 U21486 ( .A1(n18353), .A2(n18444), .ZN(n18329) );
  AOI22_X1 U21487 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18358), .B1(n18399), .B2(
        n18324), .ZN(n18328) );
  INV_X1 U21488 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18452) );
  NAND2_X1 U21489 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18353), .ZN(n18352) );
  NAND2_X1 U21490 ( .A1(n18325), .A2(n18347), .ZN(n18336) );
  NAND2_X1 U21491 ( .A1(n18415), .A2(n18336), .ZN(n18340) );
  OAI21_X1 U21492 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18372), .A(n18340), .ZN(
        n18326) );
  AOI22_X1 U21493 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18351), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n18326), .ZN(n18327) );
  OAI211_X1 U21494 ( .C1(n18330), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P3_U2713) );
  INV_X1 U21495 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18446) );
  OAI22_X1 U21496 ( .A1(n18332), .A2(n18421), .B1(n16425), .B2(n18331), .ZN(
        n18333) );
  AOI21_X1 U21497 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18351), .A(n18333), .ZN(
        n18334) );
  OAI221_X1 U21498 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18336), .C1(n18446), 
        .C2(n18340), .A(n18334), .ZN(P3_U2714) );
  AOI22_X1 U21499 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18351), .B1(n18399), .B2(
        n18335), .ZN(n18339) );
  NAND2_X1 U21500 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18347), .ZN(n18341) );
  INV_X1 U21501 ( .A(n18341), .ZN(n18337) );
  AOI22_X1 U21502 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18358), .B1(n18337), .B2(
        n18336), .ZN(n18338) );
  OAI211_X1 U21503 ( .C1(n18448), .C2(n18340), .A(n18339), .B(n18338), .ZN(
        P3_U2715) );
  AOI22_X1 U21504 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18358), .ZN(n18343) );
  OAI211_X1 U21505 ( .C1(n18347), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18415), .B(
        n18341), .ZN(n18342) );
  OAI211_X1 U21506 ( .C1(n18344), .C2(n18421), .A(n18343), .B(n18342), .ZN(
        P3_U2716) );
  AOI22_X1 U21507 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18358), .B1(n18399), .B2(
        n18345), .ZN(n18350) );
  AOI211_X1 U21508 ( .C1(n18452), .C2(n18352), .A(n18347), .B(n18346), .ZN(
        n18348) );
  INV_X1 U21509 ( .A(n18348), .ZN(n18349) );
  OAI211_X1 U21510 ( .C1(n18363), .C2(n19041), .A(n18350), .B(n18349), .ZN(
        P3_U2717) );
  AOI22_X1 U21511 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18358), .ZN(n18355) );
  OAI211_X1 U21512 ( .C1(n18353), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18415), .B(
        n18352), .ZN(n18354) );
  OAI211_X1 U21513 ( .C1(n18356), .C2(n18421), .A(n18355), .B(n18354), .ZN(
        P3_U2718) );
  AOI22_X1 U21514 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n18358), .B1(n18399), .B2(
        n18357), .ZN(n18362) );
  OAI211_X1 U21515 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18360), .A(n18415), .B(
        n18359), .ZN(n18361) );
  OAI211_X1 U21516 ( .C1(n18363), .C2(n19029), .A(n18362), .B(n18361), .ZN(
        P3_U2719) );
  NOR2_X1 U21517 ( .A1(n18364), .A2(n18365), .ZN(n18367) );
  NAND2_X1 U21518 ( .A1(n18415), .A2(n18365), .ZN(n18376) );
  INV_X1 U21519 ( .A(n18376), .ZN(n18366) );
  MUX2_X1 U21520 ( .A(n18367), .B(n18366), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n18368) );
  AOI21_X1 U21521 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n18390), .A(n18368), .ZN(
        n18369) );
  OAI21_X1 U21522 ( .B1(n18370), .B2(n18421), .A(n18369), .ZN(P3_U2720) );
  INV_X1 U21523 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18464) );
  INV_X1 U21524 ( .A(n18371), .ZN(n18373) );
  NOR3_X1 U21525 ( .A1(n18464), .A2(n18381), .A3(n18392), .ZN(n18385) );
  NAND2_X1 U21526 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18385), .ZN(n18377) );
  INV_X1 U21527 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18531) );
  AOI22_X1 U21528 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18390), .B1(n18399), .B2(
        n18374), .ZN(n18375) );
  OAI221_X1 U21529 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18377), .C1(n18531), 
        .C2(n18376), .A(n18375), .ZN(P3_U2721) );
  INV_X1 U21530 ( .A(n18377), .ZN(n18380) );
  AOI21_X1 U21531 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18415), .A(n18385), .ZN(
        n18379) );
  OAI222_X1 U21532 ( .A1(n18424), .A2(n18529), .B1(n18380), .B2(n18379), .C1(
        n18421), .C2(n18378), .ZN(P3_U2722) );
  NOR2_X1 U21533 ( .A1(n18381), .A2(n18392), .ZN(n18382) );
  AOI21_X1 U21534 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18415), .A(n18382), .ZN(
        n18384) );
  OAI222_X1 U21535 ( .A1(n18424), .A2(n18525), .B1(n18385), .B2(n18384), .C1(
        n18421), .C2(n18383), .ZN(P3_U2723) );
  INV_X1 U21536 ( .A(n18392), .ZN(n18397) );
  NAND2_X1 U21537 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18397), .ZN(n18388) );
  INV_X1 U21538 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18523) );
  INV_X1 U21539 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18467) );
  OAI21_X1 U21540 ( .B1(n18467), .B2(n18392), .A(n18415), .ZN(n18393) );
  AOI22_X1 U21541 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18390), .B1(n18399), .B2(
        n18386), .ZN(n18387) );
  OAI221_X1 U21542 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18388), .C1(n18523), 
        .C2(n18393), .A(n18387), .ZN(P3_U2724) );
  AOI22_X1 U21543 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18390), .B1(n18399), .B2(
        n18389), .ZN(n18391) );
  OAI221_X1 U21544 ( .B1(n18393), .B2(n18467), .C1(n18393), .C2(n18392), .A(
        n18391), .ZN(P3_U2725) );
  AOI21_X1 U21545 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18415), .A(n18394), .ZN(
        n18396) );
  OAI222_X1 U21546 ( .A1(n18424), .A2(n18519), .B1(n18397), .B2(n18396), .C1(
        n18421), .C2(n18395), .ZN(P3_U2726) );
  AOI22_X1 U21547 ( .A1(n18399), .A2(n18398), .B1(n18407), .B2(n18470), .ZN(
        n18402) );
  NAND3_X1 U21548 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18415), .A3(n18400), .ZN(
        n18401) );
  OAI211_X1 U21549 ( .C1(n18424), .C2(n18517), .A(n18402), .B(n18401), .ZN(
        P3_U2727) );
  INV_X1 U21550 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18474) );
  NOR2_X1 U21551 ( .A1(n18404), .A2(n18403), .ZN(n18423) );
  NAND2_X1 U21552 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18418), .ZN(n18408) );
  NOR2_X1 U21553 ( .A1(n18474), .A2(n18408), .ZN(n18411) );
  AOI21_X1 U21554 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18415), .A(n18411), .ZN(
        n18406) );
  OAI222_X1 U21555 ( .A1(n19062), .A2(n18424), .B1(n18407), .B2(n18406), .C1(
        n18421), .C2(n18405), .ZN(P3_U2728) );
  INV_X1 U21556 ( .A(n18408), .ZN(n18414) );
  AOI21_X1 U21557 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18415), .A(n18414), .ZN(
        n18410) );
  OAI222_X1 U21558 ( .A1(n21656), .A2(n18424), .B1(n18411), .B2(n18410), .C1(
        n18421), .C2(n18409), .ZN(P3_U2729) );
  AOI21_X1 U21559 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18415), .A(n18418), .ZN(
        n18413) );
  OAI222_X1 U21560 ( .A1(n19054), .A2(n18424), .B1(n18414), .B2(n18413), .C1(
        n18421), .C2(n18412), .ZN(P3_U2730) );
  AOI21_X1 U21561 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18415), .A(n18423), .ZN(
        n18417) );
  OAI222_X1 U21562 ( .A1(n19050), .A2(n18424), .B1(n18418), .B2(n18417), .C1(
        n18421), .C2(n18416), .ZN(P3_U2731) );
  AOI22_X1 U21563 ( .A1(n18419), .A2(P3_EAX_REG_2__SCAN_IN), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n18415), .ZN(n18422) );
  OAI222_X1 U21564 ( .A1(n19045), .A2(n18424), .B1(n18423), .B2(n18422), .C1(
        n18421), .C2(n18420), .ZN(P3_U2732) );
  INV_X2 U21565 ( .A(n18455), .ZN(n19623) );
  NOR2_X1 U21566 ( .A1(n18477), .A2(n18427), .ZN(P3_U2736) );
  INV_X1 U21567 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n21561) );
  AOI22_X1 U21568 ( .A1(n19623), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18429) );
  OAI21_X1 U21569 ( .B1(n21561), .B2(n18457), .A(n18429), .ZN(P3_U2737) );
  AOI22_X1 U21570 ( .A1(n19623), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18430) );
  OAI21_X1 U21571 ( .B1(n18431), .B2(n18457), .A(n18430), .ZN(P3_U2738) );
  AOI22_X1 U21572 ( .A1(n19623), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18432) );
  OAI21_X1 U21573 ( .B1(n9985), .B2(n18457), .A(n18432), .ZN(P3_U2739) );
  AOI22_X1 U21574 ( .A1(n19623), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18433) );
  OAI21_X1 U21575 ( .B1(n18434), .B2(n18457), .A(n18433), .ZN(P3_U2740) );
  INV_X1 U21576 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U21577 ( .A1(n19623), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18435) );
  OAI21_X1 U21578 ( .B1(n18436), .B2(n18457), .A(n18435), .ZN(P3_U2741) );
  AOI22_X1 U21579 ( .A1(n19623), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18437) );
  OAI21_X1 U21580 ( .B1(n18438), .B2(n18457), .A(n18437), .ZN(P3_U2742) );
  INV_X1 U21581 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18440) );
  AOI22_X1 U21582 ( .A1(n19623), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18439) );
  OAI21_X1 U21583 ( .B1(n18440), .B2(n18457), .A(n18439), .ZN(P3_U2743) );
  INV_X1 U21584 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U21585 ( .A1(n19623), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18441) );
  OAI21_X1 U21586 ( .B1(n18442), .B2(n18457), .A(n18441), .ZN(P3_U2744) );
  AOI22_X1 U21587 ( .A1(n19623), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18443) );
  OAI21_X1 U21588 ( .B1(n18444), .B2(n18457), .A(n18443), .ZN(P3_U2745) );
  AOI22_X1 U21589 ( .A1(n19623), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18445) );
  OAI21_X1 U21590 ( .B1(n18446), .B2(n18457), .A(n18445), .ZN(P3_U2746) );
  AOI22_X1 U21591 ( .A1(n19623), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18447) );
  OAI21_X1 U21592 ( .B1(n18448), .B2(n18457), .A(n18447), .ZN(P3_U2747) );
  AOI22_X1 U21593 ( .A1(n19623), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18449) );
  OAI21_X1 U21594 ( .B1(n18450), .B2(n18457), .A(n18449), .ZN(P3_U2748) );
  AOI22_X1 U21595 ( .A1(n19623), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18451) );
  OAI21_X1 U21596 ( .B1(n18452), .B2(n18457), .A(n18451), .ZN(P3_U2749) );
  INV_X1 U21597 ( .A(P3_UWORD_REG_1__SCAN_IN), .ZN(n21643) );
  INV_X1 U21598 ( .A(n18457), .ZN(n18453) );
  AOI22_X1 U21599 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18453), .B1(n18484), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18454) );
  OAI21_X1 U21600 ( .B1(n18455), .B2(n21643), .A(n18454), .ZN(P3_U2750) );
  INV_X1 U21601 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U21602 ( .A1(n19623), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18456) );
  OAI21_X1 U21603 ( .B1(n18458), .B2(n18457), .A(n18456), .ZN(P3_U2751) );
  AOI22_X1 U21604 ( .A1(n19623), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18459) );
  OAI21_X1 U21605 ( .B1(n18536), .B2(n18486), .A(n18459), .ZN(P3_U2752) );
  AOI22_X1 U21606 ( .A1(n19623), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18460) );
  OAI21_X1 U21607 ( .B1(n18531), .B2(n18486), .A(n18460), .ZN(P3_U2753) );
  INV_X1 U21608 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18462) );
  AOI22_X1 U21609 ( .A1(n19623), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18461) );
  OAI21_X1 U21610 ( .B1(n18462), .B2(n18486), .A(n18461), .ZN(P3_U2754) );
  AOI22_X1 U21611 ( .A1(n19623), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18463) );
  OAI21_X1 U21612 ( .B1(n18464), .B2(n18486), .A(n18463), .ZN(P3_U2755) );
  AOI22_X1 U21613 ( .A1(n19623), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18465) );
  OAI21_X1 U21614 ( .B1(n18523), .B2(n18486), .A(n18465), .ZN(P3_U2756) );
  AOI22_X1 U21615 ( .A1(n19623), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18466) );
  OAI21_X1 U21616 ( .B1(n18467), .B2(n18486), .A(n18466), .ZN(P3_U2757) );
  INV_X1 U21617 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n21565) );
  AOI22_X1 U21618 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18475), .B1(n19623), .B2(
        P3_LWORD_REG_9__SCAN_IN), .ZN(n18468) );
  OAI21_X1 U21619 ( .B1(n21565), .B2(n18477), .A(n18468), .ZN(P3_U2758) );
  AOI22_X1 U21620 ( .A1(n19623), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18469) );
  OAI21_X1 U21621 ( .B1(n18470), .B2(n18486), .A(n18469), .ZN(P3_U2759) );
  INV_X1 U21622 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18472) );
  AOI22_X1 U21623 ( .A1(n19623), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18471) );
  OAI21_X1 U21624 ( .B1(n18472), .B2(n18486), .A(n18471), .ZN(P3_U2760) );
  AOI22_X1 U21625 ( .A1(n19623), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18473) );
  OAI21_X1 U21626 ( .B1(n18474), .B2(n18486), .A(n18473), .ZN(P3_U2761) );
  INV_X1 U21627 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n21723) );
  AOI22_X1 U21628 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18475), .B1(n19623), .B2(
        P3_LWORD_REG_5__SCAN_IN), .ZN(n18476) );
  OAI21_X1 U21629 ( .B1(n21723), .B2(n18477), .A(n18476), .ZN(P3_U2762) );
  INV_X1 U21630 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21552) );
  AOI22_X1 U21631 ( .A1(n19623), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18478) );
  OAI21_X1 U21632 ( .B1(n21552), .B2(n18486), .A(n18478), .ZN(P3_U2763) );
  INV_X1 U21633 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18480) );
  AOI22_X1 U21634 ( .A1(n19623), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18479) );
  OAI21_X1 U21635 ( .B1(n18480), .B2(n18486), .A(n18479), .ZN(P3_U2764) );
  AOI22_X1 U21636 ( .A1(n19623), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18481) );
  OAI21_X1 U21637 ( .B1(n18482), .B2(n18486), .A(n18481), .ZN(P3_U2765) );
  INV_X1 U21638 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U21639 ( .A1(n19623), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18483) );
  OAI21_X1 U21640 ( .B1(n18509), .B2(n18486), .A(n18483), .ZN(P3_U2766) );
  INV_X1 U21641 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U21642 ( .A1(n19623), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18484), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18485) );
  OAI21_X1 U21643 ( .B1(n18487), .B2(n18486), .A(n18485), .ZN(P3_U2767) );
  AOI211_X1 U21644 ( .C1(n18490), .C2(n19529), .A(n18489), .B(n18488), .ZN(
        n18503) );
  INV_X2 U21645 ( .A(n18503), .ZN(n18532) );
  AOI22_X1 U21646 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18532), .ZN(n18491) );
  OAI21_X1 U21647 ( .B1(n19029), .B2(n18528), .A(n18491), .ZN(P3_U2768) );
  INV_X2 U21648 ( .A(n18535), .ZN(n18526) );
  AOI22_X1 U21649 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18533), .B1(
        P3_EAX_REG_17__SCAN_IN), .B2(n18526), .ZN(n18492) );
  OAI21_X1 U21650 ( .B1(n18503), .B2(n21643), .A(n18492), .ZN(P3_U2769) );
  AOI22_X1 U21651 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18532), .ZN(n18493) );
  OAI21_X1 U21652 ( .B1(n19041), .B2(n18528), .A(n18493), .ZN(P3_U2770) );
  AOI22_X1 U21653 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18532), .ZN(n18494) );
  OAI21_X1 U21654 ( .B1(n19045), .B2(n18528), .A(n18494), .ZN(P3_U2771) );
  AOI22_X1 U21655 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18532), .ZN(n18495) );
  OAI21_X1 U21656 ( .B1(n19050), .B2(n18528), .A(n18495), .ZN(P3_U2772) );
  AOI22_X1 U21657 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18532), .ZN(n18496) );
  OAI21_X1 U21658 ( .B1(n19054), .B2(n18528), .A(n18496), .ZN(P3_U2773) );
  AOI22_X1 U21659 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18532), .ZN(n18497) );
  OAI21_X1 U21660 ( .B1(n21656), .B2(n18528), .A(n18497), .ZN(P3_U2774) );
  AOI22_X1 U21661 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18532), .ZN(n18498) );
  OAI21_X1 U21662 ( .B1(n19062), .B2(n18528), .A(n18498), .ZN(P3_U2775) );
  AOI22_X1 U21663 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18532), .ZN(n18499) );
  OAI21_X1 U21664 ( .B1(n18517), .B2(n18528), .A(n18499), .ZN(P3_U2776) );
  AOI22_X1 U21665 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18532), .ZN(n18500) );
  OAI21_X1 U21666 ( .B1(n18519), .B2(n18528), .A(n18500), .ZN(P3_U2777) );
  AOI22_X1 U21667 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18532), .ZN(n18501) );
  OAI21_X1 U21668 ( .B1(n18521), .B2(n18528), .A(n18501), .ZN(P3_U2778) );
  INV_X1 U21669 ( .A(P3_UWORD_REG_11__SCAN_IN), .ZN(n21767) );
  AOI22_X1 U21670 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18533), .B1(
        P3_EAX_REG_27__SCAN_IN), .B2(n18526), .ZN(n18502) );
  OAI21_X1 U21671 ( .B1(n18503), .B2(n21767), .A(n18502), .ZN(P3_U2779) );
  AOI22_X1 U21672 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18532), .ZN(n18504) );
  OAI21_X1 U21673 ( .B1(n18525), .B2(n18528), .A(n18504), .ZN(P3_U2780) );
  AOI22_X1 U21674 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18526), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18532), .ZN(n18505) );
  OAI21_X1 U21675 ( .B1(n18529), .B2(n18528), .A(n18505), .ZN(P3_U2781) );
  AOI22_X1 U21676 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18533), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18532), .ZN(n18506) );
  OAI21_X1 U21677 ( .B1(n21561), .B2(n18535), .A(n18506), .ZN(P3_U2782) );
  AOI22_X1 U21678 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18532), .ZN(n18507) );
  OAI21_X1 U21679 ( .B1(n19029), .B2(n18528), .A(n18507), .ZN(P3_U2783) );
  AOI22_X1 U21680 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18533), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18532), .ZN(n18508) );
  OAI21_X1 U21681 ( .B1(n18509), .B2(n18535), .A(n18508), .ZN(P3_U2784) );
  AOI22_X1 U21682 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18532), .ZN(n18510) );
  OAI21_X1 U21683 ( .B1(n19041), .B2(n18528), .A(n18510), .ZN(P3_U2785) );
  AOI22_X1 U21684 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18532), .ZN(n18511) );
  OAI21_X1 U21685 ( .B1(n19045), .B2(n18528), .A(n18511), .ZN(P3_U2786) );
  AOI22_X1 U21686 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18532), .ZN(n18512) );
  OAI21_X1 U21687 ( .B1(n19050), .B2(n18528), .A(n18512), .ZN(P3_U2787) );
  AOI22_X1 U21688 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18532), .ZN(n18513) );
  OAI21_X1 U21689 ( .B1(n19054), .B2(n18528), .A(n18513), .ZN(P3_U2788) );
  AOI22_X1 U21690 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18532), .ZN(n18514) );
  OAI21_X1 U21691 ( .B1(n21656), .B2(n18528), .A(n18514), .ZN(P3_U2789) );
  AOI22_X1 U21692 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18532), .ZN(n18515) );
  OAI21_X1 U21693 ( .B1(n19062), .B2(n18528), .A(n18515), .ZN(P3_U2790) );
  AOI22_X1 U21694 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18532), .ZN(n18516) );
  OAI21_X1 U21695 ( .B1(n18517), .B2(n18528), .A(n18516), .ZN(P3_U2791) );
  AOI22_X1 U21696 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18532), .ZN(n18518) );
  OAI21_X1 U21697 ( .B1(n18519), .B2(n18528), .A(n18518), .ZN(P3_U2792) );
  AOI22_X1 U21698 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18532), .ZN(n18520) );
  OAI21_X1 U21699 ( .B1(n18521), .B2(n18528), .A(n18520), .ZN(P3_U2793) );
  AOI22_X1 U21700 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18533), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18532), .ZN(n18522) );
  OAI21_X1 U21701 ( .B1(n18523), .B2(n18535), .A(n18522), .ZN(P3_U2794) );
  AOI22_X1 U21702 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18532), .ZN(n18524) );
  OAI21_X1 U21703 ( .B1(n18525), .B2(n18528), .A(n18524), .ZN(P3_U2795) );
  AOI22_X1 U21704 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18526), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18532), .ZN(n18527) );
  OAI21_X1 U21705 ( .B1(n18529), .B2(n18528), .A(n18527), .ZN(P3_U2796) );
  AOI22_X1 U21706 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18533), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18532), .ZN(n18530) );
  OAI21_X1 U21707 ( .B1(n18531), .B2(n18535), .A(n18530), .ZN(P3_U2797) );
  AOI22_X1 U21708 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18533), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18532), .ZN(n18534) );
  OAI21_X1 U21709 ( .B1(n18536), .B2(n18535), .A(n18534), .ZN(P3_U2798) );
  OAI21_X1 U21710 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18538), .A(
        n18537), .ZN(n18819) );
  INV_X1 U21711 ( .A(n18561), .ZN(n18540) );
  AOI22_X1 U21712 ( .A1(n18694), .A2(n18540), .B1(n19409), .B2(n18539), .ZN(
        n18541) );
  OAI211_X1 U21713 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18648), .A(
        n18541), .B(n18772), .ZN(n18553) );
  NOR2_X1 U21714 ( .A1(n18593), .A2(n18539), .ZN(n18554) );
  OAI211_X1 U21715 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18554), .B(n18542), .ZN(n18543) );
  NAND2_X1 U21716 ( .A1(n9696), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18805) );
  OAI211_X1 U21717 ( .C1(n18696), .C2(n18544), .A(n18543), .B(n18805), .ZN(
        n18545) );
  AOI21_X1 U21718 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18553), .A(
        n18545), .ZN(n18550) );
  AOI22_X1 U21719 ( .A1(n9749), .A2(n18798), .B1(n18546), .B2(n9962), .ZN(
        n18816) );
  MUX2_X1 U21720 ( .A(n18547), .B(n18552), .S(n18734), .Z(n18548) );
  XNOR2_X1 U21721 ( .A(n18548), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18815) );
  AOI22_X1 U21722 ( .A1(n18792), .A2(n18816), .B1(n18760), .B2(n18815), .ZN(
        n18549) );
  OAI211_X1 U21723 ( .C1(n18700), .C2(n18819), .A(n18550), .B(n18549), .ZN(
        P3_U2805) );
  NAND2_X1 U21724 ( .A1(n18551), .A2(n18601), .ZN(n18560) );
  NOR2_X1 U21725 ( .A1(n9749), .A2(n18701), .ZN(n18574) );
  AOI21_X1 U21726 ( .B1(n18725), .B2(n18824), .A(n18574), .ZN(n18581) );
  OAI21_X1 U21727 ( .B1(n9814), .B2(n18830), .A(n18552), .ZN(n18829) );
  INV_X1 U21728 ( .A(n18553), .ZN(n18564) );
  AOI22_X1 U21729 ( .A1(n18555), .A2(n18714), .B1(n18554), .B2(n18557), .ZN(
        n18556) );
  NAND2_X1 U21730 ( .A1(n9696), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18832) );
  OAI211_X1 U21731 ( .C1(n18564), .C2(n18557), .A(n18556), .B(n18832), .ZN(
        n18558) );
  AOI21_X1 U21732 ( .B1(n18760), .B2(n18829), .A(n18558), .ZN(n18559) );
  OAI221_X1 U21733 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18560), 
        .C1(n18830), .C2(n18581), .A(n18559), .ZN(P3_U2806) );
  AND2_X1 U21734 ( .A1(n18539), .A2(n19409), .ZN(n18567) );
  INV_X1 U21735 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19579) );
  NOR2_X1 U21736 ( .A1(n10420), .A2(n19579), .ZN(n18836) );
  AOI21_X1 U21737 ( .B1(n18620), .B2(n18561), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18563) );
  OAI22_X1 U21738 ( .A1(n18564), .A2(n18563), .B1(n18696), .B2(n18562), .ZN(
        n18565) );
  AOI211_X1 U21739 ( .C1(n18567), .C2(n18566), .A(n18836), .B(n18565), .ZN(
        n18580) );
  INV_X1 U21740 ( .A(n18568), .ZN(n18571) );
  AOI21_X1 U21741 ( .B1(n18637), .B2(n18569), .A(n18582), .ZN(n18570) );
  AOI211_X1 U21742 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18734), .A(
        n18571), .B(n18570), .ZN(n18572) );
  XNOR2_X1 U21743 ( .A(n18572), .B(n18796), .ZN(n18837) );
  NOR2_X1 U21744 ( .A1(n18588), .A2(n18573), .ZN(n18578) );
  INV_X1 U21745 ( .A(n18574), .ZN(n18576) );
  NAND2_X1 U21746 ( .A1(n18725), .A2(n18824), .ZN(n18575) );
  OAI22_X1 U21747 ( .A1(n17226), .A2(n18576), .B1(n18899), .B2(n18575), .ZN(
        n18577) );
  AOI22_X1 U21748 ( .A1(n18760), .A2(n18837), .B1(n18578), .B2(n18577), .ZN(
        n18579) );
  OAI211_X1 U21749 ( .C1(n18581), .C2(n18796), .A(n18580), .B(n18579), .ZN(
        P3_U2807) );
  INV_X1 U21750 ( .A(n18842), .ZN(n18584) );
  INV_X1 U21751 ( .A(n18582), .ZN(n18583) );
  OAI21_X1 U21752 ( .B1(n18607), .B2(n18584), .A(n18583), .ZN(n18585) );
  NAND2_X1 U21753 ( .A1(n18585), .A2(n18568), .ZN(n18586) );
  XNOR2_X1 U21754 ( .A(n18586), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18859) );
  INV_X1 U21755 ( .A(n18859), .ZN(n18600) );
  NOR2_X1 U21756 ( .A1(n18588), .A2(n18587), .ZN(n18844) );
  INV_X1 U21757 ( .A(n18844), .ZN(n18622) );
  NOR2_X1 U21758 ( .A1(n18843), .A2(n18622), .ZN(n18851) );
  OAI21_X1 U21759 ( .B1(n18623), .B2(n18851), .A(n18658), .ZN(n18612) );
  OAI21_X1 U21760 ( .B1(n18590), .B2(n18648), .A(n18772), .ZN(n18591) );
  AOI21_X1 U21761 ( .B1(n18647), .B2(n18592), .A(n18591), .ZN(n18618) );
  OAI21_X1 U21762 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18615), .A(
        n18618), .ZN(n18604) );
  AOI22_X1 U21763 ( .A1(n9696), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18604), .ZN(n18596) );
  NOR2_X1 U21764 ( .A1(n18593), .A2(n18592), .ZN(n18606) );
  OAI211_X1 U21765 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18606), .B(n18594), .ZN(n18595) );
  OAI211_X1 U21766 ( .C1(n18696), .C2(n11586), .A(n18596), .B(n18595), .ZN(
        n18597) );
  AOI21_X1 U21767 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18612), .A(
        n18597), .ZN(n18599) );
  NAND3_X1 U21768 ( .A1(n18601), .A2(n18851), .A3(n18857), .ZN(n18598) );
  OAI211_X1 U21769 ( .C1(n18748), .C2(n18600), .A(n18599), .B(n18598), .ZN(
        P3_U2808) );
  INV_X1 U21770 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18858) );
  NAND2_X1 U21771 ( .A1(n18867), .A2(n18858), .ZN(n18871) );
  NAND2_X1 U21772 ( .A1(n18601), .A2(n18844), .ZN(n18642) );
  INV_X1 U21773 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18605) );
  OAI22_X1 U21774 ( .A1(n10420), .A2(n19575), .B1(n18696), .B2(n18602), .ZN(
        n18603) );
  AOI221_X1 U21775 ( .B1(n18606), .B2(n18605), .C1(n18604), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18603), .ZN(n18614) );
  INV_X1 U21776 ( .A(n18867), .ZN(n18610) );
  INV_X1 U21777 ( .A(n18607), .ZN(n18608) );
  NAND3_X1 U21778 ( .A1(n18608), .A2(n18703), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18635) );
  OAI22_X1 U21779 ( .A1(n18610), .A2(n18635), .B1(n18637), .B2(n18609), .ZN(
        n18611) );
  XOR2_X1 U21780 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18611), .Z(
        n18865) );
  AOI22_X1 U21781 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18612), .B1(
        n18760), .B2(n18865), .ZN(n18613) );
  OAI211_X1 U21782 ( .C1(n18871), .C2(n18642), .A(n18614), .B(n18613), .ZN(
        P3_U2809) );
  NAND2_X1 U21783 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18853), .ZN(
        n18880) );
  INV_X1 U21784 ( .A(n18615), .ZN(n18620) );
  AOI21_X1 U21785 ( .B1(n18616), .B2(n19409), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18617) );
  OAI22_X1 U21786 ( .A1(n18618), .A2(n18617), .B1(n10420), .B2(n21741), .ZN(
        n18619) );
  AOI221_X1 U21787 ( .B1(n18714), .B2(n18621), .C1(n18620), .C2(n18621), .A(
        n18619), .ZN(n18628) );
  NOR2_X1 U21788 ( .A1(n18887), .A2(n18622), .ZN(n18873) );
  OAI21_X1 U21789 ( .B1(n18623), .B2(n18873), .A(n18658), .ZN(n18639) );
  INV_X1 U21790 ( .A(n18636), .ZN(n18624) );
  OAI21_X1 U21791 ( .B1(n18624), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n18568), .ZN(n18625) );
  AOI21_X1 U21792 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18635), .A(
        n18625), .ZN(n18626) );
  XNOR2_X1 U21793 ( .A(n18626), .B(n18853), .ZN(n18876) );
  AOI22_X1 U21794 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18639), .B1(
        n18760), .B2(n18876), .ZN(n18627) );
  OAI211_X1 U21795 ( .C1(n18642), .C2(n18880), .A(n18628), .B(n18627), .ZN(
        P3_U2810) );
  OAI211_X1 U21796 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18630), .B(n18629), .ZN(n18631) );
  NAND2_X1 U21797 ( .A1(n9696), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18884) );
  OAI211_X1 U21798 ( .C1(n18696), .C2(n18632), .A(n18631), .B(n18884), .ZN(
        n18633) );
  AOI21_X1 U21799 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18634), .A(
        n18633), .ZN(n18641) );
  OAI21_X1 U21800 ( .B1(n18637), .B2(n18636), .A(n18635), .ZN(n18638) );
  XNOR2_X1 U21801 ( .A(n18638), .B(n18887), .ZN(n18883) );
  AOI22_X1 U21802 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18639), .B1(
        n18760), .B2(n18883), .ZN(n18640) );
  OAI211_X1 U21803 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18642), .A(
        n18641), .B(n18640), .ZN(P3_U2811) );
  INV_X1 U21804 ( .A(n18956), .ZN(n18666) );
  NAND2_X1 U21805 ( .A1(n18666), .A2(n18703), .ZN(n18749) );
  OAI22_X1 U21806 ( .A1(n18643), .A2(n18703), .B1(n18749), .B2(n18644), .ZN(
        n18645) );
  XOR2_X1 U21807 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18645), .Z(
        n18896) );
  AOI21_X1 U21808 ( .B1(n18647), .B2(n18646), .A(n17055), .ZN(n18681) );
  OAI21_X1 U21809 ( .B1(n18649), .B2(n18648), .A(n18681), .ZN(n18663) );
  AOI22_X1 U21810 ( .A1(n9696), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18663), .ZN(n18654) );
  NAND2_X1 U21811 ( .A1(n18679), .A2(n18650), .ZN(n18711) );
  NOR2_X1 U21812 ( .A1(n18651), .A2(n18711), .ZN(n18665) );
  OAI211_X1 U21813 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18665), .B(n18652), .ZN(n18653) );
  OAI211_X1 U21814 ( .C1(n18655), .C2(n18696), .A(n18654), .B(n18653), .ZN(
        n18656) );
  AOI21_X1 U21815 ( .B1(n18760), .B2(n18896), .A(n18656), .ZN(n18657) );
  OAI221_X1 U21816 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18659), 
        .C1(n18894), .C2(n18658), .A(n18657), .ZN(P3_U2814) );
  NOR2_X1 U21817 ( .A1(n18956), .A2(n18660), .ZN(n18932) );
  AND3_X1 U21818 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18932), .ZN(n18685) );
  NOR2_X1 U21819 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18685), .ZN(
        n18905) );
  NAND2_X1 U21820 ( .A1(n18725), .A2(n18899), .ZN(n18676) );
  NAND2_X1 U21821 ( .A1(n9696), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18908) );
  OAI21_X1 U21822 ( .B1(n18696), .B2(n18661), .A(n18908), .ZN(n18662) );
  AOI221_X1 U21823 ( .B1(n18665), .B2(n18664), .C1(n18663), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18662), .ZN(n18675) );
  INV_X1 U21824 ( .A(n18715), .ZN(n18943) );
  NAND3_X1 U21825 ( .A1(n18666), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n18943), .ZN(n18668) );
  OAI22_X1 U21826 ( .A1(n18703), .A2(n18947), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18913), .ZN(n18667) );
  AOI21_X1 U21827 ( .B1(n18668), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n18667), .ZN(n18669) );
  OAI21_X1 U21828 ( .B1(n18727), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n18669), .ZN(n18670) );
  XNOR2_X1 U21829 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18670), .ZN(
        n18906) );
  AND2_X1 U21830 ( .A1(n17226), .A2(n18792), .ZN(n18673) );
  OR2_X1 U21831 ( .A1(n18671), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18672) );
  AOI22_X1 U21832 ( .A1(n18760), .A2(n18906), .B1(n18673), .B2(n18672), .ZN(
        n18674) );
  OAI211_X1 U21833 ( .C1(n18905), .C2(n18676), .A(n18675), .B(n18674), .ZN(
        P3_U2815) );
  OAI21_X1 U21834 ( .B1(n18749), .B2(n18917), .A(n18677), .ZN(n18678) );
  XOR2_X1 U21835 ( .A(n18913), .B(n18678), .Z(n18929) );
  AND2_X1 U21836 ( .A1(n18679), .A2(n19409), .ZN(n18723) );
  AOI21_X1 U21837 ( .B1(n18689), .B2(n18723), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18680) );
  OAI22_X1 U21838 ( .A1(n18776), .A2(n18682), .B1(n18681), .B2(n18680), .ZN(
        n18683) );
  AOI21_X1 U21839 ( .B1(n9696), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18683), .ZN(
        n18688) );
  AOI21_X1 U21840 ( .B1(n18684), .B2(n18913), .A(n18671), .ZN(n18924) );
  NAND2_X1 U21841 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18932), .ZN(
        n18686) );
  AOI21_X1 U21842 ( .B1(n18913), .B2(n18686), .A(n18685), .ZN(n18925) );
  AOI22_X1 U21843 ( .A1(n18792), .A2(n18924), .B1(n18725), .B2(n18925), .ZN(
        n18687) );
  OAI211_X1 U21844 ( .C1(n18929), .C2(n18748), .A(n18688), .B(n18687), .ZN(
        P3_U2816) );
  NAND2_X1 U21845 ( .A1(n18911), .A2(n10164), .ZN(n18941) );
  AOI211_X1 U21846 ( .C1(n18710), .C2(n18697), .A(n18689), .B(n18711), .ZN(
        n18699) );
  OAI21_X1 U21847 ( .B1(n10099), .B2(n18691), .A(n18690), .ZN(n18692) );
  AOI21_X1 U21848 ( .B1(n18694), .B2(n18693), .A(n18692), .ZN(n18709) );
  OAI22_X1 U21849 ( .A1(n18709), .A2(n18697), .B1(n18696), .B2(n18695), .ZN(
        n18698) );
  AOI211_X1 U21850 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n9696), .A(n18699), .B(
        n18698), .ZN(n18706) );
  OAI22_X1 U21851 ( .A1(n18934), .A2(n18701), .B1(n18932), .B2(n18700), .ZN(
        n18716) );
  NOR2_X1 U21852 ( .A1(n18703), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18702) );
  OAI22_X1 U21853 ( .A1(n18727), .A2(n18703), .B1(n18932), .B2(n18702), .ZN(
        n18704) );
  XNOR2_X1 U21854 ( .A(n18704), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18930) );
  AOI22_X1 U21855 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18716), .B1(
        n18760), .B2(n18930), .ZN(n18705) );
  OAI211_X1 U21856 ( .C1(n18763), .C2(n18941), .A(n18706), .B(n18705), .ZN(
        P3_U2817) );
  INV_X1 U21857 ( .A(n18749), .ZN(n18707) );
  NAND2_X1 U21858 ( .A1(n18707), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18736) );
  NOR2_X1 U21859 ( .A1(n18970), .A2(n18736), .ZN(n18726) );
  AOI21_X1 U21860 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n18726), .A(
        n18727), .ZN(n18708) );
  XNOR2_X1 U21861 ( .A(n18708), .B(n18947), .ZN(n18954) );
  NAND2_X1 U21862 ( .A1(n9696), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18952) );
  OAI221_X1 U21863 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18711), .C1(
        n18710), .C2(n18709), .A(n18952), .ZN(n18712) );
  AOI21_X1 U21864 ( .B1(n18714), .B2(n18713), .A(n18712), .ZN(n18719) );
  OAI21_X1 U21865 ( .B1(n18715), .B2(n18763), .A(n18947), .ZN(n18717) );
  NAND2_X1 U21866 ( .A1(n18717), .A2(n18716), .ZN(n18718) );
  OAI211_X1 U21867 ( .C1(n18954), .C2(n18748), .A(n18719), .B(n18718), .ZN(
        P3_U2818) );
  NAND2_X1 U21868 ( .A1(n18958), .A2(n10248), .ZN(n18966) );
  NAND2_X1 U21869 ( .A1(n18720), .A2(n18753), .ZN(n18752) );
  NOR2_X1 U21870 ( .A1(n18740), .A2(n18752), .ZN(n18738) );
  AOI21_X1 U21871 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18764), .A(
        n18738), .ZN(n18722) );
  OAI22_X1 U21872 ( .A1(n18723), .A2(n18722), .B1(n18776), .B2(n18721), .ZN(
        n18724) );
  AOI21_X1 U21873 ( .B1(n9696), .B2(P3_REIP_REG_11__SCAN_IN), .A(n18724), .ZN(
        n18733) );
  AOI22_X1 U21874 ( .A1(n13537), .A2(n18792), .B1(n18725), .B2(n18956), .ZN(
        n18762) );
  OAI21_X1 U21875 ( .B1(n18958), .B2(n18763), .A(n18762), .ZN(n18744) );
  INV_X1 U21876 ( .A(n18726), .ZN(n18731) );
  INV_X1 U21877 ( .A(n18727), .ZN(n18730) );
  NAND3_X1 U21878 ( .A1(n18728), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18731), .ZN(n18729) );
  OAI211_X1 U21879 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n18731), .A(
        n18730), .B(n18729), .ZN(n18955) );
  AOI22_X1 U21880 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18744), .B1(
        n18760), .B2(n18955), .ZN(n18732) );
  OAI211_X1 U21881 ( .C1(n18763), .C2(n18966), .A(n18733), .B(n18732), .ZN(
        P3_U2819) );
  INV_X1 U21882 ( .A(n17139), .ZN(n18735) );
  NAND2_X1 U21883 ( .A1(n18735), .A2(n18734), .ZN(n18750) );
  OAI21_X1 U21884 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18750), .A(
        n18736), .ZN(n18737) );
  XNOR2_X1 U21885 ( .A(n18737), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18977) );
  INV_X1 U21886 ( .A(n18764), .ZN(n18739) );
  AOI211_X1 U21887 ( .C1(n18752), .C2(n18740), .A(n18739), .B(n18738), .ZN(
        n18742) );
  NOR2_X1 U21888 ( .A1(n10420), .A2(n19553), .ZN(n18741) );
  AOI211_X1 U21889 ( .C1(n18743), .C2(n18790), .A(n18742), .B(n18741), .ZN(
        n18747) );
  OAI221_X1 U21890 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n18745), .A(n18744), .ZN(
        n18746) );
  OAI211_X1 U21891 ( .C1(n18977), .C2(n18748), .A(n18747), .B(n18746), .ZN(
        P3_U2820) );
  NAND2_X1 U21892 ( .A1(n18750), .A2(n18749), .ZN(n18751) );
  XNOR2_X1 U21893 ( .A(n18751), .B(n18991), .ZN(n18988) );
  NOR2_X1 U21894 ( .A1(n10420), .A2(n21725), .ZN(n18759) );
  INV_X1 U21895 ( .A(n18752), .ZN(n18757) );
  AOI22_X1 U21896 ( .A1(n18754), .A2(n18753), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18764), .ZN(n18756) );
  OAI22_X1 U21897 ( .A1(n18757), .A2(n18756), .B1(n18776), .B2(n18755), .ZN(
        n18758) );
  AOI211_X1 U21898 ( .C1(n18760), .C2(n18988), .A(n18759), .B(n18758), .ZN(
        n18761) );
  OAI221_X1 U21899 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18763), .C1(
        n18991), .C2(n18762), .A(n18761), .ZN(P3_U2821) );
  NAND2_X1 U21900 ( .A1(n18764), .A2(n18765), .ZN(n18781) );
  OAI22_X1 U21901 ( .A1(n18766), .A2(n18786), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18765), .ZN(n18767) );
  AOI21_X1 U21902 ( .B1(n9696), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18767), .ZN(
        n18771) );
  AOI22_X1 U21903 ( .A1(n18792), .A2(n18769), .B1(n18768), .B2(n18790), .ZN(
        n18770) );
  OAI211_X1 U21904 ( .C1(n21610), .C2(n18781), .A(n18771), .B(n18770), .ZN(
        P3_U2824) );
  AOI21_X1 U21905 ( .B1(n18773), .B2(n18772), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18782) );
  OAI22_X1 U21906 ( .A1(n18776), .A2(n18775), .B1(n18786), .B2(n18774), .ZN(
        n18777) );
  AOI211_X1 U21907 ( .C1(n18792), .C2(n18779), .A(n18778), .B(n18777), .ZN(
        n18780) );
  OAI21_X1 U21908 ( .B1(n18782), .B2(n18781), .A(n18780), .ZN(P3_U2825) );
  XNOR2_X1 U21909 ( .A(n18784), .B(n18783), .ZN(n19011) );
  OAI22_X1 U21910 ( .A1(n18786), .A2(n19011), .B1(n18785), .B2(n19313), .ZN(
        n18787) );
  AOI21_X1 U21911 ( .B1(n9696), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18787), .ZN(
        n18794) );
  AOI21_X1 U21912 ( .B1(n19018), .B2(n18789), .A(n18788), .ZN(n19014) );
  AOI22_X1 U21913 ( .A1(n18792), .A2(n19014), .B1(n18791), .B2(n18790), .ZN(
        n18793) );
  OAI211_X1 U21914 ( .C1(n21640), .C2(n18795), .A(n18794), .B(n18793), .ZN(
        P3_U2826) );
  NOR3_X1 U21915 ( .A1(n18797), .A2(n19006), .A3(n18796), .ZN(n18831) );
  AOI22_X1 U21916 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18951), .B1(
        n18798), .B2(n18831), .ZN(n18803) );
  INV_X1 U21917 ( .A(n18799), .ZN(n18800) );
  AOI22_X1 U21918 ( .A1(n18800), .A2(n19002), .B1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n19008), .ZN(n18802) );
  OAI211_X1 U21919 ( .C1(n18804), .C2(n18803), .A(n18802), .B(n18801), .ZN(
        P3_U2836) );
  INV_X1 U21920 ( .A(n18805), .ZN(n18814) );
  INV_X1 U21921 ( .A(n18825), .ZN(n18807) );
  AOI221_X1 U21922 ( .B1(n18808), .B2(n10299), .C1(n18807), .C2(n10299), .A(
        n18806), .ZN(n18812) );
  NAND2_X1 U21923 ( .A1(n18810), .A2(n18809), .ZN(n18811) );
  AOI221_X1 U21924 ( .B1(n18812), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n18811), .C2(n9962), .A(n19006), .ZN(n18813) );
  AOI211_X1 U21925 ( .C1(n19008), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18814), .B(n18813), .ZN(n18818) );
  AOI22_X1 U21926 ( .A1(n19015), .A2(n18816), .B1(n19002), .B2(n18815), .ZN(
        n18817) );
  OAI211_X1 U21927 ( .C1(n18820), .C2(n18819), .A(n18818), .B(n18817), .ZN(
        P3_U2837) );
  OAI22_X1 U21928 ( .A1(n18822), .A2(n18821), .B1(n9749), .B2(n18933), .ZN(
        n18823) );
  AOI211_X1 U21929 ( .C1(n18996), .C2(n18824), .A(n19008), .B(n18823), .ZN(
        n18827) );
  OAI211_X1 U21930 ( .C1(n18825), .C2(n18889), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18827), .ZN(n18826) );
  NAND2_X1 U21931 ( .A1(n10420), .A2(n18826), .ZN(n18839) );
  INV_X1 U21932 ( .A(n18827), .ZN(n18828) );
  OAI21_X1 U21933 ( .B1(n18892), .B2(n18828), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18834) );
  AOI22_X1 U21934 ( .A1(n18831), .A2(n18830), .B1(n19002), .B2(n18829), .ZN(
        n18833) );
  OAI211_X1 U21935 ( .C1(n18839), .C2(n18834), .A(n18833), .B(n18832), .ZN(
        P3_U2838) );
  AOI21_X1 U21936 ( .B1(n18835), .B2(n18998), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18840) );
  AOI21_X1 U21937 ( .B1(n18837), .B2(n19002), .A(n18836), .ZN(n18838) );
  OAI21_X1 U21938 ( .B1(n18840), .B2(n18839), .A(n18838), .ZN(P3_U2839) );
  NOR2_X1 U21939 ( .A1(n18841), .A2(n19006), .ZN(n18864) );
  AOI22_X1 U21940 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18951), .B1(
        n18842), .B2(n18864), .ZN(n18863) );
  INV_X1 U21941 ( .A(n18843), .ZN(n18855) );
  NOR2_X1 U21942 ( .A1(n10151), .A2(n18916), .ZN(n18986) );
  NAND3_X1 U21943 ( .A1(n18888), .A2(n18844), .A3(n18986), .ZN(n18850) );
  AOI21_X1 U21944 ( .B1(n18846), .B2(n18873), .A(n18845), .ZN(n18849) );
  AOI21_X1 U21945 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18847), .A(
        n18889), .ZN(n18848) );
  AOI211_X1 U21946 ( .C1(n18978), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        n18872) );
  OAI21_X1 U21947 ( .B1(n18851), .B2(n18957), .A(n18872), .ZN(n18852) );
  AOI21_X1 U21948 ( .B1(n18981), .B2(n18853), .A(n18852), .ZN(n18866) );
  OAI211_X1 U21949 ( .C1(n18855), .C2(n18910), .A(n18854), .B(n18866), .ZN(
        n18856) );
  AOI211_X1 U21950 ( .C1(n18981), .C2(n18858), .A(n18857), .B(n18856), .ZN(
        n18862) );
  AOI22_X1 U21951 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19008), .B1(
        n19002), .B2(n18859), .ZN(n18861) );
  NAND2_X1 U21952 ( .A1(n9696), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18860) );
  OAI211_X1 U21953 ( .C1(n18863), .C2(n18862), .A(n18861), .B(n18860), .ZN(
        P3_U2840) );
  NAND2_X1 U21954 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18864), .ZN(
        n18881) );
  AOI22_X1 U21955 ( .A1(n9696), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n19002), 
        .B2(n18865), .ZN(n18870) );
  OAI21_X1 U21956 ( .B1(n18867), .B2(n18910), .A(n18866), .ZN(n18868) );
  OAI211_X1 U21957 ( .C1(n18893), .C2(n18868), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n10420), .ZN(n18869) );
  OAI211_X1 U21958 ( .C1(n18881), .C2(n18871), .A(n18870), .B(n18869), .ZN(
        P3_U2841) );
  NAND2_X1 U21959 ( .A1(n18887), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18875) );
  OAI21_X1 U21960 ( .B1(n18873), .B2(n18957), .A(n18872), .ZN(n18874) );
  OAI21_X1 U21961 ( .B1(n18893), .B2(n18874), .A(n10420), .ZN(n18886) );
  OAI21_X1 U21962 ( .B1(n18910), .B2(n18875), .A(n18886), .ZN(n18877) );
  AOI22_X1 U21963 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18877), .B1(
        n19002), .B2(n18876), .ZN(n18879) );
  NAND2_X1 U21964 ( .A1(n9696), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18878) );
  OAI211_X1 U21965 ( .C1(n18880), .C2(n18881), .A(n18879), .B(n18878), .ZN(
        P3_U2842) );
  INV_X1 U21966 ( .A(n18881), .ZN(n18882) );
  AOI22_X1 U21967 ( .A1(n19002), .A2(n18883), .B1(n18882), .B2(n18887), .ZN(
        n18885) );
  OAI211_X1 U21968 ( .C1(n18887), .C2(n18886), .A(n18885), .B(n18884), .ZN(
        P3_U2843) );
  INV_X1 U21969 ( .A(n18968), .ZN(n18937) );
  NAND2_X1 U21970 ( .A1(n18888), .A2(n18986), .ZN(n18890) );
  NOR2_X1 U21971 ( .A1(n18912), .A2(n18889), .ZN(n18979) );
  AOI211_X1 U21972 ( .C1(n18890), .C2(n18978), .A(n13199), .B(n18979), .ZN(
        n18891) );
  NAND2_X1 U21973 ( .A1(n18981), .A2(n18916), .ZN(n18967) );
  OAI211_X1 U21974 ( .C1(n18901), .C2(n18937), .A(n18891), .B(n18967), .ZN(
        n18900) );
  OAI221_X1 U21975 ( .B1(n18893), .B2(n18892), .C1(n18893), .C2(n18900), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18898) );
  AOI22_X1 U21976 ( .A1(n19002), .A2(n18896), .B1(n18895), .B2(n18894), .ZN(
        n18897) );
  OAI221_X1 U21977 ( .B1(n9696), .B2(n18898), .C1(n10420), .C2(n19566), .A(
        n18897), .ZN(P3_U2846) );
  NAND2_X1 U21978 ( .A1(n18996), .A2(n18899), .ZN(n18904) );
  OAI211_X1 U21979 ( .C1(n18671), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n19465), .B(n17226), .ZN(n18903) );
  OAI221_X1 U21980 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18901), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18945), .A(n18900), .ZN(
        n18902) );
  OAI211_X1 U21981 ( .C1(n18905), .C2(n18904), .A(n18903), .B(n18902), .ZN(
        n18907) );
  AOI22_X1 U21982 ( .A1(n18951), .A2(n18907), .B1(n19002), .B2(n18906), .ZN(
        n18909) );
  OAI211_X1 U21983 ( .C1(n18998), .C2(n13199), .A(n18909), .B(n18908), .ZN(
        P3_U2847) );
  NOR2_X1 U21984 ( .A1(n10420), .A2(n19562), .ZN(n18923) );
  INV_X1 U21985 ( .A(n18910), .ZN(n18915) );
  INV_X1 U21986 ( .A(n18917), .ZN(n18918) );
  NAND2_X1 U21987 ( .A1(n18911), .A2(n18986), .ZN(n18942) );
  NAND2_X1 U21988 ( .A1(n18978), .A2(n18942), .ZN(n18936) );
  NAND3_X1 U21989 ( .A1(n18912), .A2(n18918), .A3(n18936), .ZN(n18914) );
  AOI21_X1 U21990 ( .B1(n18915), .B2(n18914), .A(n18913), .ZN(n18921) );
  OAI21_X1 U21991 ( .B1(n18917), .B2(n18916), .A(n18981), .ZN(n18920) );
  AOI21_X1 U21992 ( .B1(n18918), .B2(n18945), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18919) );
  AOI211_X1 U21993 ( .C1(n18921), .C2(n18920), .A(n18919), .B(n19006), .ZN(
        n18922) );
  AOI211_X1 U21994 ( .C1(n19008), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18923), .B(n18922), .ZN(n18928) );
  AOI22_X1 U21995 ( .A1(n18926), .A2(n18925), .B1(n19015), .B2(n18924), .ZN(
        n18927) );
  OAI211_X1 U21996 ( .C1(n18929), .C2(n18976), .A(n18928), .B(n18927), .ZN(
        P3_U2848) );
  AOI22_X1 U21997 ( .A1(n9696), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n19002), 
        .B2(n18930), .ZN(n18940) );
  OAI21_X1 U21998 ( .B1(n18943), .B2(n18937), .A(n18967), .ZN(n18963) );
  OAI22_X1 U21999 ( .A1(n18934), .A2(n18933), .B1(n18932), .B2(n18931), .ZN(
        n18935) );
  NOR3_X1 U22000 ( .A1(n18979), .A2(n18963), .A3(n18935), .ZN(n18949) );
  OAI211_X1 U22001 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18937), .A(
        n18949), .B(n18936), .ZN(n18938) );
  OAI211_X1 U22002 ( .C1(n19006), .C2(n18938), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n10420), .ZN(n18939) );
  OAI211_X1 U22003 ( .C1(n18992), .C2(n18941), .A(n18940), .B(n18939), .ZN(
        P3_U2849) );
  OAI21_X1 U22004 ( .B1(n18947), .B2(n18978), .A(n18942), .ZN(n18948) );
  OAI21_X1 U22005 ( .B1(n18945), .B2(n18944), .A(n18943), .ZN(n18946) );
  AOI22_X1 U22006 ( .A1(n18949), .A2(n18948), .B1(n18947), .B2(n18946), .ZN(
        n18950) );
  AOI22_X1 U22007 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19008), .B1(
        n18951), .B2(n18950), .ZN(n18953) );
  OAI211_X1 U22008 ( .C1(n18954), .C2(n18976), .A(n18953), .B(n18952), .ZN(
        P3_U2850) );
  AOI22_X1 U22009 ( .A1(n9696), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19002), 
        .B2(n18955), .ZN(n18965) );
  AOI21_X1 U22010 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18986), .A(
        n18961), .ZN(n18960) );
  AOI22_X1 U22011 ( .A1(n13537), .A2(n19465), .B1(n18996), .B2(n18956), .ZN(
        n18984) );
  OAI21_X1 U22012 ( .B1(n18958), .B2(n18957), .A(n18984), .ZN(n18959) );
  NOR4_X1 U22013 ( .A1(n18960), .A2(n18979), .A3(n19006), .A4(n18959), .ZN(
        n18972) );
  OAI21_X1 U22014 ( .B1(n18961), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18972), .ZN(n18962) );
  OAI211_X1 U22015 ( .C1(n18963), .C2(n18962), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n10420), .ZN(n18964) );
  OAI211_X1 U22016 ( .C1(n18966), .C2(n18992), .A(n18965), .B(n18964), .ZN(
        P3_U2851) );
  INV_X1 U22017 ( .A(n18967), .ZN(n18969) );
  OAI21_X1 U22018 ( .B1(n18969), .B2(n18991), .A(n18968), .ZN(n18971) );
  AOI21_X1 U22019 ( .B1(n18972), .B2(n18971), .A(n18970), .ZN(n18974) );
  NOR3_X1 U22020 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18991), .A3(
        n18992), .ZN(n18973) );
  AOI221_X1 U22021 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9696), .C1(n18974), 
        .C2(n10420), .A(n18973), .ZN(n18975) );
  OAI21_X1 U22022 ( .B1(n18977), .B2(n18976), .A(n18975), .ZN(P3_U2852) );
  AOI21_X1 U22023 ( .B1(n18981), .B2(n18993), .A(n18978), .ZN(n18985) );
  AOI221_X1 U22024 ( .B1(n18982), .B2(n18981), .C1(n18980), .C2(n18981), .A(
        n18979), .ZN(n18983) );
  OAI211_X1 U22025 ( .C1(n18986), .C2(n18985), .A(n18984), .B(n18983), .ZN(
        n18987) );
  OAI21_X1 U22026 ( .B1(n19006), .B2(n18987), .A(n10420), .ZN(n18990) );
  AOI22_X1 U22027 ( .A1(n9696), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19002), .B2(
        n18988), .ZN(n18989) );
  OAI221_X1 U22028 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18992), .C1(
        n18991), .C2(n18990), .A(n18989), .ZN(P3_U2853) );
  AOI222_X1 U22029 ( .A1(n18997), .A2(n19465), .B1(n18996), .B2(n18995), .C1(
        n18994), .C2(n18993), .ZN(n19007) );
  OAI21_X1 U22030 ( .B1(n19000), .B2(n18999), .A(n18998), .ZN(n19003) );
  AOI22_X1 U22031 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n19001), .ZN(n19005) );
  OAI211_X1 U22032 ( .C1(n19007), .C2(n19006), .A(n19005), .B(n19004), .ZN(
        P3_U2854) );
  AOI21_X1 U22033 ( .B1(n19010), .B2(n19009), .A(n19008), .ZN(n19017) );
  OAI22_X1 U22034 ( .A1(n19012), .A2(n19011), .B1(n19543), .B2(n10420), .ZN(
        n19013) );
  AOI21_X1 U22035 ( .B1(n19015), .B2(n19014), .A(n19013), .ZN(n19016) );
  OAI221_X1 U22036 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19019), .C1(
        n19018), .C2(n19017), .A(n19016), .ZN(P3_U2858) );
  AOI21_X1 U22037 ( .B1(n19022), .B2(n19021), .A(n19020), .ZN(n19504) );
  OAI21_X1 U22038 ( .B1(n19504), .B2(n19069), .A(n19027), .ZN(n19023) );
  OAI221_X1 U22039 ( .B1(n19477), .B2(n19620), .C1(n19477), .C2(n19027), .A(
        n19023), .ZN(P3_U2863) );
  NOR2_X1 U22040 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19028), .ZN(
        n19200) );
  NOR2_X1 U22041 ( .A1(n19244), .A2(n19200), .ZN(n19025) );
  OAI22_X1 U22042 ( .A1(n19026), .A2(n11737), .B1(n19025), .B2(n19024), .ZN(
        P3_U2866) );
  NOR2_X1 U22043 ( .A1(n19494), .A2(n19027), .ZN(P3_U2867) );
  NOR2_X1 U22044 ( .A1(n19028), .A2(n11737), .ZN(n19346) );
  NOR2_X1 U22045 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19477), .ZN(
        n19243) );
  NAND2_X1 U22046 ( .A1(n19346), .A2(n19243), .ZN(n19452) );
  NAND2_X1 U22047 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19409), .ZN(n19379) );
  NOR2_X1 U22048 ( .A1(n11737), .A2(n19175), .ZN(n19407) );
  NAND2_X1 U22049 ( .A1(n19477), .A2(n19407), .ZN(n19080) );
  INV_X1 U22050 ( .A(n19080), .ZN(n19398) );
  NOR2_X2 U22051 ( .A1(n19313), .A2(n19815), .ZN(n19410) );
  NOR2_X2 U22052 ( .A1(n19312), .A2(n19029), .ZN(n19404) );
  NAND2_X1 U22053 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19407), .ZN(
        n19414) );
  INV_X1 U22054 ( .A(n19414), .ZN(n19458) );
  NOR2_X1 U22055 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19483) );
  NAND2_X1 U22056 ( .A1(n19483), .A2(n19487), .ZN(n19130) );
  NOR2_X1 U22057 ( .A1(n19458), .A2(n19123), .ZN(n19091) );
  NOR2_X1 U22058 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19608), .ZN(n19370) );
  NOR2_X1 U22059 ( .A1(n19091), .A2(n19370), .ZN(n19063) );
  AOI22_X1 U22060 ( .A1(n19398), .A2(n19410), .B1(n19404), .B2(n19063), .ZN(
        n19037) );
  NAND2_X1 U22061 ( .A1(n19452), .A2(n19080), .ZN(n19369) );
  AOI21_X1 U22062 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19312), .ZN(n19031) );
  INV_X1 U22063 ( .A(n19091), .ZN(n19030) );
  AOI22_X1 U22064 ( .A1(n19409), .A2(n19369), .B1(n19031), .B2(n19030), .ZN(
        n19066) );
  INV_X1 U22065 ( .A(n19032), .ZN(n19033) );
  NAND2_X1 U22066 ( .A1(n19034), .A2(n19033), .ZN(n19064) );
  NOR2_X1 U22067 ( .A1(n19035), .A2(n19064), .ZN(n19376) );
  AOI22_X1 U22068 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19376), .ZN(n19036) );
  OAI211_X1 U22069 ( .C1(n19452), .C2(n19379), .A(n19037), .B(n19036), .ZN(
        P3_U2868) );
  NAND2_X1 U22070 ( .A1(n19409), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19383) );
  INV_X1 U22071 ( .A(n19452), .ZN(n19456) );
  NAND2_X1 U22072 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19409), .ZN(n19420) );
  AND2_X1 U22073 ( .A1(n19375), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19415) );
  AOI22_X1 U22074 ( .A1(n19456), .A2(n19380), .B1(n19063), .B2(n19415), .ZN(
        n19039) );
  NOR2_X2 U22075 ( .A1(n19626), .A2(n19064), .ZN(n19417) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19417), .ZN(n19038) );
  OAI211_X1 U22077 ( .C1(n19080), .C2(n19383), .A(n19039), .B(n19038), .ZN(
        P3_U2869) );
  NAND2_X1 U22078 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19409), .ZN(n19426) );
  NOR2_X2 U22079 ( .A1(n19313), .A2(n19040), .ZN(n19422) );
  NOR2_X2 U22080 ( .A1(n19312), .A2(n19041), .ZN(n19421) );
  AOI22_X1 U22081 ( .A1(n19398), .A2(n19422), .B1(n19063), .B2(n19421), .ZN(
        n19044) );
  NOR2_X2 U22082 ( .A1(n19042), .A2(n19064), .ZN(n19423) );
  AOI22_X1 U22083 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19423), .ZN(n19043) );
  OAI211_X1 U22084 ( .C1(n19452), .C2(n19426), .A(n19044), .B(n19043), .ZN(
        P3_U2870) );
  NAND2_X1 U22085 ( .A1(n19409), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19299) );
  NOR2_X1 U22086 ( .A1(n21578), .A2(n19313), .ZN(n19296) );
  NOR2_X2 U22087 ( .A1(n19312), .A2(n19045), .ZN(n19427) );
  AOI22_X1 U22088 ( .A1(n19456), .A2(n19296), .B1(n19063), .B2(n19427), .ZN(
        n19048) );
  NOR2_X2 U22089 ( .A1(n19046), .A2(n19064), .ZN(n19429) );
  AOI22_X1 U22090 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19429), .ZN(n19047) );
  OAI211_X1 U22091 ( .C1(n19080), .C2(n19299), .A(n19048), .B(n19047), .ZN(
        P3_U2871) );
  NAND2_X1 U22092 ( .A1(n19409), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19438) );
  NOR2_X1 U22093 ( .A1(n19049), .A2(n19313), .ZN(n19433) );
  NOR2_X2 U22094 ( .A1(n19312), .A2(n19050), .ZN(n19434) );
  AOI22_X1 U22095 ( .A1(n19456), .A2(n19433), .B1(n19063), .B2(n19434), .ZN(
        n19053) );
  NOR2_X2 U22096 ( .A1(n19051), .A2(n19064), .ZN(n19435) );
  AOI22_X1 U22097 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19435), .ZN(n19052) );
  OAI211_X1 U22098 ( .C1(n19080), .C2(n19438), .A(n19053), .B(n19052), .ZN(
        P3_U2872) );
  NAND2_X1 U22099 ( .A1(n19409), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19393) );
  NAND2_X1 U22100 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19409), .ZN(n19444) );
  INV_X1 U22101 ( .A(n19444), .ZN(n19390) );
  NOR2_X2 U22102 ( .A1(n19312), .A2(n19054), .ZN(n19439) );
  AOI22_X1 U22103 ( .A1(n19456), .A2(n19390), .B1(n19063), .B2(n19439), .ZN(
        n19057) );
  NOR2_X2 U22104 ( .A1(n19055), .A2(n19064), .ZN(n19441) );
  AOI22_X1 U22105 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19441), .ZN(n19056) );
  OAI211_X1 U22106 ( .C1(n19080), .C2(n19393), .A(n19057), .B(n19056), .ZN(
        P3_U2873) );
  NAND2_X1 U22107 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19409), .ZN(n19335) );
  NAND2_X1 U22108 ( .A1(n19409), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19451) );
  INV_X1 U22109 ( .A(n19451), .ZN(n19331) );
  NOR2_X2 U22110 ( .A1(n19312), .A2(n21656), .ZN(n19445) );
  AOI22_X1 U22111 ( .A1(n19398), .A2(n19331), .B1(n19063), .B2(n19445), .ZN(
        n19060) );
  NOR2_X2 U22112 ( .A1(n19058), .A2(n19064), .ZN(n19448) );
  AOI22_X1 U22113 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19448), .ZN(n19059) );
  OAI211_X1 U22114 ( .C1(n19452), .C2(n19335), .A(n19060), .B(n19059), .ZN(
        P3_U2874) );
  NOR2_X1 U22115 ( .A1(n19313), .A2(n19061), .ZN(n19338) );
  NOR2_X2 U22116 ( .A1(n19312), .A2(n19062), .ZN(n19454) );
  AOI22_X1 U22117 ( .A1(n19456), .A2(n19338), .B1(n19063), .B2(n19454), .ZN(
        n19068) );
  NOR2_X2 U22118 ( .A1(n19065), .A2(n19064), .ZN(n19457) );
  AOI22_X1 U22119 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19066), .B1(
        n19123), .B2(n19457), .ZN(n19067) );
  OAI211_X1 U22120 ( .C1(n19080), .C2(n19342), .A(n19068), .B(n19067), .ZN(
        P3_U2875) );
  NAND2_X1 U22121 ( .A1(n19487), .A2(n19243), .ZN(n19152) );
  INV_X1 U22122 ( .A(n19379), .ZN(n19405) );
  INV_X1 U22123 ( .A(n19487), .ZN(n19089) );
  INV_X1 U22124 ( .A(n19370), .ZN(n19403) );
  NAND2_X1 U22125 ( .A1(n19478), .A2(n19403), .ZN(n19343) );
  NOR2_X1 U22126 ( .A1(n19089), .A2(n19343), .ZN(n19085) );
  AOI22_X1 U22127 ( .A1(n19405), .A2(n19398), .B1(n19404), .B2(n19085), .ZN(
        n19071) );
  NOR2_X1 U22128 ( .A1(n19312), .A2(n19069), .ZN(n19406) );
  AOI22_X1 U22129 ( .A1(n19409), .A2(n19407), .B1(n19487), .B2(n19345), .ZN(
        n19086) );
  AOI22_X1 U22130 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19086), .B1(
        n19458), .B2(n19410), .ZN(n19070) );
  OAI211_X1 U22131 ( .C1(n19413), .C2(n19152), .A(n19071), .B(n19070), .ZN(
        P3_U2876) );
  AOI22_X1 U22132 ( .A1(n19398), .A2(n19380), .B1(n19415), .B2(n19085), .ZN(
        n19073) );
  INV_X1 U22133 ( .A(n19152), .ZN(n19145) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19086), .B1(
        n19417), .B2(n19145), .ZN(n19072) );
  OAI211_X1 U22135 ( .C1(n19414), .C2(n19383), .A(n19073), .B(n19072), .ZN(
        P3_U2877) );
  AOI22_X1 U22136 ( .A1(n19458), .A2(n19422), .B1(n19421), .B2(n19085), .ZN(
        n19075) );
  AOI22_X1 U22137 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19086), .B1(
        n19423), .B2(n19145), .ZN(n19074) );
  OAI211_X1 U22138 ( .C1(n19080), .C2(n19426), .A(n19075), .B(n19074), .ZN(
        P3_U2878) );
  AOI22_X1 U22139 ( .A1(n19398), .A2(n19296), .B1(n19427), .B2(n19085), .ZN(
        n19077) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19086), .B1(
        n19429), .B2(n19145), .ZN(n19076) );
  OAI211_X1 U22141 ( .C1(n19414), .C2(n19299), .A(n19077), .B(n19076), .ZN(
        P3_U2879) );
  INV_X1 U22142 ( .A(n19438), .ZN(n19325) );
  AOI22_X1 U22143 ( .A1(n19458), .A2(n19325), .B1(n19434), .B2(n19085), .ZN(
        n19079) );
  AOI22_X1 U22144 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19086), .B1(
        n19435), .B2(n19145), .ZN(n19078) );
  OAI211_X1 U22145 ( .C1(n19080), .C2(n19328), .A(n19079), .B(n19078), .ZN(
        P3_U2880) );
  AOI22_X1 U22146 ( .A1(n19398), .A2(n19390), .B1(n19439), .B2(n19085), .ZN(
        n19082) );
  AOI22_X1 U22147 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19086), .B1(
        n19441), .B2(n19145), .ZN(n19081) );
  OAI211_X1 U22148 ( .C1(n19414), .C2(n19393), .A(n19082), .B(n19081), .ZN(
        P3_U2881) );
  INV_X1 U22149 ( .A(n19335), .ZN(n19447) );
  AOI22_X1 U22150 ( .A1(n19398), .A2(n19447), .B1(n19445), .B2(n19085), .ZN(
        n19084) );
  AOI22_X1 U22151 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19086), .B1(
        n19448), .B2(n19145), .ZN(n19083) );
  OAI211_X1 U22152 ( .C1(n19414), .C2(n19451), .A(n19084), .B(n19083), .ZN(
        P3_U2882) );
  AOI22_X1 U22153 ( .A1(n19398), .A2(n19338), .B1(n19454), .B2(n19085), .ZN(
        n19088) );
  AOI22_X1 U22154 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19086), .B1(
        n19457), .B2(n19145), .ZN(n19087) );
  OAI211_X1 U22155 ( .C1(n19414), .C2(n19342), .A(n19088), .B(n19087), .ZN(
        P3_U2883) );
  NAND2_X1 U22156 ( .A1(n19477), .A2(n19154), .ZN(n19174) );
  INV_X1 U22157 ( .A(n19174), .ZN(n19167) );
  NOR2_X1 U22158 ( .A1(n19145), .A2(n19167), .ZN(n19131) );
  NOR2_X1 U22159 ( .A1(n19370), .A2(n19131), .ZN(n19107) );
  AOI22_X1 U22160 ( .A1(n19123), .A2(n19410), .B1(n19404), .B2(n19107), .ZN(
        n19094) );
  INV_X1 U22161 ( .A(n19090), .ZN(n19372) );
  OAI21_X1 U22162 ( .B1(n19091), .B2(n19372), .A(n19131), .ZN(n19092) );
  OAI211_X1 U22163 ( .C1(n19167), .C2(n19608), .A(n19375), .B(n19092), .ZN(
        n19108) );
  AOI22_X1 U22164 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19108), .B1(
        n19376), .B2(n19167), .ZN(n19093) );
  OAI211_X1 U22165 ( .C1(n19379), .C2(n19414), .A(n19094), .B(n19093), .ZN(
        P3_U2884) );
  INV_X1 U22166 ( .A(n19383), .ZN(n19416) );
  AOI22_X1 U22167 ( .A1(n19123), .A2(n19416), .B1(n19415), .B2(n19107), .ZN(
        n19096) );
  AOI22_X1 U22168 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19108), .B1(
        n19417), .B2(n19167), .ZN(n19095) );
  OAI211_X1 U22169 ( .C1(n19414), .C2(n19420), .A(n19096), .B(n19095), .ZN(
        P3_U2885) );
  AOI22_X1 U22170 ( .A1(n19123), .A2(n19422), .B1(n19421), .B2(n19107), .ZN(
        n19098) );
  AOI22_X1 U22171 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19108), .B1(
        n19423), .B2(n19167), .ZN(n19097) );
  OAI211_X1 U22172 ( .C1(n19414), .C2(n19426), .A(n19098), .B(n19097), .ZN(
        P3_U2886) );
  INV_X1 U22173 ( .A(n19299), .ZN(n19428) );
  AOI22_X1 U22174 ( .A1(n19123), .A2(n19428), .B1(n19427), .B2(n19107), .ZN(
        n19100) );
  AOI22_X1 U22175 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19108), .B1(
        n19429), .B2(n19167), .ZN(n19099) );
  OAI211_X1 U22176 ( .C1(n19414), .C2(n19432), .A(n19100), .B(n19099), .ZN(
        P3_U2887) );
  AOI22_X1 U22177 ( .A1(n19458), .A2(n19433), .B1(n19434), .B2(n19107), .ZN(
        n19102) );
  AOI22_X1 U22178 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19108), .B1(
        n19435), .B2(n19167), .ZN(n19101) );
  OAI211_X1 U22179 ( .C1(n19130), .C2(n19438), .A(n19102), .B(n19101), .ZN(
        P3_U2888) );
  INV_X1 U22180 ( .A(n19393), .ZN(n19440) );
  AOI22_X1 U22181 ( .A1(n19123), .A2(n19440), .B1(n19439), .B2(n19107), .ZN(
        n19104) );
  AOI22_X1 U22182 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19108), .B1(
        n19441), .B2(n19167), .ZN(n19103) );
  OAI211_X1 U22183 ( .C1(n19414), .C2(n19444), .A(n19104), .B(n19103), .ZN(
        P3_U2889) );
  AOI22_X1 U22184 ( .A1(n19123), .A2(n19331), .B1(n19445), .B2(n19107), .ZN(
        n19106) );
  AOI22_X1 U22185 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19108), .B1(
        n19448), .B2(n19167), .ZN(n19105) );
  OAI211_X1 U22186 ( .C1(n19414), .C2(n19335), .A(n19106), .B(n19105), .ZN(
        P3_U2890) );
  INV_X1 U22187 ( .A(n19338), .ZN(n19463) );
  AOI22_X1 U22188 ( .A1(n19123), .A2(n19455), .B1(n19454), .B2(n19107), .ZN(
        n19110) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19108), .B1(
        n19457), .B2(n19167), .ZN(n19109) );
  OAI211_X1 U22190 ( .C1(n19414), .C2(n19463), .A(n19110), .B(n19109), .ZN(
        P3_U2891) );
  NAND2_X1 U22191 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19154), .ZN(
        n19188) );
  INV_X1 U22192 ( .A(n19188), .ZN(n19194) );
  AOI21_X1 U22193 ( .B1(n19478), .B2(n19372), .A(n19312), .ZN(n19199) );
  OAI211_X1 U22194 ( .C1(n19194), .C2(n19608), .A(n19487), .B(n19199), .ZN(
        n19127) );
  AND2_X1 U22195 ( .A1(n19403), .A2(n19154), .ZN(n19126) );
  AOI22_X1 U22196 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19127), .B1(
        n19404), .B2(n19126), .ZN(n19112) );
  AOI22_X1 U22197 ( .A1(n19376), .A2(n19194), .B1(n19410), .B2(n19145), .ZN(
        n19111) );
  OAI211_X1 U22198 ( .C1(n19379), .C2(n19130), .A(n19112), .B(n19111), .ZN(
        P3_U2892) );
  AOI22_X1 U22199 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19127), .B1(
        n19415), .B2(n19126), .ZN(n19114) );
  AOI22_X1 U22200 ( .A1(n19416), .A2(n19145), .B1(n19417), .B2(n19194), .ZN(
        n19113) );
  OAI211_X1 U22201 ( .C1(n19130), .C2(n19420), .A(n19114), .B(n19113), .ZN(
        P3_U2893) );
  INV_X1 U22202 ( .A(n19422), .ZN(n19355) );
  INV_X1 U22203 ( .A(n19426), .ZN(n19352) );
  AOI22_X1 U22204 ( .A1(n19123), .A2(n19352), .B1(n19421), .B2(n19126), .ZN(
        n19116) );
  AOI22_X1 U22205 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19127), .B1(
        n19423), .B2(n19194), .ZN(n19115) );
  OAI211_X1 U22206 ( .C1(n19355), .C2(n19152), .A(n19116), .B(n19115), .ZN(
        P3_U2894) );
  AOI22_X1 U22207 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19127), .B1(
        n19427), .B2(n19126), .ZN(n19118) );
  AOI22_X1 U22208 ( .A1(n19123), .A2(n19296), .B1(n19429), .B2(n19194), .ZN(
        n19117) );
  OAI211_X1 U22209 ( .C1(n19299), .C2(n19152), .A(n19118), .B(n19117), .ZN(
        P3_U2895) );
  AOI22_X1 U22210 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19127), .B1(
        n19434), .B2(n19126), .ZN(n19120) );
  AOI22_X1 U22211 ( .A1(n19325), .A2(n19145), .B1(n19435), .B2(n19194), .ZN(
        n19119) );
  OAI211_X1 U22212 ( .C1(n19130), .C2(n19328), .A(n19120), .B(n19119), .ZN(
        P3_U2896) );
  AOI22_X1 U22213 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19127), .B1(
        n19439), .B2(n19126), .ZN(n19122) );
  AOI22_X1 U22214 ( .A1(n19440), .A2(n19145), .B1(n19441), .B2(n19194), .ZN(
        n19121) );
  OAI211_X1 U22215 ( .C1(n19130), .C2(n19444), .A(n19122), .B(n19121), .ZN(
        P3_U2897) );
  AOI22_X1 U22216 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19127), .B1(
        n19445), .B2(n19126), .ZN(n19125) );
  AOI22_X1 U22217 ( .A1(n19123), .A2(n19447), .B1(n19448), .B2(n19194), .ZN(
        n19124) );
  OAI211_X1 U22218 ( .C1(n19451), .C2(n19152), .A(n19125), .B(n19124), .ZN(
        P3_U2898) );
  AOI22_X1 U22219 ( .A1(n19455), .A2(n19145), .B1(n19454), .B2(n19126), .ZN(
        n19129) );
  AOI22_X1 U22220 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19127), .B1(
        n19457), .B2(n19194), .ZN(n19128) );
  OAI211_X1 U22221 ( .C1(n19130), .C2(n19463), .A(n19129), .B(n19128), .ZN(
        P3_U2899) );
  NAND2_X1 U22222 ( .A1(n19483), .A2(n19200), .ZN(n19215) );
  NOR2_X1 U22223 ( .A1(n19194), .A2(n19218), .ZN(n19176) );
  NOR2_X1 U22224 ( .A1(n19370), .A2(n19176), .ZN(n19148) );
  AOI22_X1 U22225 ( .A1(n19410), .A2(n19167), .B1(n19404), .B2(n19148), .ZN(
        n19134) );
  OAI22_X1 U22226 ( .A1(n19131), .A2(n19313), .B1(n19176), .B2(n19312), .ZN(
        n19132) );
  OAI21_X1 U22227 ( .B1(n19218), .B2(n19608), .A(n19132), .ZN(n19149) );
  AOI22_X1 U22228 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19149), .B1(
        n19405), .B2(n19145), .ZN(n19133) );
  OAI211_X1 U22229 ( .C1(n19413), .C2(n19215), .A(n19134), .B(n19133), .ZN(
        P3_U2900) );
  AOI22_X1 U22230 ( .A1(n19416), .A2(n19167), .B1(n19415), .B2(n19148), .ZN(
        n19136) );
  AOI22_X1 U22231 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19149), .B1(
        n19417), .B2(n19218), .ZN(n19135) );
  OAI211_X1 U22232 ( .C1(n19420), .C2(n19152), .A(n19136), .B(n19135), .ZN(
        P3_U2901) );
  AOI22_X1 U22233 ( .A1(n19421), .A2(n19148), .B1(n19422), .B2(n19167), .ZN(
        n19138) );
  AOI22_X1 U22234 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19149), .B1(
        n19423), .B2(n19218), .ZN(n19137) );
  OAI211_X1 U22235 ( .C1(n19426), .C2(n19152), .A(n19138), .B(n19137), .ZN(
        P3_U2902) );
  AOI22_X1 U22236 ( .A1(n19428), .A2(n19167), .B1(n19427), .B2(n19148), .ZN(
        n19140) );
  AOI22_X1 U22237 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19149), .B1(
        n19429), .B2(n19218), .ZN(n19139) );
  OAI211_X1 U22238 ( .C1(n19432), .C2(n19152), .A(n19140), .B(n19139), .ZN(
        P3_U2903) );
  AOI22_X1 U22239 ( .A1(n19325), .A2(n19167), .B1(n19434), .B2(n19148), .ZN(
        n19142) );
  AOI22_X1 U22240 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19149), .B1(
        n19435), .B2(n19218), .ZN(n19141) );
  OAI211_X1 U22241 ( .C1(n19328), .C2(n19152), .A(n19142), .B(n19141), .ZN(
        P3_U2904) );
  AOI22_X1 U22242 ( .A1(n19440), .A2(n19167), .B1(n19439), .B2(n19148), .ZN(
        n19144) );
  AOI22_X1 U22243 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19149), .B1(
        n19441), .B2(n19218), .ZN(n19143) );
  OAI211_X1 U22244 ( .C1(n19444), .C2(n19152), .A(n19144), .B(n19143), .ZN(
        P3_U2905) );
  AOI22_X1 U22245 ( .A1(n19447), .A2(n19145), .B1(n19445), .B2(n19148), .ZN(
        n19147) );
  AOI22_X1 U22246 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19149), .B1(
        n19448), .B2(n19218), .ZN(n19146) );
  OAI211_X1 U22247 ( .C1(n19451), .C2(n19174), .A(n19147), .B(n19146), .ZN(
        P3_U2906) );
  AOI22_X1 U22248 ( .A1(n19455), .A2(n19167), .B1(n19454), .B2(n19148), .ZN(
        n19151) );
  AOI22_X1 U22249 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19149), .B1(
        n19457), .B2(n19218), .ZN(n19150) );
  OAI211_X1 U22250 ( .C1(n19463), .C2(n19152), .A(n19151), .B(n19150), .ZN(
        P3_U2907) );
  NAND2_X1 U22251 ( .A1(n19200), .A2(n19243), .ZN(n19231) );
  INV_X1 U22252 ( .A(n19200), .ZN(n19153) );
  NOR2_X1 U22253 ( .A1(n19153), .A2(n19343), .ZN(n19170) );
  AOI22_X1 U22254 ( .A1(n19410), .A2(n19194), .B1(n19404), .B2(n19170), .ZN(
        n19156) );
  AOI22_X1 U22255 ( .A1(n19409), .A2(n19154), .B1(n19200), .B2(n19345), .ZN(
        n19171) );
  AOI22_X1 U22256 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19171), .B1(
        n19405), .B2(n19167), .ZN(n19155) );
  OAI211_X1 U22257 ( .C1(n19413), .C2(n19231), .A(n19156), .B(n19155), .ZN(
        P3_U2908) );
  INV_X1 U22258 ( .A(n19417), .ZN(n19320) );
  AOI22_X1 U22259 ( .A1(n19415), .A2(n19170), .B1(n19380), .B2(n19167), .ZN(
        n19158) );
  AOI22_X1 U22260 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19171), .B1(
        n19416), .B2(n19194), .ZN(n19157) );
  OAI211_X1 U22261 ( .C1(n19320), .C2(n19231), .A(n19158), .B(n19157), .ZN(
        P3_U2909) );
  AOI22_X1 U22262 ( .A1(n19421), .A2(n19170), .B1(n19422), .B2(n19194), .ZN(
        n19160) );
  AOI22_X1 U22263 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19171), .B1(
        n19423), .B2(n19239), .ZN(n19159) );
  OAI211_X1 U22264 ( .C1(n19426), .C2(n19174), .A(n19160), .B(n19159), .ZN(
        P3_U2910) );
  AOI22_X1 U22265 ( .A1(n19296), .A2(n19167), .B1(n19427), .B2(n19170), .ZN(
        n19162) );
  AOI22_X1 U22266 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19171), .B1(
        n19429), .B2(n19239), .ZN(n19161) );
  OAI211_X1 U22267 ( .C1(n19299), .C2(n19188), .A(n19162), .B(n19161), .ZN(
        P3_U2911) );
  AOI22_X1 U22268 ( .A1(n19325), .A2(n19194), .B1(n19434), .B2(n19170), .ZN(
        n19164) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19171), .B1(
        n19435), .B2(n19239), .ZN(n19163) );
  OAI211_X1 U22270 ( .C1(n19328), .C2(n19174), .A(n19164), .B(n19163), .ZN(
        P3_U2912) );
  AOI22_X1 U22271 ( .A1(n19390), .A2(n19167), .B1(n19439), .B2(n19170), .ZN(
        n19166) );
  AOI22_X1 U22272 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19171), .B1(
        n19441), .B2(n19239), .ZN(n19165) );
  OAI211_X1 U22273 ( .C1(n19393), .C2(n19188), .A(n19166), .B(n19165), .ZN(
        P3_U2913) );
  AOI22_X1 U22274 ( .A1(n19447), .A2(n19167), .B1(n19445), .B2(n19170), .ZN(
        n19169) );
  AOI22_X1 U22275 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19171), .B1(
        n19448), .B2(n19239), .ZN(n19168) );
  OAI211_X1 U22276 ( .C1(n19451), .C2(n19188), .A(n19169), .B(n19168), .ZN(
        P3_U2914) );
  AOI22_X1 U22277 ( .A1(n19455), .A2(n19194), .B1(n19454), .B2(n19170), .ZN(
        n19173) );
  AOI22_X1 U22278 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19171), .B1(
        n19457), .B2(n19239), .ZN(n19172) );
  OAI211_X1 U22279 ( .C1(n19463), .C2(n19174), .A(n19173), .B(n19172), .ZN(
        P3_U2915) );
  NOR2_X2 U22280 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19198), .ZN(
        n19261) );
  NOR2_X1 U22281 ( .A1(n19239), .A2(n19261), .ZN(n19221) );
  NOR2_X1 U22282 ( .A1(n19370), .A2(n19221), .ZN(n19193) );
  AOI22_X1 U22283 ( .A1(n19410), .A2(n19218), .B1(n19404), .B2(n19193), .ZN(
        n19179) );
  OAI22_X1 U22284 ( .A1(n19176), .A2(n19313), .B1(n19221), .B2(n19312), .ZN(
        n19177) );
  OAI21_X1 U22285 ( .B1(n19261), .B2(n19608), .A(n19177), .ZN(n19195) );
  AOI22_X1 U22286 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19195), .B1(
        n19376), .B2(n19261), .ZN(n19178) );
  OAI211_X1 U22287 ( .C1(n19379), .C2(n19188), .A(n19179), .B(n19178), .ZN(
        P3_U2916) );
  AOI22_X1 U22288 ( .A1(n19416), .A2(n19218), .B1(n19415), .B2(n19193), .ZN(
        n19181) );
  AOI22_X1 U22289 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19195), .B1(
        n19417), .B2(n19261), .ZN(n19180) );
  OAI211_X1 U22290 ( .C1(n19420), .C2(n19188), .A(n19181), .B(n19180), .ZN(
        P3_U2917) );
  AOI22_X1 U22291 ( .A1(n19421), .A2(n19193), .B1(n19422), .B2(n19218), .ZN(
        n19183) );
  AOI22_X1 U22292 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19195), .B1(
        n19423), .B2(n19261), .ZN(n19182) );
  OAI211_X1 U22293 ( .C1(n19426), .C2(n19188), .A(n19183), .B(n19182), .ZN(
        P3_U2918) );
  AOI22_X1 U22294 ( .A1(n19296), .A2(n19194), .B1(n19427), .B2(n19193), .ZN(
        n19185) );
  AOI22_X1 U22295 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19195), .B1(
        n19429), .B2(n19261), .ZN(n19184) );
  OAI211_X1 U22296 ( .C1(n19299), .C2(n19215), .A(n19185), .B(n19184), .ZN(
        P3_U2919) );
  AOI22_X1 U22297 ( .A1(n19325), .A2(n19218), .B1(n19434), .B2(n19193), .ZN(
        n19187) );
  AOI22_X1 U22298 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19195), .B1(
        n19435), .B2(n19261), .ZN(n19186) );
  OAI211_X1 U22299 ( .C1(n19328), .C2(n19188), .A(n19187), .B(n19186), .ZN(
        P3_U2920) );
  AOI22_X1 U22300 ( .A1(n19390), .A2(n19194), .B1(n19439), .B2(n19193), .ZN(
        n19190) );
  AOI22_X1 U22301 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19195), .B1(
        n19441), .B2(n19261), .ZN(n19189) );
  OAI211_X1 U22302 ( .C1(n19393), .C2(n19215), .A(n19190), .B(n19189), .ZN(
        P3_U2921) );
  AOI22_X1 U22303 ( .A1(n19447), .A2(n19194), .B1(n19445), .B2(n19193), .ZN(
        n19192) );
  AOI22_X1 U22304 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19195), .B1(
        n19448), .B2(n19261), .ZN(n19191) );
  OAI211_X1 U22305 ( .C1(n19451), .C2(n19215), .A(n19192), .B(n19191), .ZN(
        P3_U2922) );
  AOI22_X1 U22306 ( .A1(n19338), .A2(n19194), .B1(n19454), .B2(n19193), .ZN(
        n19197) );
  AOI22_X1 U22307 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19195), .B1(
        n19457), .B2(n19261), .ZN(n19196) );
  OAI211_X1 U22308 ( .C1(n19342), .C2(n19215), .A(n19197), .B(n19196), .ZN(
        P3_U2923) );
  NOR2_X1 U22309 ( .A1(n19370), .A2(n19198), .ZN(n19216) );
  AOI22_X1 U22310 ( .A1(n19405), .A2(n19218), .B1(n19404), .B2(n19216), .ZN(
        n19202) );
  INV_X1 U22311 ( .A(n19282), .ZN(n19284) );
  OAI211_X1 U22312 ( .C1(n19284), .C2(n19608), .A(n19200), .B(n19199), .ZN(
        n19217) );
  AOI22_X1 U22313 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19217), .B1(
        n19410), .B2(n19239), .ZN(n19201) );
  OAI211_X1 U22314 ( .C1(n19413), .C2(n19282), .A(n19202), .B(n19201), .ZN(
        P3_U2924) );
  AOI22_X1 U22315 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19217), .B1(
        n19415), .B2(n19216), .ZN(n19204) );
  AOI22_X1 U22316 ( .A1(n19417), .A2(n19284), .B1(n19380), .B2(n19218), .ZN(
        n19203) );
  OAI211_X1 U22317 ( .C1(n19383), .C2(n19231), .A(n19204), .B(n19203), .ZN(
        P3_U2925) );
  AOI22_X1 U22318 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19217), .B1(
        n19421), .B2(n19216), .ZN(n19206) );
  AOI22_X1 U22319 ( .A1(n19423), .A2(n19284), .B1(n19422), .B2(n19239), .ZN(
        n19205) );
  OAI211_X1 U22320 ( .C1(n19426), .C2(n19215), .A(n19206), .B(n19205), .ZN(
        P3_U2926) );
  AOI22_X1 U22321 ( .A1(n19428), .A2(n19239), .B1(n19427), .B2(n19216), .ZN(
        n19208) );
  AOI22_X1 U22322 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19217), .B1(
        n19429), .B2(n19284), .ZN(n19207) );
  OAI211_X1 U22323 ( .C1(n19432), .C2(n19215), .A(n19208), .B(n19207), .ZN(
        P3_U2927) );
  AOI22_X1 U22324 ( .A1(n19325), .A2(n19239), .B1(n19434), .B2(n19216), .ZN(
        n19210) );
  AOI22_X1 U22325 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19217), .B1(
        n19435), .B2(n19284), .ZN(n19209) );
  OAI211_X1 U22326 ( .C1(n19328), .C2(n19215), .A(n19210), .B(n19209), .ZN(
        P3_U2928) );
  AOI22_X1 U22327 ( .A1(n19440), .A2(n19239), .B1(n19439), .B2(n19216), .ZN(
        n19212) );
  AOI22_X1 U22328 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19217), .B1(
        n19441), .B2(n19284), .ZN(n19211) );
  OAI211_X1 U22329 ( .C1(n19444), .C2(n19215), .A(n19212), .B(n19211), .ZN(
        P3_U2929) );
  AOI22_X1 U22330 ( .A1(n19445), .A2(n19216), .B1(n19331), .B2(n19239), .ZN(
        n19214) );
  AOI22_X1 U22331 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19217), .B1(
        n19448), .B2(n19284), .ZN(n19213) );
  OAI211_X1 U22332 ( .C1(n19335), .C2(n19215), .A(n19214), .B(n19213), .ZN(
        P3_U2930) );
  AOI22_X1 U22333 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19217), .B1(
        n19454), .B2(n19216), .ZN(n19220) );
  AOI22_X1 U22334 ( .A1(n19457), .A2(n19284), .B1(n19338), .B2(n19218), .ZN(
        n19219) );
  OAI211_X1 U22335 ( .C1(n19342), .C2(n19231), .A(n19220), .B(n19219), .ZN(
        P3_U2931) );
  NAND2_X1 U22336 ( .A1(n19483), .A2(n19244), .ZN(n19304) );
  NOR2_X1 U22337 ( .A1(n19284), .A2(n19308), .ZN(n19266) );
  NOR2_X1 U22338 ( .A1(n19370), .A2(n19266), .ZN(n19238) );
  AOI22_X1 U22339 ( .A1(n19405), .A2(n19239), .B1(n19404), .B2(n19238), .ZN(
        n19224) );
  OAI21_X1 U22340 ( .B1(n19221), .B2(n19372), .A(n19266), .ZN(n19222) );
  OAI211_X1 U22341 ( .C1(n19308), .C2(n19608), .A(n19375), .B(n19222), .ZN(
        n19240) );
  AOI22_X1 U22342 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19240), .B1(
        n19410), .B2(n19261), .ZN(n19223) );
  OAI211_X1 U22343 ( .C1(n19413), .C2(n19304), .A(n19224), .B(n19223), .ZN(
        P3_U2932) );
  AOI22_X1 U22344 ( .A1(n19415), .A2(n19238), .B1(n19380), .B2(n19239), .ZN(
        n19226) );
  AOI22_X1 U22345 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19240), .B1(
        n19416), .B2(n19261), .ZN(n19225) );
  OAI211_X1 U22346 ( .C1(n19320), .C2(n19304), .A(n19226), .B(n19225), .ZN(
        P3_U2933) );
  INV_X1 U22347 ( .A(n19261), .ZN(n19254) );
  AOI22_X1 U22348 ( .A1(n19352), .A2(n19239), .B1(n19421), .B2(n19238), .ZN(
        n19228) );
  AOI22_X1 U22349 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19240), .B1(
        n19423), .B2(n19308), .ZN(n19227) );
  OAI211_X1 U22350 ( .C1(n19355), .C2(n19254), .A(n19228), .B(n19227), .ZN(
        P3_U2934) );
  AOI22_X1 U22351 ( .A1(n19428), .A2(n19261), .B1(n19427), .B2(n19238), .ZN(
        n19230) );
  AOI22_X1 U22352 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19240), .B1(
        n19429), .B2(n19308), .ZN(n19229) );
  OAI211_X1 U22353 ( .C1(n19432), .C2(n19231), .A(n19230), .B(n19229), .ZN(
        P3_U2935) );
  AOI22_X1 U22354 ( .A1(n19434), .A2(n19238), .B1(n19433), .B2(n19239), .ZN(
        n19233) );
  AOI22_X1 U22355 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19240), .B1(
        n19435), .B2(n19308), .ZN(n19232) );
  OAI211_X1 U22356 ( .C1(n19438), .C2(n19254), .A(n19233), .B(n19232), .ZN(
        P3_U2936) );
  AOI22_X1 U22357 ( .A1(n19390), .A2(n19239), .B1(n19439), .B2(n19238), .ZN(
        n19235) );
  AOI22_X1 U22358 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19240), .B1(
        n19441), .B2(n19308), .ZN(n19234) );
  OAI211_X1 U22359 ( .C1(n19393), .C2(n19254), .A(n19235), .B(n19234), .ZN(
        P3_U2937) );
  AOI22_X1 U22360 ( .A1(n19447), .A2(n19239), .B1(n19445), .B2(n19238), .ZN(
        n19237) );
  AOI22_X1 U22361 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19240), .B1(
        n19448), .B2(n19308), .ZN(n19236) );
  OAI211_X1 U22362 ( .C1(n19451), .C2(n19254), .A(n19237), .B(n19236), .ZN(
        P3_U2938) );
  AOI22_X1 U22363 ( .A1(n19338), .A2(n19239), .B1(n19454), .B2(n19238), .ZN(
        n19242) );
  AOI22_X1 U22364 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19240), .B1(
        n19457), .B2(n19308), .ZN(n19241) );
  OAI211_X1 U22365 ( .C1(n19342), .C2(n19254), .A(n19242), .B(n19241), .ZN(
        P3_U2939) );
  NAND2_X1 U22366 ( .A1(n19244), .A2(n19243), .ZN(n19334) );
  INV_X1 U22367 ( .A(n19244), .ZN(n19265) );
  NOR2_X1 U22368 ( .A1(n19265), .A2(n19343), .ZN(n19288) );
  AOI22_X1 U22369 ( .A1(n19410), .A2(n19284), .B1(n19404), .B2(n19288), .ZN(
        n19247) );
  AOI22_X1 U22370 ( .A1(n19409), .A2(n19245), .B1(n19244), .B2(n19345), .ZN(
        n19262) );
  AOI22_X1 U22371 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19262), .B1(
        n19405), .B2(n19261), .ZN(n19246) );
  OAI211_X1 U22372 ( .C1(n19413), .C2(n19334), .A(n19247), .B(n19246), .ZN(
        P3_U2940) );
  AOI22_X1 U22373 ( .A1(n19415), .A2(n19288), .B1(n19380), .B2(n19261), .ZN(
        n19249) );
  AOI22_X1 U22374 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19262), .B1(
        n19416), .B2(n19284), .ZN(n19248) );
  OAI211_X1 U22375 ( .C1(n19320), .C2(n19334), .A(n19249), .B(n19248), .ZN(
        P3_U2941) );
  AOI22_X1 U22376 ( .A1(n19352), .A2(n19261), .B1(n19421), .B2(n19288), .ZN(
        n19251) );
  INV_X1 U22377 ( .A(n19334), .ZN(n19337) );
  AOI22_X1 U22378 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19262), .B1(
        n19423), .B2(n19337), .ZN(n19250) );
  OAI211_X1 U22379 ( .C1(n19355), .C2(n19282), .A(n19251), .B(n19250), .ZN(
        P3_U2942) );
  AOI22_X1 U22380 ( .A1(n19428), .A2(n19284), .B1(n19427), .B2(n19288), .ZN(
        n19253) );
  AOI22_X1 U22381 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19262), .B1(
        n19429), .B2(n19337), .ZN(n19252) );
  OAI211_X1 U22382 ( .C1(n19432), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P3_U2943) );
  AOI22_X1 U22383 ( .A1(n19434), .A2(n19288), .B1(n19433), .B2(n19261), .ZN(
        n19256) );
  AOI22_X1 U22384 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19262), .B1(
        n19435), .B2(n19337), .ZN(n19255) );
  OAI211_X1 U22385 ( .C1(n19438), .C2(n19282), .A(n19256), .B(n19255), .ZN(
        P3_U2944) );
  AOI22_X1 U22386 ( .A1(n19390), .A2(n19261), .B1(n19439), .B2(n19288), .ZN(
        n19258) );
  AOI22_X1 U22387 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19262), .B1(
        n19441), .B2(n19337), .ZN(n19257) );
  OAI211_X1 U22388 ( .C1(n19393), .C2(n19282), .A(n19258), .B(n19257), .ZN(
        P3_U2945) );
  AOI22_X1 U22389 ( .A1(n19447), .A2(n19261), .B1(n19445), .B2(n19288), .ZN(
        n19260) );
  AOI22_X1 U22390 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19262), .B1(
        n19448), .B2(n19337), .ZN(n19259) );
  OAI211_X1 U22391 ( .C1(n19451), .C2(n19282), .A(n19260), .B(n19259), .ZN(
        P3_U2946) );
  AOI22_X1 U22392 ( .A1(n19338), .A2(n19261), .B1(n19454), .B2(n19288), .ZN(
        n19264) );
  AOI22_X1 U22393 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19262), .B1(
        n19457), .B2(n19337), .ZN(n19263) );
  OAI211_X1 U22394 ( .C1(n19342), .C2(n19282), .A(n19264), .B(n19263), .ZN(
        P3_U2947) );
  NAND2_X1 U22395 ( .A1(n19477), .A2(n19347), .ZN(n19368) );
  INV_X1 U22396 ( .A(n19368), .ZN(n19362) );
  NOR2_X1 U22397 ( .A1(n19337), .A2(n19362), .ZN(n19314) );
  NOR2_X1 U22398 ( .A1(n19370), .A2(n19314), .ZN(n19283) );
  AOI22_X1 U22399 ( .A1(n19410), .A2(n19308), .B1(n19404), .B2(n19283), .ZN(
        n19269) );
  OAI21_X1 U22400 ( .B1(n19266), .B2(n19372), .A(n19314), .ZN(n19267) );
  OAI211_X1 U22401 ( .C1(n19362), .C2(n19608), .A(n19375), .B(n19267), .ZN(
        n19285) );
  AOI22_X1 U22402 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19285), .B1(
        n19376), .B2(n19362), .ZN(n19268) );
  OAI211_X1 U22403 ( .C1(n19379), .C2(n19282), .A(n19269), .B(n19268), .ZN(
        P3_U2948) );
  AOI22_X1 U22404 ( .A1(n19416), .A2(n19308), .B1(n19415), .B2(n19283), .ZN(
        n19271) );
  AOI22_X1 U22405 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19285), .B1(
        n19417), .B2(n19362), .ZN(n19270) );
  OAI211_X1 U22406 ( .C1(n19420), .C2(n19282), .A(n19271), .B(n19270), .ZN(
        P3_U2949) );
  AOI22_X1 U22407 ( .A1(n19421), .A2(n19283), .B1(n19422), .B2(n19308), .ZN(
        n19273) );
  AOI22_X1 U22408 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19285), .B1(
        n19423), .B2(n19362), .ZN(n19272) );
  OAI211_X1 U22409 ( .C1(n19426), .C2(n19282), .A(n19273), .B(n19272), .ZN(
        P3_U2950) );
  AOI22_X1 U22410 ( .A1(n19296), .A2(n19284), .B1(n19427), .B2(n19283), .ZN(
        n19275) );
  AOI22_X1 U22411 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19285), .B1(
        n19429), .B2(n19362), .ZN(n19274) );
  OAI211_X1 U22412 ( .C1(n19299), .C2(n19304), .A(n19275), .B(n19274), .ZN(
        P3_U2951) );
  AOI22_X1 U22413 ( .A1(n19325), .A2(n19308), .B1(n19434), .B2(n19283), .ZN(
        n19277) );
  AOI22_X1 U22414 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19285), .B1(
        n19435), .B2(n19362), .ZN(n19276) );
  OAI211_X1 U22415 ( .C1(n19328), .C2(n19282), .A(n19277), .B(n19276), .ZN(
        P3_U2952) );
  AOI22_X1 U22416 ( .A1(n19440), .A2(n19308), .B1(n19439), .B2(n19283), .ZN(
        n19279) );
  AOI22_X1 U22417 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19285), .B1(
        n19441), .B2(n19362), .ZN(n19278) );
  OAI211_X1 U22418 ( .C1(n19444), .C2(n19282), .A(n19279), .B(n19278), .ZN(
        P3_U2953) );
  AOI22_X1 U22419 ( .A1(n19445), .A2(n19283), .B1(n19331), .B2(n19308), .ZN(
        n19281) );
  AOI22_X1 U22420 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19285), .B1(
        n19448), .B2(n19362), .ZN(n19280) );
  OAI211_X1 U22421 ( .C1(n19335), .C2(n19282), .A(n19281), .B(n19280), .ZN(
        P3_U2954) );
  AOI22_X1 U22422 ( .A1(n19338), .A2(n19284), .B1(n19454), .B2(n19283), .ZN(
        n19287) );
  AOI22_X1 U22423 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19285), .B1(
        n19457), .B2(n19362), .ZN(n19286) );
  OAI211_X1 U22424 ( .C1(n19342), .C2(n19304), .A(n19287), .B(n19286), .ZN(
        P3_U2955) );
  AOI22_X1 U22425 ( .A1(n19409), .A2(n19288), .B1(n19406), .B2(n19347), .ZN(
        n19309) );
  INV_X1 U22426 ( .A(n19309), .ZN(n19291) );
  AND2_X1 U22427 ( .A1(n19403), .A2(n19347), .ZN(n19307) );
  AOI22_X1 U22428 ( .A1(n19410), .A2(n19337), .B1(n19404), .B2(n19307), .ZN(
        n19290) );
  NAND2_X1 U22429 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19347), .ZN(
        n19402) );
  INV_X1 U22430 ( .A(n19402), .ZN(n19394) );
  AOI22_X1 U22431 ( .A1(n19405), .A2(n19308), .B1(n19376), .B2(n19394), .ZN(
        n19289) );
  OAI211_X1 U22432 ( .C1(n21580), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P3_U2956) );
  AOI22_X1 U22433 ( .A1(n19415), .A2(n19307), .B1(n19380), .B2(n19308), .ZN(
        n19293) );
  AOI22_X1 U22434 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19309), .B1(
        n19417), .B2(n19394), .ZN(n19292) );
  OAI211_X1 U22435 ( .C1(n19383), .C2(n19334), .A(n19293), .B(n19292), .ZN(
        P3_U2957) );
  AOI22_X1 U22436 ( .A1(n19421), .A2(n19307), .B1(n19422), .B2(n19337), .ZN(
        n19295) );
  AOI22_X1 U22437 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19309), .B1(
        n19423), .B2(n19394), .ZN(n19294) );
  OAI211_X1 U22438 ( .C1(n19426), .C2(n19304), .A(n19295), .B(n19294), .ZN(
        P3_U2958) );
  AOI22_X1 U22439 ( .A1(n19296), .A2(n19308), .B1(n19427), .B2(n19307), .ZN(
        n19298) );
  AOI22_X1 U22440 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19309), .B1(
        n19429), .B2(n19394), .ZN(n19297) );
  OAI211_X1 U22441 ( .C1(n19299), .C2(n19334), .A(n19298), .B(n19297), .ZN(
        P3_U2959) );
  AOI22_X1 U22442 ( .A1(n19434), .A2(n19307), .B1(n19433), .B2(n19308), .ZN(
        n19301) );
  AOI22_X1 U22443 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19309), .B1(
        n19435), .B2(n19394), .ZN(n19300) );
  OAI211_X1 U22444 ( .C1(n19438), .C2(n19334), .A(n19301), .B(n19300), .ZN(
        P3_U2960) );
  AOI22_X1 U22445 ( .A1(n19440), .A2(n19337), .B1(n19439), .B2(n19307), .ZN(
        n19303) );
  AOI22_X1 U22446 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19309), .B1(
        n19441), .B2(n19394), .ZN(n19302) );
  OAI211_X1 U22447 ( .C1(n19444), .C2(n19304), .A(n19303), .B(n19302), .ZN(
        P3_U2961) );
  AOI22_X1 U22448 ( .A1(n19447), .A2(n19308), .B1(n19445), .B2(n19307), .ZN(
        n19306) );
  AOI22_X1 U22449 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19309), .B1(
        n19448), .B2(n19394), .ZN(n19305) );
  OAI211_X1 U22450 ( .C1(n19451), .C2(n19334), .A(n19306), .B(n19305), .ZN(
        P3_U2962) );
  AOI22_X1 U22451 ( .A1(n19338), .A2(n19308), .B1(n19454), .B2(n19307), .ZN(
        n19311) );
  AOI22_X1 U22452 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19309), .B1(
        n19457), .B2(n19394), .ZN(n19310) );
  OAI211_X1 U22453 ( .C1(n19342), .C2(n19334), .A(n19311), .B(n19310), .ZN(
        P3_U2963) );
  INV_X1 U22454 ( .A(n19462), .ZN(n19446) );
  NOR2_X1 U22455 ( .A1(n19394), .A2(n19446), .ZN(n19373) );
  NOR2_X1 U22456 ( .A1(n19370), .A2(n19373), .ZN(n19336) );
  AOI22_X1 U22457 ( .A1(n19405), .A2(n19337), .B1(n19404), .B2(n19336), .ZN(
        n19317) );
  OAI22_X1 U22458 ( .A1(n19314), .A2(n19313), .B1(n19373), .B2(n19312), .ZN(
        n19315) );
  OAI21_X1 U22459 ( .B1(n19446), .B2(n19608), .A(n19315), .ZN(n19339) );
  AOI22_X1 U22460 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19339), .B1(
        n19410), .B2(n19362), .ZN(n19316) );
  OAI211_X1 U22461 ( .C1(n19413), .C2(n19462), .A(n19317), .B(n19316), .ZN(
        P3_U2964) );
  AOI22_X1 U22462 ( .A1(n19415), .A2(n19336), .B1(n19380), .B2(n19337), .ZN(
        n19319) );
  AOI22_X1 U22463 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19339), .B1(
        n19416), .B2(n19362), .ZN(n19318) );
  OAI211_X1 U22464 ( .C1(n19320), .C2(n19462), .A(n19319), .B(n19318), .ZN(
        P3_U2965) );
  AOI22_X1 U22465 ( .A1(n19421), .A2(n19336), .B1(n19422), .B2(n19362), .ZN(
        n19322) );
  AOI22_X1 U22466 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19339), .B1(
        n19423), .B2(n19446), .ZN(n19321) );
  OAI211_X1 U22467 ( .C1(n19426), .C2(n19334), .A(n19322), .B(n19321), .ZN(
        P3_U2966) );
  AOI22_X1 U22468 ( .A1(n19428), .A2(n19362), .B1(n19427), .B2(n19336), .ZN(
        n19324) );
  AOI22_X1 U22469 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19339), .B1(
        n19429), .B2(n19446), .ZN(n19323) );
  OAI211_X1 U22470 ( .C1(n19432), .C2(n19334), .A(n19324), .B(n19323), .ZN(
        P3_U2967) );
  AOI22_X1 U22471 ( .A1(n19325), .A2(n19362), .B1(n19434), .B2(n19336), .ZN(
        n19327) );
  AOI22_X1 U22472 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19339), .B1(
        n19435), .B2(n19446), .ZN(n19326) );
  OAI211_X1 U22473 ( .C1(n19328), .C2(n19334), .A(n19327), .B(n19326), .ZN(
        P3_U2968) );
  AOI22_X1 U22474 ( .A1(n19440), .A2(n19362), .B1(n19439), .B2(n19336), .ZN(
        n19330) );
  AOI22_X1 U22475 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19339), .B1(
        n19441), .B2(n19446), .ZN(n19329) );
  OAI211_X1 U22476 ( .C1(n19444), .C2(n19334), .A(n19330), .B(n19329), .ZN(
        P3_U2969) );
  AOI22_X1 U22477 ( .A1(n19445), .A2(n19336), .B1(n19331), .B2(n19362), .ZN(
        n19333) );
  AOI22_X1 U22478 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19339), .B1(
        n19448), .B2(n19446), .ZN(n19332) );
  OAI211_X1 U22479 ( .C1(n19335), .C2(n19334), .A(n19333), .B(n19332), .ZN(
        P3_U2970) );
  AOI22_X1 U22480 ( .A1(n19338), .A2(n19337), .B1(n19454), .B2(n19336), .ZN(
        n19341) );
  AOI22_X1 U22481 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19339), .B1(
        n19457), .B2(n19446), .ZN(n19340) );
  OAI211_X1 U22482 ( .C1(n19342), .C2(n19368), .A(n19341), .B(n19340), .ZN(
        P3_U2971) );
  INV_X1 U22483 ( .A(n19346), .ZN(n19344) );
  NOR2_X1 U22484 ( .A1(n19344), .A2(n19343), .ZN(n19408) );
  AOI22_X1 U22485 ( .A1(n19410), .A2(n19394), .B1(n19404), .B2(n19408), .ZN(
        n19349) );
  AOI22_X1 U22486 ( .A1(n19409), .A2(n19347), .B1(n19346), .B2(n19345), .ZN(
        n19365) );
  AOI22_X1 U22487 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19376), .ZN(n19348) );
  OAI211_X1 U22488 ( .C1(n19379), .C2(n19368), .A(n19349), .B(n19348), .ZN(
        P3_U2972) );
  AOI22_X1 U22489 ( .A1(n19416), .A2(n19394), .B1(n19415), .B2(n19408), .ZN(
        n19351) );
  AOI22_X1 U22490 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19417), .ZN(n19350) );
  OAI211_X1 U22491 ( .C1(n19420), .C2(n19368), .A(n19351), .B(n19350), .ZN(
        P3_U2973) );
  AOI22_X1 U22492 ( .A1(n19352), .A2(n19362), .B1(n19421), .B2(n19408), .ZN(
        n19354) );
  AOI22_X1 U22493 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19423), .ZN(n19353) );
  OAI211_X1 U22494 ( .C1(n19355), .C2(n19402), .A(n19354), .B(n19353), .ZN(
        P3_U2974) );
  AOI22_X1 U22495 ( .A1(n19428), .A2(n19394), .B1(n19427), .B2(n19408), .ZN(
        n19357) );
  AOI22_X1 U22496 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19429), .ZN(n19356) );
  OAI211_X1 U22497 ( .C1(n19432), .C2(n19368), .A(n19357), .B(n19356), .ZN(
        P3_U2975) );
  AOI22_X1 U22498 ( .A1(n19434), .A2(n19408), .B1(n19433), .B2(n19362), .ZN(
        n19359) );
  AOI22_X1 U22499 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19435), .ZN(n19358) );
  OAI211_X1 U22500 ( .C1(n19438), .C2(n19402), .A(n19359), .B(n19358), .ZN(
        P3_U2976) );
  AOI22_X1 U22501 ( .A1(n19440), .A2(n19394), .B1(n19439), .B2(n19408), .ZN(
        n19361) );
  AOI22_X1 U22502 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19441), .ZN(n19360) );
  OAI211_X1 U22503 ( .C1(n19444), .C2(n19368), .A(n19361), .B(n19360), .ZN(
        P3_U2977) );
  AOI22_X1 U22504 ( .A1(n19447), .A2(n19362), .B1(n19445), .B2(n19408), .ZN(
        n19364) );
  AOI22_X1 U22505 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19448), .ZN(n19363) );
  OAI211_X1 U22506 ( .C1(n19451), .C2(n19402), .A(n19364), .B(n19363), .ZN(
        P3_U2978) );
  AOI22_X1 U22507 ( .A1(n19455), .A2(n19394), .B1(n19454), .B2(n19408), .ZN(
        n19367) );
  AOI22_X1 U22508 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19365), .B1(
        n19456), .B2(n19457), .ZN(n19366) );
  OAI211_X1 U22509 ( .C1(n19463), .C2(n19368), .A(n19367), .B(n19366), .ZN(
        P3_U2979) );
  INV_X1 U22510 ( .A(n19369), .ZN(n19371) );
  NOR2_X1 U22511 ( .A1(n19371), .A2(n19370), .ZN(n19397) );
  AOI22_X1 U22512 ( .A1(n19410), .A2(n19446), .B1(n19404), .B2(n19397), .ZN(
        n19378) );
  OAI21_X1 U22513 ( .B1(n19373), .B2(n19372), .A(n19371), .ZN(n19374) );
  OAI211_X1 U22514 ( .C1(n19398), .C2(n19608), .A(n19375), .B(n19374), .ZN(
        n19399) );
  AOI22_X1 U22515 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19376), .ZN(n19377) );
  OAI211_X1 U22516 ( .C1(n19379), .C2(n19402), .A(n19378), .B(n19377), .ZN(
        P3_U2980) );
  AOI22_X1 U22517 ( .A1(n19415), .A2(n19397), .B1(n19380), .B2(n19394), .ZN(
        n19382) );
  AOI22_X1 U22518 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19417), .ZN(n19381) );
  OAI211_X1 U22519 ( .C1(n19383), .C2(n19462), .A(n19382), .B(n19381), .ZN(
        P3_U2981) );
  AOI22_X1 U22520 ( .A1(n19421), .A2(n19397), .B1(n19422), .B2(n19446), .ZN(
        n19385) );
  AOI22_X1 U22521 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19423), .ZN(n19384) );
  OAI211_X1 U22522 ( .C1(n19426), .C2(n19402), .A(n19385), .B(n19384), .ZN(
        P3_U2982) );
  AOI22_X1 U22523 ( .A1(n19428), .A2(n19446), .B1(n19427), .B2(n19397), .ZN(
        n19387) );
  AOI22_X1 U22524 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19429), .ZN(n19386) );
  OAI211_X1 U22525 ( .C1(n19432), .C2(n19402), .A(n19387), .B(n19386), .ZN(
        P3_U2983) );
  AOI22_X1 U22526 ( .A1(n19434), .A2(n19397), .B1(n19433), .B2(n19394), .ZN(
        n19389) );
  AOI22_X1 U22527 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19435), .ZN(n19388) );
  OAI211_X1 U22528 ( .C1(n19438), .C2(n19462), .A(n19389), .B(n19388), .ZN(
        P3_U2984) );
  AOI22_X1 U22529 ( .A1(n19390), .A2(n19394), .B1(n19439), .B2(n19397), .ZN(
        n19392) );
  AOI22_X1 U22530 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19441), .ZN(n19391) );
  OAI211_X1 U22531 ( .C1(n19393), .C2(n19462), .A(n19392), .B(n19391), .ZN(
        P3_U2985) );
  AOI22_X1 U22532 ( .A1(n19447), .A2(n19394), .B1(n19445), .B2(n19397), .ZN(
        n19396) );
  AOI22_X1 U22533 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19448), .ZN(n19395) );
  OAI211_X1 U22534 ( .C1(n19451), .C2(n19462), .A(n19396), .B(n19395), .ZN(
        P3_U2986) );
  AOI22_X1 U22535 ( .A1(n19455), .A2(n19446), .B1(n19454), .B2(n19397), .ZN(
        n19401) );
  AOI22_X1 U22536 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19457), .ZN(n19400) );
  OAI211_X1 U22537 ( .C1(n19463), .C2(n19402), .A(n19401), .B(n19400), .ZN(
        P3_U2987) );
  AND2_X1 U22538 ( .A1(n19403), .A2(n19407), .ZN(n19453) );
  AOI22_X1 U22539 ( .A1(n19405), .A2(n19446), .B1(n19404), .B2(n19453), .ZN(
        n19412) );
  AOI22_X1 U22540 ( .A1(n19409), .A2(n19408), .B1(n19407), .B2(n19406), .ZN(
        n19459) );
  AOI22_X1 U22541 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19459), .B1(
        n19456), .B2(n19410), .ZN(n19411) );
  OAI211_X1 U22542 ( .C1(n19414), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P3_U2988) );
  AOI22_X1 U22543 ( .A1(n19456), .A2(n19416), .B1(n19415), .B2(n19453), .ZN(
        n19419) );
  AOI22_X1 U22544 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19417), .ZN(n19418) );
  OAI211_X1 U22545 ( .C1(n19420), .C2(n19462), .A(n19419), .B(n19418), .ZN(
        P3_U2989) );
  AOI22_X1 U22546 ( .A1(n19456), .A2(n19422), .B1(n19421), .B2(n19453), .ZN(
        n19425) );
  AOI22_X1 U22547 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19423), .ZN(n19424) );
  OAI211_X1 U22548 ( .C1(n19426), .C2(n19462), .A(n19425), .B(n19424), .ZN(
        P3_U2990) );
  AOI22_X1 U22549 ( .A1(n19456), .A2(n19428), .B1(n19427), .B2(n19453), .ZN(
        n19431) );
  AOI22_X1 U22550 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19429), .ZN(n19430) );
  OAI211_X1 U22551 ( .C1(n19432), .C2(n19462), .A(n19431), .B(n19430), .ZN(
        P3_U2991) );
  AOI22_X1 U22552 ( .A1(n19434), .A2(n19453), .B1(n19433), .B2(n19446), .ZN(
        n19437) );
  AOI22_X1 U22553 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19435), .ZN(n19436) );
  OAI211_X1 U22554 ( .C1(n19452), .C2(n19438), .A(n19437), .B(n19436), .ZN(
        P3_U2992) );
  AOI22_X1 U22555 ( .A1(n19456), .A2(n19440), .B1(n19439), .B2(n19453), .ZN(
        n19443) );
  AOI22_X1 U22556 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19441), .ZN(n19442) );
  OAI211_X1 U22557 ( .C1(n19444), .C2(n19462), .A(n19443), .B(n19442), .ZN(
        P3_U2993) );
  AOI22_X1 U22558 ( .A1(n19447), .A2(n19446), .B1(n19445), .B2(n19453), .ZN(
        n19450) );
  AOI22_X1 U22559 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19448), .ZN(n19449) );
  OAI211_X1 U22560 ( .C1(n19452), .C2(n19451), .A(n19450), .B(n19449), .ZN(
        P3_U2994) );
  AOI22_X1 U22561 ( .A1(n19456), .A2(n19455), .B1(n19454), .B2(n19453), .ZN(
        n19461) );
  AOI22_X1 U22562 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19459), .B1(
        n19458), .B2(n19457), .ZN(n19460) );
  OAI211_X1 U22563 ( .C1(n19463), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P3_U2995) );
  INV_X1 U22564 ( .A(n19464), .ZN(n19471) );
  NOR2_X1 U22565 ( .A1(n10299), .A2(n19465), .ZN(n19467) );
  OAI222_X1 U22566 ( .A1(n19471), .A2(n19470), .B1(n19469), .B2(n19468), .C1(
        n19467), .C2(n19466), .ZN(n19619) );
  OAI211_X1 U22567 ( .C1(P3_MORE_REG_SCAN_IN), .C2(P3_FLUSH_REG_SCAN_IN), .A(
        n19473), .B(n19472), .ZN(n19475) );
  OAI211_X1 U22568 ( .C1(n19490), .C2(n21648), .A(n19475), .B(n19474), .ZN(
        n19500) );
  MUX2_X1 U22569 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19476), .S(
        n19490), .Z(n19493) );
  INV_X1 U22570 ( .A(n19493), .ZN(n19486) );
  NOR3_X1 U22571 ( .A1(n19479), .A2(n19478), .A3(n19477), .ZN(n19482) );
  INV_X1 U22572 ( .A(n19479), .ZN(n19480) );
  OAI22_X1 U22573 ( .A1(n19482), .A2(n19481), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19480), .ZN(n19484) );
  AOI21_X1 U22574 ( .B1(n19484), .B2(n19490), .A(n19483), .ZN(n19485) );
  AOI21_X1 U22575 ( .B1(n19486), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n19485), .ZN(n19495) );
  AOI22_X1 U22576 ( .A1(n19487), .A2(n19493), .B1(n19495), .B2(n11737), .ZN(
        n19498) );
  AOI21_X1 U22577 ( .B1(n19489), .B2(n19490), .A(n19488), .ZN(n19491) );
  OAI22_X1 U22578 ( .A1(n19492), .A2(n19491), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19490), .ZN(n19497) );
  AOI221_X1 U22579 ( .B1(n19495), .B2(n19494), .C1(n11737), .C2(n19494), .A(
        n19493), .ZN(n19496) );
  OAI22_X1 U22580 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19496), .ZN(n19499) );
  NOR4_X1 U22581 ( .A1(n19501), .A2(n19619), .A3(n19500), .A4(n19499), .ZN(
        n19505) );
  OAI211_X1 U22582 ( .C1(n19503), .C2(n19502), .A(n19509), .B(n19505), .ZN(
        n19607) );
  OAI21_X1 U22583 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19627), .A(n19607), 
        .ZN(n19519) );
  AOI211_X1 U22584 ( .C1(n19630), .C2(P3_STATE2_REG_3__SCAN_IN), .A(n19504), 
        .B(n19519), .ZN(n19511) );
  INV_X1 U22585 ( .A(n19505), .ZN(n19508) );
  AOI22_X1 U22586 ( .A1(n19506), .A2(n19630), .B1(n19529), .B2(n19623), .ZN(
        n19507) );
  AOI22_X1 U22587 ( .A1(n19509), .A2(n19508), .B1(n19507), .B2(n19515), .ZN(
        n19510) );
  OAI21_X1 U22588 ( .B1(n19511), .B2(n19515), .A(n19510), .ZN(P3_U2996) );
  NAND2_X1 U22589 ( .A1(n19529), .A2(n19512), .ZN(n19514) );
  OAI21_X1 U22590 ( .B1(n19515), .B2(n19514), .A(n19513), .ZN(n19520) );
  AOI22_X1 U22591 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19520), .B1(n19529), 
        .B2(n19623), .ZN(n19516) );
  OAI221_X1 U22592 ( .B1(n19519), .B2(n19518), .C1(n19519), .C2(n19517), .A(
        n19516), .ZN(P3_U2997) );
  INV_X1 U22593 ( .A(n19606), .ZN(n19521) );
  NOR3_X1 U22594 ( .A1(n19630), .A2(n19521), .A3(n19520), .ZN(P3_U2998) );
  INV_X1 U22595 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21616) );
  NOR2_X1 U22596 ( .A1(n21616), .A2(n19605), .ZN(P3_U2999) );
  AND2_X1 U22597 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19602), .ZN(
        P3_U3000) );
  AND2_X1 U22598 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19602), .ZN(
        P3_U3001) );
  AND2_X1 U22599 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19602), .ZN(
        P3_U3002) );
  AND2_X1 U22600 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19602), .ZN(
        P3_U3003) );
  AND2_X1 U22601 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19602), .ZN(
        P3_U3004) );
  AND2_X1 U22602 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19602), .ZN(
        P3_U3005) );
  AND2_X1 U22603 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19602), .ZN(
        P3_U3006) );
  AND2_X1 U22604 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19602), .ZN(
        P3_U3007) );
  AND2_X1 U22605 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19602), .ZN(
        P3_U3008) );
  AND2_X1 U22606 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19602), .ZN(
        P3_U3009) );
  AND2_X1 U22607 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19602), .ZN(
        P3_U3010) );
  AND2_X1 U22608 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19602), .ZN(
        P3_U3011) );
  AND2_X1 U22609 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19602), .ZN(
        P3_U3012) );
  AND2_X1 U22610 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19602), .ZN(
        P3_U3013) );
  AND2_X1 U22611 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19602), .ZN(
        P3_U3014) );
  INV_X1 U22612 ( .A(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21692) );
  NOR2_X1 U22613 ( .A1(n21692), .A2(n19605), .ZN(P3_U3015) );
  AND2_X1 U22614 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19602), .ZN(
        P3_U3016) );
  AND2_X1 U22615 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19602), .ZN(
        P3_U3017) );
  AND2_X1 U22616 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19602), .ZN(
        P3_U3018) );
  AND2_X1 U22617 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19602), .ZN(
        P3_U3019) );
  AND2_X1 U22618 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19602), .ZN(
        P3_U3020) );
  AND2_X1 U22619 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19602), .ZN(P3_U3021) );
  INV_X1 U22620 ( .A(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21691) );
  NOR2_X1 U22621 ( .A1(n21691), .A2(n19605), .ZN(P3_U3022) );
  AND2_X1 U22622 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19602), .ZN(P3_U3023) );
  AND2_X1 U22623 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19602), .ZN(P3_U3024) );
  AND2_X1 U22624 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19602), .ZN(P3_U3025) );
  INV_X1 U22625 ( .A(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21568) );
  NOR2_X1 U22626 ( .A1(n21568), .A2(n19605), .ZN(P3_U3026) );
  AND2_X1 U22627 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19602), .ZN(P3_U3027) );
  AND2_X1 U22628 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19602), .ZN(P3_U3028) );
  INV_X1 U22629 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19526) );
  AOI21_X1 U22630 ( .B1(HOLD), .B2(n19522), .A(n19526), .ZN(n19525) );
  NAND2_X1 U22631 ( .A1(n19529), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19532) );
  AND2_X1 U22632 ( .A1(n19532), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19536) );
  INV_X1 U22633 ( .A(NA), .ZN(n21377) );
  OAI21_X1 U22634 ( .B1(n21377), .B2(n19523), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19535) );
  INV_X1 U22635 ( .A(n19535), .ZN(n19524) );
  OAI22_X1 U22636 ( .A1(n19635), .A2(n19525), .B1(n19536), .B2(n19524), .ZN(
        P3_U3029) );
  AOI21_X1 U22637 ( .B1(HOLD), .B2(n19527), .A(n19526), .ZN(n19528) );
  AOI22_X1 U22638 ( .A1(n19529), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19528), .ZN(n19531) );
  NAND3_X1 U22639 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n19537), .ZN(
        n19530) );
  NAND3_X1 U22640 ( .A1(n19531), .A2(n19624), .A3(n19530), .ZN(P3_U3030) );
  OAI222_X1 U22641 ( .A1(n21372), .A2(n19537), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n19532), .C2(NA), .ZN(n19533)
         );
  OAI211_X1 U22642 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n19533), .ZN(n19534) );
  OAI21_X1 U22643 ( .B1(n19536), .B2(n19535), .A(n19534), .ZN(P3_U3031) );
  INV_X1 U22644 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19539) );
  NAND2_X2 U22645 ( .A1(n19635), .A2(n19537), .ZN(n19590) );
  OAI222_X1 U22646 ( .A1(n19609), .A2(n19593), .B1(n19538), .B2(n19635), .C1(
        n19539), .C2(n19590), .ZN(P3_U3032) );
  OAI222_X1 U22647 ( .A1(n19590), .A2(n19541), .B1(n19540), .B2(n19635), .C1(
        n19539), .C2(n19593), .ZN(P3_U3033) );
  OAI222_X1 U22648 ( .A1(n19590), .A2(n19543), .B1(n19542), .B2(n19635), .C1(
        n19541), .C2(n19593), .ZN(P3_U3034) );
  OAI222_X1 U22649 ( .A1(n19590), .A2(n21593), .B1(n19544), .B2(n19635), .C1(
        n19543), .C2(n19593), .ZN(P3_U3035) );
  OAI222_X1 U22650 ( .A1(n19590), .A2(n19546), .B1(n19545), .B2(n19635), .C1(
        n21593), .C2(n19593), .ZN(P3_U3036) );
  OAI222_X1 U22651 ( .A1(n19590), .A2(n19548), .B1(n19547), .B2(n19635), .C1(
        n19546), .C2(n19593), .ZN(P3_U3037) );
  OAI222_X1 U22652 ( .A1(n19590), .A2(n19551), .B1(n19549), .B2(n19635), .C1(
        n19548), .C2(n19593), .ZN(P3_U3038) );
  OAI222_X1 U22653 ( .A1(n19551), .A2(n19593), .B1(n19550), .B2(n19635), .C1(
        n21725), .C2(n19590), .ZN(P3_U3039) );
  OAI222_X1 U22654 ( .A1(n21725), .A2(n19593), .B1(n19552), .B2(n19635), .C1(
        n19553), .C2(n19590), .ZN(P3_U3040) );
  INV_X1 U22655 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19555) );
  OAI222_X1 U22656 ( .A1(n19590), .A2(n19555), .B1(n19554), .B2(n19635), .C1(
        n19553), .C2(n19593), .ZN(P3_U3041) );
  OAI222_X1 U22657 ( .A1(n19590), .A2(n19558), .B1(n19556), .B2(n19635), .C1(
        n19555), .C2(n19593), .ZN(P3_U3042) );
  OAI222_X1 U22658 ( .A1(n19558), .A2(n19593), .B1(n19557), .B2(n19635), .C1(
        n19559), .C2(n19590), .ZN(P3_U3043) );
  OAI222_X1 U22659 ( .A1(n19590), .A2(n19562), .B1(n19560), .B2(n19635), .C1(
        n19559), .C2(n19593), .ZN(P3_U3044) );
  OAI222_X1 U22660 ( .A1(n19562), .A2(n19593), .B1(n19561), .B2(n19635), .C1(
        n19563), .C2(n19590), .ZN(P3_U3045) );
  OAI222_X1 U22661 ( .A1(n19590), .A2(n19566), .B1(n19564), .B2(n19635), .C1(
        n19563), .C2(n19593), .ZN(P3_U3046) );
  OAI222_X1 U22662 ( .A1(n19566), .A2(n19593), .B1(n19565), .B2(n19635), .C1(
        n19567), .C2(n19590), .ZN(P3_U3047) );
  OAI222_X1 U22663 ( .A1(n19590), .A2(n19569), .B1(n19568), .B2(n19635), .C1(
        n19567), .C2(n19593), .ZN(P3_U3048) );
  OAI222_X1 U22664 ( .A1(n19590), .A2(n19571), .B1(n19570), .B2(n19635), .C1(
        n19569), .C2(n19593), .ZN(P3_U3049) );
  OAI222_X1 U22665 ( .A1(n19590), .A2(n21741), .B1(n19572), .B2(n19635), .C1(
        n19571), .C2(n19593), .ZN(P3_U3050) );
  OAI222_X1 U22666 ( .A1(n19590), .A2(n19575), .B1(n19573), .B2(n19635), .C1(
        n21741), .C2(n19593), .ZN(P3_U3051) );
  OAI222_X1 U22667 ( .A1(n19575), .A2(n19593), .B1(n19574), .B2(n19635), .C1(
        n19576), .C2(n19590), .ZN(P3_U3052) );
  OAI222_X1 U22668 ( .A1(n19590), .A2(n19579), .B1(n19577), .B2(n19635), .C1(
        n19576), .C2(n19593), .ZN(P3_U3053) );
  OAI222_X1 U22669 ( .A1(n19579), .A2(n19593), .B1(n19578), .B2(n19635), .C1(
        n19580), .C2(n19590), .ZN(P3_U3054) );
  OAI222_X1 U22670 ( .A1(n19590), .A2(n21627), .B1(n19581), .B2(n19635), .C1(
        n19580), .C2(n19593), .ZN(P3_U3055) );
  OAI222_X1 U22671 ( .A1(n19590), .A2(n19583), .B1(n19582), .B2(n19635), .C1(
        n21627), .C2(n19593), .ZN(P3_U3056) );
  OAI222_X1 U22672 ( .A1(n19590), .A2(n19585), .B1(n19584), .B2(n19635), .C1(
        n19583), .C2(n19593), .ZN(P3_U3057) );
  INV_X1 U22673 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19587) );
  OAI222_X1 U22674 ( .A1(n19590), .A2(n19587), .B1(n21710), .B2(n19635), .C1(
        n19585), .C2(n19593), .ZN(P3_U3058) );
  OAI222_X1 U22675 ( .A1(n19587), .A2(n19593), .B1(n19586), .B2(n19635), .C1(
        n19588), .C2(n19590), .ZN(P3_U3059) );
  OAI222_X1 U22676 ( .A1(n19590), .A2(n21720), .B1(n19589), .B2(n19635), .C1(
        n19588), .C2(n19593), .ZN(P3_U3060) );
  OAI222_X1 U22677 ( .A1(n19593), .A2(n21720), .B1(n19592), .B2(n19635), .C1(
        n19591), .C2(n19590), .ZN(P3_U3061) );
  INV_X1 U22678 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19594) );
  AOI22_X1 U22679 ( .A1(n19635), .A2(n19595), .B1(n19594), .B2(n19616), .ZN(
        P3_U3274) );
  INV_X1 U22680 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19612) );
  INV_X1 U22681 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19596) );
  AOI22_X1 U22682 ( .A1(n19635), .A2(n19612), .B1(n19596), .B2(n19616), .ZN(
        P3_U3275) );
  INV_X1 U22683 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19597) );
  AOI22_X1 U22684 ( .A1(n19635), .A2(n19598), .B1(n19597), .B2(n19616), .ZN(
        P3_U3276) );
  INV_X1 U22685 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21786) );
  INV_X1 U22686 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19599) );
  AOI22_X1 U22687 ( .A1(n19635), .A2(n21786), .B1(n19599), .B2(n19616), .ZN(
        P3_U3277) );
  INV_X1 U22688 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19601) );
  INV_X1 U22689 ( .A(n19603), .ZN(n19600) );
  AOI21_X1 U22690 ( .B1(n19602), .B2(n19601), .A(n19600), .ZN(P3_U3280) );
  OAI21_X1 U22691 ( .B1(n19605), .B2(n19604), .A(n19603), .ZN(P3_U3281) );
  OAI221_X1 U22692 ( .B1(n19608), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19608), 
        .C2(n19607), .A(n19606), .ZN(P3_U3282) );
  AOI21_X1 U22693 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19610) );
  AOI22_X1 U22694 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19610), .B2(n19609), .ZN(n19613) );
  AOI22_X1 U22695 ( .A1(n19615), .A2(n19613), .B1(n19612), .B2(n19611), .ZN(
        P3_U3292) );
  OAI21_X1 U22696 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19615), .ZN(n19614) );
  OAI21_X1 U22697 ( .B1(n19615), .B2(n21786), .A(n19614), .ZN(P3_U3293) );
  INV_X1 U22698 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19617) );
  AOI22_X1 U22699 ( .A1(n19635), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19617), 
        .B2(n19616), .ZN(P3_U3294) );
  MUX2_X1 U22700 ( .A(P3_MORE_REG_SCAN_IN), .B(n19619), .S(n19618), .Z(
        P3_U3295) );
  OAI21_X1 U22701 ( .B1(n19621), .B2(n19620), .A(n19638), .ZN(n19622) );
  AOI21_X1 U22702 ( .B1(n19623), .B2(n19627), .A(n19622), .ZN(n19634) );
  AOI21_X1 U22703 ( .B1(n19626), .B2(n19625), .A(n19624), .ZN(n19628) );
  OAI211_X1 U22704 ( .C1(n19629), .C2(n19628), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19627), .ZN(n19631) );
  AOI21_X1 U22705 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19631), .A(n19630), 
        .ZN(n19633) );
  NAND2_X1 U22706 ( .A1(n19634), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19632) );
  OAI21_X1 U22707 ( .B1(n19634), .B2(n19633), .A(n19632), .ZN(P3_U3296) );
  MUX2_X1 U22708 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n19635), .Z(P3_U3297) );
  OAI21_X1 U22709 ( .B1(n19639), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19638), 
        .ZN(n19636) );
  OAI21_X1 U22710 ( .B1(n19638), .B2(n19637), .A(n19636), .ZN(P3_U3298) );
  NOR2_X1 U22711 ( .A1(n19639), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19641)
         );
  OAI21_X1 U22712 ( .B1(n19642), .B2(n19641), .A(n19640), .ZN(P3_U3299) );
  INV_X1 U22713 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19643) );
  NAND2_X1 U22714 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21644), .ZN(n20403) );
  NAND2_X1 U22715 ( .A1(n20395), .A2(n20394), .ZN(n20400) );
  OAI21_X1 U22716 ( .B1(n20395), .B2(n20403), .A(n20400), .ZN(n20475) );
  OAI21_X1 U22717 ( .B1(n20395), .B2(n19643), .A(n20393), .ZN(P2_U2815) );
  AOI22_X1 U22718 ( .A1(n20462), .A2(n19644), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20526), .ZN(n19645) );
  OAI21_X1 U22719 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20400), .A(n19645), 
        .ZN(P2_U2817) );
  INV_X1 U22720 ( .A(n20407), .ZN(n19646) );
  OAI21_X1 U22721 ( .B1(n19646), .B2(BS16), .A(n20475), .ZN(n20473) );
  OAI21_X1 U22722 ( .B1(n20475), .B2(n20512), .A(n20473), .ZN(P2_U2818) );
  NOR4_X1 U22723 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19656) );
  NOR4_X1 U22724 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19655) );
  AOI211_X1 U22725 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19647) );
  INV_X1 U22726 ( .A(P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21743) );
  INV_X1 U22727 ( .A(P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n21662) );
  NAND3_X1 U22728 ( .A1(n19647), .A2(n21743), .A3(n21662), .ZN(n19653) );
  NOR4_X1 U22729 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19651) );
  NOR4_X1 U22730 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19650) );
  NOR4_X1 U22731 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19649) );
  NOR4_X1 U22732 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19648) );
  NAND4_X1 U22733 ( .A1(n19651), .A2(n19650), .A3(n19649), .A4(n19648), .ZN(
        n19652) );
  NOR4_X1 U22734 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n19653), .A4(n19652), .ZN(n19654) );
  NAND3_X1 U22735 ( .A1(n19656), .A2(n19655), .A3(n19654), .ZN(n19662) );
  NOR2_X1 U22736 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19662), .ZN(n19657) );
  INV_X1 U22737 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20471) );
  AOI22_X1 U22738 ( .A1(n19657), .A2(n10758), .B1(n19662), .B2(n20471), .ZN(
        P2_U2820) );
  OR3_X1 U22739 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19661) );
  INV_X1 U22740 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20469) );
  AOI22_X1 U22741 ( .A1(n19657), .A2(n19661), .B1(n19662), .B2(n20469), .ZN(
        P2_U2821) );
  INV_X1 U22742 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20474) );
  NAND2_X1 U22743 ( .A1(n19657), .A2(n20474), .ZN(n19660) );
  INV_X1 U22744 ( .A(n19662), .ZN(n19663) );
  OAI21_X1 U22745 ( .B1(n20412), .B2(n10758), .A(n19663), .ZN(n19658) );
  OAI21_X1 U22746 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19663), .A(n19658), 
        .ZN(n19659) );
  OAI221_X1 U22747 ( .B1(n19660), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19660), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19659), .ZN(P2_U2822) );
  INV_X1 U22748 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20466) );
  OAI221_X1 U22749 ( .B1(n19663), .B2(n20466), .C1(n19662), .C2(n19661), .A(
        n19660), .ZN(P2_U2823) );
  OAI22_X1 U22750 ( .A1(n19667), .A2(n19666), .B1(n19665), .B2(n19664), .ZN(
        n19668) );
  INV_X1 U22751 ( .A(n19668), .ZN(n19688) );
  AOI22_X1 U22752 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19669), .ZN(n19687) );
  INV_X1 U22753 ( .A(n19672), .ZN(n19679) );
  INV_X1 U22754 ( .A(n19673), .ZN(n19675) );
  AOI222_X1 U22755 ( .A1(n19679), .A2(n19678), .B1(n19677), .B2(n19676), .C1(
        n19675), .C2(n19674), .ZN(n19686) );
  INV_X1 U22756 ( .A(n19680), .ZN(n19682) );
  OAI211_X1 U22757 ( .C1(n19684), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        n19685) );
  NAND4_X1 U22758 ( .A1(n19688), .A2(n19687), .A3(n19686), .A4(n19685), .ZN(
        P2_U2835) );
  INV_X1 U22759 ( .A(n19689), .ZN(n19690) );
  AOI22_X1 U22760 ( .A1(n19690), .A2(n19705), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n16451), .ZN(n19695) );
  XNOR2_X1 U22761 ( .A(n19692), .B(n19691), .ZN(n19693) );
  NAND2_X1 U22762 ( .A1(n19693), .A2(n19709), .ZN(n19694) );
  OAI211_X1 U22763 ( .C1(n19696), .C2(n19713), .A(n19695), .B(n19694), .ZN(
        P2_U2915) );
  AOI22_X1 U22764 ( .A1(n19705), .A2(n20485), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n16451), .ZN(n19702) );
  OAI21_X1 U22765 ( .B1(n19699), .B2(n19698), .A(n19697), .ZN(n19700) );
  NAND2_X1 U22766 ( .A1(n19700), .A2(n19709), .ZN(n19701) );
  OAI211_X1 U22767 ( .C1(n19703), .C2(n19713), .A(n19702), .B(n19701), .ZN(
        P2_U2916) );
  AOI22_X1 U22768 ( .A1(n19705), .A2(n19704), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n16451), .ZN(n19712) );
  OAI21_X1 U22769 ( .B1(n19708), .B2(n19707), .A(n19706), .ZN(n19710) );
  NAND2_X1 U22770 ( .A1(n19710), .A2(n19709), .ZN(n19711) );
  OAI211_X1 U22771 ( .C1(n19714), .C2(n19713), .A(n19712), .B(n19711), .ZN(
        P2_U2918) );
  NOR2_X1 U22772 ( .A1(n19747), .A2(n19715), .ZN(P2_U2920) );
  AOI22_X1 U22773 ( .A1(n19744), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19716) );
  OAI21_X1 U22774 ( .B1(n13937), .B2(n19742), .A(n19716), .ZN(P2_U2936) );
  AOI22_X1 U22775 ( .A1(n19744), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19717) );
  OAI21_X1 U22776 ( .B1(n19718), .B2(n19742), .A(n19717), .ZN(P2_U2937) );
  AOI22_X1 U22777 ( .A1(n19744), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19719) );
  OAI21_X1 U22778 ( .B1(n19720), .B2(n19742), .A(n19719), .ZN(P2_U2938) );
  AOI22_X1 U22779 ( .A1(n19744), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19721) );
  OAI21_X1 U22780 ( .B1(n19722), .B2(n19742), .A(n19721), .ZN(P2_U2939) );
  AOI22_X1 U22781 ( .A1(n19744), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19723) );
  OAI21_X1 U22782 ( .B1(n19724), .B2(n19742), .A(n19723), .ZN(P2_U2940) );
  AOI22_X1 U22783 ( .A1(n19744), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19725) );
  OAI21_X1 U22784 ( .B1(n19726), .B2(n19742), .A(n19725), .ZN(P2_U2941) );
  AOI22_X1 U22785 ( .A1(n19744), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19727) );
  OAI21_X1 U22786 ( .B1(n19728), .B2(n19742), .A(n19727), .ZN(P2_U2942) );
  AOI22_X1 U22787 ( .A1(n19744), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19729) );
  OAI21_X1 U22788 ( .B1(n19730), .B2(n19742), .A(n19729), .ZN(P2_U2943) );
  AOI22_X1 U22789 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n19739), .B1(n19744), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19731) );
  OAI21_X1 U22790 ( .B1(n21790), .B2(n19742), .A(n19731), .ZN(P2_U2944) );
  AOI22_X1 U22791 ( .A1(n19744), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19732) );
  OAI21_X1 U22792 ( .B1(n19733), .B2(n19742), .A(n19732), .ZN(P2_U2945) );
  INV_X1 U22793 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19735) );
  AOI22_X1 U22794 ( .A1(n19744), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19734) );
  OAI21_X1 U22795 ( .B1(n19735), .B2(n19742), .A(n19734), .ZN(P2_U2946) );
  INV_X1 U22796 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n21740) );
  AOI22_X1 U22797 ( .A1(n19744), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19736) );
  OAI21_X1 U22798 ( .B1(n21740), .B2(n19742), .A(n19736), .ZN(P2_U2947) );
  INV_X1 U22799 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U22800 ( .A1(n19744), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19737) );
  OAI21_X1 U22801 ( .B1(n19738), .B2(n19742), .A(n19737), .ZN(P2_U2948) );
  INV_X1 U22802 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n21611) );
  AOI22_X1 U22803 ( .A1(n19744), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19740) );
  OAI21_X1 U22804 ( .B1(n21611), .B2(n19742), .A(n19740), .ZN(P2_U2949) );
  INV_X1 U22805 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U22806 ( .A1(n19744), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19739), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19741) );
  OAI21_X1 U22807 ( .B1(n19743), .B2(n19742), .A(n19741), .ZN(P2_U2950) );
  AOI22_X1 U22808 ( .A1(P2_EAX_REG_0__SCAN_IN), .A2(n19745), .B1(n19744), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n19746) );
  OAI21_X1 U22809 ( .B1(n21641), .B2(n19747), .A(n19746), .ZN(P2_U2951) );
  AOI22_X1 U22810 ( .A1(n19779), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19748), .ZN(n19756) );
  NAND2_X1 U22811 ( .A1(n19749), .A2(n19781), .ZN(n19752) );
  NAND2_X1 U22812 ( .A1(n19750), .A2(n19763), .ZN(n19751) );
  OAI211_X1 U22813 ( .C1(n19774), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        n19754) );
  INV_X1 U22814 ( .A(n19754), .ZN(n19755) );
  OAI211_X1 U22815 ( .C1(n19758), .C2(n19757), .A(n19756), .B(n19755), .ZN(
        P2_U3010) );
  OAI21_X1 U22816 ( .B1(n19761), .B2(n19760), .A(n19759), .ZN(n19762) );
  INV_X1 U22817 ( .A(n19762), .ZN(n19793) );
  AOI22_X1 U22818 ( .A1(n19793), .A2(n19763), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19779), .ZN(n19777) );
  INV_X1 U22819 ( .A(n19764), .ZN(n19765) );
  NAND2_X1 U22820 ( .A1(n19766), .A2(n19765), .ZN(n19767) );
  AND2_X1 U22821 ( .A1(n19768), .A2(n19767), .ZN(n19795) );
  NAND2_X1 U22822 ( .A1(n19795), .A2(n19781), .ZN(n19773) );
  OR2_X1 U22823 ( .A1(n11468), .A2(n20414), .ZN(n19799) );
  INV_X1 U22824 ( .A(n19799), .ZN(n19770) );
  AOI21_X1 U22825 ( .B1(n19771), .B2(n9845), .A(n19770), .ZN(n19772) );
  OAI211_X1 U22826 ( .C1(n19802), .C2(n19774), .A(n19773), .B(n19772), .ZN(
        n19775) );
  INV_X1 U22827 ( .A(n19775), .ZN(n19776) );
  NAND2_X1 U22828 ( .A1(n19777), .A2(n19776), .ZN(P2_U3012) );
  NOR2_X1 U22829 ( .A1(n19779), .A2(n19778), .ZN(n19791) );
  INV_X1 U22830 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19790) );
  NAND2_X1 U22831 ( .A1(n19781), .A2(n19780), .ZN(n19783) );
  OAI211_X1 U22832 ( .C1(n19785), .C2(n19784), .A(n19783), .B(n19782), .ZN(
        n19786) );
  AOI21_X1 U22833 ( .B1(n19788), .B2(n19787), .A(n19786), .ZN(n19789) );
  OAI21_X1 U22834 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(P2_U3014) );
  AOI22_X1 U22835 ( .A1(n11071), .A2(n19793), .B1(n19792), .B2(n20490), .ZN(
        n19813) );
  AOI22_X1 U22836 ( .A1(n19796), .A2(n19795), .B1(n19807), .B2(n19794), .ZN(
        n19812) );
  NOR2_X1 U22837 ( .A1(n19798), .A2(n19797), .ZN(n19800) );
  OAI21_X1 U22838 ( .B1(n19801), .B2(n19800), .A(n19799), .ZN(n19805) );
  NOR2_X1 U22839 ( .A1(n19803), .A2(n19802), .ZN(n19804) );
  NOR2_X1 U22840 ( .A1(n19805), .A2(n19804), .ZN(n19811) );
  OAI21_X1 U22841 ( .B1(n19808), .B2(n19807), .A(n19806), .ZN(n19809) );
  NAND2_X1 U22842 ( .A1(n19809), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19810) );
  NAND4_X1 U22843 ( .A1(n19813), .A2(n19812), .A3(n19811), .A4(n19810), .ZN(
        P2_U3044) );
  AOI22_X1 U22844 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19844), .ZN(n20302) );
  INV_X1 U22845 ( .A(n20302), .ZN(n20340) );
  OR2_X1 U22846 ( .A1(n19847), .A2(n20510), .ZN(n19991) );
  AOI22_X1 U22847 ( .A1(n20389), .A2(n20340), .B1(n19848), .B2(n20338), .ZN(
        n19818) );
  AOI22_X1 U22848 ( .A1(n20339), .A2(n19853), .B1(n19880), .B2(n20341), .ZN(
        n19817) );
  OAI211_X1 U22849 ( .C1(n19857), .C2(n19819), .A(n19818), .B(n19817), .ZN(
        P2_U3048) );
  AOI22_X1 U22850 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19844), .ZN(n20305) );
  INV_X1 U22851 ( .A(n20305), .ZN(n20346) );
  OR2_X1 U22852 ( .A1(n19847), .A2(n11051), .ZN(n20002) );
  AOI22_X1 U22853 ( .A1(n20389), .A2(n20346), .B1(n19848), .B2(n20344), .ZN(
        n19823) );
  OAI22_X2 U22854 ( .A1(n19821), .A2(n19851), .B1(n16454), .B2(n19850), .ZN(
        n20347) );
  AOI22_X1 U22855 ( .A1(n20345), .A2(n19853), .B1(n19880), .B2(n20347), .ZN(
        n19822) );
  OAI211_X1 U22856 ( .C1(n19857), .C2(n19824), .A(n19823), .B(n19822), .ZN(
        P2_U3049) );
  AOI22_X1 U22857 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19844), .ZN(n20311) );
  INV_X1 U22858 ( .A(n20311), .ZN(n20359) );
  OR2_X1 U22859 ( .A1(n19847), .A2(n10101), .ZN(n20009) );
  AOI22_X1 U22860 ( .A1(n20389), .A2(n20359), .B1(n19848), .B2(n20357), .ZN(
        n19828) );
  AOI22_X1 U22861 ( .A1(n20358), .A2(n19853), .B1(n19880), .B2(n20360), .ZN(
        n19827) );
  OAI211_X1 U22862 ( .C1(n19857), .C2(n19829), .A(n19828), .B(n19827), .ZN(
        P2_U3051) );
  AOI22_X2 U22863 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19844), .ZN(n20314) );
  INV_X1 U22864 ( .A(n20314), .ZN(n20366) );
  NOR2_X2 U22865 ( .A1(n19847), .A2(n10739), .ZN(n20364) );
  AOI22_X1 U22866 ( .A1(n20389), .A2(n20366), .B1(n19848), .B2(n20364), .ZN(
        n19833) );
  OAI22_X2 U22867 ( .A1(n19831), .A2(n19851), .B1(n16434), .B2(n19850), .ZN(
        n20367) );
  AOI22_X1 U22868 ( .A1(n20365), .A2(n19853), .B1(n19880), .B2(n20367), .ZN(
        n19832) );
  OAI211_X1 U22869 ( .C1(n19857), .C2(n14152), .A(n19833), .B(n19832), .ZN(
        P2_U3052) );
  AOI22_X2 U22870 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19844), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19845), .ZN(n20317) );
  INV_X1 U22871 ( .A(n20317), .ZN(n20372) );
  OR2_X1 U22872 ( .A1(n19847), .A2(n9700), .ZN(n19942) );
  AOI22_X1 U22873 ( .A1(n20389), .A2(n20372), .B1(n19848), .B2(n20370), .ZN(
        n19838) );
  OAI22_X2 U22874 ( .A1(n19836), .A2(n19851), .B1(n16425), .B2(n19850), .ZN(
        n20373) );
  AOI22_X1 U22875 ( .A1(n20371), .A2(n19853), .B1(n19880), .B2(n20373), .ZN(
        n19837) );
  OAI211_X1 U22876 ( .C1(n19857), .C2(n14428), .A(n19838), .B(n19837), .ZN(
        P2_U3053) );
  INV_X1 U22877 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19843) );
  AOI22_X2 U22878 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19844), .ZN(n20320) );
  INV_X1 U22879 ( .A(n20320), .ZN(n20378) );
  OR2_X1 U22880 ( .A1(n19847), .A2(n19839), .ZN(n20018) );
  AOI22_X1 U22881 ( .A1(n20389), .A2(n20378), .B1(n19848), .B2(n20376), .ZN(
        n19842) );
  AOI22_X1 U22882 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19844), .ZN(n20210) );
  AOI22_X1 U22883 ( .A1(n20377), .A2(n19853), .B1(n19880), .B2(n20379), .ZN(
        n19841) );
  OAI211_X1 U22884 ( .C1(n19857), .C2(n19843), .A(n19842), .B(n19841), .ZN(
        P2_U3054) );
  INV_X1 U22885 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19856) );
  AOI22_X2 U22886 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19845), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19844), .ZN(n20327) );
  INV_X1 U22887 ( .A(n20327), .ZN(n20386) );
  OR2_X1 U22888 ( .A1(n19847), .A2(n19846), .ZN(n20022) );
  AOI22_X1 U22889 ( .A1(n20389), .A2(n20386), .B1(n19848), .B2(n20382), .ZN(
        n19855) );
  OAI22_X2 U22890 ( .A1(n19852), .A2(n19851), .B1(n16410), .B2(n19850), .ZN(
        n20388) );
  AOI22_X1 U22891 ( .A1(n20384), .A2(n19853), .B1(n19880), .B2(n20388), .ZN(
        n19854) );
  OAI211_X1 U22892 ( .C1(n19857), .C2(n19856), .A(n19855), .B(n19854), .ZN(
        P2_U3055) );
  OR2_X1 U22893 ( .A1(n19919), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19862) );
  INV_X1 U22894 ( .A(n19859), .ZN(n20256) );
  AND2_X1 U22895 ( .A1(n20252), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20253) );
  INV_X1 U22896 ( .A(n19919), .ZN(n19922) );
  NAND2_X1 U22897 ( .A1(n20253), .A2(n19922), .ZN(n19863) );
  NAND2_X1 U22898 ( .A1(n19863), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19860) );
  AOI211_X2 U22899 ( .C1(n19862), .C2(n20508), .A(n20256), .B(n19861), .ZN(
        n19884) );
  AOI22_X1 U22900 ( .A1(n19884), .A2(n20339), .B1(n20338), .B2(n19883), .ZN(
        n19868) );
  NOR2_X1 U22901 ( .A1(n20486), .A2(n20512), .ZN(n20066) );
  INV_X1 U22902 ( .A(n20066), .ZN(n19993) );
  OAI21_X1 U22903 ( .B1(n19993), .B2(n20125), .A(n19862), .ZN(n19866) );
  NAND2_X1 U22904 ( .A1(n19863), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19864) );
  NAND4_X1 U22905 ( .A1(n19866), .A2(n20298), .A3(n19865), .A4(n19864), .ZN(
        n19885) );
  AOI22_X1 U22906 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19885), .B1(
        n19880), .B2(n20340), .ZN(n19867) );
  OAI211_X1 U22907 ( .C1(n20265), .C2(n19918), .A(n19868), .B(n19867), .ZN(
        P2_U3056) );
  AOI22_X1 U22908 ( .A1(n19884), .A2(n20345), .B1(n20344), .B2(n19883), .ZN(
        n19870) );
  AOI22_X1 U22909 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19885), .B1(
        n19880), .B2(n20346), .ZN(n19869) );
  OAI211_X1 U22910 ( .C1(n20268), .C2(n19918), .A(n19870), .B(n19869), .ZN(
        P2_U3057) );
  AOI22_X1 U22911 ( .A1(n19884), .A2(n20352), .B1(n20351), .B2(n19883), .ZN(
        n19873) );
  INV_X1 U22912 ( .A(n20308), .ZN(n20353) );
  AOI22_X1 U22913 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19885), .B1(
        n19880), .B2(n20353), .ZN(n19872) );
  OAI211_X1 U22914 ( .C1(n20271), .C2(n19918), .A(n19873), .B(n19872), .ZN(
        P2_U3058) );
  AOI22_X1 U22915 ( .A1(n19884), .A2(n20358), .B1(n20357), .B2(n19883), .ZN(
        n19875) );
  AOI22_X1 U22916 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19885), .B1(
        n19880), .B2(n20359), .ZN(n19874) );
  OAI211_X1 U22917 ( .C1(n20274), .C2(n19918), .A(n19875), .B(n19874), .ZN(
        P2_U3059) );
  INV_X1 U22918 ( .A(n19880), .ZN(n19888) );
  AOI22_X1 U22919 ( .A1(n19884), .A2(n20365), .B1(n20364), .B2(n19883), .ZN(
        n19877) );
  INV_X1 U22920 ( .A(n19918), .ZN(n19894) );
  AOI22_X1 U22921 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19885), .B1(
        n19894), .B2(n20367), .ZN(n19876) );
  OAI211_X1 U22922 ( .C1(n20314), .C2(n19888), .A(n19877), .B(n19876), .ZN(
        P2_U3060) );
  INV_X1 U22923 ( .A(n20373), .ZN(n20207) );
  AOI22_X1 U22924 ( .A1(n19884), .A2(n20371), .B1(n20370), .B2(n19883), .ZN(
        n19879) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19885), .B1(
        n19880), .B2(n20372), .ZN(n19878) );
  OAI211_X1 U22926 ( .C1(n20207), .C2(n19918), .A(n19879), .B(n19878), .ZN(
        P2_U3061) );
  AOI22_X1 U22927 ( .A1(n19884), .A2(n20377), .B1(n20376), .B2(n19883), .ZN(
        n19882) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19885), .B1(
        n19880), .B2(n20378), .ZN(n19881) );
  OAI211_X1 U22929 ( .C1(n20210), .C2(n19918), .A(n19882), .B(n19881), .ZN(
        P2_U3062) );
  AOI22_X1 U22930 ( .A1(n19884), .A2(n20384), .B1(n20382), .B2(n19883), .ZN(
        n19887) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19885), .B1(
        n19894), .B2(n20388), .ZN(n19886) );
  OAI211_X1 U22932 ( .C1(n20327), .C2(n19888), .A(n19887), .B(n19886), .ZN(
        P2_U3063) );
  AND2_X1 U22933 ( .A1(n19889), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20154) );
  OAI21_X1 U22934 ( .B1(n19892), .B2(n19913), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19891) );
  INV_X1 U22935 ( .A(n20290), .ZN(n19890) );
  NAND2_X1 U22936 ( .A1(n19890), .A2(n19922), .ZN(n19895) );
  NAND2_X1 U22937 ( .A1(n19891), .A2(n19895), .ZN(n19914) );
  AOI22_X1 U22938 ( .A1(n19914), .A2(n20339), .B1(n19913), .B2(n20338), .ZN(
        n19900) );
  INV_X1 U22939 ( .A(n19892), .ZN(n19893) );
  AOI21_X1 U22940 ( .B1(n19893), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19898) );
  OAI21_X1 U22941 ( .B1(n19932), .B2(n19894), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19896) );
  NAND3_X1 U22942 ( .A1(n19896), .A2(n20484), .A3(n19895), .ZN(n19897) );
  AOI22_X1 U22943 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20341), .ZN(n19899) );
  OAI211_X1 U22944 ( .C1(n20302), .C2(n19918), .A(n19900), .B(n19899), .ZN(
        P2_U3064) );
  AOI22_X1 U22945 ( .A1(n19914), .A2(n20345), .B1(n19913), .B2(n20344), .ZN(
        n19902) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20347), .ZN(n19901) );
  OAI211_X1 U22947 ( .C1(n20305), .C2(n19918), .A(n19902), .B(n19901), .ZN(
        P2_U3065) );
  AOI22_X1 U22948 ( .A1(n19914), .A2(n20352), .B1(n19913), .B2(n20351), .ZN(
        n19904) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20354), .ZN(n19903) );
  OAI211_X1 U22950 ( .C1(n20308), .C2(n19918), .A(n19904), .B(n19903), .ZN(
        P2_U3066) );
  AOI22_X1 U22951 ( .A1(n19914), .A2(n20358), .B1(n19913), .B2(n20357), .ZN(
        n19906) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20360), .ZN(n19905) );
  OAI211_X1 U22953 ( .C1(n20311), .C2(n19918), .A(n19906), .B(n19905), .ZN(
        P2_U3067) );
  AOI22_X1 U22954 ( .A1(n19914), .A2(n20365), .B1(n19913), .B2(n20364), .ZN(
        n19908) );
  AOI22_X1 U22955 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20367), .ZN(n19907) );
  OAI211_X1 U22956 ( .C1(n20314), .C2(n19918), .A(n19908), .B(n19907), .ZN(
        P2_U3068) );
  AOI22_X1 U22957 ( .A1(n19914), .A2(n20371), .B1(n19913), .B2(n20370), .ZN(
        n19910) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20373), .ZN(n19909) );
  OAI211_X1 U22959 ( .C1(n20317), .C2(n19918), .A(n19910), .B(n19909), .ZN(
        P2_U3069) );
  AOI22_X1 U22960 ( .A1(n19914), .A2(n20377), .B1(n19913), .B2(n20376), .ZN(
        n19912) );
  AOI22_X1 U22961 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20379), .ZN(n19911) );
  OAI211_X1 U22962 ( .C1(n20320), .C2(n19918), .A(n19912), .B(n19911), .ZN(
        P2_U3070) );
  AOI22_X1 U22963 ( .A1(n19914), .A2(n20384), .B1(n19913), .B2(n20382), .ZN(
        n19917) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19915), .B1(
        n19932), .B2(n20388), .ZN(n19916) );
  OAI211_X1 U22965 ( .C1(n20327), .C2(n19918), .A(n19917), .B(n19916), .ZN(
        P2_U3071) );
  NOR2_X1 U22966 ( .A1(n19920), .A2(n19919), .ZN(n19951) );
  INV_X1 U22967 ( .A(n19951), .ZN(n19946) );
  OAI22_X1 U22968 ( .A1(n19947), .A2(n20302), .B1(n19946), .B2(n19991), .ZN(
        n19921) );
  INV_X1 U22969 ( .A(n19921), .ZN(n19931) );
  OAI21_X1 U22970 ( .B1(n19993), .B2(n20190), .A(n20484), .ZN(n19929) );
  AND2_X1 U22971 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19922), .ZN(
        n19925) );
  INV_X1 U22972 ( .A(n19926), .ZN(n19923) );
  OAI211_X1 U22973 ( .C1(n19923), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20478), 
        .B(n19946), .ZN(n19924) );
  OAI211_X1 U22974 ( .C1(n19929), .C2(n19925), .A(n20298), .B(n19924), .ZN(
        n19953) );
  INV_X1 U22975 ( .A(n19925), .ZN(n19928) );
  OAI21_X1 U22976 ( .B1(n19926), .B2(n19951), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19927) );
  AOI22_X1 U22977 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19953), .B1(
        n20339), .B2(n19952), .ZN(n19930) );
  OAI211_X1 U22978 ( .C1(n20265), .C2(n19990), .A(n19931), .B(n19930), .ZN(
        P2_U3072) );
  AOI22_X1 U22979 ( .A1(n20347), .A2(n19968), .B1(n19951), .B2(n20344), .ZN(
        n19934) );
  AOI22_X1 U22980 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19953), .B1(
        n20345), .B2(n19952), .ZN(n19933) );
  OAI211_X1 U22981 ( .C1(n20305), .C2(n19947), .A(n19934), .B(n19933), .ZN(
        P2_U3073) );
  AOI22_X1 U22982 ( .A1(n20354), .A2(n19968), .B1(n20351), .B2(n19951), .ZN(
        n19936) );
  AOI22_X1 U22983 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19953), .B1(
        n20352), .B2(n19952), .ZN(n19935) );
  OAI211_X1 U22984 ( .C1(n20308), .C2(n19947), .A(n19936), .B(n19935), .ZN(
        P2_U3074) );
  OAI22_X1 U22985 ( .A1(n19947), .A2(n20311), .B1(n19946), .B2(n20009), .ZN(
        n19937) );
  INV_X1 U22986 ( .A(n19937), .ZN(n19939) );
  AOI22_X1 U22987 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19953), .B1(
        n20358), .B2(n19952), .ZN(n19938) );
  OAI211_X1 U22988 ( .C1(n20274), .C2(n19990), .A(n19939), .B(n19938), .ZN(
        P2_U3075) );
  AOI22_X1 U22989 ( .A1(n20367), .A2(n19968), .B1(n19951), .B2(n20364), .ZN(
        n19941) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19953), .B1(
        n20365), .B2(n19952), .ZN(n19940) );
  OAI211_X1 U22991 ( .C1(n20314), .C2(n19947), .A(n19941), .B(n19940), .ZN(
        P2_U3076) );
  OAI22_X1 U22992 ( .A1(n19947), .A2(n20317), .B1(n19946), .B2(n19942), .ZN(
        n19943) );
  INV_X1 U22993 ( .A(n19943), .ZN(n19945) );
  AOI22_X1 U22994 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19953), .B1(
        n20371), .B2(n19952), .ZN(n19944) );
  OAI211_X1 U22995 ( .C1(n20207), .C2(n19990), .A(n19945), .B(n19944), .ZN(
        P2_U3077) );
  OAI22_X1 U22996 ( .A1(n19947), .A2(n20320), .B1(n19946), .B2(n20018), .ZN(
        n19948) );
  INV_X1 U22997 ( .A(n19948), .ZN(n19950) );
  AOI22_X1 U22998 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19953), .B1(
        n20377), .B2(n19952), .ZN(n19949) );
  OAI211_X1 U22999 ( .C1(n20210), .C2(n19990), .A(n19950), .B(n19949), .ZN(
        P2_U3078) );
  AOI22_X1 U23000 ( .A1(n20388), .A2(n19968), .B1(n19951), .B2(n20382), .ZN(
        n19955) );
  AOI22_X1 U23001 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19953), .B1(
        n20384), .B2(n19952), .ZN(n19954) );
  OAI211_X1 U23002 ( .C1(n20327), .C2(n19947), .A(n19955), .B(n19954), .ZN(
        P2_U3079) );
  NAND2_X1 U23003 ( .A1(n10864), .A2(n12673), .ZN(n19956) );
  NOR2_X1 U23004 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20497), .ZN(
        n20060) );
  INV_X1 U23005 ( .A(n20060), .ZN(n20031) );
  OR2_X1 U23006 ( .A1(n20219), .A2(n20031), .ZN(n19965) );
  NAND3_X1 U23007 ( .A1(n19956), .A2(n20478), .A3(n19965), .ZN(n19963) );
  INV_X1 U23008 ( .A(n20219), .ZN(n19959) );
  OAI21_X1 U23009 ( .B1(n19959), .B2(n20184), .A(n19958), .ZN(n20224) );
  NOR2_X1 U23010 ( .A1(n20224), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19964) );
  AOI221_X1 U23011 ( .B1(n19968), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20006), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19964), .ZN(n19960) );
  INV_X1 U23012 ( .A(n19960), .ZN(n19961) );
  AND2_X1 U23013 ( .A1(n20298), .A2(n19961), .ZN(n19962) );
  INV_X1 U23014 ( .A(n19964), .ZN(n19967) );
  INV_X1 U23015 ( .A(n19965), .ZN(n19985) );
  OAI21_X1 U23016 ( .B1(n10864), .B2(n19985), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19966) );
  AOI22_X1 U23017 ( .A1(n19986), .A2(n20339), .B1(n20338), .B2(n19985), .ZN(
        n19970) );
  AOI22_X1 U23018 ( .A1(n20006), .A2(n20341), .B1(n19968), .B2(n20340), .ZN(
        n19969) );
  OAI211_X1 U23019 ( .C1(n19972), .C2(n19971), .A(n19970), .B(n19969), .ZN(
        P2_U3080) );
  AOI22_X1 U23020 ( .A1(n19986), .A2(n20345), .B1(n20344), .B2(n19985), .ZN(
        n19974) );
  AOI22_X1 U23021 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20347), .ZN(n19973) );
  OAI211_X1 U23022 ( .C1(n20305), .C2(n19990), .A(n19974), .B(n19973), .ZN(
        P2_U3081) );
  AOI22_X1 U23023 ( .A1(n19986), .A2(n20352), .B1(n20351), .B2(n19985), .ZN(
        n19976) );
  AOI22_X1 U23024 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20354), .ZN(n19975) );
  OAI211_X1 U23025 ( .C1(n20308), .C2(n19990), .A(n19976), .B(n19975), .ZN(
        P2_U3082) );
  AOI22_X1 U23026 ( .A1(n19986), .A2(n20358), .B1(n20357), .B2(n19985), .ZN(
        n19978) );
  AOI22_X1 U23027 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20360), .ZN(n19977) );
  OAI211_X1 U23028 ( .C1(n20311), .C2(n19990), .A(n19978), .B(n19977), .ZN(
        P2_U3083) );
  AOI22_X1 U23029 ( .A1(n19986), .A2(n20365), .B1(n20364), .B2(n19985), .ZN(
        n19980) );
  AOI22_X1 U23030 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20367), .ZN(n19979) );
  OAI211_X1 U23031 ( .C1(n20314), .C2(n19990), .A(n19980), .B(n19979), .ZN(
        P2_U3084) );
  AOI22_X1 U23032 ( .A1(n19986), .A2(n20371), .B1(n20370), .B2(n19985), .ZN(
        n19982) );
  AOI22_X1 U23033 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20373), .ZN(n19981) );
  OAI211_X1 U23034 ( .C1(n20317), .C2(n19990), .A(n19982), .B(n19981), .ZN(
        P2_U3085) );
  AOI22_X1 U23035 ( .A1(n19986), .A2(n20377), .B1(n20376), .B2(n19985), .ZN(
        n19984) );
  AOI22_X1 U23036 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20379), .ZN(n19983) );
  OAI211_X1 U23037 ( .C1(n20320), .C2(n19990), .A(n19984), .B(n19983), .ZN(
        P2_U3086) );
  AOI22_X1 U23038 ( .A1(n19986), .A2(n20384), .B1(n20382), .B2(n19985), .ZN(
        n19989) );
  AOI22_X1 U23039 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19987), .B1(
        n20006), .B2(n20388), .ZN(n19988) );
  OAI211_X1 U23040 ( .C1(n20327), .C2(n19990), .A(n19989), .B(n19988), .ZN(
        P2_U3087) );
  AND2_X1 U23041 ( .A1(n20253), .A2(n20060), .ZN(n20033) );
  INV_X1 U23042 ( .A(n20033), .ZN(n20023) );
  OAI22_X1 U23043 ( .A1(n20024), .A2(n20302), .B1(n20023), .B2(n19991), .ZN(
        n19992) );
  INV_X1 U23044 ( .A(n19992), .ZN(n20001) );
  OAI21_X1 U23045 ( .B1(n19993), .B2(n20257), .A(n20484), .ZN(n19999) );
  NOR2_X1 U23046 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20031), .ZN(
        n19996) );
  INV_X1 U23047 ( .A(n10877), .ZN(n19994) );
  OAI211_X1 U23048 ( .C1(n19994), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20478), 
        .B(n20023), .ZN(n19995) );
  OAI211_X1 U23049 ( .C1(n19999), .C2(n19996), .A(n20298), .B(n19995), .ZN(
        n20027) );
  INV_X1 U23050 ( .A(n19996), .ZN(n19998) );
  OAI21_X1 U23051 ( .B1(n10877), .B2(n20033), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19997) );
  AOI22_X1 U23052 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20027), .B1(
        n20339), .B2(n20026), .ZN(n20000) );
  OAI211_X1 U23053 ( .C1(n20265), .C2(n20058), .A(n20001), .B(n20000), .ZN(
        P2_U3088) );
  OAI22_X1 U23054 ( .A1(n20024), .A2(n20305), .B1(n20023), .B2(n20002), .ZN(
        n20003) );
  INV_X1 U23055 ( .A(n20003), .ZN(n20005) );
  AOI22_X1 U23056 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20027), .B1(
        n20345), .B2(n20026), .ZN(n20004) );
  OAI211_X1 U23057 ( .C1(n20268), .C2(n20058), .A(n20005), .B(n20004), .ZN(
        P2_U3089) );
  INV_X1 U23058 ( .A(n20058), .ZN(n20015) );
  AOI22_X1 U23059 ( .A1(n20354), .A2(n20015), .B1(n20351), .B2(n20033), .ZN(
        n20008) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20027), .B1(
        n20352), .B2(n20026), .ZN(n20007) );
  OAI211_X1 U23061 ( .C1(n20308), .C2(n20024), .A(n20008), .B(n20007), .ZN(
        P2_U3090) );
  OAI22_X1 U23062 ( .A1(n20024), .A2(n20311), .B1(n20023), .B2(n20009), .ZN(
        n20010) );
  INV_X1 U23063 ( .A(n20010), .ZN(n20012) );
  AOI22_X1 U23064 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20027), .B1(
        n20358), .B2(n20026), .ZN(n20011) );
  OAI211_X1 U23065 ( .C1(n20274), .C2(n20058), .A(n20012), .B(n20011), .ZN(
        P2_U3091) );
  AOI22_X1 U23066 ( .A1(n20367), .A2(n20015), .B1(n20033), .B2(n20364), .ZN(
        n20014) );
  AOI22_X1 U23067 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20027), .B1(
        n20365), .B2(n20026), .ZN(n20013) );
  OAI211_X1 U23068 ( .C1(n20314), .C2(n20024), .A(n20014), .B(n20013), .ZN(
        P2_U3092) );
  AOI22_X1 U23069 ( .A1(n20373), .A2(n20015), .B1(n20033), .B2(n20370), .ZN(
        n20017) );
  AOI22_X1 U23070 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20027), .B1(
        n20371), .B2(n20026), .ZN(n20016) );
  OAI211_X1 U23071 ( .C1(n20317), .C2(n20024), .A(n20017), .B(n20016), .ZN(
        P2_U3093) );
  OAI22_X1 U23072 ( .A1(n20024), .A2(n20320), .B1(n20023), .B2(n20018), .ZN(
        n20019) );
  INV_X1 U23073 ( .A(n20019), .ZN(n20021) );
  AOI22_X1 U23074 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20027), .B1(
        n20377), .B2(n20026), .ZN(n20020) );
  OAI211_X1 U23075 ( .C1(n20210), .C2(n20058), .A(n20021), .B(n20020), .ZN(
        P2_U3094) );
  INV_X1 U23076 ( .A(n20388), .ZN(n20217) );
  OAI22_X1 U23077 ( .A1(n20024), .A2(n20327), .B1(n20023), .B2(n20022), .ZN(
        n20025) );
  INV_X1 U23078 ( .A(n20025), .ZN(n20029) );
  AOI22_X1 U23079 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20027), .B1(
        n20384), .B2(n20026), .ZN(n20028) );
  OAI211_X1 U23080 ( .C1(n20217), .C2(n20058), .A(n20029), .B(n20028), .ZN(
        P2_U3095) );
  NAND2_X1 U23081 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20060), .ZN(
        n20067) );
  OAI21_X1 U23082 ( .B1(n10876), .B2(n20053), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20030) );
  OAI21_X1 U23083 ( .B1(n20031), .B2(n20290), .A(n20030), .ZN(n20054) );
  AOI22_X1 U23084 ( .A1(n20054), .A2(n20339), .B1(n20338), .B2(n20053), .ZN(
        n20040) );
  AOI21_X1 U23085 ( .B1(n20058), .B2(n20038), .A(n20512), .ZN(n20034) );
  NOR2_X1 U23086 ( .A1(n20034), .A2(n20033), .ZN(n20035) );
  AOI211_X1 U23087 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20036), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20035), .ZN(n20037) );
  OAI21_X1 U23088 ( .B1(n20037), .B2(n20053), .A(n20298), .ZN(n20055) );
  AOI22_X1 U23089 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20341), .ZN(n20039) );
  OAI211_X1 U23090 ( .C1(n20302), .C2(n20058), .A(n20040), .B(n20039), .ZN(
        P2_U3096) );
  AOI22_X1 U23091 ( .A1(n20054), .A2(n20345), .B1(n20344), .B2(n20053), .ZN(
        n20042) );
  AOI22_X1 U23092 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20347), .ZN(n20041) );
  OAI211_X1 U23093 ( .C1(n20305), .C2(n20058), .A(n20042), .B(n20041), .ZN(
        P2_U3097) );
  AOI22_X1 U23094 ( .A1(n20054), .A2(n20352), .B1(n20351), .B2(n20053), .ZN(
        n20044) );
  AOI22_X1 U23095 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20354), .ZN(n20043) );
  OAI211_X1 U23096 ( .C1(n20308), .C2(n20058), .A(n20044), .B(n20043), .ZN(
        P2_U3098) );
  AOI22_X1 U23097 ( .A1(n20054), .A2(n20358), .B1(n20357), .B2(n20053), .ZN(
        n20046) );
  AOI22_X1 U23098 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20360), .ZN(n20045) );
  OAI211_X1 U23099 ( .C1(n20311), .C2(n20058), .A(n20046), .B(n20045), .ZN(
        P2_U3099) );
  AOI22_X1 U23100 ( .A1(n20054), .A2(n20365), .B1(n20364), .B2(n20053), .ZN(
        n20048) );
  AOI22_X1 U23101 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20367), .ZN(n20047) );
  OAI211_X1 U23102 ( .C1(n20314), .C2(n20058), .A(n20048), .B(n20047), .ZN(
        P2_U3100) );
  AOI22_X1 U23103 ( .A1(n20054), .A2(n20371), .B1(n20370), .B2(n20053), .ZN(
        n20050) );
  AOI22_X1 U23104 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20373), .ZN(n20049) );
  OAI211_X1 U23105 ( .C1(n20317), .C2(n20058), .A(n20050), .B(n20049), .ZN(
        P2_U3101) );
  AOI22_X1 U23106 ( .A1(n20054), .A2(n20377), .B1(n20376), .B2(n20053), .ZN(
        n20052) );
  AOI22_X1 U23107 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20379), .ZN(n20051) );
  OAI211_X1 U23108 ( .C1(n20320), .C2(n20058), .A(n20052), .B(n20051), .ZN(
        P2_U3102) );
  AOI22_X1 U23109 ( .A1(n20054), .A2(n20384), .B1(n20382), .B2(n20053), .ZN(
        n20057) );
  AOI22_X1 U23110 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20055), .B1(
        n20086), .B2(n20388), .ZN(n20056) );
  OAI211_X1 U23111 ( .C1(n20327), .C2(n20058), .A(n20057), .B(n20056), .ZN(
        P2_U3103) );
  NAND2_X1 U23112 ( .A1(n20184), .A2(n20060), .ZN(n20095) );
  NOR3_X1 U23113 ( .A1(n20061), .A2(n20098), .A3(n20508), .ZN(n20064) );
  INV_X1 U23114 ( .A(n20067), .ZN(n20062) );
  AOI21_X1 U23115 ( .B1(n12673), .B2(n20062), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20063) );
  AOI22_X1 U23116 ( .A1(n20085), .A2(n20339), .B1(n20098), .B2(n20338), .ZN(
        n20071) );
  INV_X1 U23117 ( .A(n20064), .ZN(n20069) );
  NAND2_X1 U23118 ( .A1(n20066), .A2(n20065), .ZN(n20482) );
  AOI22_X1 U23119 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20095), .B1(n20067), 
        .B2(n20482), .ZN(n20068) );
  NAND3_X1 U23120 ( .A1(n20069), .A2(n20068), .A3(n20298), .ZN(n20087) );
  AOI22_X1 U23121 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n20340), .ZN(n20070) );
  OAI211_X1 U23122 ( .C1(n20265), .C2(n20121), .A(n20071), .B(n20070), .ZN(
        P2_U3104) );
  AOI22_X1 U23123 ( .A1(n20085), .A2(n20345), .B1(n20098), .B2(n20344), .ZN(
        n20073) );
  AOI22_X1 U23124 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n20346), .ZN(n20072) );
  OAI211_X1 U23125 ( .C1(n20268), .C2(n20121), .A(n20073), .B(n20072), .ZN(
        P2_U3105) );
  AOI22_X1 U23126 ( .A1(n20085), .A2(n20352), .B1(n20351), .B2(n20098), .ZN(
        n20075) );
  AOI22_X1 U23127 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n20353), .ZN(n20074) );
  OAI211_X1 U23128 ( .C1(n20271), .C2(n20121), .A(n20075), .B(n20074), .ZN(
        P2_U3106) );
  AOI22_X1 U23129 ( .A1(n20085), .A2(n20358), .B1(n20098), .B2(n20357), .ZN(
        n20077) );
  AOI22_X1 U23130 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n20359), .ZN(n20076) );
  OAI211_X1 U23131 ( .C1(n20274), .C2(n20121), .A(n20077), .B(n20076), .ZN(
        P2_U3107) );
  AOI22_X1 U23132 ( .A1(n20085), .A2(n20365), .B1(n20098), .B2(n20364), .ZN(
        n20079) );
  INV_X1 U23133 ( .A(n20121), .ZN(n20082) );
  AOI22_X1 U23134 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20087), .B1(
        n20082), .B2(n20367), .ZN(n20078) );
  OAI211_X1 U23135 ( .C1(n20314), .C2(n20038), .A(n20079), .B(n20078), .ZN(
        P2_U3108) );
  AOI22_X1 U23136 ( .A1(n20085), .A2(n20371), .B1(n20098), .B2(n20370), .ZN(
        n20081) );
  AOI22_X1 U23137 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20087), .B1(
        n20082), .B2(n20373), .ZN(n20080) );
  OAI211_X1 U23138 ( .C1(n20317), .C2(n20038), .A(n20081), .B(n20080), .ZN(
        P2_U3109) );
  AOI22_X1 U23139 ( .A1(n20085), .A2(n20377), .B1(n20098), .B2(n20376), .ZN(
        n20084) );
  AOI22_X1 U23140 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20087), .B1(
        n20082), .B2(n20379), .ZN(n20083) );
  OAI211_X1 U23141 ( .C1(n20320), .C2(n20038), .A(n20084), .B(n20083), .ZN(
        P2_U3110) );
  AOI22_X1 U23142 ( .A1(n20085), .A2(n20384), .B1(n20098), .B2(n20382), .ZN(
        n20089) );
  AOI22_X1 U23143 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n20386), .ZN(n20088) );
  OAI211_X1 U23144 ( .C1(n20217), .C2(n20121), .A(n20089), .B(n20088), .ZN(
        P2_U3111) );
  NAND2_X1 U23145 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20497), .ZN(
        n20189) );
  NOR2_X1 U23146 ( .A1(n20219), .A2(n20189), .ZN(n20116) );
  AOI22_X1 U23147 ( .A1(n20341), .A2(n20145), .B1(n20116), .B2(n20338), .ZN(
        n20103) );
  NAND2_X1 U23148 ( .A1(n20484), .A2(n20121), .ZN(n20093) );
  INV_X1 U23149 ( .A(n20091), .ZN(n20092) );
  OAI21_X1 U23150 ( .B1(n20145), .B2(n20093), .A(n20092), .ZN(n20097) );
  OAI21_X1 U23151 ( .B1(n20099), .B2(n20508), .A(n12673), .ZN(n20094) );
  AOI21_X1 U23152 ( .B1(n20097), .B2(n20095), .A(n20094), .ZN(n20096) );
  OAI21_X1 U23153 ( .B1(n20116), .B2(n20098), .A(n20097), .ZN(n20101) );
  OAI21_X1 U23154 ( .B1(n20099), .B2(n20116), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20100) );
  AOI22_X1 U23155 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20118), .B1(
        n20339), .B2(n20117), .ZN(n20102) );
  OAI211_X1 U23156 ( .C1(n20302), .C2(n20121), .A(n20103), .B(n20102), .ZN(
        P2_U3112) );
  AOI22_X1 U23157 ( .A1(n20347), .A2(n20145), .B1(n20116), .B2(n20344), .ZN(
        n20105) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20345), .ZN(n20104) );
  OAI211_X1 U23159 ( .C1(n20305), .C2(n20121), .A(n20105), .B(n20104), .ZN(
        P2_U3113) );
  AOI22_X1 U23160 ( .A1(n20354), .A2(n20145), .B1(n20351), .B2(n20116), .ZN(
        n20107) );
  AOI22_X1 U23161 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20352), .ZN(n20106) );
  OAI211_X1 U23162 ( .C1(n20308), .C2(n20121), .A(n20107), .B(n20106), .ZN(
        P2_U3114) );
  AOI22_X1 U23163 ( .A1(n20360), .A2(n20145), .B1(n20116), .B2(n20357), .ZN(
        n20109) );
  AOI22_X1 U23164 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20358), .ZN(n20108) );
  OAI211_X1 U23165 ( .C1(n20311), .C2(n20121), .A(n20109), .B(n20108), .ZN(
        P2_U3115) );
  AOI22_X1 U23166 ( .A1(n20367), .A2(n20145), .B1(n20116), .B2(n20364), .ZN(
        n20111) );
  AOI22_X1 U23167 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20365), .ZN(n20110) );
  OAI211_X1 U23168 ( .C1(n20314), .C2(n20121), .A(n20111), .B(n20110), .ZN(
        P2_U3116) );
  AOI22_X1 U23169 ( .A1(n20373), .A2(n20145), .B1(n20116), .B2(n20370), .ZN(
        n20113) );
  AOI22_X1 U23170 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20371), .ZN(n20112) );
  OAI211_X1 U23171 ( .C1(n20317), .C2(n20121), .A(n20113), .B(n20112), .ZN(
        P2_U3117) );
  AOI22_X1 U23172 ( .A1(n20145), .A2(n20379), .B1(n20116), .B2(n20376), .ZN(
        n20115) );
  AOI22_X1 U23173 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20377), .ZN(n20114) );
  OAI211_X1 U23174 ( .C1(n20320), .C2(n20121), .A(n20115), .B(n20114), .ZN(
        P2_U3118) );
  AOI22_X1 U23175 ( .A1(n20388), .A2(n20145), .B1(n20116), .B2(n20382), .ZN(
        n20120) );
  AOI22_X1 U23176 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20118), .B1(
        n20117), .B2(n20384), .ZN(n20119) );
  OAI211_X1 U23177 ( .C1(n20327), .C2(n20121), .A(n20120), .B(n20119), .ZN(
        P2_U3119) );
  INV_X1 U23178 ( .A(n20189), .ZN(n20183) );
  AOI22_X1 U23179 ( .A1(n20145), .A2(n20340), .B1(n20158), .B2(n20338), .ZN(
        n20134) );
  OR2_X1 U23180 ( .A1(n20124), .A2(n20512), .ZN(n20332) );
  OAI21_X1 U23181 ( .B1(n20332), .B2(n20125), .A(n20484), .ZN(n20132) );
  NOR2_X1 U23182 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20189), .ZN(
        n20128) );
  INV_X1 U23183 ( .A(n20158), .ZN(n20126) );
  OAI211_X1 U23184 ( .C1(n10868), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20478), 
        .B(n20126), .ZN(n20127) );
  OAI211_X1 U23185 ( .C1(n20132), .C2(n20128), .A(n20298), .B(n20127), .ZN(
        n20150) );
  INV_X1 U23186 ( .A(n20128), .ZN(n20131) );
  INV_X1 U23187 ( .A(n10868), .ZN(n20129) );
  OAI21_X1 U23188 ( .B1(n20129), .B2(n20158), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20130) );
  AOI22_X1 U23189 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20150), .B1(
        n20339), .B2(n20149), .ZN(n20133) );
  OAI211_X1 U23190 ( .C1(n20265), .C2(n20182), .A(n20134), .B(n20133), .ZN(
        P2_U3120) );
  AOI22_X1 U23191 ( .A1(n20145), .A2(n20346), .B1(n20158), .B2(n20344), .ZN(
        n20136) );
  AOI22_X1 U23192 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20150), .B1(
        n20345), .B2(n20149), .ZN(n20135) );
  OAI211_X1 U23193 ( .C1(n20268), .C2(n20182), .A(n20136), .B(n20135), .ZN(
        P2_U3121) );
  AOI22_X1 U23194 ( .A1(n20145), .A2(n20353), .B1(n20158), .B2(n20351), .ZN(
        n20138) );
  AOI22_X1 U23195 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20150), .B1(
        n20352), .B2(n20149), .ZN(n20137) );
  OAI211_X1 U23196 ( .C1(n20271), .C2(n20182), .A(n20138), .B(n20137), .ZN(
        P2_U3122) );
  AOI22_X1 U23197 ( .A1(n20145), .A2(n20359), .B1(n20158), .B2(n20357), .ZN(
        n20140) );
  AOI22_X1 U23198 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20150), .B1(
        n20358), .B2(n20149), .ZN(n20139) );
  OAI211_X1 U23199 ( .C1(n20274), .C2(n20182), .A(n20140), .B(n20139), .ZN(
        P2_U3123) );
  INV_X1 U23200 ( .A(n20145), .ZN(n20153) );
  INV_X1 U23201 ( .A(n20182), .ZN(n20148) );
  AOI22_X1 U23202 ( .A1(n20367), .A2(n20148), .B1(n20158), .B2(n20364), .ZN(
        n20142) );
  AOI22_X1 U23203 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20150), .B1(
        n20365), .B2(n20149), .ZN(n20141) );
  OAI211_X1 U23204 ( .C1(n20314), .C2(n20153), .A(n20142), .B(n20141), .ZN(
        P2_U3124) );
  AOI22_X1 U23205 ( .A1(n20373), .A2(n20148), .B1(n20158), .B2(n20370), .ZN(
        n20144) );
  AOI22_X1 U23206 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20150), .B1(
        n20371), .B2(n20149), .ZN(n20143) );
  OAI211_X1 U23207 ( .C1(n20317), .C2(n20153), .A(n20144), .B(n20143), .ZN(
        P2_U3125) );
  AOI22_X1 U23208 ( .A1(n20145), .A2(n20378), .B1(n20158), .B2(n20376), .ZN(
        n20147) );
  AOI22_X1 U23209 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20150), .B1(
        n20377), .B2(n20149), .ZN(n20146) );
  OAI211_X1 U23210 ( .C1(n20210), .C2(n20182), .A(n20147), .B(n20146), .ZN(
        P2_U3126) );
  AOI22_X1 U23211 ( .A1(n20388), .A2(n20148), .B1(n20158), .B2(n20382), .ZN(
        n20152) );
  AOI22_X1 U23212 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20150), .B1(
        n20384), .B2(n20149), .ZN(n20151) );
  OAI211_X1 U23213 ( .C1(n20327), .C2(n20153), .A(n20152), .B(n20151), .ZN(
        P2_U3127) );
  OAI21_X1 U23214 ( .B1(n20156), .B2(n20177), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20155) );
  OAI21_X1 U23215 ( .B1(n20189), .B2(n20290), .A(n20155), .ZN(n20178) );
  AOI22_X1 U23216 ( .A1(n20178), .A2(n20339), .B1(n20177), .B2(n20338), .ZN(
        n20164) );
  INV_X1 U23217 ( .A(n20156), .ZN(n20161) );
  NOR2_X4 U23218 ( .A1(n20292), .A2(n20190), .ZN(n20213) );
  INV_X1 U23219 ( .A(n20213), .ZN(n20157) );
  AOI21_X1 U23220 ( .B1(n20157), .B2(n20182), .A(n20512), .ZN(n20159) );
  NOR2_X1 U23221 ( .A1(n20159), .A2(n20158), .ZN(n20160) );
  AOI211_X1 U23222 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20161), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20160), .ZN(n20162) );
  OAI21_X1 U23223 ( .B1(n20162), .B2(n20177), .A(n20298), .ZN(n20179) );
  AOI22_X1 U23224 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20341), .ZN(n20163) );
  OAI211_X1 U23225 ( .C1(n20302), .C2(n20182), .A(n20164), .B(n20163), .ZN(
        P2_U3128) );
  AOI22_X1 U23226 ( .A1(n20178), .A2(n20345), .B1(n20177), .B2(n20344), .ZN(
        n20166) );
  AOI22_X1 U23227 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20347), .ZN(n20165) );
  OAI211_X1 U23228 ( .C1(n20305), .C2(n20182), .A(n20166), .B(n20165), .ZN(
        P2_U3129) );
  AOI22_X1 U23229 ( .A1(n20178), .A2(n20352), .B1(n20351), .B2(n20177), .ZN(
        n20168) );
  AOI22_X1 U23230 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20354), .ZN(n20167) );
  OAI211_X1 U23231 ( .C1(n20308), .C2(n20182), .A(n20168), .B(n20167), .ZN(
        P2_U3130) );
  AOI22_X1 U23232 ( .A1(n20178), .A2(n20358), .B1(n20177), .B2(n20357), .ZN(
        n20170) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20360), .ZN(n20169) );
  OAI211_X1 U23234 ( .C1(n20311), .C2(n20182), .A(n20170), .B(n20169), .ZN(
        P2_U3131) );
  AOI22_X1 U23235 ( .A1(n20178), .A2(n20365), .B1(n20177), .B2(n20364), .ZN(
        n20172) );
  AOI22_X1 U23236 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20367), .ZN(n20171) );
  OAI211_X1 U23237 ( .C1(n20314), .C2(n20182), .A(n20172), .B(n20171), .ZN(
        P2_U3132) );
  AOI22_X1 U23238 ( .A1(n20178), .A2(n20371), .B1(n20177), .B2(n20370), .ZN(
        n20174) );
  AOI22_X1 U23239 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20373), .ZN(n20173) );
  OAI211_X1 U23240 ( .C1(n20317), .C2(n20182), .A(n20174), .B(n20173), .ZN(
        P2_U3133) );
  AOI22_X1 U23241 ( .A1(n20178), .A2(n20377), .B1(n20177), .B2(n20376), .ZN(
        n20176) );
  AOI22_X1 U23242 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20379), .ZN(n20175) );
  OAI211_X1 U23243 ( .C1(n20320), .C2(n20182), .A(n20176), .B(n20175), .ZN(
        P2_U3134) );
  AOI22_X1 U23244 ( .A1(n20178), .A2(n20384), .B1(n20177), .B2(n20382), .ZN(
        n20181) );
  AOI22_X1 U23245 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20179), .B1(
        n20213), .B2(n20388), .ZN(n20180) );
  OAI211_X1 U23246 ( .C1(n20327), .C2(n20182), .A(n20181), .B(n20180), .ZN(
        P2_U3135) );
  NAND3_X1 U23247 ( .A1(n12673), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n20183), .ZN(n20188) );
  NAND2_X1 U23248 ( .A1(n20184), .A2(n20183), .ZN(n20191) );
  AND2_X1 U23249 ( .A1(n20191), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20185) );
  NAND2_X1 U23250 ( .A1(n20186), .A2(n20185), .ZN(n20193) );
  INV_X1 U23251 ( .A(n20193), .ZN(n20187) );
  INV_X1 U23252 ( .A(n20191), .ZN(n20211) );
  AOI22_X1 U23253 ( .A1(n20212), .A2(n20339), .B1(n20338), .B2(n20211), .ZN(
        n20196) );
  OAI22_X1 U23254 ( .A1(n20332), .A2(n20190), .B1(n20189), .B2(n20252), .ZN(
        n20194) );
  NAND2_X1 U23255 ( .A1(n20191), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20192) );
  NAND4_X1 U23256 ( .A1(n20194), .A2(n20298), .A3(n20193), .A4(n20192), .ZN(
        n20214) );
  AOI22_X1 U23257 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20340), .ZN(n20195) );
  OAI211_X1 U23258 ( .C1(n20265), .C2(n20249), .A(n20196), .B(n20195), .ZN(
        P2_U3136) );
  AOI22_X1 U23259 ( .A1(n20212), .A2(n20345), .B1(n20344), .B2(n20211), .ZN(
        n20198) );
  AOI22_X1 U23260 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20346), .ZN(n20197) );
  OAI211_X1 U23261 ( .C1(n20268), .C2(n20249), .A(n20198), .B(n20197), .ZN(
        P2_U3137) );
  AOI22_X1 U23262 ( .A1(n20212), .A2(n20352), .B1(n20351), .B2(n20211), .ZN(
        n20200) );
  AOI22_X1 U23263 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20353), .ZN(n20199) );
  OAI211_X1 U23264 ( .C1(n20271), .C2(n20249), .A(n20200), .B(n20199), .ZN(
        P2_U3138) );
  AOI22_X1 U23265 ( .A1(n20212), .A2(n20358), .B1(n20357), .B2(n20211), .ZN(
        n20202) );
  AOI22_X1 U23266 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20359), .ZN(n20201) );
  OAI211_X1 U23267 ( .C1(n20274), .C2(n20249), .A(n20202), .B(n20201), .ZN(
        P2_U3139) );
  AOI22_X1 U23268 ( .A1(n20212), .A2(n20365), .B1(n20364), .B2(n20211), .ZN(
        n20204) );
  INV_X1 U23269 ( .A(n20249), .ZN(n20222) );
  AOI22_X1 U23270 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20214), .B1(
        n20222), .B2(n20367), .ZN(n20203) );
  OAI211_X1 U23271 ( .C1(n20314), .C2(n20157), .A(n20204), .B(n20203), .ZN(
        P2_U3140) );
  AOI22_X1 U23272 ( .A1(n20212), .A2(n20371), .B1(n20370), .B2(n20211), .ZN(
        n20206) );
  AOI22_X1 U23273 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20372), .ZN(n20205) );
  OAI211_X1 U23274 ( .C1(n20207), .C2(n20249), .A(n20206), .B(n20205), .ZN(
        P2_U3141) );
  AOI22_X1 U23275 ( .A1(n20212), .A2(n20377), .B1(n20376), .B2(n20211), .ZN(
        n20209) );
  AOI22_X1 U23276 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20378), .ZN(n20208) );
  OAI211_X1 U23277 ( .C1(n20210), .C2(n20249), .A(n20209), .B(n20208), .ZN(
        P2_U3142) );
  AOI22_X1 U23278 ( .A1(n20212), .A2(n20384), .B1(n20382), .B2(n20211), .ZN(
        n20216) );
  AOI22_X1 U23279 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20214), .B1(
        n20213), .B2(n20386), .ZN(n20215) );
  OAI211_X1 U23280 ( .C1(n20217), .C2(n20249), .A(n20216), .B(n20215), .ZN(
        P2_U3143) );
  INV_X1 U23281 ( .A(n20218), .ZN(n20221) );
  INV_X1 U23282 ( .A(n20288), .ZN(n20291) );
  OR2_X1 U23283 ( .A1(n20219), .A2(n20291), .ZN(n20226) );
  INV_X1 U23284 ( .A(n20226), .ZN(n20244) );
  OAI21_X1 U23285 ( .B1(n20225), .B2(n20244), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20220) );
  AOI22_X1 U23286 ( .A1(n20245), .A2(n20339), .B1(n20244), .B2(n20338), .ZN(
        n20231) );
  NOR2_X2 U23287 ( .A1(n20292), .A2(n20257), .ZN(n20275) );
  OAI21_X1 U23288 ( .B1(n20222), .B2(n20275), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20223) );
  OAI21_X1 U23289 ( .B1(n21570), .B2(n20224), .A(n20223), .ZN(n20229) );
  INV_X1 U23290 ( .A(n20225), .ZN(n20227) );
  OAI211_X1 U23291 ( .C1(n20227), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20478), 
        .B(n20226), .ZN(n20228) );
  NAND3_X1 U23292 ( .A1(n20229), .A2(n20298), .A3(n20228), .ZN(n20246) );
  AOI22_X1 U23293 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20341), .ZN(n20230) );
  OAI211_X1 U23294 ( .C1(n20302), .C2(n20249), .A(n20231), .B(n20230), .ZN(
        P2_U3144) );
  AOI22_X1 U23295 ( .A1(n20245), .A2(n20345), .B1(n20244), .B2(n20344), .ZN(
        n20233) );
  AOI22_X1 U23296 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20347), .ZN(n20232) );
  OAI211_X1 U23297 ( .C1(n20305), .C2(n20249), .A(n20233), .B(n20232), .ZN(
        P2_U3145) );
  AOI22_X1 U23298 ( .A1(n20245), .A2(n20352), .B1(n20244), .B2(n20351), .ZN(
        n20235) );
  AOI22_X1 U23299 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20354), .ZN(n20234) );
  OAI211_X1 U23300 ( .C1(n20308), .C2(n20249), .A(n20235), .B(n20234), .ZN(
        P2_U3146) );
  AOI22_X1 U23301 ( .A1(n20245), .A2(n20358), .B1(n20244), .B2(n20357), .ZN(
        n20237) );
  AOI22_X1 U23302 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20360), .ZN(n20236) );
  OAI211_X1 U23303 ( .C1(n20311), .C2(n20249), .A(n20237), .B(n20236), .ZN(
        P2_U3147) );
  AOI22_X1 U23304 ( .A1(n20245), .A2(n20365), .B1(n20244), .B2(n20364), .ZN(
        n20239) );
  AOI22_X1 U23305 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20367), .ZN(n20238) );
  OAI211_X1 U23306 ( .C1(n20314), .C2(n20249), .A(n20239), .B(n20238), .ZN(
        P2_U3148) );
  AOI22_X1 U23307 ( .A1(n20245), .A2(n20371), .B1(n20244), .B2(n20370), .ZN(
        n20241) );
  AOI22_X1 U23308 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20373), .ZN(n20240) );
  OAI211_X1 U23309 ( .C1(n20317), .C2(n20249), .A(n20241), .B(n20240), .ZN(
        P2_U3149) );
  AOI22_X1 U23310 ( .A1(n20245), .A2(n20377), .B1(n20244), .B2(n20376), .ZN(
        n20243) );
  AOI22_X1 U23311 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20379), .ZN(n20242) );
  OAI211_X1 U23312 ( .C1(n20320), .C2(n20249), .A(n20243), .B(n20242), .ZN(
        P2_U3150) );
  AOI22_X1 U23313 ( .A1(n20245), .A2(n20384), .B1(n20244), .B2(n20382), .ZN(
        n20248) );
  AOI22_X1 U23314 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20246), .B1(
        n20275), .B2(n20388), .ZN(n20247) );
  OAI211_X1 U23315 ( .C1(n20327), .C2(n20249), .A(n20248), .B(n20247), .ZN(
        P2_U3151) );
  NAND2_X1 U23316 ( .A1(n20252), .A2(n20288), .ZN(n20258) );
  INV_X1 U23317 ( .A(n20294), .ZN(n20254) );
  NAND3_X1 U23318 ( .A1(n10870), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20254), 
        .ZN(n20260) );
  INV_X1 U23319 ( .A(n20260), .ZN(n20255) );
  AOI211_X2 U23320 ( .C1(n20508), .C2(n20258), .A(n20256), .B(n20255), .ZN(
        n20282) );
  AOI22_X1 U23321 ( .A1(n20282), .A2(n20339), .B1(n20294), .B2(n20338), .ZN(
        n20264) );
  NOR3_X1 U23322 ( .A1(n20332), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n20257), 
        .ZN(n20262) );
  NOR2_X1 U23323 ( .A1(n20259), .A2(n20258), .ZN(n20261) );
  OAI211_X1 U23324 ( .C1(n20262), .C2(n20261), .A(n20298), .B(n20260), .ZN(
        n20284) );
  AOI22_X1 U23325 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20284), .B1(
        n20275), .B2(n20340), .ZN(n20263) );
  OAI211_X1 U23326 ( .C1(n20265), .C2(n20326), .A(n20264), .B(n20263), .ZN(
        P2_U3152) );
  AOI22_X1 U23327 ( .A1(n20282), .A2(n20345), .B1(n20294), .B2(n20344), .ZN(
        n20267) );
  AOI22_X1 U23328 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20284), .B1(
        n20275), .B2(n20346), .ZN(n20266) );
  OAI211_X1 U23329 ( .C1(n20268), .C2(n20326), .A(n20267), .B(n20266), .ZN(
        P2_U3153) );
  AOI22_X1 U23330 ( .A1(n20282), .A2(n20352), .B1(n20351), .B2(n20294), .ZN(
        n20270) );
  AOI22_X1 U23331 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20284), .B1(
        n20275), .B2(n20353), .ZN(n20269) );
  OAI211_X1 U23332 ( .C1(n20271), .C2(n20326), .A(n20270), .B(n20269), .ZN(
        P2_U3154) );
  AOI22_X1 U23333 ( .A1(n20282), .A2(n20358), .B1(n20294), .B2(n20357), .ZN(
        n20273) );
  AOI22_X1 U23334 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20284), .B1(
        n20275), .B2(n20359), .ZN(n20272) );
  OAI211_X1 U23335 ( .C1(n20274), .C2(n20326), .A(n20273), .B(n20272), .ZN(
        P2_U3155) );
  INV_X1 U23336 ( .A(n20275), .ZN(n20287) );
  AOI22_X1 U23337 ( .A1(n20282), .A2(n20365), .B1(n20294), .B2(n20364), .ZN(
        n20277) );
  INV_X1 U23338 ( .A(n20326), .ZN(n20283) );
  AOI22_X1 U23339 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20367), .ZN(n20276) );
  OAI211_X1 U23340 ( .C1(n20314), .C2(n20287), .A(n20277), .B(n20276), .ZN(
        P2_U3156) );
  AOI22_X1 U23341 ( .A1(n20282), .A2(n20371), .B1(n20294), .B2(n20370), .ZN(
        n20279) );
  AOI22_X1 U23342 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20373), .ZN(n20278) );
  OAI211_X1 U23343 ( .C1(n20317), .C2(n20287), .A(n20279), .B(n20278), .ZN(
        P2_U3157) );
  AOI22_X1 U23344 ( .A1(n20282), .A2(n20377), .B1(n20294), .B2(n20376), .ZN(
        n20281) );
  AOI22_X1 U23345 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20379), .ZN(n20280) );
  OAI211_X1 U23346 ( .C1(n20320), .C2(n20287), .A(n20281), .B(n20280), .ZN(
        P2_U3158) );
  AOI22_X1 U23347 ( .A1(n20282), .A2(n20384), .B1(n20294), .B2(n20382), .ZN(
        n20286) );
  AOI22_X1 U23348 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20388), .ZN(n20285) );
  OAI211_X1 U23349 ( .C1(n20327), .C2(n20287), .A(n20286), .B(n20285), .ZN(
        P2_U3159) );
  NAND2_X1 U23350 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20288), .ZN(
        n20334) );
  OAI21_X1 U23351 ( .B1(n10866), .B2(n20321), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20289) );
  OAI21_X1 U23352 ( .B1(n20291), .B2(n20290), .A(n20289), .ZN(n20322) );
  AOI22_X1 U23353 ( .A1(n20322), .A2(n20339), .B1(n20338), .B2(n20321), .ZN(
        n20301) );
  INV_X1 U23354 ( .A(n10866), .ZN(n20297) );
  NOR2_X4 U23355 ( .A1(n20292), .A2(n20333), .ZN(n20387) );
  INV_X1 U23356 ( .A(n20387), .ZN(n20293) );
  AOI21_X1 U23357 ( .B1(n20293), .B2(n20326), .A(n20512), .ZN(n20295) );
  NOR2_X1 U23358 ( .A1(n20295), .A2(n20294), .ZN(n20296) );
  AOI211_X1 U23359 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20297), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20296), .ZN(n20299) );
  OAI21_X1 U23360 ( .B1(n20299), .B2(n20321), .A(n20298), .ZN(n20323) );
  AOI22_X1 U23361 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20341), .ZN(n20300) );
  OAI211_X1 U23362 ( .C1(n20302), .C2(n20326), .A(n20301), .B(n20300), .ZN(
        P2_U3160) );
  AOI22_X1 U23363 ( .A1(n20322), .A2(n20345), .B1(n20344), .B2(n20321), .ZN(
        n20304) );
  AOI22_X1 U23364 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20347), .ZN(n20303) );
  OAI211_X1 U23365 ( .C1(n20305), .C2(n20326), .A(n20304), .B(n20303), .ZN(
        P2_U3161) );
  AOI22_X1 U23366 ( .A1(n20322), .A2(n20352), .B1(n20351), .B2(n20321), .ZN(
        n20307) );
  AOI22_X1 U23367 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20354), .ZN(n20306) );
  OAI211_X1 U23368 ( .C1(n20308), .C2(n20326), .A(n20307), .B(n20306), .ZN(
        P2_U3162) );
  AOI22_X1 U23369 ( .A1(n20322), .A2(n20358), .B1(n20357), .B2(n20321), .ZN(
        n20310) );
  AOI22_X1 U23370 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20360), .ZN(n20309) );
  OAI211_X1 U23371 ( .C1(n20311), .C2(n20326), .A(n20310), .B(n20309), .ZN(
        P2_U3163) );
  AOI22_X1 U23372 ( .A1(n20322), .A2(n20365), .B1(n20364), .B2(n20321), .ZN(
        n20313) );
  AOI22_X1 U23373 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20367), .ZN(n20312) );
  OAI211_X1 U23374 ( .C1(n20314), .C2(n20326), .A(n20313), .B(n20312), .ZN(
        P2_U3164) );
  AOI22_X1 U23375 ( .A1(n20322), .A2(n20371), .B1(n20370), .B2(n20321), .ZN(
        n20316) );
  AOI22_X1 U23376 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20373), .ZN(n20315) );
  OAI211_X1 U23377 ( .C1(n20317), .C2(n20326), .A(n20316), .B(n20315), .ZN(
        P2_U3165) );
  AOI22_X1 U23378 ( .A1(n20322), .A2(n20377), .B1(n20376), .B2(n20321), .ZN(
        n20319) );
  AOI22_X1 U23379 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20379), .ZN(n20318) );
  OAI211_X1 U23380 ( .C1(n20320), .C2(n20326), .A(n20319), .B(n20318), .ZN(
        P2_U3166) );
  AOI22_X1 U23381 ( .A1(n20322), .A2(n20384), .B1(n20382), .B2(n20321), .ZN(
        n20325) );
  AOI22_X1 U23382 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20323), .B1(
        n20387), .B2(n20388), .ZN(n20324) );
  OAI211_X1 U23383 ( .C1(n20327), .C2(n20326), .A(n20325), .B(n20324), .ZN(
        P2_U3167) );
  INV_X1 U23384 ( .A(n20328), .ZN(n20383) );
  NOR3_X1 U23385 ( .A1(n20329), .A2(n20383), .A3(n20508), .ZN(n20337) );
  INV_X1 U23386 ( .A(n20337), .ZN(n20330) );
  OAI211_X1 U23387 ( .C1(n20383), .C2(n12673), .A(n20330), .B(n20298), .ZN(
        n20331) );
  INV_X1 U23388 ( .A(n20334), .ZN(n20335) );
  AOI21_X1 U23389 ( .B1(n12673), .B2(n20335), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20336) );
  AOI22_X1 U23390 ( .A1(n20385), .A2(n20339), .B1(n20383), .B2(n20338), .ZN(
        n20343) );
  AOI22_X1 U23391 ( .A1(n20389), .A2(n20341), .B1(n20387), .B2(n20340), .ZN(
        n20342) );
  OAI211_X1 U23392 ( .C1(n20392), .C2(n12705), .A(n20343), .B(n20342), .ZN(
        P2_U3168) );
  INV_X1 U23393 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20350) );
  AOI22_X1 U23394 ( .A1(n20385), .A2(n20345), .B1(n20383), .B2(n20344), .ZN(
        n20349) );
  AOI22_X1 U23395 ( .A1(n20389), .A2(n20347), .B1(n20387), .B2(n20346), .ZN(
        n20348) );
  OAI211_X1 U23396 ( .C1(n20392), .C2(n20350), .A(n20349), .B(n20348), .ZN(
        P2_U3169) );
  AOI22_X1 U23397 ( .A1(n20385), .A2(n20352), .B1(n20383), .B2(n20351), .ZN(
        n20356) );
  AOI22_X1 U23398 ( .A1(n20389), .A2(n20354), .B1(n20387), .B2(n20353), .ZN(
        n20355) );
  OAI211_X1 U23399 ( .C1(n20392), .C2(n12739), .A(n20356), .B(n20355), .ZN(
        P2_U3170) );
  INV_X1 U23400 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20363) );
  AOI22_X1 U23401 ( .A1(n20385), .A2(n20358), .B1(n20383), .B2(n20357), .ZN(
        n20362) );
  AOI22_X1 U23402 ( .A1(n20389), .A2(n20360), .B1(n20387), .B2(n20359), .ZN(
        n20361) );
  OAI211_X1 U23403 ( .C1(n20392), .C2(n20363), .A(n20362), .B(n20361), .ZN(
        P2_U3171) );
  AOI22_X1 U23404 ( .A1(n20385), .A2(n20365), .B1(n20383), .B2(n20364), .ZN(
        n20369) );
  AOI22_X1 U23405 ( .A1(n20389), .A2(n20367), .B1(n20387), .B2(n20366), .ZN(
        n20368) );
  OAI211_X1 U23406 ( .C1(n20392), .C2(n12773), .A(n20369), .B(n20368), .ZN(
        P2_U3172) );
  AOI22_X1 U23407 ( .A1(n20385), .A2(n20371), .B1(n20383), .B2(n20370), .ZN(
        n20375) );
  AOI22_X1 U23408 ( .A1(n20389), .A2(n20373), .B1(n20387), .B2(n20372), .ZN(
        n20374) );
  OAI211_X1 U23409 ( .C1(n20392), .C2(n12807), .A(n20375), .B(n20374), .ZN(
        P2_U3173) );
  AOI22_X1 U23410 ( .A1(n20385), .A2(n20377), .B1(n20383), .B2(n20376), .ZN(
        n20381) );
  AOI22_X1 U23411 ( .A1(n20389), .A2(n20379), .B1(n20387), .B2(n20378), .ZN(
        n20380) );
  OAI211_X1 U23412 ( .C1(n20392), .C2(n12790), .A(n20381), .B(n20380), .ZN(
        P2_U3174) );
  AOI22_X1 U23413 ( .A1(n20385), .A2(n20384), .B1(n20383), .B2(n20382), .ZN(
        n20391) );
  AOI22_X1 U23414 ( .A1(n20389), .A2(n20388), .B1(n20387), .B2(n20386), .ZN(
        n20390) );
  OAI211_X1 U23415 ( .C1(n20392), .C2(n12992), .A(n20391), .B(n20390), .ZN(
        P2_U3175) );
  AND2_X1 U23416 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20393), .ZN(
        P2_U3179) );
  NOR2_X1 U23417 ( .A1(n21743), .A2(n20475), .ZN(P2_U3180) );
  AND2_X1 U23418 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20393), .ZN(
        P2_U3181) );
  AND2_X1 U23419 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20393), .ZN(
        P2_U3182) );
  AND2_X1 U23420 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20393), .ZN(
        P2_U3183) );
  AND2_X1 U23421 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20393), .ZN(
        P2_U3184) );
  AND2_X1 U23422 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20393), .ZN(
        P2_U3185) );
  AND2_X1 U23423 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20393), .ZN(
        P2_U3186) );
  AND2_X1 U23424 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20393), .ZN(
        P2_U3187) );
  AND2_X1 U23425 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20393), .ZN(
        P2_U3188) );
  AND2_X1 U23426 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20393), .ZN(
        P2_U3189) );
  AND2_X1 U23427 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20393), .ZN(
        P2_U3190) );
  AND2_X1 U23428 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20393), .ZN(
        P2_U3191) );
  AND2_X1 U23429 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20393), .ZN(
        P2_U3192) );
  AND2_X1 U23430 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20393), .ZN(
        P2_U3193) );
  AND2_X1 U23431 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20393), .ZN(
        P2_U3194) );
  AND2_X1 U23432 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20393), .ZN(
        P2_U3195) );
  NOR2_X1 U23433 ( .A1(n21662), .A2(n20475), .ZN(P2_U3196) );
  AND2_X1 U23434 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20393), .ZN(
        P2_U3197) );
  AND2_X1 U23435 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20393), .ZN(
        P2_U3198) );
  AND2_X1 U23436 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20393), .ZN(
        P2_U3199) );
  AND2_X1 U23437 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20393), .ZN(
        P2_U3200) );
  AND2_X1 U23438 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20393), .ZN(P2_U3201) );
  AND2_X1 U23439 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20393), .ZN(P2_U3202) );
  INV_X1 U23440 ( .A(P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n21759) );
  NOR2_X1 U23441 ( .A1(n21759), .A2(n20475), .ZN(P2_U3203) );
  AND2_X1 U23442 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20393), .ZN(P2_U3204) );
  AND2_X1 U23443 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20393), .ZN(P2_U3205) );
  AND2_X1 U23444 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20393), .ZN(P2_U3206) );
  AND2_X1 U23445 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20393), .ZN(P2_U3207) );
  AND2_X1 U23446 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20393), .ZN(P2_U3208) );
  NOR2_X1 U23447 ( .A1(n20394), .A2(n20520), .ZN(n20405) );
  INV_X1 U23448 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20399) );
  NOR3_X1 U23449 ( .A1(n20405), .A2(n20399), .A3(n20395), .ZN(n20398) );
  OAI211_X1 U23450 ( .C1(HOLD), .C2(n20399), .A(n20526), .B(n20407), .ZN(
        n20397) );
  NOR2_X1 U23451 ( .A1(n21377), .A2(n20400), .ZN(n20411) );
  INV_X1 U23452 ( .A(n20411), .ZN(n20396) );
  OAI211_X1 U23453 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20398), .A(n20397), 
        .B(n20396), .ZN(P2_U3209) );
  AOI21_X1 U23454 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21372), .A(n21644), 
        .ZN(n20404) );
  NOR2_X1 U23455 ( .A1(n20399), .A2(n20404), .ZN(n20401) );
  AOI21_X1 U23456 ( .B1(n20401), .B2(n20400), .A(n20405), .ZN(n20402) );
  OAI211_X1 U23457 ( .C1(n21372), .C2(n20403), .A(n20402), .B(n20513), .ZN(
        P2_U3210) );
  AOI21_X1 U23458 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20405), .A(n20404), 
        .ZN(n20410) );
  INV_X1 U23459 ( .A(n20405), .ZN(n20406) );
  OAI22_X1 U23460 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20407), .B1(NA), 
        .B2(n20406), .ZN(n20408) );
  OAI211_X1 U23461 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20408), .ZN(n20409) );
  OAI21_X1 U23462 ( .B1(n20411), .B2(n20410), .A(n20409), .ZN(P2_U3211) );
  NAND2_X2 U23463 ( .A1(n20462), .A2(n21644), .ZN(n20464) );
  OAI222_X1 U23464 ( .A1(n20464), .A2(n20414), .B1(n20413), .B2(n20462), .C1(
        n20412), .C2(n20458), .ZN(P2_U3212) );
  CLKBUF_X1 U23465 ( .A(n20458), .Z(n20461) );
  OAI222_X1 U23466 ( .A1(n20464), .A2(n10772), .B1(n20415), .B2(n20462), .C1(
        n20414), .C2(n20461), .ZN(P2_U3213) );
  OAI222_X1 U23467 ( .A1(n20464), .A2(n20417), .B1(n20416), .B2(n20462), .C1(
        n10772), .C2(n20461), .ZN(P2_U3214) );
  OAI222_X1 U23468 ( .A1(n20464), .A2(n16206), .B1(n20418), .B2(n20462), .C1(
        n20417), .C2(n20461), .ZN(P2_U3215) );
  OAI222_X1 U23469 ( .A1(n20464), .A2(n20420), .B1(n20419), .B2(n20462), .C1(
        n16206), .C2(n20461), .ZN(P2_U3216) );
  OAI222_X1 U23470 ( .A1(n20464), .A2(n21760), .B1(n20421), .B2(n20462), .C1(
        n20420), .C2(n20461), .ZN(P2_U3217) );
  OAI222_X1 U23471 ( .A1(n20464), .A2(n16671), .B1(n20422), .B2(n20462), .C1(
        n21760), .C2(n20461), .ZN(P2_U3218) );
  OAI222_X1 U23472 ( .A1(n20464), .A2(n20424), .B1(n20423), .B2(n20462), .C1(
        n16671), .C2(n20461), .ZN(P2_U3219) );
  OAI222_X1 U23473 ( .A1(n20464), .A2(n20426), .B1(n20425), .B2(n20462), .C1(
        n20424), .C2(n20461), .ZN(P2_U3220) );
  OAI222_X1 U23474 ( .A1(n20464), .A2(n20428), .B1(n20427), .B2(n20462), .C1(
        n20426), .C2(n20461), .ZN(P2_U3221) );
  OAI222_X1 U23475 ( .A1(n20464), .A2(n20430), .B1(n20429), .B2(n20462), .C1(
        n20428), .C2(n20461), .ZN(P2_U3222) );
  OAI222_X1 U23476 ( .A1(n20464), .A2(n21718), .B1(n20431), .B2(n20462), .C1(
        n20430), .C2(n20461), .ZN(P2_U3223) );
  OAI222_X1 U23477 ( .A1(n20464), .A2(n20433), .B1(n20432), .B2(n20462), .C1(
        n21718), .C2(n20461), .ZN(P2_U3224) );
  OAI222_X1 U23478 ( .A1(n20464), .A2(n20435), .B1(n20434), .B2(n20462), .C1(
        n20433), .C2(n20461), .ZN(P2_U3225) );
  OAI222_X1 U23479 ( .A1(n20464), .A2(n20437), .B1(n20436), .B2(n20462), .C1(
        n20435), .C2(n20461), .ZN(P2_U3226) );
  OAI222_X1 U23480 ( .A1(n20464), .A2(n20439), .B1(n20438), .B2(n20462), .C1(
        n20437), .C2(n20461), .ZN(P2_U3227) );
  OAI222_X1 U23481 ( .A1(n20464), .A2(n13325), .B1(n20440), .B2(n20462), .C1(
        n20439), .C2(n20461), .ZN(P2_U3228) );
  OAI222_X1 U23482 ( .A1(n20464), .A2(n20442), .B1(n20441), .B2(n20462), .C1(
        n13325), .C2(n20461), .ZN(P2_U3229) );
  OAI222_X1 U23483 ( .A1(n20464), .A2(n19665), .B1(n21600), .B2(n20462), .C1(
        n20442), .C2(n20461), .ZN(P2_U3230) );
  OAI222_X1 U23484 ( .A1(n20464), .A2(n20444), .B1(n20443), .B2(n20462), .C1(
        n19665), .C2(n20461), .ZN(P2_U3231) );
  OAI222_X1 U23485 ( .A1(n20464), .A2(n20446), .B1(n20445), .B2(n20462), .C1(
        n20444), .C2(n20461), .ZN(P2_U3232) );
  OAI222_X1 U23486 ( .A1(n20464), .A2(n20448), .B1(n20447), .B2(n20462), .C1(
        n20446), .C2(n20461), .ZN(P2_U3233) );
  OAI222_X1 U23487 ( .A1(n20464), .A2(n15985), .B1(n20449), .B2(n20462), .C1(
        n20448), .C2(n20461), .ZN(P2_U3234) );
  OAI222_X1 U23488 ( .A1(n20464), .A2(n20451), .B1(n20450), .B2(n20462), .C1(
        n15985), .C2(n20458), .ZN(P2_U3235) );
  OAI222_X1 U23489 ( .A1(n20464), .A2(n20452), .B1(n21738), .B2(n20462), .C1(
        n20451), .C2(n20458), .ZN(P2_U3236) );
  OAI222_X1 U23490 ( .A1(n20464), .A2(n20455), .B1(n20453), .B2(n20462), .C1(
        n20452), .C2(n20458), .ZN(P2_U3237) );
  OAI222_X1 U23491 ( .A1(n20461), .A2(n20455), .B1(n20454), .B2(n20462), .C1(
        n20456), .C2(n20464), .ZN(P2_U3238) );
  OAI222_X1 U23492 ( .A1(n20464), .A2(n20459), .B1(n20457), .B2(n20462), .C1(
        n20456), .C2(n20458), .ZN(P2_U3239) );
  OAI222_X1 U23493 ( .A1(n20464), .A2(n11480), .B1(n20460), .B2(n20462), .C1(
        n20459), .C2(n20458), .ZN(P2_U3240) );
  OAI222_X1 U23494 ( .A1(n20464), .A2(n21704), .B1(n20463), .B2(n20462), .C1(
        n11480), .C2(n20461), .ZN(P2_U3241) );
  INV_X1 U23495 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20465) );
  AOI22_X1 U23496 ( .A1(n20462), .A2(n20466), .B1(n20465), .B2(n20526), .ZN(
        P2_U3585) );
  INV_X1 U23497 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20467) );
  AOI22_X1 U23498 ( .A1(n20462), .A2(n20467), .B1(n21773), .B2(n20526), .ZN(
        P2_U3586) );
  INV_X1 U23499 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20468) );
  AOI22_X1 U23500 ( .A1(n20462), .A2(n20469), .B1(n20468), .B2(n20526), .ZN(
        P2_U3587) );
  INV_X1 U23501 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20470) );
  AOI22_X1 U23502 ( .A1(n20462), .A2(n20471), .B1(n20470), .B2(n20526), .ZN(
        P2_U3588) );
  OAI21_X1 U23503 ( .B1(n20475), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20473), 
        .ZN(n20472) );
  INV_X1 U23504 ( .A(n20472), .ZN(P2_U3591) );
  OAI21_X1 U23505 ( .B1(n20475), .B2(n20474), .A(n20473), .ZN(P2_U3592) );
  NAND2_X1 U23506 ( .A1(n20477), .A2(n20476), .ZN(n20494) );
  OR2_X1 U23507 ( .A1(n20479), .A2(n20478), .ZN(n20481) );
  AND2_X1 U23508 ( .A1(n20481), .A2(n20480), .ZN(n20489) );
  NAND2_X1 U23509 ( .A1(n20494), .A2(n20489), .ZN(n20487) );
  INV_X1 U23510 ( .A(n20482), .ZN(n20483) );
  AOI222_X1 U23511 ( .A1(n20487), .A2(n20486), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20485), .C1(n20484), .C2(n20483), .ZN(n20488) );
  AOI22_X1 U23512 ( .A1(n20498), .A2(n21570), .B1(n20488), .B2(n20495), .ZN(
        P2_U3602) );
  INV_X1 U23513 ( .A(n20489), .ZN(n20492) );
  AOI22_X1 U23514 ( .A1(n20492), .A2(n20491), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20490), .ZN(n20493) );
  AND2_X1 U23515 ( .A1(n20494), .A2(n20493), .ZN(n20496) );
  AOI22_X1 U23516 ( .A1(n20498), .A2(n20497), .B1(n20496), .B2(n20495), .ZN(
        P2_U3603) );
  AOI22_X1 U23517 ( .A1(n20462), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20499), 
        .B2(n20526), .ZN(P2_U3608) );
  INV_X1 U23518 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n21647) );
  AOI22_X1 U23519 ( .A1(n20503), .A2(n20502), .B1(n20501), .B2(n20500), .ZN(
        n20506) );
  NOR2_X1 U23520 ( .A1(n20507), .A2(n20504), .ZN(n20505) );
  AOI22_X1 U23521 ( .A1(n21647), .A2(n20507), .B1(n20506), .B2(n20505), .ZN(
        P2_U3609) );
  NOR2_X1 U23522 ( .A1(n20509), .A2(n20508), .ZN(n20518) );
  NAND3_X1 U23523 ( .A1(n20513), .A2(n20510), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20515) );
  OAI21_X1 U23524 ( .B1(n20513), .B2(n20512), .A(n20511), .ZN(n20514) );
  MUX2_X1 U23525 ( .A(n20515), .B(n20514), .S(n11051), .Z(n20516) );
  OAI21_X1 U23526 ( .B1(n20518), .B2(n20517), .A(n20516), .ZN(n20525) );
  INV_X1 U23527 ( .A(n20519), .ZN(n20523) );
  AND2_X1 U23528 ( .A1(n20520), .A2(n19744), .ZN(n20522) );
  AOI211_X1 U23529 ( .C1(n12673), .C2(n20523), .A(n20522), .B(n20521), .ZN(
        n20524) );
  MUX2_X1 U23530 ( .A(n20525), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n20524), 
        .Z(P2_U3610) );
  INV_X1 U23531 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20527) );
  AOI22_X1 U23532 ( .A1(n20462), .A2(n20528), .B1(n20527), .B2(n20526), .ZN(
        P2_U3611) );
  OAI21_X1 U23533 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20529), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n21379) );
  NAND2_X1 U23534 ( .A1(n21379), .A2(n21494), .ZN(n21448) );
  OAI21_X1 U23535 ( .B1(n21439), .B2(n21567), .A(n21448), .ZN(P1_U2802) );
  INV_X1 U23536 ( .A(n20530), .ZN(n20534) );
  OAI21_X1 U23537 ( .B1(n20532), .B2(n20531), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20533) );
  OAI21_X1 U23538 ( .B1(n20534), .B2(n21369), .A(n20533), .ZN(P1_U2803) );
  NOR2_X1 U23539 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20536) );
  OAI21_X1 U23540 ( .B1(n20536), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21494), .ZN(
        n20535) );
  OAI21_X1 U23541 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21494), .A(n20535), 
        .ZN(P1_U2804) );
  OAI21_X1 U23542 ( .B1(BS16), .B2(n20536), .A(n21452), .ZN(n21450) );
  OAI21_X1 U23543 ( .B1(n21452), .B2(n20830), .A(n21450), .ZN(P1_U2805) );
  OAI21_X1 U23544 ( .B1(n20539), .B2(n20538), .A(n20537), .ZN(P1_U2806) );
  NOR4_X1 U23545 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20543) );
  NOR4_X1 U23546 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20542) );
  NOR4_X1 U23547 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20541) );
  NOR4_X1 U23548 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20540) );
  NAND4_X1 U23549 ( .A1(n20543), .A2(n20542), .A3(n20541), .A4(n20540), .ZN(
        n20549) );
  NOR4_X1 U23550 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20547) );
  AOI211_X1 U23551 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_11__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20546) );
  NOR4_X1 U23552 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20545) );
  NOR4_X1 U23553 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20544) );
  NAND4_X1 U23554 ( .A1(n20547), .A2(n20546), .A3(n20545), .A4(n20544), .ZN(
        n20548) );
  NOR2_X1 U23555 ( .A1(n20549), .A2(n20548), .ZN(n21483) );
  INV_X1 U23556 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21446) );
  NOR3_X1 U23557 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20551) );
  OAI21_X1 U23558 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20551), .A(n21483), .ZN(
        n20550) );
  OAI21_X1 U23559 ( .B1(n21483), .B2(n21446), .A(n20550), .ZN(P1_U2807) );
  INV_X1 U23560 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21476) );
  INV_X1 U23561 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21451) );
  AOI21_X1 U23562 ( .B1(n21476), .B2(n21451), .A(n20551), .ZN(n20552) );
  INV_X1 U23563 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21444) );
  INV_X1 U23564 ( .A(n21483), .ZN(n21478) );
  AOI22_X1 U23565 ( .A1(n21483), .A2(n20552), .B1(n21444), .B2(n21478), .ZN(
        P1_U2808) );
  AOI22_X1 U23566 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20622), .B1(n20608), .B2(
        n20639), .ZN(n20556) );
  NOR2_X1 U23567 ( .A1(n20553), .A2(n21402), .ZN(n20554) );
  AOI211_X1 U23568 ( .C1(n20625), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20718), .B(n20554), .ZN(n20555) );
  OAI211_X1 U23569 ( .C1(n20557), .C2(n20620), .A(n20556), .B(n20555), .ZN(
        n20558) );
  AOI21_X1 U23570 ( .B1(n20640), .B2(n20582), .A(n20558), .ZN(n20559) );
  OAI21_X1 U23571 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20560), .A(n20559), .ZN(
        P1_U2831) );
  OAI21_X1 U23572 ( .B1(n20595), .B2(n20596), .A(n20561), .ZN(n20594) );
  AOI21_X1 U23573 ( .B1(n20612), .B2(n20562), .A(n20594), .ZN(n20585) );
  NAND2_X1 U23574 ( .A1(n20563), .A2(n20586), .ZN(n20564) );
  NOR2_X1 U23575 ( .A1(n20564), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n20569) );
  INV_X1 U23576 ( .A(n20565), .ZN(n20566) );
  NAND2_X1 U23577 ( .A1(n20623), .A2(n20566), .ZN(n20567) );
  OAI211_X1 U23578 ( .C1(n12329), .C2(n20588), .A(n20567), .B(n20576), .ZN(
        n20568) );
  NOR2_X1 U23579 ( .A1(n20569), .A2(n20568), .ZN(n20571) );
  AOI22_X1 U23580 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20622), .B1(n20608), .B2(
        n20643), .ZN(n20570) );
  NAND2_X1 U23581 ( .A1(n20571), .A2(n20570), .ZN(n20572) );
  AOI21_X1 U23582 ( .B1(n20644), .B2(n20582), .A(n20572), .ZN(n20573) );
  OAI21_X1 U23583 ( .B1(n20585), .B2(n21398), .A(n20573), .ZN(P1_U2833) );
  INV_X1 U23584 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21680) );
  AOI22_X1 U23585 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20625), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(n20622), .ZN(n20575) );
  NAND3_X1 U23586 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20586), .A3(n21680), 
        .ZN(n20574) );
  NAND3_X1 U23587 ( .A1(n20576), .A2(n20575), .A3(n20574), .ZN(n20577) );
  AOI21_X1 U23588 ( .B1(n20608), .B2(n20578), .A(n20577), .ZN(n20579) );
  OAI21_X1 U23589 ( .B1(n20620), .B2(n20580), .A(n20579), .ZN(n20581) );
  AOI21_X1 U23590 ( .B1(n20583), .B2(n20582), .A(n20581), .ZN(n20584) );
  OAI21_X1 U23591 ( .B1(n20585), .B2(n21680), .A(n20584), .ZN(P1_U2834) );
  INV_X1 U23592 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21396) );
  AOI22_X1 U23593 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20622), .B1(n20586), .B2(
        n21396), .ZN(n20593) );
  OAI22_X1 U23594 ( .A1(n20589), .A2(n20588), .B1(n20587), .B2(n20620), .ZN(
        n20590) );
  AOI211_X1 U23595 ( .C1(n20608), .C2(n20647), .A(n20718), .B(n20590), .ZN(
        n20592) );
  AOI22_X1 U23596 ( .A1(n20650), .A2(n20633), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20594), .ZN(n20591) );
  NAND3_X1 U23597 ( .A1(n20593), .A2(n20592), .A3(n20591), .ZN(P1_U2835) );
  INV_X1 U23598 ( .A(n20594), .ZN(n20606) );
  AOI22_X1 U23599 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(n20622), .B1(n20608), .B2(
        n20719), .ZN(n20603) );
  NOR3_X1 U23600 ( .A1(n20597), .A2(n20596), .A3(n20595), .ZN(n20598) );
  AOI21_X1 U23601 ( .B1(n20599), .B2(n20626), .A(n20598), .ZN(n20600) );
  INV_X1 U23602 ( .A(n20600), .ZN(n20601) );
  AOI211_X1 U23603 ( .C1(n20625), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20718), .B(n20601), .ZN(n20602) );
  OAI211_X1 U23604 ( .C1(n20620), .C2(n20713), .A(n20603), .B(n20602), .ZN(
        n20604) );
  AOI21_X1 U23605 ( .B1(n20708), .B2(n20633), .A(n20604), .ZN(n20605) );
  OAI21_X1 U23606 ( .B1(n20606), .B2(n21393), .A(n20605), .ZN(P1_U2836) );
  INV_X1 U23607 ( .A(n20607), .ZN(n20621) );
  AOI22_X1 U23608 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(n20622), .B1(n20608), .B2(
        n20728), .ZN(n20619) );
  INV_X1 U23609 ( .A(n20609), .ZN(n20617) );
  NOR2_X1 U23610 ( .A1(n20611), .A2(n20610), .ZN(n20631) );
  INV_X1 U23611 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21392) );
  AOI22_X1 U23612 ( .A1(n20626), .A2(n21464), .B1(n20625), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20615) );
  AND2_X1 U23613 ( .A1(n20612), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20628) );
  OR2_X1 U23614 ( .A1(n21392), .A2(n20627), .ZN(n20613) );
  OAI211_X1 U23615 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20628), .B(n20613), .ZN(n20614) );
  OAI211_X1 U23616 ( .C1(n20631), .C2(n21392), .A(n20615), .B(n20614), .ZN(
        n20616) );
  AOI21_X1 U23617 ( .B1(n20617), .B2(n20633), .A(n20616), .ZN(n20618) );
  OAI211_X1 U23618 ( .C1(n20621), .C2(n20620), .A(n20619), .B(n20618), .ZN(
        P1_U2837) );
  AOI22_X1 U23619 ( .A1(n20624), .A2(n20623), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n20622), .ZN(n20636) );
  INV_X1 U23620 ( .A(n13843), .ZN(n20780) );
  AOI22_X1 U23621 ( .A1(n20626), .A2(n20780), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20625), .ZN(n20630) );
  NAND2_X1 U23622 ( .A1(n20628), .A2(n20627), .ZN(n20629) );
  OAI211_X1 U23623 ( .C1(n20631), .C2(n20627), .A(n20630), .B(n20629), .ZN(
        n20632) );
  AOI21_X1 U23624 ( .B1(n20634), .B2(n20633), .A(n20632), .ZN(n20635) );
  OAI211_X1 U23625 ( .C1(n20638), .C2(n20637), .A(n20636), .B(n20635), .ZN(
        P1_U2838) );
  AOI22_X1 U23626 ( .A1(n20640), .A2(n20649), .B1(n20648), .B2(n20639), .ZN(
        n20641) );
  OAI21_X1 U23627 ( .B1(n20653), .B2(n20642), .A(n20641), .ZN(P1_U2863) );
  AOI22_X1 U23628 ( .A1(n20644), .A2(n20649), .B1(n20648), .B2(n20643), .ZN(
        n20645) );
  OAI21_X1 U23629 ( .B1(n20653), .B2(n20646), .A(n20645), .ZN(P1_U2865) );
  AOI22_X1 U23630 ( .A1(n20650), .A2(n20649), .B1(n20648), .B2(n20647), .ZN(
        n20651) );
  OAI21_X1 U23631 ( .B1(n20653), .B2(n20652), .A(n20651), .ZN(P1_U2867) );
  INV_X1 U23632 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n21694) );
  AOI22_X1 U23633 ( .A1(n20658), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20662), .ZN(n20655) );
  OAI21_X1 U23634 ( .B1(n21694), .B2(n20675), .A(n20655), .ZN(P1_U2907) );
  AOI22_X1 U23635 ( .A1(n20658), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20662), .ZN(n20656) );
  OAI21_X1 U23636 ( .B1(n21594), .B2(n20675), .A(n20656), .ZN(P1_U2911) );
  AOI22_X1 U23637 ( .A1(n20658), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20662), .ZN(n20657) );
  OAI21_X1 U23638 ( .B1(n21744), .B2(n20675), .A(n20657), .ZN(P1_U2918) );
  INV_X1 U23639 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n21665) );
  AOI22_X1 U23640 ( .A1(n20681), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n20658), .ZN(n20659) );
  OAI21_X1 U23641 ( .B1(n21665), .B2(n20674), .A(n20659), .ZN(P1_U2920) );
  AOI22_X1 U23642 ( .A1(n20662), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20660) );
  OAI21_X1 U23643 ( .B1(n20661), .B2(n20683), .A(n20660), .ZN(P1_U2921) );
  AOI22_X1 U23644 ( .A1(n20662), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20663) );
  OAI21_X1 U23645 ( .B1(n15468), .B2(n20683), .A(n20663), .ZN(P1_U2922) );
  AOI22_X1 U23646 ( .A1(n20662), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20664) );
  OAI21_X1 U23647 ( .B1(n15471), .B2(n20683), .A(n20664), .ZN(P1_U2923) );
  AOI22_X1 U23648 ( .A1(n20662), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20665) );
  OAI21_X1 U23649 ( .B1(n15472), .B2(n20683), .A(n20665), .ZN(P1_U2924) );
  AOI22_X1 U23650 ( .A1(n20662), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20666) );
  OAI21_X1 U23651 ( .B1(n15475), .B2(n20683), .A(n20666), .ZN(P1_U2925) );
  INV_X1 U23652 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n20667) );
  OAI222_X1 U23653 ( .A1(n20675), .A2(n21586), .B1(n20683), .B2(n14248), .C1(
        n20674), .C2(n20667), .ZN(P1_U2926) );
  AOI22_X1 U23654 ( .A1(n20662), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20668) );
  OAI21_X1 U23655 ( .B1(n15483), .B2(n20683), .A(n20668), .ZN(P1_U2927) );
  AOI22_X1 U23656 ( .A1(n20662), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20669) );
  OAI21_X1 U23657 ( .B1(n20670), .B2(n20683), .A(n20669), .ZN(P1_U2928) );
  AOI22_X1 U23658 ( .A1(n20662), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20671) );
  OAI21_X1 U23659 ( .B1(n14260), .B2(n20683), .A(n20671), .ZN(P1_U2929) );
  AOI22_X1 U23660 ( .A1(n20662), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20672) );
  OAI21_X1 U23661 ( .B1(n15488), .B2(n20683), .A(n20672), .ZN(P1_U2930) );
  INV_X1 U23662 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n20673) );
  OAI222_X1 U23663 ( .A1(n20675), .A2(n21754), .B1(n20683), .B2(n14256), .C1(
        n20674), .C2(n20673), .ZN(P1_U2931) );
  AOI22_X1 U23664 ( .A1(n20662), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20676) );
  OAI21_X1 U23665 ( .B1(n14252), .B2(n20683), .A(n20676), .ZN(P1_U2932) );
  AOI22_X1 U23666 ( .A1(n20662), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20677) );
  OAI21_X1 U23667 ( .B1(n14277), .B2(n20683), .A(n20677), .ZN(P1_U2933) );
  AOI22_X1 U23668 ( .A1(n20662), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20678) );
  OAI21_X1 U23669 ( .B1(n20679), .B2(n20683), .A(n20678), .ZN(P1_U2934) );
  AOI22_X1 U23670 ( .A1(n20662), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20680) );
  OAI21_X1 U23671 ( .B1(n14280), .B2(n20683), .A(n20680), .ZN(P1_U2935) );
  AOI22_X1 U23672 ( .A1(n20662), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20681), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20682) );
  OAI21_X1 U23673 ( .B1(n20684), .B2(n20683), .A(n20682), .ZN(P1_U2936) );
  AOI22_X1 U23674 ( .A1(n20700), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n21497), .ZN(n20687) );
  INV_X1 U23675 ( .A(n20685), .ZN(n20686) );
  NAND2_X1 U23676 ( .A1(n20690), .A2(n20686), .ZN(n20692) );
  NAND2_X1 U23677 ( .A1(n20687), .A2(n20692), .ZN(P1_U2946) );
  AOI22_X1 U23678 ( .A1(n20700), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n21497), .ZN(n20691) );
  INV_X1 U23679 ( .A(n20688), .ZN(n20689) );
  NAND2_X1 U23680 ( .A1(n20690), .A2(n20689), .ZN(n20698) );
  NAND2_X1 U23681 ( .A1(n20691), .A2(n20698), .ZN(P1_U2950) );
  AOI22_X1 U23682 ( .A1(n20700), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21497), .ZN(n20693) );
  NAND2_X1 U23683 ( .A1(n20693), .A2(n20692), .ZN(P1_U2961) );
  AOI22_X1 U23684 ( .A1(n20700), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n21497), .ZN(n20695) );
  NAND2_X1 U23685 ( .A1(n20695), .A2(n20694), .ZN(P1_U2963) );
  AOI22_X1 U23686 ( .A1(n20700), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21497), .ZN(n20697) );
  NAND2_X1 U23687 ( .A1(n20697), .A2(n20696), .ZN(P1_U2964) );
  AOI22_X1 U23688 ( .A1(n20700), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n21497), .ZN(n20699) );
  NAND2_X1 U23689 ( .A1(n20699), .A2(n20698), .ZN(P1_U2965) );
  AOI22_X1 U23690 ( .A1(n20700), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21497), .ZN(n20702) );
  NAND2_X1 U23691 ( .A1(n20702), .A2(n20701), .ZN(P1_U2966) );
  AOI22_X1 U23692 ( .A1(n20703), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20718), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20712) );
  AOI21_X1 U23693 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14573), .A(
        n20704), .ZN(n20707) );
  XNOR2_X1 U23694 ( .A(n20705), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20706) );
  XNOR2_X1 U23695 ( .A(n20707), .B(n20706), .ZN(n20722) );
  AOI22_X1 U23696 ( .A1(n20722), .A2(n20710), .B1(n20709), .B2(n20708), .ZN(
        n20711) );
  OAI211_X1 U23697 ( .C1(n20714), .C2(n20713), .A(n20712), .B(n20711), .ZN(
        P1_U2995) );
  AOI21_X1 U23698 ( .B1(n20716), .B2(n12123), .A(n20715), .ZN(n20717) );
  INV_X1 U23699 ( .A(n20717), .ZN(n20725) );
  AOI22_X1 U23700 ( .A1(n20742), .A2(n20719), .B1(n20718), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20724) );
  NAND2_X1 U23701 ( .A1(n20736), .A2(n20720), .ZN(n20745) );
  NAND3_X1 U23702 ( .A1(n20750), .A2(n20721), .A3(n20745), .ZN(n20729) );
  AOI22_X1 U23703 ( .A1(n20722), .A2(n20738), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20729), .ZN(n20723) );
  OAI211_X1 U23704 ( .C1(n20733), .C2(n20725), .A(n20724), .B(n20723), .ZN(
        P1_U3027) );
  INV_X1 U23705 ( .A(n20726), .ZN(n20727) );
  AOI21_X1 U23706 ( .B1(n20742), .B2(n20728), .A(n20727), .ZN(n20732) );
  AOI22_X1 U23707 ( .A1(n20730), .A2(n20738), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20729), .ZN(n20731) );
  OAI211_X1 U23708 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20733), .A(
        n20732), .B(n20731), .ZN(P1_U3028) );
  NOR2_X1 U23709 ( .A1(n20734), .A2(n20767), .ZN(n20737) );
  AOI22_X1 U23710 ( .A1(n20737), .A2(n20736), .B1(n20767), .B2(n20735), .ZN(
        n20749) );
  NAND3_X1 U23711 ( .A1(n20739), .A2(n14631), .A3(n20738), .ZN(n20747) );
  AOI21_X1 U23712 ( .B1(n20742), .B2(n20741), .A(n20740), .ZN(n20746) );
  OR3_X1 U23713 ( .A1(n20743), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n20767), .ZN(n20744) );
  AND4_X1 U23714 ( .A1(n20747), .A2(n20746), .A3(n20745), .A4(n20744), .ZN(
        n20748) );
  OAI221_X1 U23715 ( .B1(n20751), .B2(n20750), .C1(n20751), .C2(n20749), .A(
        n20748), .ZN(P1_U3029) );
  NOR3_X1 U23716 ( .A1(n20755), .A2(n20754), .A3(n20753), .ZN(n20764) );
  AND3_X1 U23717 ( .A1(n20757), .A2(n20767), .A3(n20756), .ZN(n20762) );
  INV_X1 U23718 ( .A(n20758), .ZN(n20759) );
  NOR2_X1 U23719 ( .A1(n20760), .A2(n20759), .ZN(n20761) );
  NOR4_X1 U23720 ( .A1(n20764), .A2(n20763), .A3(n20762), .A4(n20761), .ZN(
        n20765) );
  OAI221_X1 U23721 ( .B1(n20767), .B2(n20766), .C1(n20767), .C2(n15895), .A(
        n20765), .ZN(P1_U3030) );
  NOR2_X1 U23722 ( .A1(n20768), .A2(n21475), .ZN(P1_U3032) );
  AOI22_X2 U23723 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20816), .B1(DATAI_16_), 
        .B2(n20817), .ZN(n21266) );
  INV_X1 U23724 ( .A(n21065), .ZN(n20772) );
  AOI22_X1 U23725 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20816), .B1(DATAI_24_), 
        .B2(n20817), .ZN(n21320) );
  INV_X1 U23726 ( .A(n21320), .ZN(n21263) );
  NAND2_X1 U23727 ( .A1(n21474), .A2(n21066), .ZN(n20892) );
  OR2_X1 U23728 ( .A1(n21198), .A2(n20892), .ZN(n20781) );
  INV_X1 U23729 ( .A(n20781), .ZN(n20820) );
  NAND2_X1 U23730 ( .A1(n20819), .A2(n20776), .ZN(n21116) );
  AOI22_X1 U23731 ( .A1(n21362), .A2(n21263), .B1(n20820), .B2(n21310), .ZN(
        n20791) );
  INV_X1 U23732 ( .A(n21120), .ZN(n20777) );
  NOR2_X1 U23733 ( .A1(n20777), .A2(n21067), .ZN(n20787) );
  OR2_X1 U23734 ( .A1(n20785), .A2(n21306), .ZN(n21254) );
  INV_X1 U23735 ( .A(n21254), .ZN(n20778) );
  NAND2_X1 U23736 ( .A1(n20854), .A2(n9694), .ZN(n20779) );
  NAND2_X1 U23737 ( .A1(n9694), .A2(n20830), .ZN(n21199) );
  OAI21_X1 U23738 ( .B1(n20779), .B2(n21362), .A(n21199), .ZN(n20784) );
  OR2_X1 U23739 ( .A1(n21464), .A2(n20780), .ZN(n20895) );
  AOI22_X1 U23740 ( .A1(n20784), .A2(n20788), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20781), .ZN(n20782) );
  NOR2_X2 U23741 ( .A1(n20945), .A2(n20783), .ZN(n21309) );
  INV_X1 U23742 ( .A(n20784), .ZN(n20789) );
  INV_X1 U23743 ( .A(n20785), .ZN(n20786) );
  NOR2_X1 U23744 ( .A1(n20786), .A2(n21306), .ZN(n20946) );
  INV_X1 U23745 ( .A(n20946), .ZN(n21126) );
  INV_X1 U23746 ( .A(n20787), .ZN(n20940) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20823), .B1(
        n21309), .B2(n20822), .ZN(n20790) );
  OAI211_X1 U23748 ( .C1(n21266), .C2(n20854), .A(n20791), .B(n20790), .ZN(
        P1_U3033) );
  AOI22_X1 U23749 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20816), .B1(DATAI_17_), 
        .B2(n20817), .ZN(n21270) );
  INV_X1 U23750 ( .A(n21326), .ZN(n21267) );
  NAND2_X1 U23751 ( .A1(n20819), .A2(n20792), .ZN(n21131) );
  AOI22_X1 U23752 ( .A1(n21362), .A2(n21267), .B1(n20820), .B2(n21322), .ZN(
        n20795) );
  NOR2_X2 U23753 ( .A1(n20945), .A2(n20793), .ZN(n21321) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20823), .B1(
        n21321), .B2(n20822), .ZN(n20794) );
  OAI211_X1 U23755 ( .C1(n21270), .C2(n20854), .A(n20795), .B(n20794), .ZN(
        P1_U3034) );
  AOI22_X1 U23756 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20816), .B1(DATAI_26_), 
        .B2(n20817), .ZN(n21332) );
  INV_X1 U23757 ( .A(n21332), .ZN(n21271) );
  NAND2_X1 U23758 ( .A1(n20819), .A2(n20796), .ZN(n21135) );
  AOI22_X1 U23759 ( .A1(n21362), .A2(n21271), .B1(n20820), .B2(n21328), .ZN(
        n20799) );
  NOR2_X2 U23760 ( .A1(n20945), .A2(n20797), .ZN(n21327) );
  AOI22_X1 U23761 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20823), .B1(
        n21327), .B2(n20822), .ZN(n20798) );
  OAI211_X1 U23762 ( .C1(n21274), .C2(n20854), .A(n20799), .B(n20798), .ZN(
        P1_U3035) );
  AOI22_X1 U23763 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20816), .B1(DATAI_27_), 
        .B2(n20817), .ZN(n21338) );
  INV_X1 U23764 ( .A(n21338), .ZN(n21275) );
  NAND2_X1 U23765 ( .A1(n20819), .A2(n20800), .ZN(n21139) );
  AOI22_X1 U23766 ( .A1(n21362), .A2(n21275), .B1(n20820), .B2(n21334), .ZN(
        n20803) );
  NOR2_X2 U23767 ( .A1(n20945), .A2(n20801), .ZN(n21333) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20823), .B1(
        n21333), .B2(n20822), .ZN(n20802) );
  OAI211_X1 U23769 ( .C1(n21278), .C2(n20854), .A(n20803), .B(n20802), .ZN(
        P1_U3036) );
  AOI22_X1 U23770 ( .A1(DATAI_20_), .A2(n20817), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20816), .ZN(n21282) );
  AOI22_X1 U23771 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20816), .B1(DATAI_28_), 
        .B2(n20817), .ZN(n21344) );
  INV_X1 U23772 ( .A(n21344), .ZN(n21279) );
  NAND2_X1 U23773 ( .A1(n20819), .A2(n20804), .ZN(n21143) );
  AOI22_X1 U23774 ( .A1(n21362), .A2(n21279), .B1(n20820), .B2(n21340), .ZN(
        n20807) );
  NOR2_X2 U23775 ( .A1(n20945), .A2(n20805), .ZN(n21339) );
  AOI22_X1 U23776 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20823), .B1(
        n21339), .B2(n20822), .ZN(n20806) );
  OAI211_X1 U23777 ( .C1(n21282), .C2(n20854), .A(n20807), .B(n20806), .ZN(
        P1_U3037) );
  AOI22_X1 U23778 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20816), .B1(DATAI_21_), 
        .B2(n20817), .ZN(n21286) );
  INV_X1 U23779 ( .A(n21350), .ZN(n21283) );
  NAND2_X1 U23780 ( .A1(n20819), .A2(n20808), .ZN(n21147) );
  AOI22_X1 U23781 ( .A1(n21362), .A2(n21283), .B1(n20820), .B2(n21346), .ZN(
        n20811) );
  NOR2_X2 U23782 ( .A1(n20945), .A2(n20809), .ZN(n21345) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20823), .B1(
        n21345), .B2(n20822), .ZN(n20810) );
  OAI211_X1 U23784 ( .C1(n21286), .C2(n20854), .A(n20811), .B(n20810), .ZN(
        P1_U3038) );
  AOI22_X1 U23785 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20816), .B1(DATAI_22_), 
        .B2(n20817), .ZN(n21290) );
  AOI22_X1 U23786 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20816), .B1(DATAI_30_), 
        .B2(n20817), .ZN(n21356) );
  INV_X1 U23787 ( .A(n21356), .ZN(n21287) );
  NAND2_X1 U23788 ( .A1(n20819), .A2(n20812), .ZN(n21151) );
  AOI22_X1 U23789 ( .A1(n21362), .A2(n21287), .B1(n20820), .B2(n21352), .ZN(
        n20815) );
  NOR2_X2 U23790 ( .A1(n20945), .A2(n20813), .ZN(n21351) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20823), .B1(
        n21351), .B2(n20822), .ZN(n20814) );
  OAI211_X1 U23792 ( .C1(n21290), .C2(n20854), .A(n20815), .B(n20814), .ZN(
        P1_U3039) );
  AOI22_X1 U23793 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20816), .B1(DATAI_23_), 
        .B2(n20817), .ZN(n21298) );
  AOI22_X1 U23794 ( .A1(DATAI_31_), .A2(n20817), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20816), .ZN(n21367) );
  INV_X1 U23795 ( .A(n21367), .ZN(n21293) );
  NAND2_X1 U23796 ( .A1(n20819), .A2(n20818), .ZN(n21156) );
  AOI22_X1 U23797 ( .A1(n21362), .A2(n21293), .B1(n20820), .B2(n21360), .ZN(
        n20825) );
  NOR2_X2 U23798 ( .A1(n20945), .A2(n20821), .ZN(n21358) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20823), .B1(
        n21358), .B2(n20822), .ZN(n20824) );
  OAI211_X1 U23800 ( .C1(n21298), .C2(n20854), .A(n20825), .B(n20824), .ZN(
        P1_U3040) );
  INV_X1 U23801 ( .A(n20895), .ZN(n20827) );
  INV_X1 U23802 ( .A(n20826), .ZN(n21091) );
  NOR3_X2 U23803 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21677), .A3(
        n20892), .ZN(n20848) );
  AOI21_X1 U23804 ( .B1(n20827), .B2(n21091), .A(n20848), .ZN(n20829) );
  NOR2_X1 U23805 ( .A1(n20892), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20832) );
  INV_X1 U23806 ( .A(n20832), .ZN(n20828) );
  OAI22_X1 U23807 ( .A1(n20829), .A2(n21304), .B1(n20828), .B2(n21306), .ZN(
        n20849) );
  AOI22_X1 U23808 ( .A1(n20849), .A2(n21309), .B1(n21310), .B2(n20848), .ZN(
        n20834) );
  INV_X1 U23809 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20830) );
  OAI211_X1 U23810 ( .C1(n20897), .C2(n20830), .A(n9694), .B(n20829), .ZN(
        n20831) );
  OAI211_X1 U23811 ( .C1(n9694), .C2(n20832), .A(n21314), .B(n20831), .ZN(
        n20851) );
  INV_X1 U23812 ( .A(n20854), .ZN(n20839) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20851), .B1(
        n20839), .B2(n21263), .ZN(n20833) );
  OAI211_X1 U23814 ( .C1(n21266), .C2(n20883), .A(n20834), .B(n20833), .ZN(
        P1_U3041) );
  AOI22_X1 U23815 ( .A1(n20849), .A2(n21321), .B1(n21322), .B2(n20848), .ZN(
        n20836) );
  INV_X1 U23816 ( .A(n20883), .ZN(n20850) );
  INV_X1 U23817 ( .A(n21270), .ZN(n21323) );
  AOI22_X1 U23818 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20851), .B1(
        n20850), .B2(n21323), .ZN(n20835) );
  OAI211_X1 U23819 ( .C1(n21326), .C2(n20854), .A(n20836), .B(n20835), .ZN(
        P1_U3042) );
  AOI22_X1 U23820 ( .A1(n20849), .A2(n21327), .B1(n21328), .B2(n20848), .ZN(
        n20838) );
  AOI22_X1 U23821 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20851), .B1(
        n20839), .B2(n21271), .ZN(n20837) );
  OAI211_X1 U23822 ( .C1(n21274), .C2(n20883), .A(n20838), .B(n20837), .ZN(
        P1_U3043) );
  AOI22_X1 U23823 ( .A1(n20849), .A2(n21333), .B1(n21334), .B2(n20848), .ZN(
        n20841) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20851), .B1(
        n20839), .B2(n21275), .ZN(n20840) );
  OAI211_X1 U23825 ( .C1(n21278), .C2(n20883), .A(n20841), .B(n20840), .ZN(
        P1_U3044) );
  AOI22_X1 U23826 ( .A1(n20849), .A2(n21339), .B1(n21340), .B2(n20848), .ZN(
        n20843) );
  INV_X1 U23827 ( .A(n21282), .ZN(n21341) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20851), .B1(
        n20850), .B2(n21341), .ZN(n20842) );
  OAI211_X1 U23829 ( .C1(n21344), .C2(n20854), .A(n20843), .B(n20842), .ZN(
        P1_U3045) );
  AOI22_X1 U23830 ( .A1(n20849), .A2(n21345), .B1(n21346), .B2(n20848), .ZN(
        n20845) );
  INV_X1 U23831 ( .A(n21286), .ZN(n21347) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20851), .B1(
        n20850), .B2(n21347), .ZN(n20844) );
  OAI211_X1 U23833 ( .C1(n21350), .C2(n20854), .A(n20845), .B(n20844), .ZN(
        P1_U3046) );
  AOI22_X1 U23834 ( .A1(n20849), .A2(n21351), .B1(n21352), .B2(n20848), .ZN(
        n20847) );
  INV_X1 U23835 ( .A(n21290), .ZN(n21353) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20851), .B1(
        n20850), .B2(n21353), .ZN(n20846) );
  OAI211_X1 U23837 ( .C1(n21356), .C2(n20854), .A(n20847), .B(n20846), .ZN(
        P1_U3047) );
  AOI22_X1 U23838 ( .A1(n20849), .A2(n21358), .B1(n21360), .B2(n20848), .ZN(
        n20853) );
  INV_X1 U23839 ( .A(n21298), .ZN(n21361) );
  AOI22_X1 U23840 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20851), .B1(
        n20850), .B2(n21361), .ZN(n20852) );
  OAI211_X1 U23841 ( .C1(n21367), .C2(n20854), .A(n20853), .B(n20852), .ZN(
        P1_U3048) );
  NAND2_X1 U23842 ( .A1(n20971), .A2(n20855), .ZN(n20996) );
  OR3_X1 U23843 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21302), .A3(
        n20892), .ZN(n20882) );
  OAI22_X1 U23844 ( .A1(n20932), .A2(n21266), .B1(n21116), .B2(n20882), .ZN(
        n20856) );
  INV_X1 U23845 ( .A(n20856), .ZN(n20863) );
  NAND3_X1 U23846 ( .A1(n20932), .A2(n20883), .A3(n9694), .ZN(n20857) );
  NAND2_X1 U23847 ( .A1(n20857), .A2(n21199), .ZN(n20859) );
  OR2_X1 U23848 ( .A1(n20895), .A2(n13858), .ZN(n20860) );
  AOI22_X1 U23849 ( .A1(n20859), .A2(n20860), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20882), .ZN(n20858) );
  OR2_X1 U23850 ( .A1(n21120), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21004) );
  NAND2_X1 U23851 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21004), .ZN(n21001) );
  NAND3_X1 U23852 ( .A1(n21123), .A2(n20858), .A3(n21001), .ZN(n20886) );
  INV_X1 U23853 ( .A(n20859), .ZN(n20861) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20886), .B1(
        n21309), .B2(n20885), .ZN(n20862) );
  OAI211_X1 U23855 ( .C1(n21320), .C2(n20883), .A(n20863), .B(n20862), .ZN(
        P1_U3049) );
  OAI22_X1 U23856 ( .A1(n20932), .A2(n21270), .B1(n21131), .B2(n20882), .ZN(
        n20864) );
  INV_X1 U23857 ( .A(n20864), .ZN(n20866) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20886), .B1(
        n21321), .B2(n20885), .ZN(n20865) );
  OAI211_X1 U23859 ( .C1(n21326), .C2(n20883), .A(n20866), .B(n20865), .ZN(
        P1_U3050) );
  OAI22_X1 U23860 ( .A1(n20883), .A2(n21332), .B1(n21135), .B2(n20882), .ZN(
        n20867) );
  INV_X1 U23861 ( .A(n20867), .ZN(n20869) );
  AOI22_X1 U23862 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20886), .B1(
        n21327), .B2(n20885), .ZN(n20868) );
  OAI211_X1 U23863 ( .C1(n21274), .C2(n20932), .A(n20869), .B(n20868), .ZN(
        P1_U3051) );
  OAI22_X1 U23864 ( .A1(n20932), .A2(n21278), .B1(n21139), .B2(n20882), .ZN(
        n20870) );
  INV_X1 U23865 ( .A(n20870), .ZN(n20872) );
  AOI22_X1 U23866 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20886), .B1(
        n21333), .B2(n20885), .ZN(n20871) );
  OAI211_X1 U23867 ( .C1(n21338), .C2(n20883), .A(n20872), .B(n20871), .ZN(
        P1_U3052) );
  OAI22_X1 U23868 ( .A1(n20932), .A2(n21282), .B1(n21143), .B2(n20882), .ZN(
        n20873) );
  INV_X1 U23869 ( .A(n20873), .ZN(n20875) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20886), .B1(
        n21339), .B2(n20885), .ZN(n20874) );
  OAI211_X1 U23871 ( .C1(n21344), .C2(n20883), .A(n20875), .B(n20874), .ZN(
        P1_U3053) );
  OAI22_X1 U23872 ( .A1(n20932), .A2(n21286), .B1(n21147), .B2(n20882), .ZN(
        n20876) );
  INV_X1 U23873 ( .A(n20876), .ZN(n20878) );
  AOI22_X1 U23874 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20886), .B1(
        n21345), .B2(n20885), .ZN(n20877) );
  OAI211_X1 U23875 ( .C1(n21350), .C2(n20883), .A(n20878), .B(n20877), .ZN(
        P1_U3054) );
  OAI22_X1 U23876 ( .A1(n20883), .A2(n21356), .B1(n21151), .B2(n20882), .ZN(
        n20879) );
  INV_X1 U23877 ( .A(n20879), .ZN(n20881) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20886), .B1(
        n21351), .B2(n20885), .ZN(n20880) );
  OAI211_X1 U23879 ( .C1(n21290), .C2(n20932), .A(n20881), .B(n20880), .ZN(
        P1_U3055) );
  OAI22_X1 U23880 ( .A1(n20883), .A2(n21367), .B1(n21156), .B2(n20882), .ZN(
        n20884) );
  INV_X1 U23881 ( .A(n20884), .ZN(n20888) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20886), .B1(
        n21358), .B2(n20885), .ZN(n20887) );
  OAI211_X1 U23883 ( .C1(n21298), .C2(n20932), .A(n20888), .B(n20887), .ZN(
        P1_U3056) );
  INV_X1 U23884 ( .A(n21163), .ZN(n20889) );
  INV_X1 U23885 ( .A(n20892), .ZN(n20890) );
  NAND2_X1 U23886 ( .A1(n21300), .A2(n20890), .ZN(n20926) );
  OAI22_X1 U23887 ( .A1(n20932), .A2(n21320), .B1(n21116), .B2(n20926), .ZN(
        n20891) );
  INV_X1 U23888 ( .A(n20891), .ZN(n20907) );
  NOR2_X1 U23889 ( .A1(n21302), .A2(n20892), .ZN(n20902) );
  AND2_X1 U23890 ( .A1(n20894), .A2(n20893), .ZN(n21167) );
  INV_X1 U23891 ( .A(n21167), .ZN(n21307) );
  OR2_X1 U23892 ( .A1(n20895), .A2(n21307), .ZN(n20896) );
  INV_X1 U23893 ( .A(n20897), .ZN(n20899) );
  OAI21_X1 U23894 ( .B1(n20899), .B2(n21304), .A(n20898), .ZN(n20903) );
  NAND2_X1 U23895 ( .A1(n20901), .A2(n20903), .ZN(n20900) );
  OAI211_X1 U23896 ( .C1(n9694), .C2(n20902), .A(n21314), .B(n20900), .ZN(
        n20929) );
  INV_X1 U23897 ( .A(n20901), .ZN(n20904) );
  AOI22_X1 U23898 ( .A1(n20904), .A2(n20903), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20902), .ZN(n20905) );
  AOI22_X1 U23899 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20929), .B1(
        n21309), .B2(n20928), .ZN(n20906) );
  OAI211_X1 U23900 ( .C1(n21266), .C2(n20942), .A(n20907), .B(n20906), .ZN(
        P1_U3057) );
  OAI22_X1 U23901 ( .A1(n20932), .A2(n21326), .B1(n21131), .B2(n20926), .ZN(
        n20908) );
  INV_X1 U23902 ( .A(n20908), .ZN(n20910) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20929), .B1(
        n21321), .B2(n20928), .ZN(n20909) );
  OAI211_X1 U23904 ( .C1(n21270), .C2(n20942), .A(n20910), .B(n20909), .ZN(
        P1_U3058) );
  OAI22_X1 U23905 ( .A1(n20942), .A2(n21274), .B1(n21135), .B2(n20926), .ZN(
        n20911) );
  INV_X1 U23906 ( .A(n20911), .ZN(n20913) );
  AOI22_X1 U23907 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20929), .B1(
        n21327), .B2(n20928), .ZN(n20912) );
  OAI211_X1 U23908 ( .C1(n21332), .C2(n20932), .A(n20913), .B(n20912), .ZN(
        P1_U3059) );
  OAI22_X1 U23909 ( .A1(n20932), .A2(n21338), .B1(n21139), .B2(n20926), .ZN(
        n20914) );
  INV_X1 U23910 ( .A(n20914), .ZN(n20916) );
  AOI22_X1 U23911 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20929), .B1(
        n21333), .B2(n20928), .ZN(n20915) );
  OAI211_X1 U23912 ( .C1(n21278), .C2(n20942), .A(n20916), .B(n20915), .ZN(
        P1_U3060) );
  OAI22_X1 U23913 ( .A1(n20942), .A2(n21282), .B1(n21143), .B2(n20926), .ZN(
        n20917) );
  INV_X1 U23914 ( .A(n20917), .ZN(n20919) );
  AOI22_X1 U23915 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20929), .B1(
        n21339), .B2(n20928), .ZN(n20918) );
  OAI211_X1 U23916 ( .C1(n21344), .C2(n20932), .A(n20919), .B(n20918), .ZN(
        P1_U3061) );
  OAI22_X1 U23917 ( .A1(n20942), .A2(n21286), .B1(n21147), .B2(n20926), .ZN(
        n20920) );
  INV_X1 U23918 ( .A(n20920), .ZN(n20922) );
  AOI22_X1 U23919 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20929), .B1(
        n21345), .B2(n20928), .ZN(n20921) );
  OAI211_X1 U23920 ( .C1(n21350), .C2(n20932), .A(n20922), .B(n20921), .ZN(
        P1_U3062) );
  OAI22_X1 U23921 ( .A1(n20942), .A2(n21290), .B1(n21151), .B2(n20926), .ZN(
        n20923) );
  INV_X1 U23922 ( .A(n20923), .ZN(n20925) );
  AOI22_X1 U23923 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20929), .B1(
        n21351), .B2(n20928), .ZN(n20924) );
  OAI211_X1 U23924 ( .C1(n21356), .C2(n20932), .A(n20925), .B(n20924), .ZN(
        P1_U3063) );
  OAI22_X1 U23925 ( .A1(n20942), .A2(n21298), .B1(n21156), .B2(n20926), .ZN(
        n20927) );
  INV_X1 U23926 ( .A(n20927), .ZN(n20931) );
  AOI22_X1 U23927 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20929), .B1(
        n21358), .B2(n20928), .ZN(n20930) );
  OAI211_X1 U23928 ( .C1(n21367), .C2(n20932), .A(n20931), .B(n20930), .ZN(
        P1_U3064) );
  INV_X1 U23929 ( .A(n20933), .ZN(n20934) );
  AND2_X1 U23930 ( .A1(n20935), .A2(n20934), .ZN(n20937) );
  OR2_X1 U23931 ( .A1(n13843), .A2(n20939), .ZN(n21000) );
  NAND2_X1 U23932 ( .A1(n13858), .A2(n9694), .ZN(n20941) );
  OAI22_X1 U23933 ( .A1(n21000), .A2(n20941), .B1(n20940), .B2(n21254), .ZN(
        n20962) );
  AOI22_X1 U23934 ( .A1(n21310), .A2(n9828), .B1(n21309), .B2(n20962), .ZN(
        n20949) );
  INV_X1 U23935 ( .A(n20995), .ZN(n20943) );
  OAI21_X1 U23936 ( .B1(n20963), .B2(n20943), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20944) );
  OAI21_X1 U23937 ( .B1(n21256), .B2(n21000), .A(n20944), .ZN(n20947) );
  AOI22_X1 U23938 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21263), .ZN(n20948) );
  OAI211_X1 U23939 ( .C1(n21266), .C2(n20995), .A(n20949), .B(n20948), .ZN(
        P1_U3065) );
  AOI22_X1 U23940 ( .A1(n21322), .A2(n9828), .B1(n21321), .B2(n20962), .ZN(
        n20951) );
  AOI22_X1 U23941 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21267), .ZN(n20950) );
  OAI211_X1 U23942 ( .C1(n21270), .C2(n20995), .A(n20951), .B(n20950), .ZN(
        P1_U3066) );
  AOI22_X1 U23943 ( .A1(n21328), .A2(n9828), .B1(n21327), .B2(n20962), .ZN(
        n20953) );
  AOI22_X1 U23944 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21271), .ZN(n20952) );
  OAI211_X1 U23945 ( .C1(n21274), .C2(n20995), .A(n20953), .B(n20952), .ZN(
        P1_U3067) );
  AOI22_X1 U23946 ( .A1(n21334), .A2(n9828), .B1(n21333), .B2(n20962), .ZN(
        n20955) );
  AOI22_X1 U23947 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21275), .ZN(n20954) );
  OAI211_X1 U23948 ( .C1(n21278), .C2(n20995), .A(n20955), .B(n20954), .ZN(
        P1_U3068) );
  AOI22_X1 U23949 ( .A1(n21340), .A2(n9828), .B1(n21339), .B2(n20962), .ZN(
        n20957) );
  AOI22_X1 U23950 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21279), .ZN(n20956) );
  OAI211_X1 U23951 ( .C1(n21282), .C2(n20995), .A(n20957), .B(n20956), .ZN(
        P1_U3069) );
  AOI22_X1 U23952 ( .A1(n21346), .A2(n9828), .B1(n21345), .B2(n20962), .ZN(
        n20959) );
  AOI22_X1 U23953 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21283), .ZN(n20958) );
  OAI211_X1 U23954 ( .C1(n21286), .C2(n20995), .A(n20959), .B(n20958), .ZN(
        P1_U3070) );
  AOI22_X1 U23955 ( .A1(n21352), .A2(n9828), .B1(n21351), .B2(n20962), .ZN(
        n20961) );
  AOI22_X1 U23956 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21287), .ZN(n20960) );
  OAI211_X1 U23957 ( .C1(n21290), .C2(n20995), .A(n20961), .B(n20960), .ZN(
        P1_U3071) );
  AOI22_X1 U23958 ( .A1(n21360), .A2(n9828), .B1(n21358), .B2(n20962), .ZN(
        n20966) );
  AOI22_X1 U23959 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20964), .B1(
        n20963), .B2(n21293), .ZN(n20965) );
  OAI211_X1 U23960 ( .C1(n21298), .C2(n20995), .A(n20966), .B(n20965), .ZN(
        P1_U3072) );
  NOR2_X1 U23961 ( .A1(n20997), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20972) );
  INV_X1 U23962 ( .A(n20972), .ZN(n20967) );
  NOR2_X1 U23963 ( .A1(n21677), .A2(n20967), .ZN(n20990) );
  INV_X1 U23964 ( .A(n21000), .ZN(n21036) );
  AOI21_X1 U23965 ( .B1(n21036), .B2(n21091), .A(n20990), .ZN(n20968) );
  OAI22_X1 U23966 ( .A1(n20968), .A2(n21304), .B1(n20967), .B2(n21306), .ZN(
        n20989) );
  AOI22_X1 U23967 ( .A1(n21310), .A2(n20990), .B1(n21309), .B2(n20989), .ZN(
        n20976) );
  INV_X1 U23968 ( .A(n20969), .ZN(n20970) );
  NOR2_X1 U23969 ( .A1(n20971), .A2(n20970), .ZN(n21230) );
  AND2_X1 U23970 ( .A1(n21034), .A2(n21230), .ZN(n20973) );
  INV_X1 U23971 ( .A(n21266), .ZN(n21317) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21317), .ZN(n20975) );
  OAI211_X1 U23973 ( .C1(n21320), .C2(n20995), .A(n20976), .B(n20975), .ZN(
        P1_U3073) );
  AOI22_X1 U23974 ( .A1(n21322), .A2(n20990), .B1(n21321), .B2(n20989), .ZN(
        n20978) );
  AOI22_X1 U23975 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21323), .ZN(n20977) );
  OAI211_X1 U23976 ( .C1(n21326), .C2(n20995), .A(n20978), .B(n20977), .ZN(
        P1_U3074) );
  AOI22_X1 U23977 ( .A1(n21328), .A2(n20990), .B1(n21327), .B2(n20989), .ZN(
        n20980) );
  INV_X1 U23978 ( .A(n21274), .ZN(n21329) );
  AOI22_X1 U23979 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21329), .ZN(n20979) );
  OAI211_X1 U23980 ( .C1(n21332), .C2(n20995), .A(n20980), .B(n20979), .ZN(
        P1_U3075) );
  AOI22_X1 U23981 ( .A1(n21334), .A2(n20990), .B1(n21333), .B2(n20989), .ZN(
        n20982) );
  INV_X1 U23982 ( .A(n21278), .ZN(n21335) );
  AOI22_X1 U23983 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21335), .ZN(n20981) );
  OAI211_X1 U23984 ( .C1(n21338), .C2(n20995), .A(n20982), .B(n20981), .ZN(
        P1_U3076) );
  AOI22_X1 U23985 ( .A1(n21340), .A2(n20990), .B1(n21339), .B2(n20989), .ZN(
        n20984) );
  AOI22_X1 U23986 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21341), .ZN(n20983) );
  OAI211_X1 U23987 ( .C1(n21344), .C2(n20995), .A(n20984), .B(n20983), .ZN(
        P1_U3077) );
  AOI22_X1 U23988 ( .A1(n21346), .A2(n20990), .B1(n21345), .B2(n20989), .ZN(
        n20986) );
  AOI22_X1 U23989 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21347), .ZN(n20985) );
  OAI211_X1 U23990 ( .C1(n21350), .C2(n20995), .A(n20986), .B(n20985), .ZN(
        P1_U3078) );
  AOI22_X1 U23991 ( .A1(n21352), .A2(n20990), .B1(n21351), .B2(n20989), .ZN(
        n20988) );
  AOI22_X1 U23992 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21353), .ZN(n20987) );
  OAI211_X1 U23993 ( .C1(n21356), .C2(n20995), .A(n20988), .B(n20987), .ZN(
        P1_U3079) );
  AOI22_X1 U23994 ( .A1(n21360), .A2(n20990), .B1(n21358), .B2(n20989), .ZN(
        n20994) );
  AOI22_X1 U23995 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20992), .B1(
        n20991), .B2(n21361), .ZN(n20993) );
  OAI211_X1 U23996 ( .C1(n21367), .C2(n20995), .A(n20994), .B(n20993), .ZN(
        P1_U3080) );
  NOR2_X1 U23997 ( .A1(n21302), .A2(n20997), .ZN(n21042) );
  INV_X1 U23998 ( .A(n21042), .ZN(n21037) );
  OAI22_X1 U23999 ( .A1(n21028), .A2(n21320), .B1(n21116), .B2(n21027), .ZN(
        n20998) );
  INV_X1 U24000 ( .A(n20998), .ZN(n21008) );
  NAND3_X1 U24001 ( .A1(n21064), .A2(n21028), .A3(n9694), .ZN(n20999) );
  NAND2_X1 U24002 ( .A1(n20999), .A2(n21199), .ZN(n21003) );
  OR2_X1 U24003 ( .A1(n21000), .A2(n13858), .ZN(n21005) );
  AOI22_X1 U24004 ( .A1(n21003), .A2(n21005), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21027), .ZN(n21002) );
  NAND3_X1 U24005 ( .A1(n21260), .A2(n21002), .A3(n21001), .ZN(n21031) );
  INV_X1 U24006 ( .A(n21003), .ZN(n21006) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21031), .B1(
        n21309), .B2(n21030), .ZN(n21007) );
  OAI211_X1 U24008 ( .C1(n21266), .C2(n21064), .A(n21008), .B(n21007), .ZN(
        P1_U3081) );
  OAI22_X1 U24009 ( .A1(n21028), .A2(n21326), .B1(n21131), .B2(n21027), .ZN(
        n21009) );
  INV_X1 U24010 ( .A(n21009), .ZN(n21011) );
  AOI22_X1 U24011 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21031), .B1(
        n21321), .B2(n21030), .ZN(n21010) );
  OAI211_X1 U24012 ( .C1(n21270), .C2(n21064), .A(n21011), .B(n21010), .ZN(
        P1_U3082) );
  OAI22_X1 U24013 ( .A1(n21064), .A2(n21274), .B1(n21135), .B2(n21027), .ZN(
        n21012) );
  INV_X1 U24014 ( .A(n21012), .ZN(n21014) );
  AOI22_X1 U24015 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21031), .B1(
        n21327), .B2(n21030), .ZN(n21013) );
  OAI211_X1 U24016 ( .C1(n21332), .C2(n21028), .A(n21014), .B(n21013), .ZN(
        P1_U3083) );
  OAI22_X1 U24017 ( .A1(n21064), .A2(n21278), .B1(n21139), .B2(n21027), .ZN(
        n21015) );
  INV_X1 U24018 ( .A(n21015), .ZN(n21017) );
  AOI22_X1 U24019 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21031), .B1(
        n21333), .B2(n21030), .ZN(n21016) );
  OAI211_X1 U24020 ( .C1(n21338), .C2(n21028), .A(n21017), .B(n21016), .ZN(
        P1_U3084) );
  OAI22_X1 U24021 ( .A1(n21064), .A2(n21282), .B1(n21143), .B2(n21027), .ZN(
        n21018) );
  INV_X1 U24022 ( .A(n21018), .ZN(n21020) );
  AOI22_X1 U24023 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21031), .B1(
        n21339), .B2(n21030), .ZN(n21019) );
  OAI211_X1 U24024 ( .C1(n21344), .C2(n21028), .A(n21020), .B(n21019), .ZN(
        P1_U3085) );
  OAI22_X1 U24025 ( .A1(n21028), .A2(n21350), .B1(n21147), .B2(n21027), .ZN(
        n21021) );
  INV_X1 U24026 ( .A(n21021), .ZN(n21023) );
  AOI22_X1 U24027 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21031), .B1(
        n21345), .B2(n21030), .ZN(n21022) );
  OAI211_X1 U24028 ( .C1(n21286), .C2(n21064), .A(n21023), .B(n21022), .ZN(
        P1_U3086) );
  OAI22_X1 U24029 ( .A1(n21028), .A2(n21356), .B1(n21151), .B2(n21027), .ZN(
        n21024) );
  INV_X1 U24030 ( .A(n21024), .ZN(n21026) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21031), .B1(
        n21351), .B2(n21030), .ZN(n21025) );
  OAI211_X1 U24032 ( .C1(n21290), .C2(n21064), .A(n21026), .B(n21025), .ZN(
        P1_U3087) );
  OAI22_X1 U24033 ( .A1(n21028), .A2(n21367), .B1(n21156), .B2(n21027), .ZN(
        n21029) );
  INV_X1 U24034 ( .A(n21029), .ZN(n21033) );
  AOI22_X1 U24035 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21031), .B1(
        n21358), .B2(n21030), .ZN(n21032) );
  OAI211_X1 U24036 ( .C1(n21298), .C2(n21064), .A(n21033), .B(n21032), .ZN(
        P1_U3088) );
  NAND2_X1 U24037 ( .A1(n21034), .A2(n21163), .ZN(n21050) );
  AOI21_X1 U24038 ( .B1(n21036), .B2(n21167), .A(n21060), .ZN(n21040) );
  OAI22_X1 U24039 ( .A1(n21040), .A2(n21304), .B1(n21037), .B2(n21306), .ZN(
        n21059) );
  AOI22_X1 U24040 ( .A1(n21060), .A2(n21310), .B1(n21059), .B2(n21309), .ZN(
        n21044) );
  OR2_X1 U24041 ( .A1(n21039), .A2(n21038), .ZN(n21462) );
  NAND2_X1 U24042 ( .A1(n21040), .A2(n21462), .ZN(n21041) );
  OAI221_X1 U24043 ( .B1(n9694), .B2(n21042), .C1(n21304), .C2(n21041), .A(
        n21314), .ZN(n21061) );
  INV_X1 U24044 ( .A(n21064), .ZN(n21047) );
  AOI22_X1 U24045 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21061), .B1(
        n21047), .B2(n21263), .ZN(n21043) );
  OAI211_X1 U24046 ( .C1(n21266), .C2(n21050), .A(n21044), .B(n21043), .ZN(
        P1_U3089) );
  AOI22_X1 U24047 ( .A1(n21060), .A2(n21322), .B1(n21059), .B2(n21321), .ZN(
        n21046) );
  AOI22_X1 U24048 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21061), .B1(
        n21087), .B2(n21323), .ZN(n21045) );
  OAI211_X1 U24049 ( .C1(n21326), .C2(n21064), .A(n21046), .B(n21045), .ZN(
        P1_U3090) );
  AOI22_X1 U24050 ( .A1(n21060), .A2(n21328), .B1(n21059), .B2(n21327), .ZN(
        n21049) );
  AOI22_X1 U24051 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21061), .B1(
        n21047), .B2(n21271), .ZN(n21048) );
  OAI211_X1 U24052 ( .C1(n21274), .C2(n21050), .A(n21049), .B(n21048), .ZN(
        P1_U3091) );
  AOI22_X1 U24053 ( .A1(n21060), .A2(n21334), .B1(n21059), .B2(n21333), .ZN(
        n21052) );
  AOI22_X1 U24054 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21061), .B1(
        n21087), .B2(n21335), .ZN(n21051) );
  OAI211_X1 U24055 ( .C1(n21338), .C2(n21064), .A(n21052), .B(n21051), .ZN(
        P1_U3092) );
  AOI22_X1 U24056 ( .A1(n21060), .A2(n21340), .B1(n21059), .B2(n21339), .ZN(
        n21054) );
  AOI22_X1 U24057 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21061), .B1(
        n21087), .B2(n21341), .ZN(n21053) );
  OAI211_X1 U24058 ( .C1(n21344), .C2(n21064), .A(n21054), .B(n21053), .ZN(
        P1_U3093) );
  AOI22_X1 U24059 ( .A1(n21060), .A2(n21346), .B1(n21059), .B2(n21345), .ZN(
        n21056) );
  AOI22_X1 U24060 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21061), .B1(
        n21087), .B2(n21347), .ZN(n21055) );
  OAI211_X1 U24061 ( .C1(n21350), .C2(n21064), .A(n21056), .B(n21055), .ZN(
        P1_U3094) );
  AOI22_X1 U24062 ( .A1(n21060), .A2(n21352), .B1(n21059), .B2(n21351), .ZN(
        n21058) );
  AOI22_X1 U24063 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21061), .B1(
        n21087), .B2(n21353), .ZN(n21057) );
  OAI211_X1 U24064 ( .C1(n21356), .C2(n21064), .A(n21058), .B(n21057), .ZN(
        P1_U3095) );
  AOI22_X1 U24065 ( .A1(n21060), .A2(n21360), .B1(n21059), .B2(n21358), .ZN(
        n21063) );
  AOI22_X1 U24066 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21061), .B1(
        n21087), .B2(n21361), .ZN(n21062) );
  OAI211_X1 U24067 ( .C1(n21367), .C2(n21064), .A(n21063), .B(n21062), .ZN(
        P1_U3096) );
  AND2_X1 U24068 ( .A1(n21464), .A2(n13843), .ZN(n21168) );
  NAND2_X1 U24069 ( .A1(n21066), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21165) );
  AOI21_X1 U24070 ( .B1(n21168), .B2(n13858), .A(n10408), .ZN(n21069) );
  NAND2_X1 U24071 ( .A1(n21067), .A2(n21120), .ZN(n21204) );
  OAI22_X1 U24072 ( .A1(n21069), .A2(n21304), .B1(n21126), .B2(n21204), .ZN(
        n21086) );
  AOI22_X1 U24073 ( .A1(n21086), .A2(n21309), .B1(n21310), .B2(n10408), .ZN(
        n21073) );
  INV_X1 U24074 ( .A(n21115), .ZN(n21068) );
  OAI21_X1 U24075 ( .B1(n21068), .B2(n21087), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21070) );
  NAND2_X1 U24076 ( .A1(n21070), .A2(n21069), .ZN(n21071) );
  AOI22_X1 U24077 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21263), .ZN(n21072) );
  OAI211_X1 U24078 ( .C1(n21266), .C2(n21115), .A(n21073), .B(n21072), .ZN(
        P1_U3097) );
  AOI22_X1 U24079 ( .A1(n21086), .A2(n21321), .B1(n21322), .B2(n10408), .ZN(
        n21075) );
  AOI22_X1 U24080 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21267), .ZN(n21074) );
  OAI211_X1 U24081 ( .C1(n21270), .C2(n21115), .A(n21075), .B(n21074), .ZN(
        P1_U3098) );
  AOI22_X1 U24082 ( .A1(n21086), .A2(n21327), .B1(n21328), .B2(n10408), .ZN(
        n21077) );
  AOI22_X1 U24083 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21271), .ZN(n21076) );
  OAI211_X1 U24084 ( .C1(n21274), .C2(n21115), .A(n21077), .B(n21076), .ZN(
        P1_U3099) );
  AOI22_X1 U24085 ( .A1(n21086), .A2(n21333), .B1(n21334), .B2(n10408), .ZN(
        n21079) );
  AOI22_X1 U24086 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21275), .ZN(n21078) );
  OAI211_X1 U24087 ( .C1(n21278), .C2(n21115), .A(n21079), .B(n21078), .ZN(
        P1_U3100) );
  AOI22_X1 U24088 ( .A1(n21086), .A2(n21339), .B1(n21340), .B2(n10408), .ZN(
        n21081) );
  AOI22_X1 U24089 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21279), .ZN(n21080) );
  OAI211_X1 U24090 ( .C1(n21282), .C2(n21115), .A(n21081), .B(n21080), .ZN(
        P1_U3101) );
  AOI22_X1 U24091 ( .A1(n21086), .A2(n21345), .B1(n21346), .B2(n10408), .ZN(
        n21083) );
  AOI22_X1 U24092 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21283), .ZN(n21082) );
  OAI211_X1 U24093 ( .C1(n21286), .C2(n21115), .A(n21083), .B(n21082), .ZN(
        P1_U3102) );
  AOI22_X1 U24094 ( .A1(n21086), .A2(n21351), .B1(n21352), .B2(n10408), .ZN(
        n21085) );
  AOI22_X1 U24095 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21287), .ZN(n21084) );
  OAI211_X1 U24096 ( .C1(n21290), .C2(n21115), .A(n21085), .B(n21084), .ZN(
        P1_U3103) );
  AOI22_X1 U24097 ( .A1(n21086), .A2(n21358), .B1(n21360), .B2(n10408), .ZN(
        n21090) );
  AOI22_X1 U24098 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21088), .B1(
        n21087), .B2(n21293), .ZN(n21089) );
  OAI211_X1 U24099 ( .C1(n21298), .C2(n21115), .A(n21090), .B(n21089), .ZN(
        P1_U3104) );
  NOR2_X1 U24100 ( .A1(n21165), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21095) );
  INV_X1 U24101 ( .A(n21095), .ZN(n21092) );
  NOR2_X1 U24102 ( .A1(n21677), .A2(n21092), .ZN(n21110) );
  AOI21_X1 U24103 ( .B1(n21168), .B2(n21091), .A(n21110), .ZN(n21093) );
  OAI22_X1 U24104 ( .A1(n21093), .A2(n21304), .B1(n21092), .B2(n21306), .ZN(
        n21111) );
  AOI22_X1 U24105 ( .A1(n21111), .A2(n21309), .B1(n21310), .B2(n21110), .ZN(
        n21097) );
  NAND2_X1 U24106 ( .A1(n21164), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21172) );
  NAND3_X1 U24107 ( .A1(n21172), .A2(n21093), .A3(n9694), .ZN(n21094) );
  OAI211_X1 U24108 ( .C1(n9694), .C2(n21095), .A(n21314), .B(n21094), .ZN(
        n21112) );
  AOI22_X1 U24109 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21317), .ZN(n21096) );
  OAI211_X1 U24110 ( .C1(n21320), .C2(n21115), .A(n21097), .B(n21096), .ZN(
        P1_U3105) );
  AOI22_X1 U24111 ( .A1(n21111), .A2(n21321), .B1(n21322), .B2(n21110), .ZN(
        n21099) );
  AOI22_X1 U24112 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21323), .ZN(n21098) );
  OAI211_X1 U24113 ( .C1(n21326), .C2(n21115), .A(n21099), .B(n21098), .ZN(
        P1_U3106) );
  AOI22_X1 U24114 ( .A1(n21111), .A2(n21327), .B1(n21328), .B2(n21110), .ZN(
        n21101) );
  AOI22_X1 U24115 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21329), .ZN(n21100) );
  OAI211_X1 U24116 ( .C1(n21332), .C2(n21115), .A(n21101), .B(n21100), .ZN(
        P1_U3107) );
  AOI22_X1 U24117 ( .A1(n21111), .A2(n21333), .B1(n21334), .B2(n21110), .ZN(
        n21103) );
  AOI22_X1 U24118 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21335), .ZN(n21102) );
  OAI211_X1 U24119 ( .C1(n21338), .C2(n21115), .A(n21103), .B(n21102), .ZN(
        P1_U3108) );
  AOI22_X1 U24120 ( .A1(n21111), .A2(n21339), .B1(n21340), .B2(n21110), .ZN(
        n21105) );
  AOI22_X1 U24121 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21341), .ZN(n21104) );
  OAI211_X1 U24122 ( .C1(n21344), .C2(n21115), .A(n21105), .B(n21104), .ZN(
        P1_U3109) );
  AOI22_X1 U24123 ( .A1(n21111), .A2(n21345), .B1(n21346), .B2(n21110), .ZN(
        n21107) );
  AOI22_X1 U24124 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21347), .ZN(n21106) );
  OAI211_X1 U24125 ( .C1(n21350), .C2(n21115), .A(n21107), .B(n21106), .ZN(
        P1_U3110) );
  AOI22_X1 U24126 ( .A1(n21111), .A2(n21351), .B1(n21352), .B2(n21110), .ZN(
        n21109) );
  AOI22_X1 U24127 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21353), .ZN(n21108) );
  OAI211_X1 U24128 ( .C1(n21356), .C2(n21115), .A(n21109), .B(n21108), .ZN(
        P1_U3111) );
  AOI22_X1 U24129 ( .A1(n21111), .A2(n21358), .B1(n21360), .B2(n21110), .ZN(
        n21114) );
  AOI22_X1 U24130 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21112), .B1(
        n21118), .B2(n21361), .ZN(n21113) );
  OAI211_X1 U24131 ( .C1(n21367), .C2(n21115), .A(n21114), .B(n21113), .ZN(
        P1_U3112) );
  NOR2_X1 U24132 ( .A1(n21302), .A2(n21165), .ZN(n21174) );
  INV_X1 U24133 ( .A(n21174), .ZN(n21169) );
  NOR2_X1 U24134 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21169), .ZN(
        n21121) );
  INV_X1 U24135 ( .A(n21121), .ZN(n21155) );
  OAI22_X1 U24136 ( .A1(n21157), .A2(n21320), .B1(n21116), .B2(n21155), .ZN(
        n21117) );
  INV_X1 U24137 ( .A(n21117), .ZN(n21130) );
  OAI21_X1 U24138 ( .B1(n21193), .B2(n21118), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21119) );
  NAND2_X1 U24139 ( .A1(n21119), .A2(n9694), .ZN(n21128) );
  AND2_X1 U24140 ( .A1(n21168), .A2(n21256), .ZN(n21125) );
  OR2_X1 U24141 ( .A1(n21120), .A2(n21474), .ZN(n21253) );
  NAND2_X1 U24142 ( .A1(n21253), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21259) );
  OAI21_X1 U24143 ( .B1(n21660), .B2(n21121), .A(n21259), .ZN(n21122) );
  INV_X1 U24144 ( .A(n21122), .ZN(n21124) );
  INV_X1 U24145 ( .A(n21125), .ZN(n21127) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21160), .B1(
        n21309), .B2(n21159), .ZN(n21129) );
  OAI211_X1 U24147 ( .C1(n21266), .C2(n21188), .A(n21130), .B(n21129), .ZN(
        P1_U3113) );
  OAI22_X1 U24148 ( .A1(n21157), .A2(n21326), .B1(n21131), .B2(n21155), .ZN(
        n21132) );
  INV_X1 U24149 ( .A(n21132), .ZN(n21134) );
  AOI22_X1 U24150 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21160), .B1(
        n21321), .B2(n21159), .ZN(n21133) );
  OAI211_X1 U24151 ( .C1(n21270), .C2(n21188), .A(n21134), .B(n21133), .ZN(
        P1_U3114) );
  OAI22_X1 U24152 ( .A1(n21188), .A2(n21274), .B1(n21135), .B2(n21155), .ZN(
        n21136) );
  INV_X1 U24153 ( .A(n21136), .ZN(n21138) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21160), .B1(
        n21327), .B2(n21159), .ZN(n21137) );
  OAI211_X1 U24155 ( .C1(n21332), .C2(n21157), .A(n21138), .B(n21137), .ZN(
        P1_U3115) );
  OAI22_X1 U24156 ( .A1(n21188), .A2(n21278), .B1(n21139), .B2(n21155), .ZN(
        n21140) );
  INV_X1 U24157 ( .A(n21140), .ZN(n21142) );
  AOI22_X1 U24158 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21160), .B1(
        n21333), .B2(n21159), .ZN(n21141) );
  OAI211_X1 U24159 ( .C1(n21338), .C2(n21157), .A(n21142), .B(n21141), .ZN(
        P1_U3116) );
  OAI22_X1 U24160 ( .A1(n21188), .A2(n21282), .B1(n21143), .B2(n21155), .ZN(
        n21144) );
  INV_X1 U24161 ( .A(n21144), .ZN(n21146) );
  AOI22_X1 U24162 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21160), .B1(
        n21339), .B2(n21159), .ZN(n21145) );
  OAI211_X1 U24163 ( .C1(n21344), .C2(n21157), .A(n21146), .B(n21145), .ZN(
        P1_U3117) );
  OAI22_X1 U24164 ( .A1(n21157), .A2(n21350), .B1(n21147), .B2(n21155), .ZN(
        n21148) );
  INV_X1 U24165 ( .A(n21148), .ZN(n21150) );
  AOI22_X1 U24166 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21160), .B1(
        n21345), .B2(n21159), .ZN(n21149) );
  OAI211_X1 U24167 ( .C1(n21286), .C2(n21188), .A(n21150), .B(n21149), .ZN(
        P1_U3118) );
  OAI22_X1 U24168 ( .A1(n21157), .A2(n21356), .B1(n21151), .B2(n21155), .ZN(
        n21152) );
  INV_X1 U24169 ( .A(n21152), .ZN(n21154) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21160), .B1(
        n21351), .B2(n21159), .ZN(n21153) );
  OAI211_X1 U24171 ( .C1(n21290), .C2(n21188), .A(n21154), .B(n21153), .ZN(
        P1_U3119) );
  OAI22_X1 U24172 ( .A1(n21157), .A2(n21367), .B1(n21156), .B2(n21155), .ZN(
        n21158) );
  INV_X1 U24173 ( .A(n21158), .ZN(n21162) );
  AOI22_X1 U24174 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21160), .B1(
        n21358), .B2(n21159), .ZN(n21161) );
  OAI211_X1 U24175 ( .C1(n21298), .C2(n21188), .A(n21162), .B(n21161), .ZN(
        P1_U3120) );
  NOR2_X1 U24176 ( .A1(n21166), .A2(n21165), .ZN(n21191) );
  AOI21_X1 U24177 ( .B1(n21168), .B2(n21167), .A(n21191), .ZN(n21170) );
  OAI22_X1 U24178 ( .A1(n21170), .A2(n21304), .B1(n21169), .B2(n21306), .ZN(
        n21192) );
  AOI22_X1 U24179 ( .A1(n21192), .A2(n21309), .B1(n21310), .B2(n21191), .ZN(
        n21176) );
  OAI211_X1 U24180 ( .C1(n21172), .C2(n21171), .A(n9694), .B(n21170), .ZN(
        n21173) );
  OAI211_X1 U24181 ( .C1(n9694), .C2(n21174), .A(n21314), .B(n21173), .ZN(
        n21194) );
  AOI22_X1 U24182 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21263), .ZN(n21175) );
  OAI211_X1 U24183 ( .C1(n21266), .C2(n21225), .A(n21176), .B(n21175), .ZN(
        P1_U3121) );
  AOI22_X1 U24184 ( .A1(n21192), .A2(n21321), .B1(n21322), .B2(n21191), .ZN(
        n21178) );
  INV_X1 U24185 ( .A(n21225), .ZN(n21185) );
  AOI22_X1 U24186 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21194), .B1(
        n21185), .B2(n21323), .ZN(n21177) );
  OAI211_X1 U24187 ( .C1(n21326), .C2(n21188), .A(n21178), .B(n21177), .ZN(
        P1_U3122) );
  AOI22_X1 U24188 ( .A1(n21192), .A2(n21327), .B1(n21328), .B2(n21191), .ZN(
        n21180) );
  AOI22_X1 U24189 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21194), .B1(
        n21185), .B2(n21329), .ZN(n21179) );
  OAI211_X1 U24190 ( .C1(n21332), .C2(n21188), .A(n21180), .B(n21179), .ZN(
        P1_U3123) );
  AOI22_X1 U24191 ( .A1(n21192), .A2(n21333), .B1(n21334), .B2(n21191), .ZN(
        n21182) );
  AOI22_X1 U24192 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21275), .ZN(n21181) );
  OAI211_X1 U24193 ( .C1(n21278), .C2(n21225), .A(n21182), .B(n21181), .ZN(
        P1_U3124) );
  AOI22_X1 U24194 ( .A1(n21192), .A2(n21339), .B1(n21340), .B2(n21191), .ZN(
        n21184) );
  AOI22_X1 U24195 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21279), .ZN(n21183) );
  OAI211_X1 U24196 ( .C1(n21282), .C2(n21225), .A(n21184), .B(n21183), .ZN(
        P1_U3125) );
  AOI22_X1 U24197 ( .A1(n21192), .A2(n21345), .B1(n21346), .B2(n21191), .ZN(
        n21187) );
  AOI22_X1 U24198 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21194), .B1(
        n21185), .B2(n21347), .ZN(n21186) );
  OAI211_X1 U24199 ( .C1(n21350), .C2(n21188), .A(n21187), .B(n21186), .ZN(
        P1_U3126) );
  AOI22_X1 U24200 ( .A1(n21192), .A2(n21351), .B1(n21352), .B2(n21191), .ZN(
        n21190) );
  AOI22_X1 U24201 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21287), .ZN(n21189) );
  OAI211_X1 U24202 ( .C1(n21290), .C2(n21225), .A(n21190), .B(n21189), .ZN(
        P1_U3127) );
  AOI22_X1 U24203 ( .A1(n21192), .A2(n21358), .B1(n21360), .B2(n21191), .ZN(
        n21196) );
  AOI22_X1 U24204 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21293), .ZN(n21195) );
  OAI211_X1 U24205 ( .C1(n21298), .C2(n21225), .A(n21196), .B(n21195), .ZN(
        P1_U3128) );
  NAND2_X1 U24206 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21301) );
  AOI22_X1 U24207 ( .A1(n21248), .A2(n21317), .B1(n21310), .B2(n9829), .ZN(
        n21208) );
  NAND2_X1 U24208 ( .A1(n21225), .A2(n9694), .ZN(n21200) );
  OAI21_X1 U24209 ( .B1(n21200), .B2(n21248), .A(n21199), .ZN(n21203) );
  OR2_X1 U24210 ( .A1(n13843), .A2(n21201), .ZN(n21227) );
  OR2_X1 U24211 ( .A1(n21227), .A2(n21256), .ZN(n21205) );
  AOI22_X1 U24212 ( .A1(n21203), .A2(n21205), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21204), .ZN(n21202) );
  INV_X1 U24213 ( .A(n21203), .ZN(n21206) );
  AOI22_X1 U24214 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21222), .B1(
        n21309), .B2(n21221), .ZN(n21207) );
  OAI211_X1 U24215 ( .C1(n21320), .C2(n21225), .A(n21208), .B(n21207), .ZN(
        P1_U3129) );
  AOI22_X1 U24216 ( .A1(n21248), .A2(n21323), .B1(n9829), .B2(n21322), .ZN(
        n21210) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21222), .B1(
        n21321), .B2(n21221), .ZN(n21209) );
  OAI211_X1 U24218 ( .C1(n21326), .C2(n21225), .A(n21210), .B(n21209), .ZN(
        P1_U3130) );
  AOI22_X1 U24219 ( .A1(n21248), .A2(n21329), .B1(n9829), .B2(n21328), .ZN(
        n21212) );
  AOI22_X1 U24220 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21222), .B1(
        n21327), .B2(n21221), .ZN(n21211) );
  OAI211_X1 U24221 ( .C1(n21332), .C2(n21225), .A(n21212), .B(n21211), .ZN(
        P1_U3131) );
  AOI22_X1 U24222 ( .A1(n21248), .A2(n21335), .B1(n9829), .B2(n21334), .ZN(
        n21214) );
  AOI22_X1 U24223 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21222), .B1(
        n21333), .B2(n21221), .ZN(n21213) );
  OAI211_X1 U24224 ( .C1(n21338), .C2(n21225), .A(n21214), .B(n21213), .ZN(
        P1_U3132) );
  AOI22_X1 U24225 ( .A1(n21248), .A2(n21341), .B1(n9829), .B2(n21340), .ZN(
        n21216) );
  AOI22_X1 U24226 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21222), .B1(
        n21339), .B2(n21221), .ZN(n21215) );
  OAI211_X1 U24227 ( .C1(n21344), .C2(n21225), .A(n21216), .B(n21215), .ZN(
        P1_U3133) );
  AOI22_X1 U24228 ( .A1(n21248), .A2(n21347), .B1(n9829), .B2(n21346), .ZN(
        n21218) );
  AOI22_X1 U24229 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21222), .B1(
        n21345), .B2(n21221), .ZN(n21217) );
  OAI211_X1 U24230 ( .C1(n21350), .C2(n21225), .A(n21218), .B(n21217), .ZN(
        P1_U3134) );
  AOI22_X1 U24231 ( .A1(n21248), .A2(n21353), .B1(n9829), .B2(n21352), .ZN(
        n21220) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21222), .B1(
        n21351), .B2(n21221), .ZN(n21219) );
  OAI211_X1 U24233 ( .C1(n21356), .C2(n21225), .A(n21220), .B(n21219), .ZN(
        P1_U3135) );
  AOI22_X1 U24234 ( .A1(n21248), .A2(n21361), .B1(n9829), .B2(n21360), .ZN(
        n21224) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21222), .B1(
        n21358), .B2(n21221), .ZN(n21223) );
  OAI211_X1 U24236 ( .C1(n21367), .C2(n21225), .A(n21224), .B(n21223), .ZN(
        P1_U3136) );
  NOR3_X2 U24237 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21677), .A3(
        n21301), .ZN(n21246) );
  INV_X1 U24238 ( .A(n21246), .ZN(n21229) );
  NOR2_X1 U24239 ( .A1(n21301), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21231) );
  INV_X1 U24240 ( .A(n21231), .ZN(n21228) );
  INV_X1 U24241 ( .A(n21227), .ZN(n21257) );
  NAND2_X1 U24242 ( .A1(n21257), .A2(n9694), .ZN(n21308) );
  OAI222_X1 U24243 ( .A1(n21229), .A2(n21304), .B1(n21306), .B2(n21228), .C1(
        n20826), .C2(n21308), .ZN(n21247) );
  AOI22_X1 U24244 ( .A1(n21309), .A2(n21247), .B1(n21310), .B2(n21246), .ZN(
        n21233) );
  AND2_X1 U24245 ( .A1(n21311), .A2(n21230), .ZN(n21467) );
  AOI22_X1 U24246 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21263), .ZN(n21232) );
  OAI211_X1 U24247 ( .C1(n21266), .C2(n21262), .A(n21233), .B(n21232), .ZN(
        P1_U3137) );
  AOI22_X1 U24248 ( .A1(n21321), .A2(n21247), .B1(n21322), .B2(n21246), .ZN(
        n21235) );
  AOI22_X1 U24249 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21267), .ZN(n21234) );
  OAI211_X1 U24250 ( .C1(n21270), .C2(n21262), .A(n21235), .B(n21234), .ZN(
        P1_U3138) );
  AOI22_X1 U24251 ( .A1(n21327), .A2(n21247), .B1(n21328), .B2(n21246), .ZN(
        n21237) );
  AOI22_X1 U24252 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21271), .ZN(n21236) );
  OAI211_X1 U24253 ( .C1(n21274), .C2(n21262), .A(n21237), .B(n21236), .ZN(
        P1_U3139) );
  AOI22_X1 U24254 ( .A1(n21333), .A2(n21247), .B1(n21334), .B2(n21246), .ZN(
        n21239) );
  AOI22_X1 U24255 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21275), .ZN(n21238) );
  OAI211_X1 U24256 ( .C1(n21278), .C2(n21262), .A(n21239), .B(n21238), .ZN(
        P1_U3140) );
  AOI22_X1 U24257 ( .A1(n21339), .A2(n21247), .B1(n21340), .B2(n21246), .ZN(
        n21241) );
  AOI22_X1 U24258 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21279), .ZN(n21240) );
  OAI211_X1 U24259 ( .C1(n21282), .C2(n21262), .A(n21241), .B(n21240), .ZN(
        P1_U3141) );
  AOI22_X1 U24260 ( .A1(n21345), .A2(n21247), .B1(n21346), .B2(n21246), .ZN(
        n21243) );
  AOI22_X1 U24261 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21283), .ZN(n21242) );
  OAI211_X1 U24262 ( .C1(n21286), .C2(n21262), .A(n21243), .B(n21242), .ZN(
        P1_U3142) );
  AOI22_X1 U24263 ( .A1(n21351), .A2(n21247), .B1(n21352), .B2(n21246), .ZN(
        n21245) );
  AOI22_X1 U24264 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21287), .ZN(n21244) );
  OAI211_X1 U24265 ( .C1(n21290), .C2(n21262), .A(n21245), .B(n21244), .ZN(
        P1_U3143) );
  AOI22_X1 U24266 ( .A1(n21358), .A2(n21247), .B1(n21360), .B2(n21246), .ZN(
        n21251) );
  AOI22_X1 U24267 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21249), .B1(
        n21248), .B2(n21293), .ZN(n21250) );
  OAI211_X1 U24268 ( .C1(n21298), .C2(n21262), .A(n21251), .B(n21250), .ZN(
        P1_U3144) );
  NOR3_X2 U24269 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21302), .A3(
        n21301), .ZN(n21292) );
  OAI22_X1 U24270 ( .A1(n21308), .A2(n13858), .B1(n21254), .B2(n21253), .ZN(
        n21291) );
  AOI22_X1 U24271 ( .A1(n21310), .A2(n21292), .B1(n21309), .B2(n21291), .ZN(
        n21265) );
  AOI21_X1 U24272 ( .B1(n21262), .B2(n21366), .A(n20830), .ZN(n21255) );
  AOI21_X1 U24273 ( .B1(n21257), .B2(n21256), .A(n21255), .ZN(n21258) );
  NOR2_X1 U24274 ( .A1(n21258), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21261) );
  AOI22_X1 U24275 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21263), .ZN(n21264) );
  OAI211_X1 U24276 ( .C1(n21266), .C2(n21366), .A(n21265), .B(n21264), .ZN(
        P1_U3145) );
  AOI22_X1 U24277 ( .A1(n21322), .A2(n21292), .B1(n21321), .B2(n21291), .ZN(
        n21269) );
  AOI22_X1 U24278 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21267), .ZN(n21268) );
  OAI211_X1 U24279 ( .C1(n21270), .C2(n21366), .A(n21269), .B(n21268), .ZN(
        P1_U3146) );
  AOI22_X1 U24280 ( .A1(n21328), .A2(n21292), .B1(n21327), .B2(n21291), .ZN(
        n21273) );
  AOI22_X1 U24281 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21271), .ZN(n21272) );
  OAI211_X1 U24282 ( .C1(n21274), .C2(n21366), .A(n21273), .B(n21272), .ZN(
        P1_U3147) );
  AOI22_X1 U24283 ( .A1(n21334), .A2(n21292), .B1(n21333), .B2(n21291), .ZN(
        n21277) );
  AOI22_X1 U24284 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21275), .ZN(n21276) );
  OAI211_X1 U24285 ( .C1(n21278), .C2(n21366), .A(n21277), .B(n21276), .ZN(
        P1_U3148) );
  AOI22_X1 U24286 ( .A1(n21340), .A2(n21292), .B1(n21339), .B2(n21291), .ZN(
        n21281) );
  AOI22_X1 U24287 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21279), .ZN(n21280) );
  OAI211_X1 U24288 ( .C1(n21282), .C2(n21366), .A(n21281), .B(n21280), .ZN(
        P1_U3149) );
  AOI22_X1 U24289 ( .A1(n21346), .A2(n21292), .B1(n21345), .B2(n21291), .ZN(
        n21285) );
  AOI22_X1 U24290 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21283), .ZN(n21284) );
  OAI211_X1 U24291 ( .C1(n21286), .C2(n21366), .A(n21285), .B(n21284), .ZN(
        P1_U3150) );
  AOI22_X1 U24292 ( .A1(n21352), .A2(n21292), .B1(n21351), .B2(n21291), .ZN(
        n21289) );
  AOI22_X1 U24293 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21287), .ZN(n21288) );
  OAI211_X1 U24294 ( .C1(n21290), .C2(n21366), .A(n21289), .B(n21288), .ZN(
        P1_U3151) );
  AOI22_X1 U24295 ( .A1(n21360), .A2(n21292), .B1(n21358), .B2(n21291), .ZN(
        n21297) );
  AOI22_X1 U24296 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21295), .B1(
        n21294), .B2(n21293), .ZN(n21296) );
  OAI211_X1 U24297 ( .C1(n21298), .C2(n21366), .A(n21297), .B(n21296), .ZN(
        P1_U3152) );
  INV_X1 U24298 ( .A(n21301), .ZN(n21299) );
  NAND2_X1 U24299 ( .A1(n21300), .A2(n21299), .ZN(n21303) );
  INV_X1 U24300 ( .A(n21303), .ZN(n21359) );
  NOR2_X1 U24301 ( .A1(n21302), .A2(n21301), .ZN(n21315) );
  INV_X1 U24302 ( .A(n21315), .ZN(n21305) );
  OAI222_X1 U24303 ( .A1(n21308), .A2(n21307), .B1(n21306), .B2(n21305), .C1(
        n21304), .C2(n21303), .ZN(n21357) );
  AOI22_X1 U24304 ( .A1(n21310), .A2(n21359), .B1(n21309), .B2(n21357), .ZN(
        n21319) );
  INV_X1 U24305 ( .A(n21311), .ZN(n21313) );
  NOR2_X1 U24306 ( .A1(n21313), .A2(n21312), .ZN(n21316) );
  AOI22_X1 U24307 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21317), .ZN(n21318) );
  OAI211_X1 U24308 ( .C1(n21320), .C2(n21366), .A(n21319), .B(n21318), .ZN(
        P1_U3153) );
  AOI22_X1 U24309 ( .A1(n21322), .A2(n21359), .B1(n21321), .B2(n21357), .ZN(
        n21325) );
  AOI22_X1 U24310 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21323), .ZN(n21324) );
  OAI211_X1 U24311 ( .C1(n21326), .C2(n21366), .A(n21325), .B(n21324), .ZN(
        P1_U3154) );
  AOI22_X1 U24312 ( .A1(n21328), .A2(n21359), .B1(n21327), .B2(n21357), .ZN(
        n21331) );
  AOI22_X1 U24313 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21329), .ZN(n21330) );
  OAI211_X1 U24314 ( .C1(n21332), .C2(n21366), .A(n21331), .B(n21330), .ZN(
        P1_U3155) );
  AOI22_X1 U24315 ( .A1(n21334), .A2(n21359), .B1(n21333), .B2(n21357), .ZN(
        n21337) );
  AOI22_X1 U24316 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21335), .ZN(n21336) );
  OAI211_X1 U24317 ( .C1(n21338), .C2(n21366), .A(n21337), .B(n21336), .ZN(
        P1_U3156) );
  AOI22_X1 U24318 ( .A1(n21340), .A2(n21359), .B1(n21339), .B2(n21357), .ZN(
        n21343) );
  AOI22_X1 U24319 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21341), .ZN(n21342) );
  OAI211_X1 U24320 ( .C1(n21344), .C2(n21366), .A(n21343), .B(n21342), .ZN(
        P1_U3157) );
  AOI22_X1 U24321 ( .A1(n21346), .A2(n21359), .B1(n21345), .B2(n21357), .ZN(
        n21349) );
  AOI22_X1 U24322 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21347), .ZN(n21348) );
  OAI211_X1 U24323 ( .C1(n21350), .C2(n21366), .A(n21349), .B(n21348), .ZN(
        P1_U3158) );
  AOI22_X1 U24324 ( .A1(n21352), .A2(n21359), .B1(n21351), .B2(n21357), .ZN(
        n21355) );
  AOI22_X1 U24325 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21353), .ZN(n21354) );
  OAI211_X1 U24326 ( .C1(n21356), .C2(n21366), .A(n21355), .B(n21354), .ZN(
        P1_U3159) );
  AOI22_X1 U24327 ( .A1(n21360), .A2(n21359), .B1(n21358), .B2(n21357), .ZN(
        n21365) );
  AOI22_X1 U24328 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21363), .B1(
        n21362), .B2(n21361), .ZN(n21364) );
  OAI211_X1 U24329 ( .C1(n21367), .C2(n21366), .A(n21365), .B(n21364), .ZN(
        P1_U3160) );
  AOI21_X1 U24330 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21369), .A(n21368), 
        .ZN(n21371) );
  NAND2_X1 U24331 ( .A1(n21371), .A2(n21370), .ZN(P1_U3163) );
  AND2_X1 U24332 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21448), .ZN(
        P1_U3164) );
  AND2_X1 U24333 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21448), .ZN(
        P1_U3165) );
  AND2_X1 U24334 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21448), .ZN(
        P1_U3166) );
  AND2_X1 U24335 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21448), .ZN(
        P1_U3167) );
  AND2_X1 U24336 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21448), .ZN(
        P1_U3168) );
  AND2_X1 U24337 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21448), .ZN(
        P1_U3169) );
  AND2_X1 U24338 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21448), .ZN(
        P1_U3170) );
  AND2_X1 U24339 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21448), .ZN(
        P1_U3171) );
  AND2_X1 U24340 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21448), .ZN(
        P1_U3172) );
  AND2_X1 U24341 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21448), .ZN(
        P1_U3173) );
  AND2_X1 U24342 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21448), .ZN(
        P1_U3174) );
  AND2_X1 U24343 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21448), .ZN(
        P1_U3175) );
  AND2_X1 U24344 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21448), .ZN(
        P1_U3176) );
  AND2_X1 U24345 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21448), .ZN(
        P1_U3177) );
  AND2_X1 U24346 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21448), .ZN(
        P1_U3178) );
  AND2_X1 U24347 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21448), .ZN(
        P1_U3179) );
  AND2_X1 U24348 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21448), .ZN(
        P1_U3180) );
  AND2_X1 U24349 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21448), .ZN(
        P1_U3181) );
  AND2_X1 U24350 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21448), .ZN(
        P1_U3182) );
  AND2_X1 U24351 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21448), .ZN(
        P1_U3183) );
  INV_X1 U24352 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21753) );
  NOR2_X1 U24353 ( .A1(n21452), .A2(n21753), .ZN(P1_U3184) );
  AND2_X1 U24354 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21448), .ZN(
        P1_U3185) );
  INV_X1 U24355 ( .A(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21613) );
  NOR2_X1 U24356 ( .A1(n21452), .A2(n21613), .ZN(P1_U3186) );
  AND2_X1 U24357 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21448), .ZN(P1_U3187) );
  AND2_X1 U24358 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21448), .ZN(P1_U3188) );
  AND2_X1 U24359 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21448), .ZN(P1_U3189) );
  AND2_X1 U24360 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21448), .ZN(P1_U3190) );
  AND2_X1 U24361 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21448), .ZN(P1_U3191) );
  AND2_X1 U24362 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21448), .ZN(P1_U3192) );
  INV_X1 U24363 ( .A(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21774) );
  NOR2_X1 U24364 ( .A1(n21452), .A2(n21774), .ZN(P1_U3193) );
  AOI21_X1 U24365 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21378), .A(n21380), 
        .ZN(n21387) );
  OAI22_X1 U24366 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21377), .B1(n21388), 
        .B2(n21372), .ZN(n21373) );
  NOR3_X1 U24367 ( .A1(n21374), .A2(n21383), .A3(n21373), .ZN(n21375) );
  OAI22_X1 U24368 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21387), .B1(n21439), 
        .B2(n21375), .ZN(P1_U3194) );
  OAI21_X1 U24369 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21376), .A(n21377), 
        .ZN(n21386) );
  NAND2_X1 U24370 ( .A1(n21378), .A2(n21377), .ZN(n21381) );
  OAI21_X1 U24371 ( .B1(n21381), .B2(n21380), .A(n21379), .ZN(n21382) );
  OAI211_X1 U24372 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21383), .A(HOLD), .B(
        n21382), .ZN(n21384) );
  OAI221_X1 U24373 ( .B1(n21387), .B2(n21386), .C1(n21387), .C2(n21385), .A(
        n21384), .ZN(P1_U3196) );
  INV_X1 U24374 ( .A(n21436), .ZN(n21420) );
  INV_X1 U24375 ( .A(n21420), .ZN(n21437) );
  INV_X1 U24376 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21389) );
  INV_X2 U24377 ( .A(n21423), .ZN(n21442) );
  OAI222_X1 U24378 ( .A1(n21437), .A2(n20627), .B1(n21389), .B2(n21439), .C1(
        n21476), .C2(n21442), .ZN(P1_U3197) );
  INV_X1 U24379 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21390) );
  OAI222_X1 U24380 ( .A1(n21442), .A2(n20627), .B1(n21390), .B2(n21439), .C1(
        n21392), .C2(n21436), .ZN(P1_U3198) );
  INV_X1 U24381 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21391) );
  OAI222_X1 U24382 ( .A1(n21442), .A2(n21392), .B1(n21391), .B2(n21439), .C1(
        n21393), .C2(n21437), .ZN(P1_U3199) );
  INV_X1 U24383 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21394) );
  OAI222_X1 U24384 ( .A1(n21437), .A2(n21396), .B1(n21394), .B2(n21439), .C1(
        n21393), .C2(n21442), .ZN(P1_U3200) );
  INV_X1 U24385 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21395) );
  OAI222_X1 U24386 ( .A1(n21442), .A2(n21396), .B1(n21395), .B2(n21439), .C1(
        n21680), .C2(n21436), .ZN(P1_U3201) );
  INV_X1 U24387 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21397) );
  OAI222_X1 U24388 ( .A1(n21442), .A2(n21680), .B1(n21397), .B2(n21439), .C1(
        n21398), .C2(n21436), .ZN(P1_U3202) );
  INV_X1 U24389 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21562) );
  OAI222_X1 U24390 ( .A1(n21442), .A2(n21398), .B1(n21562), .B2(n21439), .C1(
        n21399), .C2(n21436), .ZN(P1_U3203) );
  INV_X1 U24391 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21400) );
  OAI222_X1 U24392 ( .A1(n21436), .A2(n21402), .B1(n21400), .B2(n21439), .C1(
        n21399), .C2(n21442), .ZN(P1_U3204) );
  INV_X1 U24393 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21401) );
  OAI222_X1 U24394 ( .A1(n21442), .A2(n21402), .B1(n21401), .B2(n21439), .C1(
        n21403), .C2(n21436), .ZN(P1_U3205) );
  INV_X1 U24395 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21404) );
  OAI222_X1 U24396 ( .A1(n21436), .A2(n21406), .B1(n21404), .B2(n21439), .C1(
        n21403), .C2(n21442), .ZN(P1_U3206) );
  INV_X1 U24397 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21405) );
  OAI222_X1 U24398 ( .A1(n21442), .A2(n21406), .B1(n21405), .B2(n21439), .C1(
        n21407), .C2(n21436), .ZN(P1_U3207) );
  INV_X1 U24399 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21775) );
  OAI222_X1 U24400 ( .A1(n21442), .A2(n21407), .B1(n21775), .B2(n21439), .C1(
        n21408), .C2(n21436), .ZN(P1_U3208) );
  INV_X1 U24401 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21657) );
  OAI222_X1 U24402 ( .A1(n21442), .A2(n21408), .B1(n21657), .B2(n21439), .C1(
        n21409), .C2(n21437), .ZN(P1_U3209) );
  INV_X1 U24403 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21410) );
  OAI222_X1 U24404 ( .A1(n21436), .A2(n21766), .B1(n21410), .B2(n21439), .C1(
        n21409), .C2(n21442), .ZN(P1_U3210) );
  INV_X1 U24405 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21411) );
  OAI222_X1 U24406 ( .A1(n21436), .A2(n21413), .B1(n21411), .B2(n21439), .C1(
        n21766), .C2(n21442), .ZN(P1_U3211) );
  INV_X1 U24407 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21412) );
  OAI222_X1 U24408 ( .A1(n21442), .A2(n21413), .B1(n21412), .B2(n21439), .C1(
        n21415), .C2(n21437), .ZN(P1_U3212) );
  INV_X1 U24409 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21414) );
  OAI222_X1 U24410 ( .A1(n21442), .A2(n21415), .B1(n21414), .B2(n21439), .C1(
        n21417), .C2(n21436), .ZN(P1_U3213) );
  AOI22_X1 U24411 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21494), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21420), .ZN(n21416) );
  OAI21_X1 U24412 ( .B1(n21417), .B2(n21442), .A(n21416), .ZN(P1_U3214) );
  AOI22_X1 U24413 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21494), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21423), .ZN(n21418) );
  OAI21_X1 U24414 ( .B1(n21419), .B2(n21437), .A(n21418), .ZN(P1_U3215) );
  INV_X1 U24415 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21749) );
  OAI222_X1 U24416 ( .A1(n21442), .A2(n21419), .B1(n21749), .B2(n21439), .C1(
        n15559), .C2(n21437), .ZN(P1_U3216) );
  INV_X1 U24417 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21682) );
  OAI222_X1 U24418 ( .A1(n21442), .A2(n15559), .B1(n21682), .B2(n21439), .C1(
        n21422), .C2(n21437), .ZN(P1_U3217) );
  AOI22_X1 U24419 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21494), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21420), .ZN(n21421) );
  OAI21_X1 U24420 ( .B1(n21422), .B2(n21442), .A(n21421), .ZN(P1_U3218) );
  AOI22_X1 U24421 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21494), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21423), .ZN(n21424) );
  OAI21_X1 U24422 ( .B1(n21426), .B2(n21437), .A(n21424), .ZN(P1_U3219) );
  INV_X1 U24423 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21425) );
  OAI222_X1 U24424 ( .A1(n21442), .A2(n21426), .B1(n21425), .B2(n21439), .C1(
        n15125), .C2(n21437), .ZN(P1_U3220) );
  INV_X1 U24425 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21427) );
  OAI222_X1 U24426 ( .A1(n21442), .A2(n15125), .B1(n21427), .B2(n21439), .C1(
        n21429), .C2(n21437), .ZN(P1_U3221) );
  INV_X1 U24427 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21428) );
  OAI222_X1 U24428 ( .A1(n21442), .A2(n21429), .B1(n21428), .B2(n21439), .C1(
        n21431), .C2(n21437), .ZN(P1_U3222) );
  INV_X1 U24429 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21430) );
  OAI222_X1 U24430 ( .A1(n21442), .A2(n21431), .B1(n21430), .B2(n21439), .C1(
        n21433), .C2(n21437), .ZN(P1_U3223) );
  INV_X1 U24431 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21432) );
  OAI222_X1 U24432 ( .A1(n21442), .A2(n21433), .B1(n21432), .B2(n21439), .C1(
        n21434), .C2(n21437), .ZN(P1_U3224) );
  INV_X1 U24433 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21441) );
  INV_X1 U24434 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21435) );
  OAI222_X1 U24435 ( .A1(n21436), .A2(n21441), .B1(n21435), .B2(n21439), .C1(
        n21434), .C2(n21442), .ZN(P1_U3225) );
  INV_X1 U24436 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21440) );
  OAI222_X1 U24437 ( .A1(n21442), .A2(n21441), .B1(n21440), .B2(n21439), .C1(
        n21438), .C2(n21437), .ZN(P1_U3226) );
  INV_X1 U24438 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21443) );
  AOI22_X1 U24439 ( .A1(n21439), .A2(n21444), .B1(n21443), .B2(n21494), .ZN(
        P1_U3458) );
  INV_X1 U24440 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21479) );
  AOI22_X1 U24441 ( .A1(n21439), .A2(n21479), .B1(n21549), .B2(n21494), .ZN(
        P1_U3459) );
  AOI22_X1 U24442 ( .A1(n21439), .A2(n21446), .B1(n21445), .B2(n21494), .ZN(
        P1_U3460) );
  INV_X1 U24443 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21482) );
  AOI22_X1 U24444 ( .A1(n21439), .A2(n21482), .B1(n21789), .B2(n21494), .ZN(
        P1_U3461) );
  INV_X1 U24445 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21449) );
  INV_X1 U24446 ( .A(n21450), .ZN(n21447) );
  AOI21_X1 U24447 ( .B1(n21449), .B2(n21448), .A(n21447), .ZN(P1_U3464) );
  OAI21_X1 U24448 ( .B1(n21452), .B2(n21451), .A(n21450), .ZN(P1_U3465) );
  INV_X1 U24449 ( .A(n21453), .ZN(n21455) );
  OAI21_X1 U24450 ( .B1(n21455), .B2(n21454), .A(n21457), .ZN(n21456) );
  OAI21_X1 U24451 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21457), .A(
        n21456), .ZN(n21458) );
  OAI21_X1 U24452 ( .B1(n21460), .B2(n21459), .A(n21458), .ZN(P1_U3469) );
  OAI211_X1 U24453 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21463), .A(n21462), 
        .B(n21461), .ZN(n21469) );
  INV_X1 U24454 ( .A(n21464), .ZN(n21466) );
  NOR2_X1 U24455 ( .A1(n21466), .A2(n21465), .ZN(n21468) );
  AOI211_X1 U24456 ( .C1(n9694), .C2(n21469), .A(n21468), .B(n21467), .ZN(
        n21471) );
  OR2_X1 U24457 ( .A1(n21472), .A2(n21471), .ZN(n21473) );
  OAI21_X1 U24458 ( .B1(n21475), .B2(n21474), .A(n21473), .ZN(P1_U3475) );
  AOI21_X1 U24459 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21477) );
  AOI22_X1 U24460 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21477), .B2(n21476), .ZN(n21480) );
  AOI22_X1 U24461 ( .A1(n21483), .A2(n21480), .B1(n21479), .B2(n21478), .ZN(
        P1_U3481) );
  OAI21_X1 U24462 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21483), .ZN(n21481) );
  OAI21_X1 U24463 ( .B1(n21483), .B2(n21482), .A(n21481), .ZN(P1_U3482) );
  INV_X1 U24464 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21484) );
  AOI22_X1 U24465 ( .A1(n21439), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21484), 
        .B2(n21494), .ZN(P1_U3483) );
  AOI211_X1 U24466 ( .C1(n20662), .C2(n21487), .A(n21486), .B(n21485), .ZN(
        n21493) );
  OAI211_X1 U24467 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11957), .A(n21488), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21490) );
  AOI21_X1 U24468 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21490), .A(n21489), 
        .ZN(n21492) );
  NAND2_X1 U24469 ( .A1(n21493), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21491) );
  OAI21_X1 U24470 ( .B1(n21493), .B2(n21492), .A(n21491), .ZN(P1_U3485) );
  OAI22_X1 U24471 ( .A1(n21494), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n21439), .ZN(n21495) );
  INV_X1 U24472 ( .A(n21495), .ZN(P1_U3486) );
  AOI21_X1 U24473 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21497), .A(n21496), 
        .ZN(n21498) );
  OAI21_X1 U24474 ( .B1(n14041), .B2(n21499), .A(n21498), .ZN(n21806) );
  NOR4_X1 U24475 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(
        BUF1_REG_8__SCAN_IN), .A3(P3_ADDRESS_REG_26__SCAN_IN), .A4(n21704), 
        .ZN(n21500) );
  NAND3_X1 U24476 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_DATAO_REG_5__SCAN_IN), 
        .A3(n21500), .ZN(n21510) );
  INV_X1 U24477 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21571) );
  NAND4_X1 U24478 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(P3_DATAO_REG_9__SCAN_IN), 
        .A3(P1_ADS_N_REG_SCAN_IN), .A4(n21571), .ZN(n21501) );
  NOR3_X1 U24479 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n21564), .A3(n21501), 
        .ZN(n21508) );
  INV_X1 U24480 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21550) );
  NAND4_X1 U24481 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(n21550), .A3(n10871), 
        .A4(n14248), .ZN(n21506) );
  NAND4_X1 U24482 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .A3(n21586), .A4(n21587), .ZN(n21505) );
  NAND4_X1 U24483 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A4(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n21504) );
  NAND4_X1 U24484 ( .A1(n21502), .A2(n15125), .A3(P1_EBX_REG_14__SCAN_IN), 
        .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n21503) );
  NOR4_X1 U24485 ( .A1(n21506), .A2(n21505), .A3(n21504), .A4(n21503), .ZN(
        n21507) );
  NAND4_X1 U24486 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        BUF2_REG_27__SCAN_IN), .A3(n21508), .A4(n21507), .ZN(n21509) );
  NOR4_X1 U24487 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n21510), .A4(n21509), .ZN(
        n21545) );
  NAND4_X1 U24488 ( .A1(n21512), .A2(n21511), .A3(P3_EBX_REG_12__SCAN_IN), 
        .A4(P3_EBX_REG_11__SCAN_IN), .ZN(n21543) );
  INV_X1 U24489 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n21513) );
  NAND4_X1 U24490 ( .A1(n21513), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_13__1__SCAN_IN), .A4(n21787), .ZN(n21514) );
  NOR3_X1 U24491 ( .A1(n21514), .A2(P2_DATAWIDTH_REG_14__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21520) );
  NAND4_X1 U24492 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_DATAO_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        n21657), .ZN(n21518) );
  INV_X1 U24493 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21553) );
  NAND4_X1 U24494 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_5__2__SCAN_IN), .A3(P1_INSTQUEUE_REG_13__7__SCAN_IN), 
        .A4(n21553), .ZN(n21517) );
  NAND4_X1 U24495 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(
        P1_DATAO_REG_18__SCAN_IN), .A3(n21736), .A4(n16206), .ZN(n21516) );
  NAND4_X1 U24496 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(n21751), .A4(n21760), .ZN(n21515) );
  NOR4_X1 U24497 ( .A1(n21518), .A2(n21517), .A3(n21516), .A4(n21515), .ZN(
        n21519) );
  NAND4_X1 U24498 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_1__0__SCAN_IN), .A3(n21520), .A4(n21519), .ZN(n21542)
         );
  NAND4_X1 U24499 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_DATAO_REG_29__SCAN_IN), .A3(n21680), .A4(n21676), .ZN(n21524) );
  NAND4_X1 U24500 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_15__5__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), 
        .A4(n21692), .ZN(n21523) );
  NAND4_X1 U24501 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(BUF1_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(n21717), .ZN(n21522) );
  NAND4_X1 U24502 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .A3(P2_EBX_REG_24__SCAN_IN), .A4(P3_REIP_REG_30__SCAN_IN), .ZN(n21521)
         );
  NOR4_X1 U24503 ( .A1(n21524), .A2(n21523), .A3(n21522), .A4(n21521), .ZN(
        n21540) );
  NAND4_X1 U24504 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P2_EAX_REG_7__SCAN_IN), 
        .A3(P3_BYTEENABLE_REG_0__SCAN_IN), .A4(n21774), .ZN(n21528) );
  INV_X1 U24505 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21781) );
  NAND4_X1 U24506 ( .A1(n21740), .A2(n21781), .A3(n21780), .A4(n21741), .ZN(
        n21527) );
  NAND4_X1 U24507 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(
        P1_REIP_REG_15__SCAN_IN), .A3(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), 
        .A4(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21526) );
  NAND4_X1 U24508 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(
        P2_BE_N_REG_2__SCAN_IN), .A3(P3_UWORD_REG_11__SCAN_IN), .A4(n14256), 
        .ZN(n21525) );
  NOR4_X1 U24509 ( .A1(n21528), .A2(n21527), .A3(n21526), .A4(n21525), .ZN(
        n21539) );
  NAND4_X1 U24510 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_MORE_REG_SCAN_IN), .A3(n21646), .A4(n21641), .ZN(n21532) );
  NAND4_X1 U24511 ( .A1(DATAI_25_), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A3(
        n10545), .A4(n21627), .ZN(n21531) );
  NAND4_X1 U24512 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(BUF1_REG_24__SCAN_IN), 
        .A3(BUF1_REG_1__SCAN_IN), .A4(n21659), .ZN(n21530) );
  NAND4_X1 U24513 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        P2_STATE_REG_2__SCAN_IN), .A3(BUF2_REG_6__SCAN_IN), .A4(n21643), .ZN(
        n21529) );
  NOR4_X1 U24514 ( .A1(n21532), .A2(n21531), .A3(n21530), .A4(n21529), .ZN(
        n21538) );
  NAND4_X1 U24515 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(P1_EAX_REG_6__SCAN_IN), 
        .A3(BUF1_REG_18__SCAN_IN), .A4(n21613), .ZN(n21536) );
  NAND4_X1 U24516 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .A3(P3_REIP_REG_5__SCAN_IN), .A4(
        n21598), .ZN(n21535) );
  INV_X1 U24517 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21617) );
  NAND4_X1 U24518 ( .A1(BUF2_REG_30__SCAN_IN), .A2(READY22_REG_SCAN_IN), .A3(
        P3_LWORD_REG_14__SCAN_IN), .A4(n21617), .ZN(n21534) );
  NAND4_X1 U24519 ( .A1(n21611), .A2(n12123), .A3(n21610), .A4(n21616), .ZN(
        n21533) );
  NOR4_X1 U24520 ( .A1(n21536), .A2(n21535), .A3(n21534), .A4(n21533), .ZN(
        n21537) );
  NAND4_X1 U24521 ( .A1(n21540), .A2(n21539), .A3(n21538), .A4(n21537), .ZN(
        n21541) );
  NOR4_X1 U24522 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21543), .A3(n21542), 
        .A4(n21541), .ZN(n21544) );
  AOI21_X1 U24523 ( .B1(n21545), .B2(n21544), .A(P1_ADDRESS_REG_19__SCAN_IN), 
        .ZN(n21804) );
  INV_X1 U24524 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21547) );
  AOI22_X1 U24525 ( .A1(n21547), .A2(keyinput35), .B1(keyinput17), .B2(n15125), 
        .ZN(n21546) );
  OAI221_X1 U24526 ( .B1(n21547), .B2(keyinput35), .C1(n15125), .C2(keyinput17), .A(n21546), .ZN(n21559) );
  AOI22_X1 U24527 ( .A1(n21550), .A2(keyinput95), .B1(keyinput81), .B2(n21549), 
        .ZN(n21548) );
  OAI221_X1 U24528 ( .B1(n21550), .B2(keyinput95), .C1(n21549), .C2(keyinput81), .A(n21548), .ZN(n21558) );
  AOI22_X1 U24529 ( .A1(n21553), .A2(keyinput27), .B1(keyinput75), .B2(n21552), 
        .ZN(n21551) );
  OAI221_X1 U24530 ( .B1(n21553), .B2(keyinput27), .C1(n21552), .C2(keyinput75), .A(n21551), .ZN(n21557) );
  XNOR2_X1 U24531 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput87), .ZN(
        n21555) );
  XNOR2_X1 U24532 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput96), .ZN(n21554) );
  NAND2_X1 U24533 ( .A1(n21555), .A2(n21554), .ZN(n21556) );
  NOR4_X1 U24534 ( .A1(n21559), .A2(n21558), .A3(n21557), .A4(n21556), .ZN(
        n21608) );
  AOI22_X1 U24535 ( .A1(n21562), .A2(keyinput42), .B1(keyinput47), .B2(n21561), 
        .ZN(n21560) );
  OAI221_X1 U24536 ( .B1(n21562), .B2(keyinput42), .C1(n21561), .C2(keyinput47), .A(n21560), .ZN(n21575) );
  AOI22_X1 U24537 ( .A1(n21565), .A2(keyinput117), .B1(n21564), .B2(keyinput49), .ZN(n21563) );
  OAI221_X1 U24538 ( .B1(n21565), .B2(keyinput117), .C1(n21564), .C2(
        keyinput49), .A(n21563), .ZN(n21574) );
  AOI22_X1 U24539 ( .A1(n21568), .A2(keyinput26), .B1(keyinput3), .B2(n21567), 
        .ZN(n21566) );
  OAI221_X1 U24540 ( .B1(n21568), .B2(keyinput26), .C1(n21567), .C2(keyinput3), 
        .A(n21566), .ZN(n21573) );
  AOI22_X1 U24541 ( .A1(n21571), .A2(keyinput33), .B1(n21570), .B2(keyinput8), 
        .ZN(n21569) );
  OAI221_X1 U24542 ( .B1(n21571), .B2(keyinput33), .C1(n21570), .C2(keyinput8), 
        .A(n21569), .ZN(n21572) );
  NOR4_X1 U24543 ( .A1(n21575), .A2(n21574), .A3(n21573), .A4(n21572), .ZN(
        n21607) );
  AOI22_X1 U24544 ( .A1(n21578), .A2(keyinput102), .B1(keyinput46), .B2(n21577), .ZN(n21576) );
  OAI221_X1 U24545 ( .B1(n21578), .B2(keyinput102), .C1(n21577), .C2(
        keyinput46), .A(n21576), .ZN(n21591) );
  AOI22_X1 U24546 ( .A1(n21581), .A2(keyinput103), .B1(n21580), .B2(
        keyinput113), .ZN(n21579) );
  OAI221_X1 U24547 ( .B1(n21581), .B2(keyinput103), .C1(n21580), .C2(
        keyinput113), .A(n21579), .ZN(n21590) );
  AOI22_X1 U24548 ( .A1(n21584), .A2(keyinput63), .B1(n21583), .B2(keyinput34), 
        .ZN(n21582) );
  OAI221_X1 U24549 ( .B1(n21584), .B2(keyinput63), .C1(n21583), .C2(keyinput34), .A(n21582), .ZN(n21589) );
  AOI22_X1 U24550 ( .A1(n21587), .A2(keyinput98), .B1(keyinput36), .B2(n21586), 
        .ZN(n21585) );
  OAI221_X1 U24551 ( .B1(n21587), .B2(keyinput98), .C1(n21586), .C2(keyinput36), .A(n21585), .ZN(n21588) );
  NOR4_X1 U24552 ( .A1(n21591), .A2(n21590), .A3(n21589), .A4(n21588), .ZN(
        n21606) );
  AOI22_X1 U24553 ( .A1(n21594), .A2(keyinput92), .B1(n21593), .B2(keyinput31), 
        .ZN(n21592) );
  OAI221_X1 U24554 ( .B1(n21594), .B2(keyinput92), .C1(n21593), .C2(keyinput31), .A(n21592), .ZN(n21604) );
  AOI22_X1 U24555 ( .A1(n13937), .A2(keyinput105), .B1(n10469), .B2(
        keyinput107), .ZN(n21595) );
  OAI221_X1 U24556 ( .B1(n13937), .B2(keyinput105), .C1(n10469), .C2(
        keyinput107), .A(n21595), .ZN(n21603) );
  AOI22_X1 U24557 ( .A1(n21598), .A2(keyinput70), .B1(keyinput97), .B2(n21597), 
        .ZN(n21596) );
  OAI221_X1 U24558 ( .B1(n21598), .B2(keyinput70), .C1(n21597), .C2(keyinput97), .A(n21596), .ZN(n21602) );
  AOI22_X1 U24559 ( .A1(n15488), .A2(keyinput2), .B1(n21600), .B2(keyinput39), 
        .ZN(n21599) );
  OAI221_X1 U24560 ( .B1(n15488), .B2(keyinput2), .C1(n21600), .C2(keyinput39), 
        .A(n21599), .ZN(n21601) );
  NOR4_X1 U24561 ( .A1(n21604), .A2(n21603), .A3(n21602), .A4(n21601), .ZN(
        n21605) );
  NAND4_X1 U24562 ( .A1(n21608), .A2(n21607), .A3(n21606), .A4(n21605), .ZN(
        n21802) );
  AOI22_X1 U24563 ( .A1(n21611), .A2(keyinput52), .B1(keyinput28), .B2(n21610), 
        .ZN(n21609) );
  OAI221_X1 U24564 ( .B1(n21611), .B2(keyinput52), .C1(n21610), .C2(keyinput28), .A(n21609), .ZN(n21623) );
  INV_X1 U24565 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21614) );
  AOI22_X1 U24566 ( .A1(n21614), .A2(keyinput118), .B1(keyinput54), .B2(n21613), .ZN(n21612) );
  OAI221_X1 U24567 ( .B1(n21614), .B2(keyinput118), .C1(n21613), .C2(
        keyinput54), .A(n21612), .ZN(n21622) );
  AOI22_X1 U24568 ( .A1(n21616), .A2(keyinput24), .B1(n12123), .B2(keyinput91), 
        .ZN(n21615) );
  OAI221_X1 U24569 ( .B1(n21616), .B2(keyinput24), .C1(n12123), .C2(keyinput91), .A(n21615), .ZN(n21621) );
  XOR2_X1 U24570 ( .A(n21617), .B(keyinput11), .Z(n21619) );
  XNOR2_X1 U24571 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B(keyinput38), .ZN(
        n21618) );
  NAND2_X1 U24572 ( .A1(n21619), .A2(n21618), .ZN(n21620) );
  NOR4_X1 U24573 ( .A1(n21623), .A2(n21622), .A3(n21621), .A4(n21620), .ZN(
        n21674) );
  AOI22_X1 U24574 ( .A1(n21625), .A2(keyinput61), .B1(n10545), .B2(keyinput44), 
        .ZN(n21624) );
  OAI221_X1 U24575 ( .B1(n21625), .B2(keyinput61), .C1(n10545), .C2(keyinput44), .A(n21624), .ZN(n21638) );
  INV_X1 U24576 ( .A(DATAI_25_), .ZN(n21628) );
  AOI22_X1 U24577 ( .A1(n21628), .A2(keyinput10), .B1(keyinput60), .B2(n21627), 
        .ZN(n21626) );
  OAI221_X1 U24578 ( .B1(n21628), .B2(keyinput10), .C1(n21627), .C2(keyinput60), .A(n21626), .ZN(n21637) );
  INV_X1 U24579 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n21631) );
  AOI22_X1 U24580 ( .A1(n21631), .A2(keyinput79), .B1(n21630), .B2(keyinput59), 
        .ZN(n21629) );
  OAI221_X1 U24581 ( .B1(n21631), .B2(keyinput79), .C1(n21630), .C2(keyinput59), .A(n21629), .ZN(n21636) );
  INV_X1 U24582 ( .A(READY22_REG_SCAN_IN), .ZN(n21632) );
  XOR2_X1 U24583 ( .A(keyinput18), .B(n21632), .Z(n21634) );
  XNOR2_X1 U24584 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B(keyinput67), .ZN(
        n21633) );
  NAND2_X1 U24585 ( .A1(n21634), .A2(n21633), .ZN(n21635) );
  NOR4_X1 U24586 ( .A1(n21638), .A2(n21637), .A3(n21636), .A4(n21635), .ZN(
        n21673) );
  AOI22_X1 U24587 ( .A1(n21641), .A2(keyinput125), .B1(n21640), .B2(keyinput71), .ZN(n21639) );
  OAI221_X1 U24588 ( .B1(n21641), .B2(keyinput125), .C1(n21640), .C2(
        keyinput71), .A(n21639), .ZN(n21654) );
  AOI22_X1 U24589 ( .A1(n21644), .A2(keyinput127), .B1(keyinput78), .B2(n21643), .ZN(n21642) );
  OAI221_X1 U24590 ( .B1(n21644), .B2(keyinput127), .C1(n21643), .C2(
        keyinput78), .A(n21642), .ZN(n21653) );
  AOI22_X1 U24591 ( .A1(n21647), .A2(keyinput45), .B1(n21646), .B2(keyinput9), 
        .ZN(n21645) );
  OAI221_X1 U24592 ( .B1(n21647), .B2(keyinput45), .C1(n21646), .C2(keyinput9), 
        .A(n21645), .ZN(n21652) );
  XOR2_X1 U24593 ( .A(n21648), .B(keyinput66), .Z(n21650) );
  XNOR2_X1 U24594 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B(keyinput65), .ZN(
        n21649) );
  NAND2_X1 U24595 ( .A1(n21650), .A2(n21649), .ZN(n21651) );
  NOR4_X1 U24596 ( .A1(n21654), .A2(n21653), .A3(n21652), .A4(n21651), .ZN(
        n21672) );
  AOI22_X1 U24597 ( .A1(n21657), .A2(keyinput68), .B1(keyinput55), .B2(n21656), 
        .ZN(n21655) );
  OAI221_X1 U24598 ( .B1(n21657), .B2(keyinput68), .C1(n21656), .C2(keyinput55), .A(n21655), .ZN(n21670) );
  AOI22_X1 U24599 ( .A1(n21660), .A2(keyinput109), .B1(keyinput77), .B2(n21659), .ZN(n21658) );
  OAI221_X1 U24600 ( .B1(n21660), .B2(keyinput109), .C1(n21659), .C2(
        keyinput77), .A(n21658), .ZN(n21669) );
  AOI22_X1 U24601 ( .A1(n21663), .A2(keyinput29), .B1(keyinput86), .B2(n21662), 
        .ZN(n21661) );
  OAI221_X1 U24602 ( .B1(n21663), .B2(keyinput29), .C1(n21662), .C2(keyinput86), .A(n21661), .ZN(n21668) );
  AOI22_X1 U24603 ( .A1(n21666), .A2(keyinput101), .B1(keyinput88), .B2(n21665), .ZN(n21664) );
  OAI221_X1 U24604 ( .B1(n21666), .B2(keyinput101), .C1(n21665), .C2(
        keyinput88), .A(n21664), .ZN(n21667) );
  NOR4_X1 U24605 ( .A1(n21670), .A2(n21669), .A3(n21668), .A4(n21667), .ZN(
        n21671) );
  NAND4_X1 U24606 ( .A1(n21674), .A2(n21673), .A3(n21672), .A4(n21671), .ZN(
        n21801) );
  AOI22_X1 U24607 ( .A1(n21677), .A2(keyinput51), .B1(keyinput25), .B2(n21676), 
        .ZN(n21675) );
  OAI221_X1 U24608 ( .B1(n21677), .B2(keyinput51), .C1(n21676), .C2(keyinput25), .A(n21675), .ZN(n21689) );
  AOI22_X1 U24609 ( .A1(n21680), .A2(keyinput115), .B1(n21679), .B2(keyinput56), .ZN(n21678) );
  OAI221_X1 U24610 ( .B1(n21680), .B2(keyinput115), .C1(n21679), .C2(
        keyinput56), .A(n21678), .ZN(n21688) );
  INV_X1 U24611 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n21683) );
  AOI22_X1 U24612 ( .A1(n21683), .A2(keyinput0), .B1(keyinput4), .B2(n21682), 
        .ZN(n21681) );
  OAI221_X1 U24613 ( .B1(n21683), .B2(keyinput0), .C1(n21682), .C2(keyinput4), 
        .A(n21681), .ZN(n21687) );
  INV_X1 U24614 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n21685) );
  AOI22_X1 U24615 ( .A1(n21685), .A2(keyinput93), .B1(keyinput15), .B2(n15979), 
        .ZN(n21684) );
  OAI221_X1 U24616 ( .B1(n21685), .B2(keyinput93), .C1(n15979), .C2(keyinput15), .A(n21684), .ZN(n21686) );
  NOR4_X1 U24617 ( .A1(n21689), .A2(n21688), .A3(n21687), .A4(n21686), .ZN(
        n21734) );
  AOI22_X1 U24618 ( .A1(n21692), .A2(keyinput89), .B1(keyinput112), .B2(n21691), .ZN(n21690) );
  OAI221_X1 U24619 ( .B1(n21692), .B2(keyinput89), .C1(n21691), .C2(
        keyinput112), .A(n21690), .ZN(n21701) );
  AOI22_X1 U24620 ( .A1(n17968), .A2(keyinput90), .B1(keyinput94), .B2(n21694), 
        .ZN(n21693) );
  OAI221_X1 U24621 ( .B1(n17968), .B2(keyinput90), .C1(n21694), .C2(keyinput94), .A(n21693), .ZN(n21700) );
  XNOR2_X1 U24622 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput6), 
        .ZN(n21698) );
  XNOR2_X1 U24623 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B(keyinput30), 
        .ZN(n21697) );
  XNOR2_X1 U24624 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B(keyinput116), .ZN(
        n21696) );
  XNOR2_X1 U24625 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(keyinput7), .ZN(
        n21695) );
  NAND4_X1 U24626 ( .A1(n21698), .A2(n21697), .A3(n21696), .A4(n21695), .ZN(
        n21699) );
  NOR3_X1 U24627 ( .A1(n21701), .A2(n21700), .A3(n21699), .ZN(n21733) );
  AOI22_X1 U24628 ( .A1(n21704), .A2(keyinput84), .B1(n21703), .B2(keyinput41), 
        .ZN(n21702) );
  OAI221_X1 U24629 ( .B1(n21704), .B2(keyinput84), .C1(n21703), .C2(keyinput41), .A(n21702), .ZN(n21715) );
  AOI22_X1 U24630 ( .A1(n21707), .A2(keyinput37), .B1(keyinput108), .B2(n21706), .ZN(n21705) );
  OAI221_X1 U24631 ( .B1(n21707), .B2(keyinput37), .C1(n21706), .C2(
        keyinput108), .A(n21705), .ZN(n21714) );
  AOI22_X1 U24632 ( .A1(n14248), .A2(keyinput32), .B1(n10871), .B2(keyinput104), .ZN(n21708) );
  OAI221_X1 U24633 ( .B1(n14248), .B2(keyinput32), .C1(n10871), .C2(
        keyinput104), .A(n21708), .ZN(n21713) );
  AOI22_X1 U24634 ( .A1(n21711), .A2(keyinput22), .B1(keyinput110), .B2(n21710), .ZN(n21709) );
  OAI221_X1 U24635 ( .B1(n21711), .B2(keyinput22), .C1(n21710), .C2(
        keyinput110), .A(n21709), .ZN(n21712) );
  NOR4_X1 U24636 ( .A1(n21715), .A2(n21714), .A3(n21713), .A4(n21712), .ZN(
        n21732) );
  AOI22_X1 U24637 ( .A1(n21718), .A2(keyinput111), .B1(keyinput19), .B2(n21717), .ZN(n21716) );
  OAI221_X1 U24638 ( .B1(n21718), .B2(keyinput111), .C1(n21717), .C2(
        keyinput19), .A(n21716), .ZN(n21730) );
  AOI22_X1 U24639 ( .A1(n21720), .A2(keyinput82), .B1(keyinput83), .B2(n14292), 
        .ZN(n21719) );
  OAI221_X1 U24640 ( .B1(n21720), .B2(keyinput82), .C1(n14292), .C2(keyinput83), .A(n21719), .ZN(n21729) );
  INV_X1 U24641 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n21722) );
  AOI22_X1 U24642 ( .A1(n21723), .A2(keyinput73), .B1(n21722), .B2(keyinput106), .ZN(n21721) );
  OAI221_X1 U24643 ( .B1(n21723), .B2(keyinput73), .C1(n21722), .C2(
        keyinput106), .A(n21721), .ZN(n21728) );
  AOI22_X1 U24644 ( .A1(n21726), .A2(keyinput58), .B1(keyinput114), .B2(n21725), .ZN(n21724) );
  OAI221_X1 U24645 ( .B1(n21726), .B2(keyinput58), .C1(n21725), .C2(
        keyinput114), .A(n21724), .ZN(n21727) );
  NOR4_X1 U24646 ( .A1(n21730), .A2(n21729), .A3(n21728), .A4(n21727), .ZN(
        n21731) );
  NAND4_X1 U24647 ( .A1(n21734), .A2(n21733), .A3(n21732), .A4(n21731), .ZN(
        n21800) );
  AOI22_X1 U24648 ( .A1(n16206), .A2(keyinput12), .B1(keyinput64), .B2(n21736), 
        .ZN(n21735) );
  OAI221_X1 U24649 ( .B1(n16206), .B2(keyinput12), .C1(n21736), .C2(keyinput64), .A(n21735), .ZN(n21748) );
  AOI22_X1 U24650 ( .A1(n21738), .A2(keyinput23), .B1(n11282), .B2(keyinput14), 
        .ZN(n21737) );
  OAI221_X1 U24651 ( .B1(n21738), .B2(keyinput23), .C1(n11282), .C2(keyinput14), .A(n21737), .ZN(n21747) );
  AOI22_X1 U24652 ( .A1(n21741), .A2(keyinput126), .B1(n21740), .B2(keyinput69), .ZN(n21739) );
  OAI221_X1 U24653 ( .B1(n21741), .B2(keyinput126), .C1(n21740), .C2(
        keyinput69), .A(n21739), .ZN(n21746) );
  AOI22_X1 U24654 ( .A1(n21744), .A2(keyinput119), .B1(n21743), .B2(keyinput13), .ZN(n21742) );
  OAI221_X1 U24655 ( .B1(n21744), .B2(keyinput119), .C1(n21743), .C2(
        keyinput13), .A(n21742), .ZN(n21745) );
  NOR4_X1 U24656 ( .A1(n21748), .A2(n21747), .A3(n21746), .A4(n21745), .ZN(
        n21798) );
  AOI22_X1 U24657 ( .A1(keyinput72), .A2(n21751), .B1(keyinput123), .B2(n21749), .ZN(n21750) );
  OAI21_X1 U24658 ( .B1(n21751), .B2(keyinput72), .A(n21750), .ZN(n21764) );
  AOI22_X1 U24659 ( .A1(n21754), .A2(keyinput16), .B1(keyinput50), .B2(n21753), 
        .ZN(n21752) );
  OAI221_X1 U24660 ( .B1(n21754), .B2(keyinput16), .C1(n21753), .C2(keyinput50), .A(n21752), .ZN(n21763) );
  INV_X1 U24661 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n21757) );
  AOI22_X1 U24662 ( .A1(n21757), .A2(keyinput76), .B1(keyinput62), .B2(n21756), 
        .ZN(n21755) );
  OAI221_X1 U24663 ( .B1(n21757), .B2(keyinput76), .C1(n21756), .C2(keyinput62), .A(n21755), .ZN(n21762) );
  AOI22_X1 U24664 ( .A1(n21760), .A2(keyinput21), .B1(keyinput74), .B2(n21759), 
        .ZN(n21758) );
  OAI221_X1 U24665 ( .B1(n21760), .B2(keyinput21), .C1(n21759), .C2(keyinput74), .A(n21758), .ZN(n21761) );
  NOR4_X1 U24666 ( .A1(n21764), .A2(n21763), .A3(n21762), .A4(n21761), .ZN(
        n21797) );
  AOI22_X1 U24667 ( .A1(n14256), .A2(keyinput120), .B1(keyinput124), .B2(
        n21766), .ZN(n21765) );
  OAI221_X1 U24668 ( .B1(n14256), .B2(keyinput120), .C1(n21766), .C2(
        keyinput124), .A(n21765), .ZN(n21771) );
  XNOR2_X1 U24669 ( .A(n21767), .B(keyinput100), .ZN(n21770) );
  XOR2_X1 U24670 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B(keyinput48), .Z(
        n21769) );
  XOR2_X1 U24671 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B(keyinput80), .Z(
        n21768) );
  OR4_X1 U24672 ( .A1(n21771), .A2(n21770), .A3(n21769), .A4(n21768), .ZN(
        n21778) );
  AOI22_X1 U24673 ( .A1(n21774), .A2(keyinput57), .B1(keyinput43), .B2(n21773), 
        .ZN(n21772) );
  OAI221_X1 U24674 ( .B1(n21774), .B2(keyinput57), .C1(n21773), .C2(keyinput43), .A(n21772), .ZN(n21777) );
  XNOR2_X1 U24675 ( .A(n21775), .B(keyinput122), .ZN(n21776) );
  NOR3_X1 U24676 ( .A1(n21778), .A2(n21777), .A3(n21776), .ZN(n21796) );
  AOI22_X1 U24677 ( .A1(n21781), .A2(keyinput121), .B1(keyinput53), .B2(n21780), .ZN(n21779) );
  OAI221_X1 U24678 ( .B1(n21781), .B2(keyinput121), .C1(n21780), .C2(
        keyinput53), .A(n21779), .ZN(n21794) );
  INV_X1 U24679 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n21784) );
  AOI22_X1 U24680 ( .A1(n21784), .A2(keyinput20), .B1(keyinput40), .B2(n21783), 
        .ZN(n21782) );
  OAI221_X1 U24681 ( .B1(n21784), .B2(keyinput20), .C1(n21783), .C2(keyinput40), .A(n21782), .ZN(n21793) );
  AOI22_X1 U24682 ( .A1(n21787), .A2(keyinput5), .B1(keyinput99), .B2(n21786), 
        .ZN(n21785) );
  OAI221_X1 U24683 ( .B1(n21787), .B2(keyinput5), .C1(n21786), .C2(keyinput99), 
        .A(n21785), .ZN(n21792) );
  AOI22_X1 U24684 ( .A1(n21790), .A2(keyinput1), .B1(keyinput85), .B2(n21789), 
        .ZN(n21788) );
  OAI221_X1 U24685 ( .B1(n21790), .B2(keyinput1), .C1(n21789), .C2(keyinput85), 
        .A(n21788), .ZN(n21791) );
  NOR4_X1 U24686 ( .A1(n21794), .A2(n21793), .A3(n21792), .A4(n21791), .ZN(
        n21795) );
  NAND4_X1 U24687 ( .A1(n21798), .A2(n21797), .A3(n21796), .A4(n21795), .ZN(
        n21799) );
  NOR4_X1 U24688 ( .A1(n21802), .A2(n21801), .A3(n21800), .A4(n21799), .ZN(
        n21803) );
  OAI21_X1 U24689 ( .B1(keyinput123), .B2(n21804), .A(n21803), .ZN(n21805) );
  XNOR2_X1 U24690 ( .A(n21806), .B(n21805), .ZN(P1_U2947) );
  NAND2_X1 U11365 ( .A1(n16246), .A2(n10786), .ZN(n10870) );
  NOR2_X2 U13115 ( .A1(n10803), .A2(n12681), .ZN(n20099) );
  AND2_X1 U13095 ( .A1(n10809), .A2(n10806), .ZN(n20061) );
  AND2_X1 U13097 ( .A1(n10809), .A2(n10799), .ZN(n10877) );
  AND2_X1 U14060 ( .A1(n10809), .A2(n10808), .ZN(n10876) );
  BUF_X2 U11156 ( .A(n14760), .Z(n16643) );
  CLKBUF_X2 U11189 ( .A(n11975), .Z(n14784) );
  CLKBUF_X1 U11211 ( .A(n11093), .Z(n11094) );
  CLKBUF_X1 U11289 ( .A(n11940), .Z(n20796) );
  CLKBUF_X2 U11531 ( .A(n11130), .Z(n10980) );
  AND2_X1 U11791 ( .A1(n14070), .A2(n10810), .ZN(n10807) );
  AND2_X1 U12531 ( .A1(n10809), .A2(n10796), .ZN(n10864) );
  CLKBUF_X1 U12897 ( .A(n12293), .Z(n21463) );
  CLKBUF_X1 U12953 ( .A(n16485), .Z(n16486) );
  NAND2_X1 U13060 ( .A1(n16643), .A2(n11563), .ZN(n9836) );
  CLKBUF_X1 U13297 ( .A(n10755), .Z(n14514) );
  CLKBUF_X1 U14053 ( .A(n12009), .Z(n11973) );
endmodule

