

module b15_C_AntiSAT_k_128_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3011, n3012, n3013, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802;

  CLKBUF_X2 U3441 ( .A(n4077), .Z(n4686) );
  AOI21_X1 U3443 ( .B1(n4329), .B2(n6599), .A(n3228), .ZN(n3230) );
  CLKBUF_X2 U3444 ( .A(n3141), .Z(n3837) );
  CLKBUF_X2 U34450 ( .A(n3072), .Z(n3775) );
  CLKBUF_X2 U34460 ( .A(n3824), .Z(n3013) );
  CLKBUF_X2 U34470 ( .A(n3123), .Z(n3840) );
  CLKBUF_X1 U34480 ( .A(n3073), .Z(n3800) );
  CLKBUF_X2 U3449 ( .A(n3096), .Z(n3730) );
  CLKBUF_X1 U3450 ( .A(n3452), .Z(n3848) );
  CLKBUF_X1 U34510 ( .A(n3780), .Z(n3007) );
  NOR2_X1 U34520 ( .A1(n3926), .A2(n5072), .ZN(n4218) );
  OR2_X1 U34530 ( .A1(n3187), .A2(n3935), .ZN(n3179) );
  AND4_X1 U3454 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3084)
         );
  AND2_X1 U34550 ( .A1(n4212), .A2(n4561), .ZN(n3072) );
  AND2_X1 U34560 ( .A1(n3033), .A2(n4212), .ZN(n3073) );
  AND2_X1 U3457 ( .A1(n4216), .A2(n3033), .ZN(n3824) );
  AND2_X2 U3458 ( .A1(n3042), .A2(n4561), .ZN(n3118) );
  AND2_X1 U34590 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4211) );
  CLKBUF_X1 U34600 ( .A(n6129), .Z(n2993) );
  NOR2_X1 U34610 ( .A1(n5075), .A2(n5074), .ZN(n6129) );
  AND4_X1 U34630 ( .A1(n3032), .A2(n3031), .A3(n3030), .A4(n3029), .ZN(n3050)
         );
  AND4_X1 U34640 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n3021)
         );
  NAND2_X1 U34650 ( .A1(n3299), .A2(n3281), .ZN(n3290) );
  BUF_X1 U3466 ( .A(n4161), .Z(n5723) );
  AND4_X1 U3467 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3135)
         );
  AND2_X1 U34680 ( .A1(n5279), .A2(n3286), .ZN(n3198) );
  NAND2_X1 U34700 ( .A1(n3313), .A2(n4303), .ZN(n4310) );
  INV_X4 U34710 ( .A(n5824), .ZN(n5720) );
  INV_X1 U34720 ( .A(n6102), .ZN(n6135) );
  CLKBUF_X1 U34730 ( .A(n3097), .Z(n2994) );
  INV_X1 U34740 ( .A(n3158), .ZN(n3061) );
  NOR2_X2 U3475 ( .A1(n5703), .A2(n5463), .ZN(n5480) );
  NAND2_X2 U3476 ( .A1(n5462), .A2(n5461), .ZN(n5703) );
  OAI21_X2 U3477 ( .B1(n5547), .B2(n5271), .A(n5444), .ZN(n5470) );
  NOR2_X2 U3478 ( .A1(n5438), .A2(n5466), .ZN(n5481) );
  AND2_X1 U3479 ( .A1(n4216), .A2(n4542), .ZN(n3780) );
  AND2_X2 U3481 ( .A1(n3026), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3033)
         );
  AND2_X1 U3482 ( .A1(n5656), .A2(n4050), .ZN(n4053) );
  NAND2_X1 U3483 ( .A1(n5270), .A2(n5271), .ZN(n5444) );
  OR2_X1 U3485 ( .A1(n3411), .A2(n3410), .ZN(n4126) );
  NAND2_X2 U3486 ( .A1(n4286), .A2(n4285), .ZN(n4284) );
  NAND2_X1 U3487 ( .A1(n3177), .A2(n3176), .ZN(n3260) );
  BUF_X1 U3488 ( .A(n3181), .Z(n4348) );
  INV_X1 U3489 ( .A(n4257), .ZN(n3109) );
  INV_X1 U3490 ( .A(n4557), .ZN(n3096) );
  CLKBUF_X2 U3492 ( .A(n3103), .Z(n3735) );
  NAND2_X1 U3493 ( .A1(n3033), .A2(n4211), .ZN(n4557) );
  CLKBUF_X2 U3494 ( .A(n3102), .Z(n3847) );
  NOR2_X4 U3495 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4561) );
  AND2_X2 U3496 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4542) );
  AND2_X1 U3497 ( .A1(n5336), .A2(n5459), .ZN(n5458) );
  CLKBUF_X1 U3498 ( .A(n4163), .Z(n5378) );
  NOR2_X1 U3499 ( .A1(n5444), .A2(n5443), .ZN(n5448) );
  AND2_X1 U3500 ( .A1(n5656), .A2(n5655), .ZN(n6147) );
  OAI21_X1 U3501 ( .B1(n5395), .B2(n5394), .A(n5645), .ZN(n5652) );
  CLKBUF_X1 U3502 ( .A(n5270), .Z(n5547) );
  OR2_X1 U3503 ( .A1(n5578), .A2(n5579), .ZN(n5654) );
  NOR2_X1 U3504 ( .A1(n5368), .A2(n5548), .ZN(n5270) );
  OAI21_X1 U3505 ( .B1(n5592), .B2(n5327), .A(n5578), .ZN(n5665) );
  OR2_X1 U3506 ( .A1(n4170), .A2(n5619), .ZN(n5610) );
  AND2_X1 U3507 ( .A1(n3509), .A2(n3508), .ZN(n5256) );
  CLKBUF_X1 U3508 ( .A(n4870), .Z(n5032) );
  NOR2_X2 U3509 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  AOI21_X1 U3510 ( .B1(n4112), .B2(n3724), .A(n3418), .ZN(n4868) );
  AOI21_X1 U3511 ( .B1(n4686), .B2(n3724), .A(n3348), .ZN(n4309) );
  AOI21_X1 U3512 ( .B1(n4094), .B2(n3724), .A(n3388), .ZN(n4414) );
  NOR2_X2 U3513 ( .A1(n5595), .A2(n5594), .ZN(n5667) );
  XNOR2_X1 U3514 ( .A(n3383), .B(n3389), .ZN(n4094) );
  AND2_X1 U3515 ( .A1(n3340), .A2(n3369), .ZN(n4077) );
  OR2_X2 U3516 ( .A1(n5267), .A2(n5266), .ZN(n5595) );
  INV_X1 U3517 ( .A(n3369), .ZN(n3392) );
  NAND2_X1 U3518 ( .A1(n3285), .A2(n3284), .ZN(n3338) );
  OAI21_X1 U3519 ( .B1(n3283), .B2(n3282), .A(n3290), .ZN(n3285) );
  XNOR2_X1 U3521 ( .A(n3230), .B(n3229), .ZN(n3314) );
  NAND2_X1 U3522 ( .A1(n3317), .A2(n3316), .ZN(n4538) );
  NAND2_X2 U3523 ( .A1(n5453), .A2(n4300), .ZN(n5917) );
  OR2_X1 U3524 ( .A1(n3301), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U3525 ( .A1(n3260), .A2(n3261), .ZN(n3264) );
  OR2_X1 U3526 ( .A1(n4195), .A2(n4059), .ZN(n5522) );
  CLKBUF_X1 U3527 ( .A(n3924), .Z(n4210) );
  AND2_X1 U3528 ( .A1(n3951), .A2(n3950), .ZN(n4307) );
  AND3_X1 U3529 ( .A1(n3184), .A2(n3183), .A3(n4205), .ZN(n3191) );
  NAND2_X1 U3530 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  CLKBUF_X1 U3531 ( .A(n3186), .Z(n4202) );
  BUF_X1 U3532 ( .A(n3945), .Z(n4028) );
  NAND2_X1 U3533 ( .A1(n3110), .A2(n3109), .ZN(n3553) );
  OR2_X1 U3534 ( .A1(n3945), .A2(EBX_REG_1__SCAN_IN), .ZN(n3943) );
  INV_X1 U3535 ( .A(n3920), .ZN(n4054) );
  AND2_X2 U3536 ( .A1(n3873), .A2(n3109), .ZN(n3903) );
  NAND2_X1 U3537 ( .A1(n3196), .A2(n4257), .ZN(n3180) );
  OR2_X1 U3538 ( .A1(n3935), .A2(n3181), .ZN(n3920) );
  NAND2_X1 U3539 ( .A1(n3927), .A2(n3926), .ZN(n3934) );
  NAND3_X1 U3540 ( .A1(n3094), .A2(n3022), .A3(n3017), .ZN(n3181) );
  AND2_X2 U3541 ( .A1(n3108), .A2(n3016), .ZN(n4257) );
  NAND4_X1 U3542 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3927)
         );
  NAND4_X2 U3543 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .ZN(n3158)
         );
  NAND2_X2 U3544 ( .A1(n3021), .A2(n3060), .ZN(n3286) );
  AND4_X1 U3545 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3156)
         );
  AND4_X1 U3546 ( .A1(n3140), .A2(n3139), .A3(n3138), .A4(n3137), .ZN(n3157)
         );
  AND4_X1 U3547 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3049)
         );
  AND4_X1 U3548 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3154)
         );
  AND4_X1 U3549 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3136)
         );
  AND4_X1 U3550 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n3060)
         );
  AND4_X1 U3551 ( .A1(n3041), .A2(n3040), .A3(n3039), .A4(n3038), .ZN(n3048)
         );
  AND4_X1 U3552 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3047)
         );
  AND4_X1 U3553 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3134)
         );
  AND4_X1 U3554 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3133)
         );
  AND4_X1 U3555 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3155)
         );
  CLKBUF_X1 U3556 ( .A(n3759), .Z(n3818) );
  AND3_X1 U3557 ( .A1(n3081), .A2(n3080), .A3(n3079), .ZN(n3083) );
  AND2_X2 U3558 ( .A1(n3042), .A2(n4542), .ZN(n3221) );
  AND2_X2 U3559 ( .A1(n4555), .A2(n4211), .ZN(n3452) );
  INV_X2 U3560 ( .A(n6535), .ZN(n6607) );
  AND2_X2 U3561 ( .A1(n4561), .A2(n4211), .ZN(n3846) );
  NOR2_X2 U3562 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5055) );
  NOR2_X1 U3563 ( .A1(n4170), .A2(n2995), .ZN(n5612) );
  OR2_X1 U3564 ( .A1(n5619), .A2(n5611), .ZN(n2995) );
  XNOR2_X1 U3565 ( .A(n5444), .B(n3869), .ZN(n5496) );
  NAND2_X2 U3567 ( .A1(n5401), .A2(n4131), .ZN(n5160) );
  NAND2_X1 U3568 ( .A1(n5160), .A2(n3000), .ZN(n2997) );
  AND2_X2 U3569 ( .A1(n2997), .A2(n2998), .ZN(n6220) );
  OR2_X1 U3570 ( .A1(n2999), .A2(n5159), .ZN(n2998) );
  INV_X1 U3571 ( .A(n5215), .ZN(n2999) );
  AND2_X1 U3572 ( .A1(n5158), .A2(n5215), .ZN(n3000) );
  AND2_X1 U3573 ( .A1(n3260), .A2(n3261), .ZN(n3001) );
  XNOR2_X1 U3574 ( .A(n3001), .B(n3233), .ZN(n4191) );
  AND2_X1 U3575 ( .A1(n5225), .A2(n3002), .ZN(n3003) );
  INV_X1 U3576 ( .A(n5185), .ZN(n3002) );
  AND2_X1 U3577 ( .A1(n5034), .A2(n3002), .ZN(n5226) );
  NAND2_X1 U3578 ( .A1(n5411), .A2(n3004), .ZN(n5617) );
  AND2_X1 U3579 ( .A1(n5621), .A2(n3005), .ZN(n3004) );
  INV_X1 U3580 ( .A(n5615), .ZN(n3005) );
  NOR2_X2 U3581 ( .A1(n5551), .A2(n5550), .ZN(n5278) );
  OR2_X1 U3582 ( .A1(n5617), .A2(n5357), .ZN(n5551) );
  AND2_X2 U3583 ( .A1(n3025), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4216)
         );
  INV_X1 U3584 ( .A(n3314), .ZN(n3339) );
  BUF_X1 U3588 ( .A(n3452), .Z(n3011) );
  AND2_X1 U3589 ( .A1(n4555), .A2(n4212), .ZN(n3089) );
  BUF_X1 U3590 ( .A(n3089), .Z(n3838) );
  AND2_X1 U3591 ( .A1(n4216), .A2(n4555), .ZN(n3012) );
  AND2_X1 U3592 ( .A1(n4216), .A2(n4555), .ZN(n3123) );
  NOR2_X4 U3593 ( .A1(n3061), .A2(n3286), .ZN(n3187) );
  NAND2_X1 U3596 ( .A1(n4030), .A2(n4262), .ZN(n5272) );
  XNOR2_X1 U3597 ( .A(n3291), .B(n3290), .ZN(n4322) );
  AND2_X1 U3598 ( .A1(n4216), .A2(n4561), .ZN(n3141) );
  AND2_X2 U3599 ( .A1(n5633), .A2(n5412), .ZN(n5411) );
  NOR2_X1 U3600 ( .A1(n5480), .A2(n5481), .ZN(n5464) );
  OR2_X2 U3601 ( .A1(n5640), .A2(n5641), .ZN(n5632) );
  AND2_X1 U3602 ( .A1(n4216), .A2(n4542), .ZN(n3015) );
  AND2_X2 U3603 ( .A1(n3003), .A2(n5034), .ZN(n5224) );
  NAND2_X1 U3604 ( .A1(n4059), .A2(n3926), .ZN(n4188) );
  INV_X1 U3605 ( .A(n3926), .ZN(n4243) );
  NAND2_X1 U3606 ( .A1(n3392), .A2(n3391), .ZN(n3411) );
  AND2_X1 U3607 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  NAND2_X1 U3608 ( .A1(n5307), .A2(n4030), .ZN(n3945) );
  AND2_X1 U3609 ( .A1(n3015), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3051) );
  OR2_X1 U3610 ( .A1(n3684), .A2(n5593), .ZN(n5635) );
  INV_X1 U3611 ( .A(n3198), .ZN(n4244) );
  INV_X1 U3612 ( .A(n3181), .ZN(n4246) );
  AND3_X1 U3613 ( .A1(n3259), .A2(n3258), .A3(n3257), .ZN(n3288) );
  OAI21_X1 U3614 ( .B1(n5993), .B2(n4580), .A(n6483), .ZN(n4331) );
  CLKBUF_X1 U3615 ( .A(n4195), .Z(n4196) );
  NAND2_X1 U3616 ( .A1(n6066), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5075) );
  AND2_X1 U3617 ( .A1(n4229), .A2(n4228), .ZN(n5514) );
  OR2_X1 U3618 ( .A1(n3711), .A2(n4169), .ZN(n3728) );
  AND2_X1 U3619 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3628), .ZN(n3627)
         );
  AND2_X1 U3620 ( .A1(n5943), .A2(n4141), .ZN(n4142) );
  AND2_X1 U3621 ( .A1(n3405), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3430)
         );
  NAND2_X1 U3622 ( .A1(n3364), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3384)
         );
  INV_X1 U3623 ( .A(n4294), .ZN(n4373) );
  NAND2_X1 U3624 ( .A1(n5458), .A2(n5705), .ZN(n5438) );
  XNOR2_X1 U3625 ( .A(n3314), .B(n3338), .ZN(n4321) );
  AND2_X1 U3626 ( .A1(n3917), .A2(n3916), .ZN(n5524) );
  NOR2_X1 U3627 ( .A1(n5485), .A2(n6145), .ZN(n5430) );
  NOR2_X1 U3628 ( .A1(n5485), .A2(n5670), .ZN(n4047) );
  XNOR2_X1 U3629 ( .A(n5448), .B(n5447), .ZN(n5529) );
  INV_X1 U3630 ( .A(n5443), .ZN(n3869) );
  INV_X1 U3631 ( .A(n5415), .ZN(n5421) );
  CLKBUF_X1 U3632 ( .A(n4324), .Z(n4888) );
  CLKBUF_X1 U3633 ( .A(n4322), .Z(n5837) );
  CLKBUF_X1 U3634 ( .A(n4321), .Z(n5841) );
  AND2_X1 U3635 ( .A1(n5072), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3873) );
  CLKBUF_X1 U3636 ( .A(n3800), .Z(n3823) );
  OR2_X1 U3637 ( .A1(n3243), .A2(n3242), .ZN(n4067) );
  NAND2_X1 U3638 ( .A1(n4257), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4123) );
  AND2_X2 U3639 ( .A1(n3027), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3042)
         );
  INV_X1 U3640 ( .A(n3180), .ZN(n3874) );
  OR2_X1 U3641 ( .A1(n5635), .A2(n5637), .ZN(n5627) );
  OR2_X1 U3642 ( .A1(n6452), .A2(n6599), .ZN(n3863) );
  OR2_X1 U3643 ( .A1(n5720), .A2(n4149), .ZN(n4150) );
  NAND2_X1 U3644 ( .A1(n5824), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4135) );
  NAND2_X1 U3645 ( .A1(n3953), .A2(n3952), .ZN(n4304) );
  INV_X1 U3646 ( .A(n4307), .ZN(n3952) );
  INV_X1 U3647 ( .A(n4306), .ZN(n3953) );
  OR2_X1 U3648 ( .A1(n3275), .A2(n3274), .ZN(n4068) );
  NAND2_X1 U3649 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  NAND2_X1 U3650 ( .A1(n3903), .A2(n4122), .ZN(n3915) );
  NAND2_X1 U3651 ( .A1(n4123), .A2(n3323), .ZN(n3911) );
  AND2_X1 U3652 ( .A1(n3910), .A2(n3909), .ZN(n3914) );
  NAND2_X1 U3653 ( .A1(n3216), .A2(n3215), .ZN(n3316) );
  XNOR2_X1 U3654 ( .A(n4538), .B(n4536), .ZN(n4327) );
  INV_X1 U3655 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4716) );
  INV_X1 U3656 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6461) );
  INV_X1 U3657 ( .A(n5075), .ZN(n5148) );
  OR2_X1 U3658 ( .A1(n3796), .A2(n5554), .ZN(n3865) );
  AND2_X1 U3659 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3556), .ZN(n3699)
         );
  AND2_X1 U3660 ( .A1(n3627), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3594)
         );
  NOR2_X1 U3661 ( .A1(n3635), .A2(n5586), .ZN(n3628) );
  NOR2_X1 U3662 ( .A1(n3669), .A2(n5601), .ZN(n3652) );
  AND2_X1 U3663 ( .A1(n3497), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3498)
         );
  NAND2_X1 U3664 ( .A1(n3498), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3712)
         );
  NAND2_X1 U3665 ( .A1(n3521), .A2(n3502), .ZN(n3508) );
  NOR2_X1 U3666 ( .A1(n3492), .A2(n3491), .ZN(n3497) );
  NAND2_X1 U3667 ( .A1(n3467), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3492)
         );
  NOR2_X1 U3668 ( .A1(n6757), .A2(n3436), .ZN(n3467) );
  CLKBUF_X1 U3669 ( .A(n5030), .Z(n5031) );
  AND2_X1 U3670 ( .A1(n3430), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3435)
         );
  AOI21_X1 U3671 ( .B1(n4102), .B2(n3724), .A(n3409), .ZN(n4619) );
  NOR2_X1 U3672 ( .A1(n3384), .A2(n5076), .ZN(n3405) );
  INV_X1 U3673 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5076) );
  AND2_X1 U3674 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3341), .ZN(n3364)
         );
  NAND2_X1 U3675 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U3676 ( .A1(n4022), .A2(n4262), .ZN(n5531) );
  OR2_X1 U3677 ( .A1(n5984), .A2(n5364), .ZN(n5831) );
  CLKBUF_X1 U3678 ( .A(n5323), .Z(n5825) );
  AND2_X1 U3679 ( .A1(n5720), .A2(n5298), .ZN(n4144) );
  OR2_X2 U3680 ( .A1(n4152), .A2(n5072), .ZN(n4263) );
  CLKBUF_X1 U3681 ( .A(n5246), .Z(n5942) );
  OR2_X1 U3682 ( .A1(n5720), .A2(n4133), .ZN(n6219) );
  OR2_X1 U3683 ( .A1(n5720), .A2(n5174), .ZN(n5159) );
  OR2_X1 U3684 ( .A1(n6579), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4156) );
  AND2_X1 U3685 ( .A1(n3969), .A2(n3968), .ZN(n4622) );
  OR2_X1 U3686 ( .A1(n5975), .A2(n5977), .ZN(n5345) );
  OAI21_X1 U3687 ( .B1(n4255), .B2(n4294), .A(n4254), .ZN(n4275) );
  NAND2_X1 U3688 ( .A1(n3263), .A2(n3262), .ZN(n3265) );
  XNOR2_X1 U3689 ( .A(n3289), .B(n3288), .ZN(n3291) );
  CLKBUF_X1 U3690 ( .A(n4191), .Z(n4192) );
  CLKBUF_X1 U3691 ( .A(n4329), .Z(n5205) );
  OR2_X1 U3692 ( .A1(n4298), .A2(n4231), .ZN(n6458) );
  INV_X1 U3693 ( .A(n5841), .ZN(n4628) );
  OR2_X1 U3694 ( .A1(n4607), .A2(n5837), .ZN(n4889) );
  NOR2_X1 U3695 ( .A1(n4714), .A2(n5837), .ZN(n4723) );
  CLKBUF_X1 U3696 ( .A(n4327), .Z(n4632) );
  INV_X1 U3697 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U3698 ( .A1(n6599), .A2(n4331), .ZN(n4572) );
  CLKBUF_X1 U3699 ( .A(n3286), .Z(n4353) );
  AND2_X1 U3700 ( .A1(n4326), .A2(n4331), .ZN(n4365) );
  AND2_X1 U3701 ( .A1(n6066), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6133) );
  AND2_X1 U3702 ( .A1(n6066), .A2(n5067), .ZN(n6102) );
  INV_X1 U3703 ( .A(n6099), .ZN(n6112) );
  AND2_X1 U3704 ( .A1(n5539), .A2(n5066), .ZN(n6079) );
  NAND2_X1 U3705 ( .A1(n3933), .A2(n5528), .ZN(n5674) );
  INV_X1 U3706 ( .A(n5670), .ZN(n5675) );
  OR2_X1 U3707 ( .A1(n5674), .A2(n5279), .ZN(n5670) );
  INV_X1 U3708 ( .A(n5496), .ZN(n5437) );
  AND2_X1 U3709 ( .A1(n5453), .A2(n4301), .ZN(n5689) );
  NOR2_X1 U3710 ( .A1(n6604), .A2(n6160), .ZN(n6175) );
  INV_X1 U3711 ( .A(n6217), .ZN(n6211) );
  INV_X1 U3712 ( .A(n4843), .ZN(n6215) );
  INV_X1 U3713 ( .A(n6196), .ZN(n6214) );
  AOI21_X1 U3714 ( .B1(n5646), .B2(n5645), .A(n5644), .ZN(n5924) );
  CLKBUF_X1 U3715 ( .A(n5297), .Z(n5300) );
  NAND2_X1 U3716 ( .A1(n5481), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5482) );
  NOR2_X1 U3717 ( .A1(n6256), .A2(n5976), .ZN(n5984) );
  INV_X1 U3718 ( .A(n6283), .ZN(n6338) );
  AND2_X1 U3719 ( .A1(n4275), .A2(n6454), .ZN(n5975) );
  AND2_X1 U3720 ( .A1(n5837), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5840) );
  INV_X1 U3721 ( .A(n5836), .ZN(n5844) );
  NOR2_X1 U3722 ( .A1(n3174), .A2(n5524), .ZN(n5500) );
  CLKBUF_X1 U3723 ( .A(n4193), .Z(n4194) );
  CLKBUF_X1 U3724 ( .A(n4639), .Z(n5141) );
  INV_X1 U3725 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6599) );
  INV_X1 U3726 ( .A(n5500), .ZN(n6483) );
  NOR2_X1 U3727 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  NOR2_X1 U3728 ( .A1(n5669), .A2(n4045), .ZN(n4046) );
  AOI21_X1 U3729 ( .B1(n5529), .B2(n6225), .A(n5451), .ZN(n5452) );
  OAI21_X1 U3730 ( .B1(n5686), .B2(n5406), .A(n4174), .ZN(n4175) );
  OAI21_X1 U3731 ( .B1(n5823), .B2(n6229), .A(n4158), .ZN(n4159) );
  AOI21_X1 U3732 ( .B1(n6224), .B2(n5315), .A(n4157), .ZN(n4158) );
  NAND2_X1 U3733 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  OR2_X2 U3734 ( .A1(n3071), .A2(n3070), .ZN(n4364) );
  NAND2_X1 U3735 ( .A1(n5265), .A2(n3729), .ZN(n4170) );
  NOR2_X1 U3736 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  INV_X1 U3737 ( .A(n4409), .ZN(n3964) );
  AND4_X1 U3738 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(n3016)
         );
  AND4_X1 U3739 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3017)
         );
  NAND2_X1 U3740 ( .A1(n5720), .A2(n4147), .ZN(n3018) );
  AND2_X1 U3741 ( .A1(n6219), .A2(n4135), .ZN(n3019) );
  NOR2_X2 U3742 ( .A1(n4889), .A2(n4888), .ZN(n3020) );
  NAND2_X1 U3743 ( .A1(n5738), .A2(n5729), .ZN(n5721) );
  AND3_X1 U3744 ( .A1(n3088), .A2(n3087), .A3(n3086), .ZN(n3022) );
  INV_X1 U3745 ( .A(n4415), .ZN(n3963) );
  INV_X1 U3746 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U3747 ( .A1(n3336), .A2(n3335), .ZN(n3337) );
  INV_X1 U3748 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6466) );
  INV_X1 U3749 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5479) );
  XOR2_X1 U3750 ( .A(n5536), .B(n5535), .Z(n3023) );
  OR2_X1 U3751 ( .A1(n3205), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3024)
         );
  INV_X1 U3752 ( .A(n3159), .ZN(n3160) );
  NOR2_X1 U3753 ( .A1(n3165), .A2(n4202), .ZN(n3169) );
  NAND2_X1 U3754 ( .A1(n3903), .A2(n3171), .ZN(n3172) );
  NAND2_X1 U3755 ( .A1(n3199), .A2(n4218), .ZN(n3185) );
  OR2_X1 U3756 ( .A1(n3358), .A2(n3357), .ZN(n4104) );
  AOI22_X1 U3757 ( .A1(n3124), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3086) );
  AOI21_X1 U3758 ( .B1(n3097), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n3051), 
        .ZN(n3055) );
  AND2_X1 U3759 ( .A1(n6455), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3884)
         );
  BUF_X1 U3761 ( .A(n3221), .Z(n3839) );
  AND2_X1 U3762 ( .A1(n3162), .A2(n5279), .ZN(n3163) );
  OR2_X1 U3763 ( .A1(n3227), .A2(n3226), .ZN(n4069) );
  NAND2_X1 U3764 ( .A1(n3204), .A2(n3024), .ZN(n3232) );
  INV_X1 U3765 ( .A(n3288), .ZN(n3282) );
  AOI22_X1 U3766 ( .A1(n3073), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3098) );
  NOR2_X1 U3767 ( .A1(n3707), .A2(n3558), .ZN(n3748) );
  OR2_X1 U3768 ( .A1(n3255), .A2(n3254), .ZN(n4121) );
  OR2_X1 U3769 ( .A1(n5072), .A2(n6599), .ZN(n3323) );
  AND4_X1 U3770 ( .A1(n3101), .A2(n3100), .A3(n3099), .A4(n3098), .ZN(n3108)
         );
  NOR2_X1 U3771 ( .A1(n3920), .A2(n3196), .ZN(n3194) );
  OR2_X1 U3772 ( .A1(n5941), .A2(n4137), .ZN(n4138) );
  NAND2_X1 U3773 ( .A1(n3085), .A2(n5279), .ZN(n4264) );
  AND2_X1 U3774 ( .A1(n3404), .A2(n3403), .ZN(n3410) );
  NAND2_X1 U3775 ( .A1(n3964), .A2(n3963), .ZN(n4416) );
  OR2_X1 U3776 ( .A1(n4296), .A2(n4244), .ZN(n4273) );
  INV_X1 U3777 ( .A(n3553), .ZN(n3554) );
  AND2_X2 U3778 ( .A1(n3028), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4555)
         );
  NAND2_X1 U3779 ( .A1(n3322), .A2(n3321), .ZN(n4536) );
  INV_X1 U3780 ( .A(n3927), .ZN(n4059) );
  INV_X1 U3781 ( .A(n3954), .ZN(n4022) );
  NOR2_X1 U3782 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  NAND2_X1 U3783 ( .A1(n3928), .A2(n4218), .ZN(n4296) );
  OR2_X1 U3784 ( .A1(n5059), .A2(n5426), .ZN(n5061) );
  OR2_X1 U3785 ( .A1(n3769), .A2(n6737), .ZN(n3794) );
  OR2_X1 U3786 ( .A1(n3712), .A2(n6038), .ZN(n3669) );
  INV_X1 U3787 ( .A(n5179), .ZN(n3466) );
  XNOR2_X1 U3788 ( .A(n4126), .B(n3413), .ZN(n4112) );
  INV_X1 U3789 ( .A(n4264), .ZN(n3300) );
  NAND2_X1 U3790 ( .A1(n4039), .A2(n5532), .ZN(n4044) );
  NAND2_X1 U3791 ( .A1(n5335), .A2(n5334), .ZN(n5457) );
  CLKBUF_X1 U3792 ( .A(n4416), .Z(n4623) );
  NAND2_X1 U3793 ( .A1(n3937), .A2(n3936), .ZN(n4236) );
  AND2_X1 U3794 ( .A1(n3926), .A2(n3196), .ZN(n4122) );
  OR2_X1 U3795 ( .A1(n3915), .A2(n4182), .ZN(n3916) );
  NAND2_X1 U3796 ( .A1(n4327), .A2(n6599), .ZN(n3336) );
  AND2_X2 U3797 ( .A1(n3280), .A2(n3279), .ZN(n3299) );
  AND2_X1 U3798 ( .A1(n2993), .A2(EBX_REG_30__SCAN_IN), .ZN(n5427) );
  INV_X1 U3799 ( .A(n3593), .ZN(n3556) );
  NAND2_X1 U3800 ( .A1(n5667), .A2(n5666), .ZN(n5580) );
  NAND2_X1 U3801 ( .A1(n3435), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3436)
         );
  NAND2_X1 U3802 ( .A1(n5148), .A2(n5064), .ZN(n6083) );
  OR2_X1 U3803 ( .A1(n5627), .A2(n3710), .ZN(n4169) );
  INV_X1 U3804 ( .A(n4868), .ZN(n3419) );
  NAND2_X1 U3805 ( .A1(n3594), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3593)
         );
  NAND2_X1 U3806 ( .A1(n4051), .A2(n5327), .ZN(n5578) );
  INV_X1 U3807 ( .A(n5031), .ZN(n5180) );
  INV_X1 U3808 ( .A(n4618), .ZN(n4867) );
  AND2_X1 U3809 ( .A1(n4044), .A2(n4043), .ZN(n5485) );
  NAND2_X1 U3810 ( .A1(n5703), .A2(n5692), .ZN(n5696) );
  INV_X1 U3811 ( .A(n5419), .ZN(n5420) );
  NOR2_X1 U3812 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5729)
         );
  AND2_X1 U3813 ( .A1(n4126), .A2(n4125), .ZN(n5824) );
  AND2_X1 U3814 ( .A1(n3981), .A2(n3980), .ZN(n5185) );
  OR2_X1 U3815 ( .A1(n5524), .A2(n6488), .ZN(n4294) );
  CLKBUF_X1 U3816 ( .A(n4211), .Z(n5499) );
  OR2_X1 U3817 ( .A1(n4574), .A2(n4722), .ZN(n4743) );
  OR2_X1 U3818 ( .A1(n5428), .A2(n5427), .ZN(n5429) );
  NAND2_X1 U3819 ( .A1(n3699), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3707)
         );
  OR2_X1 U3820 ( .A1(n6601), .A2(n5058), .ZN(n6066) );
  CLKBUF_X1 U3821 ( .A(n4874), .Z(n5035) );
  NAND2_X1 U3822 ( .A1(n4287), .A2(n4030), .ZN(n4290) );
  AND2_X1 U3823 ( .A1(n5453), .A2(n5280), .ZN(n6157) );
  INV_X1 U3824 ( .A(n5453), .ZN(n6156) );
  AND2_X1 U3825 ( .A1(n4375), .A2(n5525), .ZN(n6160) );
  AOI21_X1 U3826 ( .B1(n5548), .B2(n5368), .A(n5547), .ZN(n5701) );
  INV_X1 U3827 ( .A(n5732), .ZN(n5921) );
  INV_X1 U3828 ( .A(n6255), .ZN(n6224) );
  AOI21_X1 U3829 ( .B1(n5696), .B2(n5695), .A(n5694), .ZN(n5697) );
  AND2_X1 U3830 ( .A1(n5736), .A2(n4165), .ZN(n5738) );
  AND2_X1 U3831 ( .A1(n5360), .A2(n6331), .ZN(n6256) );
  INV_X1 U3832 ( .A(n6342), .ZN(n6324) );
  AND2_X1 U3833 ( .A1(n5345), .A2(n4678), .ZN(n6331) );
  INV_X1 U3834 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6571) );
  INV_X1 U3835 ( .A(n4930), .ZN(n4974) );
  INV_X1 U3836 ( .A(n5146), .ZN(n5089) );
  INV_X1 U3837 ( .A(n4664), .ZN(n4451) );
  INV_X1 U3838 ( .A(n4751), .ZN(n4883) );
  INV_X1 U3839 ( .A(n4978), .ZN(n5013) );
  NAND2_X1 U3840 ( .A1(n4628), .A2(n4686), .ZN(n4714) );
  INV_X1 U3841 ( .A(n4460), .ZN(n6441) );
  INV_X1 U3842 ( .A(n4743), .ZN(n4780) );
  INV_X1 U3843 ( .A(n4888), .ZN(n4722) );
  INV_X1 U3844 ( .A(n4499), .ZN(n4533) );
  NAND2_X1 U3845 ( .A1(n4187), .A2(n4186), .ZN(n6601) );
  NOR2_X1 U3846 ( .A1(n5430), .A2(n5429), .ZN(n5434) );
  INV_X1 U3847 ( .A(n6133), .ZN(n6124) );
  NAND2_X1 U3848 ( .A1(n6066), .A2(n5062), .ZN(n6099) );
  INV_X1 U3849 ( .A(n2993), .ZN(n6138) );
  INV_X1 U3850 ( .A(n6079), .ZN(n6145) );
  NAND2_X1 U3851 ( .A1(n5496), .A2(n5672), .ZN(n4049) );
  OR2_X1 U3852 ( .A1(n5639), .A2(n5638), .ZN(n5732) );
  INV_X1 U3853 ( .A(n5674), .ZN(n5669) );
  OR2_X1 U3854 ( .A1(n5630), .A2(n5629), .ZN(n5875) );
  NAND2_X1 U3855 ( .A1(n6196), .A2(n4299), .ZN(n5453) );
  INV_X1 U3856 ( .A(n6160), .ZN(n6187) );
  INV_X1 U3857 ( .A(n6210), .ZN(n4843) );
  NAND2_X1 U3858 ( .A1(n4373), .A2(n4315), .ZN(n6217) );
  INV_X1 U3859 ( .A(n4175), .ZN(n4176) );
  OR2_X1 U3860 ( .A1(n6236), .A2(n4278), .ZN(n6255) );
  XNOR2_X1 U3861 ( .A(n5464), .B(n5479), .ZN(n5478) );
  INV_X1 U3862 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6455) );
  INV_X1 U3863 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5510) );
  AND2_X1 U3864 ( .A1(n4939), .A2(n4938), .ZN(n4977) );
  OR2_X1 U3865 ( .A1(n4889), .A2(n4722), .ZN(n4919) );
  OR2_X1 U3866 ( .A1(n4607), .A2(n4638), .ZN(n6410) );
  NAND2_X1 U3867 ( .A1(n4723), .A2(n4888), .ZN(n4842) );
  OR2_X1 U3868 ( .A1(n4714), .A2(n4638), .ZN(n6450) );
  NOR2_X1 U3869 ( .A1(n4459), .A2(n4458), .ZN(n4497) );
  NAND2_X1 U3870 ( .A1(n4498), .A2(n4722), .ZN(n4782) );
  INV_X1 U3871 ( .A(n4931), .ZN(n4972) );
  NAND2_X1 U3872 ( .A1(n4049), .A2(n4048), .ZN(U2829) );
  INV_X1 U3873 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3025) );
  NAND2_X1 U3874 ( .A1(n3780), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3032)
         );
  INV_X1 U3875 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3026) );
  INV_X1 U3876 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3027) );
  AND2_X2 U3877 ( .A1(n3033), .A2(n3042), .ZN(n3097) );
  NAND2_X1 U3878 ( .A1(n3097), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3031) );
  INV_X1 U3879 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3028) );
  AND2_X2 U3880 ( .A1(n4555), .A2(n3042), .ZN(n3103) );
  NAND2_X1 U3881 ( .A1(n3103), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3030)
         );
  NOR2_X4 U3882 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U3883 ( .A1(n3073), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U3884 ( .A1(n3824), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3885 ( .A1(n3452), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3036)
         );
  NAND2_X1 U3886 ( .A1(n3096), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3035) );
  NAND2_X1 U3887 ( .A1(n3072), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3034) );
  NAND2_X1 U3888 ( .A1(n3089), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3041) );
  NAND2_X1 U3889 ( .A1(n3141), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3040) );
  NAND2_X1 U3890 ( .A1(n3118), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U3891 ( .A1(n3846), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3038) );
  NAND2_X1 U3892 ( .A1(n3123), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3046) );
  NAND2_X1 U3893 ( .A1(n3221), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3045)
         );
  AND2_X2 U3894 ( .A1(n4212), .A2(n4542), .ZN(n3102) );
  NAND2_X1 U3895 ( .A1(n3102), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3044)
         );
  AND2_X2 U3896 ( .A1(n4542), .A2(n4211), .ZN(n3074) );
  NAND2_X1 U3897 ( .A1(n3074), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3043)
         );
  AOI22_X1 U3898 ( .A1(n3452), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U3899 ( .A1(n3824), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3900 ( .A1(n3073), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3901 ( .A1(n3089), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3059) );
  AOI22_X1 U3902 ( .A1(n3123), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U3903 ( .A1(n3141), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3904 ( .A1(n3103), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3905 ( .A1(n3780), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3906 ( .A1(n3824), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3907 ( .A1(n3073), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U3908 ( .A1(n3452), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3062) );
  NAND4_X1 U3909 ( .A1(n3065), .A2(n3064), .A3(n3063), .A4(n3062), .ZN(n3071)
         );
  AOI22_X1 U3910 ( .A1(n3089), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3911 ( .A1(n3141), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U3912 ( .A1(n3103), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3913 ( .A1(n3012), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3066) );
  NAND4_X1 U3914 ( .A1(n3067), .A2(n3068), .A3(n3069), .A4(n3066), .ZN(n3070)
         );
  INV_X1 U3915 ( .A(n3286), .ZN(n3085) );
  AOI22_X1 U3916 ( .A1(n3780), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U3917 ( .A1(n3824), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U3918 ( .A1(n3073), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3076) );
  AOI22_X1 U3919 ( .A1(n3452), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3075) );
  AOI22_X1 U3920 ( .A1(n3089), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3081) );
  AOI22_X1 U3921 ( .A1(n3123), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3080) );
  AOI22_X1 U3922 ( .A1(n3141), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U3923 ( .A1(n3103), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3082) );
  NAND3_X4 U3924 ( .A1(n3084), .A2(n3083), .A3(n3082), .ZN(n5279) );
  AOI22_X1 U3925 ( .A1(n3015), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3094) );
  AOI22_X1 U3926 ( .A1(n3011), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3088) );
  AOI22_X1 U3927 ( .A1(n3073), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3087) );
  AOI22_X1 U3928 ( .A1(n3097), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3093) );
  AOI22_X1 U3929 ( .A1(n3838), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3141), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3092) );
  AOI22_X1 U3930 ( .A1(n3103), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3091) );
  AOI22_X1 U3931 ( .A1(n3221), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3932 ( .A1(n3300), .A2(n4348), .ZN(n3095) );
  AND2_X2 U3933 ( .A1(n3179), .A2(n3095), .ZN(n3113) );
  INV_X1 U3934 ( .A(n3158), .ZN(n3161) );
  AOI22_X1 U3935 ( .A1(n3198), .A2(n3161), .B1(n5279), .B2(n3181), .ZN(n3111)
         );
  INV_X1 U3936 ( .A(n4264), .ZN(n3110) );
  AOI22_X1 U3937 ( .A1(n3452), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3101) );
  AOI22_X1 U3938 ( .A1(n3824), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3100) );
  AOI22_X1 U3939 ( .A1(n3780), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3099) );
  AOI22_X1 U3940 ( .A1(n3089), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U3941 ( .A1(n3141), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3106) );
  AOI22_X1 U3942 ( .A1(n3103), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U3943 ( .A1(n3123), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U3944 ( .A1(n3111), .A2(n3553), .ZN(n3112) );
  NAND2_X2 U3945 ( .A1(n3113), .A2(n3112), .ZN(n3199) );
  NAND2_X1 U3946 ( .A1(n3780), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3117)
         );
  NAND2_X1 U3947 ( .A1(n3097), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U3948 ( .A1(n3824), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3115) );
  NAND2_X1 U3949 ( .A1(n3096), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3114) );
  NAND2_X1 U3950 ( .A1(n3103), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3122)
         );
  NAND2_X1 U3951 ( .A1(n3089), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3121) );
  NAND2_X1 U3952 ( .A1(n3118), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3120) );
  NAND2_X1 U3953 ( .A1(n3102), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3119)
         );
  BUF_X1 U3954 ( .A(n3123), .Z(n3124) );
  NAND2_X1 U3955 ( .A1(n3123), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U3956 ( .A1(n3141), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U3957 ( .A1(n3221), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3126)
         );
  NAND2_X1 U3958 ( .A1(n3846), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U3959 ( .A1(n3452), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3132)
         );
  NAND2_X1 U3960 ( .A1(n3073), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U3961 ( .A1(n3072), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U3962 ( .A1(n3074), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3129)
         );
  NAND4_X4 U3963 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n3926)
         );
  NAND2_X1 U3964 ( .A1(n3780), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U3965 ( .A1(n3097), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U3966 ( .A1(n3073), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U3967 ( .A1(n3096), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3968 ( .A1(n3141), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U3969 ( .A1(n3123), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U3970 ( .A1(n3089), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U3971 ( .A1(n3846), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U3972 ( .A1(n3452), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3149)
         );
  NAND2_X1 U3973 ( .A1(n3103), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3148)
         );
  NAND2_X1 U3974 ( .A1(n3221), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3147)
         );
  NAND2_X1 U3975 ( .A1(n3074), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3146)
         );
  NAND2_X1 U3976 ( .A1(n3824), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U3977 ( .A1(n3118), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U3978 ( .A1(n3072), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U3979 ( .A1(n3102), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3150)
         );
  INV_X1 U3980 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6497) );
  XNOR2_X1 U3981 ( .A(n6497), .B(STATE_REG_1__SCAN_IN), .ZN(n4224) );
  NOR2_X1 U3982 ( .A1(n3926), .A2(n4224), .ZN(n3200) );
  BUF_X4 U3983 ( .A(n3158), .Z(n3196) );
  OAI21_X1 U3984 ( .B1(n3200), .B2(n3196), .A(n4188), .ZN(n3159) );
  NAND2_X1 U3985 ( .A1(n4054), .A2(n3160), .ZN(n3165) );
  NAND2_X1 U3986 ( .A1(n3187), .A2(n4257), .ZN(n3164) );
  NAND2_X1 U3987 ( .A1(n3161), .A2(n3286), .ZN(n3162) );
  NAND2_X1 U3988 ( .A1(n3164), .A2(n3163), .ZN(n3186) );
  NAND2_X1 U3989 ( .A1(n3300), .A2(n4257), .ZN(n3168) );
  INV_X1 U3990 ( .A(n3180), .ZN(n3166) );
  NAND2_X1 U3991 ( .A1(n3166), .A2(n5279), .ZN(n3167) );
  AND2_X2 U3993 ( .A1(n4243), .A2(n5072), .ZN(n6592) );
  NAND2_X4 U3994 ( .A1(n4364), .A2(n3926), .ZN(n3938) );
  NOR2_X1 U3995 ( .A1(n3180), .A2(n3938), .ZN(n4197) );
  AOI21_X2 U3996 ( .B1(n3918), .B2(n6592), .A(n4197), .ZN(n3192) );
  NAND3_X1 U3997 ( .A1(n3185), .A2(n3169), .A3(n3192), .ZN(n3170) );
  NAND2_X1 U3998 ( .A1(n3170), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3173) );
  INV_X1 U3999 ( .A(n3187), .ZN(n3171) );
  NAND2_X2 U4000 ( .A1(n3173), .A2(n3172), .ZN(n3209) );
  NAND2_X1 U4001 ( .A1(n3209), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3177) );
  AND2_X1 U4002 ( .A1(n6571), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3932) );
  INV_X1 U4003 ( .A(n3932), .ZN(n3213) );
  INV_X1 U4004 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n3174) );
  NAND2_X1 U4005 ( .A1(n3174), .A2(n6571), .ZN(n6579) );
  INV_X1 U4006 ( .A(n4156), .ZN(n3214) );
  MUX2_X1 U4007 ( .A(n3213), .B(n3214), .S(n6455), .Z(n3175) );
  INV_X1 U4008 ( .A(n3175), .ZN(n3176) );
  NAND2_X1 U4009 ( .A1(n3553), .A2(n4243), .ZN(n3178) );
  INV_X1 U4010 ( .A(n4364), .ZN(n3935) );
  NAND2_X1 U4011 ( .A1(n3178), .A2(n3935), .ZN(n3184) );
  OR2_X1 U4012 ( .A1(n6579), .A2(n6599), .ZN(n6489) );
  AOI21_X1 U4013 ( .B1(n3179), .B2(n6592), .A(n6489), .ZN(n3183) );
  INV_X1 U4014 ( .A(n3874), .ZN(n4152) );
  NAND2_X1 U4015 ( .A1(n4188), .A2(n4246), .ZN(n3182) );
  NAND2_X1 U4016 ( .A1(n4263), .A2(n3182), .ZN(n4205) );
  INV_X1 U4017 ( .A(n3186), .ZN(n3189) );
  OR2_X1 U4018 ( .A1(n3187), .A2(n4257), .ZN(n3188) );
  NAND2_X1 U4019 ( .A1(n3189), .A2(n3188), .ZN(n3193) );
  NAND2_X1 U4020 ( .A1(n3193), .A2(n3926), .ZN(n3190) );
  NAND4_X1 U4021 ( .A1(n3192), .A2(n3191), .A3(n3185), .A4(n3190), .ZN(n3261)
         );
  INV_X1 U4022 ( .A(n3193), .ZN(n3195) );
  NAND2_X1 U4023 ( .A1(n3195), .A2(n3194), .ZN(n4195) );
  NOR2_X1 U4024 ( .A1(n4364), .A2(n3196), .ZN(n3197) );
  AND2_X1 U4025 ( .A1(n3197), .A2(n4246), .ZN(n3928) );
  NOR2_X2 U4026 ( .A1(n3199), .A2(n4263), .ZN(n3924) );
  NAND2_X1 U4027 ( .A1(n3924), .A2(n4243), .ZN(n4193) );
  OAI211_X1 U4028 ( .C1(n5522), .C2(n3200), .A(n4273), .B(n4193), .ZN(n3201)
         );
  NAND2_X1 U4029 ( .A1(n3201), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3207) );
  INV_X1 U4030 ( .A(n3207), .ZN(n3204) );
  XNOR2_X1 U4031 ( .A(n6461), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6350)
         );
  NAND2_X1 U4032 ( .A1(n3214), .A2(n6350), .ZN(n3203) );
  NAND2_X1 U4033 ( .A1(n3213), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4034 ( .A1(n3203), .A2(n3202), .ZN(n3205) );
  NAND2_X1 U4035 ( .A1(n3264), .A2(n3232), .ZN(n3208) );
  AOI21_X1 U4036 ( .B1(n3209), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3205), 
        .ZN(n3206) );
  NAND2_X1 U4037 ( .A1(n3207), .A2(n3206), .ZN(n3231) );
  NAND2_X1 U4038 ( .A1(n3208), .A2(n3231), .ZN(n3315) );
  NAND2_X1 U4039 ( .A1(n3209), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3216) );
  AND2_X1 U4040 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4041 ( .A1(n3210), .A2(n4716), .ZN(n4633) );
  INV_X1 U4042 ( .A(n3210), .ZN(n3211) );
  NAND2_X1 U4043 ( .A1(n3211), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4044 ( .A1(n4633), .A2(n3212), .ZN(n4423) );
  AOI22_X1 U4045 ( .A1(n3214), .A2(n4423), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3213), .ZN(n3215) );
  XNOR2_X1 U4046 ( .A(n3315), .B(n3316), .ZN(n4329) );
  AOI22_X1 U4047 ( .A1(n3006), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4048 ( .A1(n3013), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4049 ( .A1(n3823), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4050 ( .A1(n3848), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3217) );
  NAND4_X1 U4051 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3227)
         );
  AOI22_X1 U4052 ( .A1(n3818), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3225) );
  AOI22_X1 U4053 ( .A1(n3837), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4054 ( .A1(n3735), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3223) );
  BUF_X1 U4055 ( .A(n3846), .Z(n3782) );
  AOI22_X1 U4056 ( .A1(n3840), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3222) );
  NAND4_X1 U4057 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3226)
         );
  INV_X1 U4058 ( .A(n4069), .ZN(n4078) );
  NOR2_X1 U4059 ( .A1(n4123), .A2(n4078), .ZN(n3228) );
  INV_X1 U4060 ( .A(n3323), .ZN(n3256) );
  AOI22_X1 U4061 ( .A1(n3903), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3256), 
        .B2(n4069), .ZN(n3229) );
  NAND2_X1 U4062 ( .A1(n3232), .A2(n3231), .ZN(n3233) );
  AOI22_X1 U4063 ( .A1(n3848), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4064 ( .A1(n3818), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4065 ( .A1(n3006), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4066 ( .A1(n3823), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3234) );
  NAND4_X1 U4067 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3243)
         );
  AOI22_X1 U4068 ( .A1(n3013), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4070 ( .A1(n3781), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4071 ( .A1(n3847), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4072 ( .A1(n3840), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3238) );
  NAND4_X1 U4073 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3242)
         );
  INV_X1 U4074 ( .A(n4067), .ZN(n3244) );
  NOR2_X1 U4075 ( .A1(n4123), .A2(n3244), .ZN(n3245) );
  AOI21_X2 U4076 ( .B1(n4191), .B2(n6599), .A(n3245), .ZN(n3289) );
  INV_X1 U4077 ( .A(n3289), .ZN(n3283) );
  NAND2_X1 U4078 ( .A1(n3903), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4079 ( .A1(n3007), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4080 ( .A1(n3800), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4081 ( .A1(n3837), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4082 ( .A1(n3840), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4083 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3255)
         );
  AOI22_X1 U4084 ( .A1(n3735), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4085 ( .A1(n3013), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4086 ( .A1(n3452), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4087 ( .A1(n3847), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3250) );
  NAND4_X1 U4088 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3254)
         );
  OR2_X1 U4089 ( .A1(n4123), .A2(n4121), .ZN(n3258) );
  NAND2_X1 U4090 ( .A1(n3256), .A2(n4067), .ZN(n3257) );
  INV_X1 U4091 ( .A(n3260), .ZN(n3263) );
  INV_X1 U4092 ( .A(n3261), .ZN(n3262) );
  NAND2_X1 U4093 ( .A1(n3265), .A2(n3264), .ZN(n3301) );
  INV_X1 U4094 ( .A(n3903), .ZN(n3888) );
  INV_X1 U4095 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4953) );
  AOI21_X1 U4096 ( .B1(n4257), .B2(n4121), .A(n6599), .ZN(n3277) );
  AOI22_X1 U4097 ( .A1(n3013), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4098 ( .A1(n3735), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4099 ( .A1(n3847), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4100 ( .A1(n3837), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3266) );
  NAND4_X1 U4101 ( .A1(n3269), .A2(n3268), .A3(n3267), .A4(n3266), .ZN(n3275)
         );
  AOI22_X1 U4102 ( .A1(n3006), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4103 ( .A1(n3800), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4104 ( .A1(n3840), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4105 ( .A1(n3730), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3270) );
  NAND4_X1 U4106 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3274)
         );
  NAND2_X1 U4107 ( .A1(n4059), .A2(n4068), .ZN(n3276) );
  OAI211_X1 U4108 ( .C1(n3888), .C2(n4953), .A(n3277), .B(n3276), .ZN(n3297)
         );
  XNOR2_X1 U4109 ( .A(n4068), .B(n4121), .ZN(n3278) );
  NOR2_X1 U4110 ( .A1(n3278), .A2(n4123), .ZN(n3296) );
  NAND2_X1 U4111 ( .A1(n3297), .A2(n3296), .ZN(n3279) );
  INV_X1 U4112 ( .A(n4121), .ZN(n4127) );
  OR2_X1 U4113 ( .A1(n4123), .A2(n4127), .ZN(n3281) );
  NOR2_X2 U4114 ( .A1(n4353), .A2(n4987), .ZN(n3724) );
  NAND2_X1 U4115 ( .A1(n4321), .A2(n3724), .ZN(n3287) );
  NAND2_X1 U4116 ( .A1(n4987), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3561) );
  NAND2_X1 U4117 ( .A1(n3287), .A2(n3561), .ZN(n4302) );
  NAND2_X1 U4118 ( .A1(n4322), .A2(n3724), .ZN(n3295) );
  OR2_X1 U4119 ( .A1(n5279), .A2(n4987), .ZN(n3417) );
  INV_X2 U4120 ( .A(n3417), .ZN(n5446) );
  AOI22_X1 U4121 ( .A1(n5446), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4987), .ZN(n3293) );
  AND2_X1 U4122 ( .A1(n3198), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4123 ( .A1(n3305), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3292) );
  AND2_X1 U4124 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  NAND2_X1 U4125 ( .A1(n3295), .A2(n3294), .ZN(n4286) );
  OR2_X1 U4126 ( .A1(n3297), .A2(n3296), .ZN(n3298) );
  NAND2_X2 U4127 ( .A1(n3299), .A2(n3298), .ZN(n4324) );
  AOI21_X1 U4128 ( .B1(n4324), .B2(n3300), .A(n4987), .ZN(n4239) );
  INV_X1 U4129 ( .A(n3305), .ZN(n3363) );
  BUF_X1 U4130 ( .A(n3301), .Z(n4328) );
  INV_X1 U4131 ( .A(n3724), .ZN(n3495) );
  OR2_X1 U4132 ( .A1(n4328), .A2(n3495), .ZN(n3303) );
  AOI22_X1 U4133 ( .A1(n5446), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4987), .ZN(n3302) );
  OAI211_X1 U4134 ( .C1(n3363), .C2(n3304), .A(n3303), .B(n3302), .ZN(n4240)
         );
  MUX2_X1 U4135 ( .A(n5055), .B(n4239), .S(n4240), .Z(n4285) );
  NAND2_X1 U4136 ( .A1(n3305), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3310) );
  INV_X1 U4137 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3307) );
  OAI21_X1 U4138 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3342), .ZN(n6254) );
  NAND2_X1 U4139 ( .A1(n5055), .A2(n6254), .ZN(n3306) );
  OAI21_X1 U4140 ( .B1(n3561), .B2(n3307), .A(n3306), .ZN(n3308) );
  AOI21_X1 U4141 ( .B1(n5446), .B2(EAX_REG_2__SCAN_IN), .A(n3308), .ZN(n3309)
         );
  AND2_X1 U4142 ( .A1(n3310), .A2(n3309), .ZN(n3312) );
  NOR2_X1 U4143 ( .A1(n4284), .A2(n3312), .ZN(n3311) );
  OR2_X1 U4144 ( .A1(n4302), .A2(n3311), .ZN(n3313) );
  NAND2_X1 U4145 ( .A1(n4284), .A2(n3312), .ZN(n4303) );
  NAND2_X1 U4146 ( .A1(n3339), .A2(n3338), .ZN(n3334) );
  INV_X1 U4147 ( .A(n3315), .ZN(n3317) );
  NAND2_X1 U4148 ( .A1(n3209), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3322) );
  NAND3_X1 U4149 ( .A1(n6466), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6349) );
  INV_X1 U4150 ( .A(n6349), .ZN(n3318) );
  NAND2_X1 U4151 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3318), .ZN(n4605) );
  NAND2_X1 U4152 ( .A1(n6466), .A2(n4605), .ZN(n3319) );
  NOR3_X1 U4153 ( .A1(n6466), .A2(n4716), .A3(n6461), .ZN(n4501) );
  NAND2_X1 U4154 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4501), .ZN(n4368) );
  NAND2_X1 U4155 ( .A1(n3319), .A2(n4368), .ZN(n4457) );
  OAI22_X1 U4156 ( .A1(n4156), .A2(n4457), .B1(n3932), .B2(n6466), .ZN(n3320)
         );
  INV_X1 U4157 ( .A(n3320), .ZN(n3321) );
  AOI22_X1 U4158 ( .A1(n3818), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4159 ( .A1(n3013), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4160 ( .A1(n3837), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4161 ( .A1(n3775), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3324) );
  NAND4_X1 U4162 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3333)
         );
  INV_X1 U4163 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U4164 ( .A1(n3840), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4165 ( .A1(n3823), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4166 ( .A1(n3735), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4167 ( .A1(n3848), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3328) );
  NAND4_X1 U4168 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3332)
         );
  OR2_X1 U4169 ( .A1(n3333), .A2(n3332), .ZN(n4087) );
  AOI22_X1 U4170 ( .A1(n3911), .A2(n4087), .B1(n3903), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3335) );
  AND2_X1 U4171 ( .A1(n3336), .A2(n3335), .ZN(n4454) );
  NAND2_X1 U4172 ( .A1(n3334), .A2(n4454), .ZN(n3340) );
  NAND3_X2 U4173 ( .A1(n3339), .A2(n3338), .A3(n3337), .ZN(n3369) );
  INV_X1 U4174 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4558) );
  INV_X1 U4175 ( .A(n3342), .ZN(n3341) );
  INV_X1 U4176 ( .A(n3364), .ZN(n3345) );
  INV_X1 U4177 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4178 ( .A1(n3343), .A2(n3342), .ZN(n3344) );
  NAND2_X1 U4179 ( .A1(n3345), .A2(n3344), .ZN(n5149) );
  INV_X1 U4180 ( .A(n3561), .ZN(n5445) );
  AOI22_X1 U4181 ( .A1(n5149), .A2(n5055), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4182 ( .A1(n5446), .A2(EAX_REG_3__SCAN_IN), .ZN(n3346) );
  OAI211_X1 U4183 ( .C1(n3363), .C2(n4558), .A(n3347), .B(n3346), .ZN(n3348)
         );
  NOR2_X1 U4184 ( .A1(n4310), .A2(n4309), .ZN(n4404) );
  AOI22_X1 U4185 ( .A1(n3007), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4186 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3013), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4187 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3823), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4188 ( .A1(n3848), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3349) );
  NAND4_X1 U4189 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3358)
         );
  AOI22_X1 U4190 ( .A1(n3818), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4191 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3837), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4192 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3735), .B1(n3847), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4193 ( .A1(n3840), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3353) );
  NAND4_X1 U4194 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3357)
         );
  NAND2_X1 U4195 ( .A1(n3911), .A2(n4104), .ZN(n3360) );
  NAND2_X1 U4196 ( .A1(n3903), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4197 ( .A1(n3360), .A2(n3359), .ZN(n3390) );
  XNOR2_X1 U4198 ( .A(n3369), .B(n3390), .ZN(n4086) );
  NAND2_X1 U4199 ( .A1(n4086), .A2(n3724), .ZN(n3368) );
  INV_X1 U4200 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3902) );
  NAND2_X1 U4201 ( .A1(n4987), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3362)
         );
  NAND2_X1 U4202 ( .A1(n5446), .A2(EAX_REG_4__SCAN_IN), .ZN(n3361) );
  OAI211_X1 U4203 ( .C1(n3363), .C2(n3902), .A(n3362), .B(n3361), .ZN(n3366)
         );
  INV_X1 U4204 ( .A(n5055), .ZN(n3860) );
  OAI21_X1 U4205 ( .B1(n3364), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3384), 
        .ZN(n6244) );
  AND2_X1 U4206 ( .A1(n6244), .A2(n5055), .ZN(n3365) );
  AOI21_X1 U4207 ( .B1(n3366), .B2(n3860), .A(n3365), .ZN(n3367) );
  NAND2_X1 U4208 ( .A1(n3368), .A2(n3367), .ZN(n4403) );
  NAND2_X1 U4209 ( .A1(n4404), .A2(n4403), .ZN(n4402) );
  NAND2_X1 U4210 ( .A1(n3392), .A2(n3390), .ZN(n3383) );
  AOI22_X1 U4211 ( .A1(n3006), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4212 ( .A1(n3013), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4213 ( .A1(n3823), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3372) );
  INV_X1 U4214 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4215 ( .A1(n3848), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4216 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3380)
         );
  AOI22_X1 U4217 ( .A1(n3818), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4218 ( .A1(n3837), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4219 ( .A1(n3735), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4220 ( .A1(n3840), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4221 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3379)
         );
  OR2_X1 U4222 ( .A1(n3380), .A2(n3379), .ZN(n4103) );
  NAND2_X1 U4223 ( .A1(n3911), .A2(n4103), .ZN(n3382) );
  NAND2_X1 U4224 ( .A1(n3903), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4225 ( .A1(n3382), .A2(n3381), .ZN(n3389) );
  INV_X1 U4226 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4861) );
  AND2_X1 U4227 ( .A1(n3384), .A2(n5076), .ZN(n3385) );
  OR2_X1 U4228 ( .A1(n3385), .A2(n3405), .ZN(n5068) );
  NOR2_X1 U4229 ( .A1(n3561), .A2(n5076), .ZN(n3386) );
  AOI21_X1 U4230 ( .B1(n5068), .B2(n5055), .A(n3386), .ZN(n3387) );
  OAI21_X1 U4231 ( .B1(n3417), .B2(n4861), .A(n3387), .ZN(n3388) );
  OR2_X2 U4232 ( .A1(n4402), .A2(n4414), .ZN(n4620) );
  AOI22_X1 U4233 ( .A1(n3007), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4234 ( .A1(n3013), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4235 ( .A1(n3823), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4236 ( .A1(n3848), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3393) );
  NAND4_X1 U4237 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3402)
         );
  AOI22_X1 U4238 ( .A1(n3818), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4239 ( .A1(n3837), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4240 ( .A1(n3735), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4241 ( .A1(n3840), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4242 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  OR2_X1 U4243 ( .A1(n3402), .A2(n3401), .ZN(n4114) );
  NAND2_X1 U4244 ( .A1(n3911), .A2(n4114), .ZN(n3404) );
  NAND2_X1 U4245 ( .A1(n3903), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4246 ( .A1(n3411), .A2(n3410), .ZN(n4102) );
  NOR2_X1 U4247 ( .A1(n3405), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3406)
         );
  OR2_X1 U4248 ( .A1(n3430), .A2(n3406), .ZN(n6235) );
  INV_X1 U4249 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4849) );
  INV_X1 U4250 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3407) );
  OAI22_X1 U4251 ( .A1(n3417), .A2(n4849), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3407), .ZN(n3408) );
  MUX2_X1 U4252 ( .A(n6235), .B(n3408), .S(n3860), .Z(n3409) );
  INV_X1 U4253 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U4254 ( .A1(n3911), .A2(n4121), .ZN(n3412) );
  OAI21_X1 U4255 ( .B1(n4957), .B2(n3888), .A(n3412), .ZN(n3413) );
  INV_X1 U4256 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3416) );
  XNOR2_X1 U4257 ( .A(n3430), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U4258 ( .A1(n5198), .A2(n5055), .ZN(n3415) );
  NAND2_X1 U4259 ( .A1(n5445), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3414)
         );
  OAI211_X1 U4260 ( .C1(n3417), .C2(n3416), .A(n3415), .B(n3414), .ZN(n3418)
         );
  AND2_X2 U4261 ( .A1(n4618), .A2(n3419), .ZN(n4872) );
  AOI22_X1 U4262 ( .A1(n3007), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3013), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4263 ( .A1(n3730), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4264 ( .A1(n3452), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4265 ( .A1(n3837), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3420) );
  NAND4_X1 U4266 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3429)
         );
  AOI22_X1 U4267 ( .A1(n3818), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4268 ( .A1(n3840), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4269 ( .A1(n2994), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4270 ( .A1(n3735), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4271 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3428)
         );
  OAI21_X1 U4272 ( .B1(n3429), .B2(n3428), .A(n3724), .ZN(n3434) );
  NAND2_X1 U4273 ( .A1(n5446), .A2(EAX_REG_8__SCAN_IN), .ZN(n3433) );
  INV_X1 U4274 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U4275 ( .A(n3435), .B(n5405), .ZN(n6103) );
  OR2_X1 U4276 ( .A1(n6103), .A2(n3860), .ZN(n3432) );
  NAND2_X1 U4277 ( .A1(n5445), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3431)
         );
  NAND4_X1 U4278 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(n4871)
         );
  NAND2_X1 U4279 ( .A1(n4872), .A2(n4871), .ZN(n4870) );
  INV_X1 U4280 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6757) );
  AOI21_X1 U4281 ( .B1(n6757), .B2(n3436), .A(n3467), .ZN(n6088) );
  OR2_X1 U4282 ( .A1(n6088), .A2(n3860), .ZN(n3451) );
  AOI22_X1 U4283 ( .A1(n3840), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4284 ( .A1(n3730), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4285 ( .A1(n3837), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4286 ( .A1(n3848), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4287 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3446)
         );
  AOI22_X1 U4288 ( .A1(n3007), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4289 ( .A1(n3013), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4290 ( .A1(n3735), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4291 ( .A1(n3818), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4292 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  OAI21_X1 U4293 ( .B1(n3446), .B2(n3445), .A(n3724), .ZN(n3449) );
  NAND2_X1 U4294 ( .A1(n5446), .A2(EAX_REG_9__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4295 ( .A1(n5445), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3447)
         );
  AND3_X1 U4296 ( .A1(n3449), .A2(n3448), .A3(n3447), .ZN(n3450) );
  AND2_X1 U4297 ( .A1(n3451), .A2(n3450), .ZN(n5033) );
  NOR2_X1 U4298 ( .A1(n4870), .A2(n5033), .ZN(n5030) );
  INV_X1 U4299 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U4300 ( .A(n3467), .B(n5217), .ZN(n6074) );
  OR2_X1 U4301 ( .A1(n6074), .A2(n3860), .ZN(n3465) );
  AOI22_X1 U4302 ( .A1(n5446), .A2(EAX_REG_10__SCAN_IN), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4303 ( .A1(n3007), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4304 ( .A1(n3848), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4305 ( .A1(n3840), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4306 ( .A1(n3759), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4307 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3462)
         );
  AOI22_X1 U4308 ( .A1(n3013), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4309 ( .A1(n3735), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4310 ( .A1(n3775), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4311 ( .A1(n3837), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3457) );
  NAND4_X1 U4312 ( .A1(n3460), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(n3461)
         );
  OAI21_X1 U4313 ( .B1(n3462), .B2(n3461), .A(n3724), .ZN(n3463) );
  AND3_X1 U4314 ( .A1(n3465), .A2(n3464), .A3(n3463), .ZN(n5179) );
  AND2_X2 U4315 ( .A1(n5030), .A2(n3466), .ZN(n5181) );
  INV_X1 U4316 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3491) );
  XOR2_X1 U4317 ( .A(n3491), .B(n3492), .Z(n6223) );
  AOI22_X1 U4318 ( .A1(n3848), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4319 ( .A1(n3818), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4320 ( .A1(n2994), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4321 ( .A1(n3735), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4322 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3477)
         );
  AOI22_X1 U4323 ( .A1(n3006), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3013), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4324 ( .A1(n3837), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4325 ( .A1(n3730), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4326 ( .A1(n3840), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4327 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3476)
         );
  OR2_X1 U4328 ( .A1(n3477), .A2(n3476), .ZN(n3478) );
  AOI22_X1 U4329 ( .A1(n3724), .A2(n3478), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4330 ( .A1(n5446), .A2(EAX_REG_11__SCAN_IN), .ZN(n3479) );
  OAI211_X1 U4331 ( .C1(n6223), .C2(n3860), .A(n3480), .B(n3479), .ZN(n5221)
         );
  AND2_X2 U4332 ( .A1(n5181), .A2(n5221), .ZN(n5229) );
  AOI22_X1 U4333 ( .A1(n3007), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4334 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3759), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4335 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3840), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4336 ( .A1(n3847), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4337 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3490)
         );
  AOI22_X1 U4338 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3013), .B1(n2994), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4339 ( .A1(n3735), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4340 ( .A1(n3730), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4341 ( .A1(n3837), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3485) );
  NAND4_X1 U4342 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), .ZN(n3489)
         );
  NOR2_X1 U4343 ( .A1(n3490), .A2(n3489), .ZN(n3496) );
  XNOR2_X1 U4344 ( .A(n3497), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5250)
         );
  NAND2_X1 U4345 ( .A1(n5250), .A2(n5055), .ZN(n3494) );
  AOI22_X1 U4346 ( .A1(n5446), .A2(EAX_REG_12__SCAN_IN), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3493) );
  OAI211_X1 U4347 ( .C1(n3496), .C2(n3495), .A(n3494), .B(n3493), .ZN(n5230)
         );
  INV_X1 U4348 ( .A(n5230), .ZN(n3505) );
  INV_X1 U4350 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3500) );
  OAI21_X1 U4351 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3498), .A(n3712), 
        .ZN(n6056) );
  NAND2_X1 U4352 ( .A1(n6056), .A2(n5055), .ZN(n3499) );
  OAI21_X1 U4353 ( .B1(n3500), .B2(n3561), .A(n3499), .ZN(n3501) );
  AOI21_X1 U4354 ( .B1(n5446), .B2(EAX_REG_13__SCAN_IN), .A(n3501), .ZN(n3507)
         );
  INV_X1 U4355 ( .A(n3507), .ZN(n3502) );
  NAND2_X2 U4356 ( .A1(n3503), .A2(n3502), .ZN(n3521) );
  INV_X1 U4357 ( .A(n3521), .ZN(n3504) );
  NOR2_X1 U4358 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U4359 ( .A1(n5229), .A2(n3506), .ZN(n3509) );
  AOI22_X1 U4360 ( .A1(n3006), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4361 ( .A1(n3013), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4362 ( .A1(n3800), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4363 ( .A1(n3735), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3510) );
  NAND4_X1 U4364 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3519)
         );
  AOI22_X1 U4365 ( .A1(n3759), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4366 ( .A1(n3840), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4367 ( .A1(n3848), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4368 ( .A1(n3781), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U4369 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3518)
         );
  OR2_X1 U4370 ( .A1(n3519), .A2(n3518), .ZN(n3520) );
  NAND2_X1 U4371 ( .A1(n3724), .A2(n3520), .ZN(n5255) );
  OR2_X2 U4372 ( .A1(n5256), .A2(n5255), .ZN(n5258) );
  NAND2_X2 U4373 ( .A1(n5258), .A2(n3521), .ZN(n5265) );
  AOI22_X1 U4374 ( .A1(n3013), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4375 ( .A1(n3848), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4376 ( .A1(n3735), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4377 ( .A1(n3759), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3522) );
  NAND4_X1 U4378 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3531)
         );
  AOI22_X1 U4379 ( .A1(n2994), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4380 ( .A1(n3840), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4381 ( .A1(n3775), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4382 ( .A1(n3837), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4383 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3530)
         );
  NOR2_X1 U4384 ( .A1(n3531), .A2(n3530), .ZN(n3703) );
  AOI22_X1 U4385 ( .A1(n3759), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4386 ( .A1(n3007), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4387 ( .A1(n3848), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4388 ( .A1(n3221), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3532) );
  NAND4_X1 U4389 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3541)
         );
  AOI22_X1 U4390 ( .A1(n3013), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4391 ( .A1(n3840), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4392 ( .A1(n3730), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4393 ( .A1(n3103), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4394 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3540)
         );
  NOR2_X1 U4395 ( .A1(n3541), .A2(n3540), .ZN(n3702) );
  NOR2_X1 U4396 ( .A1(n3703), .A2(n3702), .ZN(n3743) );
  AOI22_X1 U4397 ( .A1(n3007), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4398 ( .A1(n3013), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4399 ( .A1(n3800), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4400 ( .A1(n3848), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3542) );
  NAND4_X1 U4401 ( .A1(n3545), .A2(n3544), .A3(n3543), .A4(n3542), .ZN(n3551)
         );
  AOI22_X1 U4402 ( .A1(n3759), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4403 ( .A1(n3837), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4404 ( .A1(n3103), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4405 ( .A1(n3840), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3546) );
  NAND4_X1 U4406 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3550)
         );
  OR2_X1 U4407 ( .A1(n3551), .A2(n3550), .ZN(n3742) );
  INV_X1 U4408 ( .A(n3742), .ZN(n3552) );
  XNOR2_X1 U4409 ( .A(n3743), .B(n3552), .ZN(n3555) );
  NAND2_X1 U4410 ( .A1(n3554), .A2(n3196), .ZN(n6452) );
  INV_X1 U4411 ( .A(n3863), .ZN(n3831) );
  NAND2_X1 U4412 ( .A1(n3555), .A2(n3831), .ZN(n3564) );
  INV_X1 U4413 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5571) );
  INV_X1 U4414 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6038) );
  INV_X1 U4415 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U4416 ( .A1(n3652), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3635)
         );
  INV_X1 U4417 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5586) );
  INV_X1 U4418 ( .A(n3707), .ZN(n3557) );
  AOI21_X1 U4419 ( .B1(n3557), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4420 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3558) );
  OR2_X1 U4421 ( .A1(n3559), .A2(n3748), .ZN(n5570) );
  NAND2_X1 U4422 ( .A1(n5570), .A2(n5055), .ZN(n3560) );
  OAI21_X1 U4423 ( .B1(n5571), .B2(n3561), .A(n3560), .ZN(n3562) );
  AOI21_X1 U4424 ( .B1(n5446), .B2(EAX_REG_24__SCAN_IN), .A(n3562), .ZN(n3563)
         );
  NAND2_X1 U4425 ( .A1(n3564), .A2(n3563), .ZN(n4171) );
  INV_X1 U4426 ( .A(n4171), .ZN(n3711) );
  AOI22_X1 U4427 ( .A1(n3006), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4428 ( .A1(n3800), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4429 ( .A1(n3759), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4430 ( .A1(n3840), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3565) );
  NAND4_X1 U4431 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n3574)
         );
  AOI22_X1 U4432 ( .A1(n3735), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4433 ( .A1(n3013), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4434 ( .A1(n3848), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4435 ( .A1(n3847), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3569) );
  NAND4_X1 U4436 ( .A1(n3572), .A2(n3571), .A3(n3570), .A4(n3569), .ZN(n3573)
         );
  NOR2_X1 U4437 ( .A1(n3574), .A2(n3573), .ZN(n3577) );
  INV_X1 U4438 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5894) );
  OAI21_X1 U4439 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5894), .A(n3860), .ZN(
        n3575) );
  AOI21_X1 U4440 ( .B1(n5446), .B2(EAX_REG_21__SCAN_IN), .A(n3575), .ZN(n3576)
         );
  OAI21_X1 U4441 ( .B1(n3863), .B2(n3577), .A(n3576), .ZN(n3579) );
  XNOR2_X1 U4442 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3593), .ZN(n5898)
         );
  NAND2_X1 U4443 ( .A1(n5055), .A2(n5898), .ZN(n3578) );
  NAND2_X1 U4444 ( .A1(n3579), .A2(n3578), .ZN(n5646) );
  INV_X1 U4445 ( .A(n5646), .ZN(n3668) );
  AOI22_X1 U4446 ( .A1(n3007), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4447 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3735), .B1(n3759), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4448 ( .A1(n3848), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4449 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3840), .B1(n3839), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3580) );
  NAND4_X1 U4450 ( .A1(n3583), .A2(n3582), .A3(n3581), .A4(n3580), .ZN(n3589)
         );
  AOI22_X1 U4451 ( .A1(n3013), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4452 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3781), .B1(n3847), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4453 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3837), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4454 ( .A1(n3775), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3584) );
  NAND4_X1 U4455 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3588)
         );
  NOR2_X1 U4456 ( .A1(n3589), .A2(n3588), .ZN(n3590) );
  OR2_X1 U4457 ( .A1(n3863), .A2(n3590), .ZN(n3597) );
  INV_X1 U4458 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6593) );
  OAI21_X1 U4459 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6593), .A(n4987), 
        .ZN(n3591) );
  INV_X1 U4460 ( .A(n3591), .ZN(n3592) );
  AOI21_X1 U4461 ( .B1(n5446), .B2(EAX_REG_20__SCAN_IN), .A(n3592), .ZN(n3596)
         );
  OAI21_X1 U4462 ( .B1(n3594), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3593), 
        .ZN(n5902) );
  NOR2_X1 U4463 ( .A1(n5902), .A2(n3860), .ZN(n3595) );
  AOI21_X1 U4464 ( .B1(n3597), .B2(n3596), .A(n3595), .ZN(n5394) );
  AOI22_X1 U4465 ( .A1(n3007), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3013), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4466 ( .A1(n3730), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4467 ( .A1(n3735), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4468 ( .A1(n3848), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3598) );
  NAND4_X1 U4469 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3607)
         );
  AOI22_X1 U4470 ( .A1(n3837), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4471 ( .A1(n2994), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4472 ( .A1(n3818), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4473 ( .A1(n3840), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3602) );
  NAND4_X1 U4474 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3606)
         );
  NOR2_X1 U4475 ( .A1(n3607), .A2(n3606), .ZN(n3610) );
  INV_X1 U4476 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5313) );
  OAI21_X1 U4477 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5313), .A(n3860), .ZN(
        n3608) );
  AOI21_X1 U4478 ( .B1(n5446), .B2(EAX_REG_19__SCAN_IN), .A(n3608), .ZN(n3609)
         );
  OAI21_X1 U4479 ( .B1(n3863), .B2(n3610), .A(n3609), .ZN(n3612) );
  XNOR2_X1 U4480 ( .A(n3627), .B(n5313), .ZN(n5315) );
  NAND2_X1 U4481 ( .A1(n5315), .A2(n5055), .ZN(n3611) );
  NAND2_X1 U4482 ( .A1(n3612), .A2(n3611), .ZN(n4050) );
  AOI22_X1 U4483 ( .A1(n3013), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4484 ( .A1(n3848), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4485 ( .A1(n3840), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4486 ( .A1(n3781), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4487 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3622)
         );
  AOI22_X1 U4488 ( .A1(n3735), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4489 ( .A1(n3006), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4490 ( .A1(n3837), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4491 ( .A1(n3823), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4492 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3621)
         );
  NOR2_X1 U4493 ( .A1(n3622), .A2(n3621), .ZN(n3626) );
  OAI21_X1 U4494 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6593), .A(n4987), 
        .ZN(n3623) );
  INV_X1 U4495 ( .A(n3623), .ZN(n3624) );
  AOI21_X1 U4496 ( .B1(n5446), .B2(EAX_REG_18__SCAN_IN), .A(n3624), .ZN(n3625)
         );
  OAI21_X1 U4497 ( .B1(n3863), .B2(n3626), .A(n3625), .ZN(n3634) );
  INV_X1 U4498 ( .A(n3627), .ZN(n3632) );
  INV_X1 U4499 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3630) );
  INV_X1 U4500 ( .A(n3628), .ZN(n3629) );
  NAND2_X1 U4501 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  NAND2_X1 U4502 ( .A1(n3632), .A2(n3631), .ZN(n6023) );
  OR2_X1 U4503 ( .A1(n6023), .A2(n3860), .ZN(n3633) );
  NAND2_X1 U4504 ( .A1(n3634), .A2(n3633), .ZN(n5653) );
  OR2_X1 U4505 ( .A1(n4050), .A2(n5653), .ZN(n3651) );
  XNOR2_X1 U4506 ( .A(n3635), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5938)
         );
  NAND2_X1 U4507 ( .A1(n5938), .A2(n5055), .ZN(n3650) );
  AOI22_X1 U4508 ( .A1(n3007), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4509 ( .A1(n3013), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4510 ( .A1(n3823), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4511 ( .A1(n3848), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3636) );
  NAND4_X1 U4512 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3645)
         );
  AOI22_X1 U4513 ( .A1(n3818), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4514 ( .A1(n3837), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4515 ( .A1(n3735), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4516 ( .A1(n3840), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3640) );
  NAND4_X1 U4517 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3644)
         );
  NOR2_X1 U4518 ( .A1(n3645), .A2(n3644), .ZN(n3648) );
  AOI21_X1 U4519 ( .B1(n5586), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3646) );
  AOI21_X1 U4520 ( .B1(n5446), .B2(EAX_REG_17__SCAN_IN), .A(n3646), .ZN(n3647)
         );
  OAI21_X1 U4521 ( .B1(n3863), .B2(n3648), .A(n3647), .ZN(n3649) );
  NAND2_X1 U4522 ( .A1(n3650), .A2(n3649), .ZN(n5579) );
  NOR2_X1 U4523 ( .A1(n3651), .A2(n5579), .ZN(n3667) );
  XOR2_X1 U4524 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3652), .Z(n6031) );
  AOI22_X1 U4525 ( .A1(n3013), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4526 ( .A1(n3818), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4527 ( .A1(n3837), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4528 ( .A1(n3823), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4529 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3662)
         );
  AOI22_X1 U4530 ( .A1(n3006), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4531 ( .A1(n3848), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4532 ( .A1(n3735), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4533 ( .A1(n3840), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3657) );
  NAND4_X1 U4534 ( .A1(n3660), .A2(n3659), .A3(n3658), .A4(n3657), .ZN(n3661)
         );
  NOR2_X1 U4535 ( .A1(n3662), .A2(n3661), .ZN(n3664) );
  AOI22_X1 U4536 ( .A1(n5446), .A2(EAX_REG_16__SCAN_IN), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3663) );
  OAI21_X1 U4537 ( .B1(n3863), .B2(n3664), .A(n3663), .ZN(n3665) );
  INV_X1 U4538 ( .A(n3665), .ZN(n3666) );
  OAI21_X1 U4539 ( .B1(n6031), .B2(n3860), .A(n3666), .ZN(n5327) );
  AND2_X1 U4540 ( .A1(n3667), .A2(n5327), .ZN(n4052) );
  AND2_X1 U4541 ( .A1(n5394), .A2(n4052), .ZN(n5393) );
  NAND2_X1 U4542 ( .A1(n3668), .A2(n5393), .ZN(n3684) );
  XNOR2_X1 U4543 ( .A(n3669), .B(n5601), .ZN(n5748) );
  AOI22_X1 U4544 ( .A1(n3006), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4545 ( .A1(n3452), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4546 ( .A1(n3730), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4547 ( .A1(n3221), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4548 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3679)
         );
  AOI22_X1 U4549 ( .A1(n3759), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4550 ( .A1(n3735), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4551 ( .A1(n3013), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4552 ( .A1(n3840), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3674) );
  NAND4_X1 U4553 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3678)
         );
  OAI21_X1 U4554 ( .B1(n3679), .B2(n3678), .A(n3724), .ZN(n3682) );
  NAND2_X1 U4555 ( .A1(n5446), .A2(EAX_REG_15__SCAN_IN), .ZN(n3681) );
  NAND2_X1 U4556 ( .A1(n5445), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3680)
         );
  NAND3_X1 U4557 ( .A1(n3682), .A2(n3681), .A3(n3680), .ZN(n3683) );
  AOI21_X1 U4558 ( .B1(n5748), .B2(n5055), .A(n3683), .ZN(n5593) );
  AOI22_X1 U4559 ( .A1(n3006), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4560 ( .A1(n3735), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4561 ( .A1(n3840), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4562 ( .A1(n3800), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4563 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3694)
         );
  AOI22_X1 U4564 ( .A1(n3013), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4565 ( .A1(n3452), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4566 ( .A1(n3837), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4567 ( .A1(n3781), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4568 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3693)
         );
  NOR2_X1 U4569 ( .A1(n3694), .A2(n3693), .ZN(n3698) );
  OAI21_X1 U4570 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6593), .A(n4987), 
        .ZN(n3695) );
  INV_X1 U4571 ( .A(n3695), .ZN(n3696) );
  AOI21_X1 U4572 ( .B1(n5446), .B2(EAX_REG_22__SCAN_IN), .A(n3696), .ZN(n3697)
         );
  OAI21_X1 U4573 ( .B1(n3863), .B2(n3698), .A(n3697), .ZN(n3701) );
  OAI21_X1 U4574 ( .B1(n3699), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3707), 
        .ZN(n5893) );
  OR2_X1 U4575 ( .A1(n5893), .A2(n3860), .ZN(n3700) );
  NAND2_X1 U4576 ( .A1(n3701), .A2(n3700), .ZN(n5637) );
  XNOR2_X1 U4577 ( .A(n3703), .B(n3702), .ZN(n3706) );
  INV_X1 U4578 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5881) );
  AOI21_X1 U4579 ( .B1(n5881), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3704) );
  AOI21_X1 U4580 ( .B1(n5446), .B2(EAX_REG_23__SCAN_IN), .A(n3704), .ZN(n3705)
         );
  OAI21_X1 U4581 ( .B1(n3863), .B2(n3706), .A(n3705), .ZN(n3709) );
  XNOR2_X1 U4582 ( .A(n3707), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5873)
         );
  NAND2_X1 U4583 ( .A1(n5873), .A2(n5055), .ZN(n3708) );
  AND2_X1 U4584 ( .A1(n3709), .A2(n3708), .ZN(n5628) );
  INV_X1 U4585 ( .A(n5628), .ZN(n3710) );
  XOR2_X1 U4586 ( .A(n6038), .B(n3712), .Z(n6041) );
  AOI22_X1 U4587 ( .A1(n3735), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4588 ( .A1(n3013), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4589 ( .A1(n3800), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4590 ( .A1(n3840), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4591 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3722)
         );
  AOI22_X1 U4592 ( .A1(n3007), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4593 ( .A1(n3759), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4594 ( .A1(n3452), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4595 ( .A1(n3781), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4596 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3721)
         );
  OR2_X1 U4597 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  AOI22_X1 U4598 ( .A1(n3724), .A2(n3723), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4599 ( .A1(n5446), .A2(EAX_REG_14__SCAN_IN), .ZN(n3725) );
  OAI211_X1 U4600 ( .C1(n6041), .C2(n3860), .A(n3726), .B(n3725), .ZN(n5264)
         );
  INV_X1 U4601 ( .A(n5264), .ZN(n3727) );
  AOI22_X1 U4602 ( .A1(n3006), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4603 ( .A1(n3013), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4604 ( .A1(n3823), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4605 ( .A1(n3848), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3731) );
  NAND4_X1 U4606 ( .A1(n3734), .A2(n3733), .A3(n3732), .A4(n3731), .ZN(n3741)
         );
  AOI22_X1 U4607 ( .A1(n3759), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3781), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4608 ( .A1(n3837), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4609 ( .A1(n3735), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4610 ( .A1(n3840), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4611 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NOR2_X1 U4612 ( .A1(n3741), .A2(n3740), .ZN(n3753) );
  NAND2_X1 U4613 ( .A1(n3743), .A2(n3742), .ZN(n3752) );
  XOR2_X1 U4614 ( .A(n3753), .B(n3752), .Z(n3744) );
  NAND2_X1 U4615 ( .A1(n3744), .A2(n3831), .ZN(n3747) );
  INV_X1 U4616 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6782) );
  OAI21_X1 U4617 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6782), .A(n3860), .ZN(
        n3745) );
  AOI21_X1 U4618 ( .B1(n5446), .B2(EAX_REG_25__SCAN_IN), .A(n3745), .ZN(n3746)
         );
  NAND2_X1 U4619 ( .A1(n3747), .A2(n3746), .ZN(n3751) );
  NAND2_X1 U4620 ( .A1(n3748), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3769)
         );
  OR2_X1 U4621 ( .A1(n3748), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3749)
         );
  AND2_X1 U4622 ( .A1(n3769), .A2(n3749), .ZN(n5862) );
  NAND2_X1 U4623 ( .A1(n5862), .A2(n5055), .ZN(n3750) );
  NAND2_X1 U4624 ( .A1(n3751), .A2(n3750), .ZN(n5619) );
  NOR2_X1 U4625 ( .A1(n3753), .A2(n3752), .ZN(n3774) );
  AOI22_X1 U4626 ( .A1(n3007), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4627 ( .A1(n3013), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4628 ( .A1(n3800), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4629 ( .A1(n3452), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3754), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3755) );
  NAND4_X1 U4630 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3765)
         );
  AOI22_X1 U4631 ( .A1(n3759), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4632 ( .A1(n3837), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4633 ( .A1(n3103), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3847), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4634 ( .A1(n3840), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4635 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3764)
         );
  OR2_X1 U4636 ( .A1(n3765), .A2(n3764), .ZN(n3773) );
  XNOR2_X1 U4637 ( .A(n3774), .B(n3773), .ZN(n3768) );
  INV_X1 U4638 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U4639 ( .B1(n6737), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3766) );
  AOI21_X1 U4640 ( .B1(n5446), .B2(EAX_REG_26__SCAN_IN), .A(n3766), .ZN(n3767)
         );
  OAI21_X1 U4641 ( .B1(n3768), .B2(n3863), .A(n3767), .ZN(n3772) );
  NAND2_X1 U4642 ( .A1(n3769), .A2(n6737), .ZN(n3770) );
  NAND2_X1 U4643 ( .A1(n3794), .A2(n3770), .ZN(n5852) );
  OR2_X1 U4644 ( .A1(n5852), .A2(n3860), .ZN(n3771) );
  NAND2_X1 U4645 ( .A1(n3772), .A2(n3771), .ZN(n5611) );
  NAND2_X1 U4646 ( .A1(n3774), .A2(n3773), .ZN(n3798) );
  AOI22_X1 U4647 ( .A1(n3103), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4648 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3840), .B1(n3221), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4649 ( .A1(n3013), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4650 ( .A1(n3848), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4651 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3788)
         );
  AOI22_X1 U4652 ( .A1(n3007), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4653 ( .A1(n3730), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4654 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3781), .B1(n3102), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4655 ( .A1(n3837), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3782), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3783) );
  NAND4_X1 U4656 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3787)
         );
  NOR2_X1 U4657 ( .A1(n3788), .A2(n3787), .ZN(n3799) );
  XOR2_X1 U4658 ( .A(n3798), .B(n3799), .Z(n3789) );
  NAND2_X1 U4659 ( .A1(n3789), .A2(n3831), .ZN(n3793) );
  INV_X1 U4660 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3790) );
  NOR2_X1 U4661 ( .A1(n3790), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3791) );
  AOI211_X1 U4662 ( .C1(n5446), .C2(EAX_REG_27__SCAN_IN), .A(n5055), .B(n3791), 
        .ZN(n3792) );
  XNOR2_X1 U4663 ( .A(n3794), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5562)
         );
  AOI22_X1 U4664 ( .A1(n3793), .A2(n3792), .B1(n5055), .B2(n5562), .ZN(n5369)
         );
  NAND2_X1 U4665 ( .A1(n5612), .A2(n5369), .ZN(n5368) );
  INV_X1 U4666 ( .A(n3794), .ZN(n3795) );
  NAND2_X1 U4667 ( .A1(n3795), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3796)
         );
  INV_X1 U4668 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U4669 ( .A1(n3796), .A2(n5554), .ZN(n3797) );
  NAND2_X1 U4670 ( .A1(n3865), .A2(n3797), .ZN(n5699) );
  NOR2_X1 U4671 ( .A1(n3799), .A2(n3798), .ZN(n3817) );
  AOI22_X1 U4672 ( .A1(n3007), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4673 ( .A1(n3013), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4674 ( .A1(n3800), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4675 ( .A1(n3848), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4676 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3811)
         );
  AOI22_X1 U4677 ( .A1(n3759), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4678 ( .A1(n3837), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4679 ( .A1(n3103), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4680 ( .A1(n3840), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4681 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3810)
         );
  OR2_X1 U4682 ( .A1(n3811), .A2(n3810), .ZN(n3816) );
  XNOR2_X1 U4683 ( .A(n3817), .B(n3816), .ZN(n3814) );
  AOI21_X1 U4684 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n4987), .A(n5055), 
        .ZN(n3813) );
  NAND2_X1 U4685 ( .A1(n5446), .A2(EAX_REG_28__SCAN_IN), .ZN(n3812) );
  OAI211_X1 U4686 ( .C1(n3814), .C2(n3863), .A(n3813), .B(n3812), .ZN(n3815)
         );
  OAI21_X1 U4687 ( .B1(n3860), .B2(n5699), .A(n3815), .ZN(n5548) );
  NAND2_X1 U4688 ( .A1(n3817), .A2(n3816), .ZN(n3855) );
  AOI22_X1 U4689 ( .A1(n3735), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4690 ( .A1(n3759), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4691 ( .A1(n3840), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4692 ( .A1(n3730), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4693 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3830)
         );
  AOI22_X1 U4694 ( .A1(n3006), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4695 ( .A1(n3452), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4696 ( .A1(n3013), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4697 ( .A1(n3847), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4698 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  NOR2_X1 U4699 ( .A1(n3830), .A2(n3829), .ZN(n3856) );
  XOR2_X1 U4700 ( .A(n3855), .B(n3856), .Z(n3832) );
  NAND2_X1 U4701 ( .A1(n3832), .A2(n3831), .ZN(n3836) );
  INV_X1 U4702 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3833) );
  AOI21_X1 U4703 ( .B1(n3833), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3834) );
  AOI21_X1 U4704 ( .B1(n5446), .B2(EAX_REG_29__SCAN_IN), .A(n3834), .ZN(n3835)
         );
  XNOR2_X1 U4705 ( .A(n3865), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5471)
         );
  AOI22_X1 U4706 ( .A1(n3836), .A2(n3835), .B1(n5055), .B2(n5471), .ZN(n5271)
         );
  AOI22_X1 U4707 ( .A1(n2994), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3730), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4708 ( .A1(n3759), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4709 ( .A1(n3735), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4710 ( .A1(n3840), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3839), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4711 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3854)
         );
  AOI22_X1 U4712 ( .A1(n3013), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3007), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4713 ( .A1(n3800), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4714 ( .A1(n3847), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4715 ( .A1(n3452), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3074), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4716 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3853)
         );
  NOR2_X1 U4717 ( .A1(n3854), .A2(n3853), .ZN(n3858) );
  NOR2_X1 U4718 ( .A1(n3856), .A2(n3855), .ZN(n3857) );
  XOR2_X1 U4719 ( .A(n3858), .B(n3857), .Z(n3864) );
  NAND2_X1 U4720 ( .A1(n4987), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3859)
         );
  NAND2_X1 U4721 ( .A1(n3860), .A2(n3859), .ZN(n3861) );
  AOI21_X1 U4722 ( .B1(n5446), .B2(EAX_REG_30__SCAN_IN), .A(n3861), .ZN(n3862)
         );
  OAI21_X1 U4723 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3868) );
  INV_X1 U4724 ( .A(n3865), .ZN(n3866) );
  NAND2_X1 U4725 ( .A1(n3866), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5059)
         );
  XNOR2_X1 U4726 ( .A(n5059), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5425)
         );
  NAND2_X1 U4727 ( .A1(n5425), .A2(n5055), .ZN(n3867) );
  NAND2_X1 U4728 ( .A1(n3868), .A2(n3867), .ZN(n5443) );
  XNOR2_X1 U4729 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3883) );
  XOR2_X1 U4730 ( .A(n3883), .B(n3884), .Z(n4180) );
  INV_X1 U4731 ( .A(n3911), .ZN(n3870) );
  OAI21_X1 U4732 ( .B1(n3870), .B2(n4243), .A(n3196), .ZN(n3880) );
  AOI21_X1 U4733 ( .B1(n4243), .B2(n3196), .A(n4218), .ZN(n3894) );
  INV_X1 U4734 ( .A(n3884), .ZN(n3872) );
  NAND2_X1 U4735 ( .A1(n3304), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4736 ( .A1(n3872), .A2(n3871), .ZN(n3875) );
  OAI21_X1 U4737 ( .B1(n3874), .B2(n3875), .A(n3873), .ZN(n3878) );
  INV_X1 U4738 ( .A(n3875), .ZN(n3876) );
  NAND2_X1 U4739 ( .A1(n3911), .A2(n3876), .ZN(n3877) );
  AOI22_X1 U4740 ( .A1(n3894), .A2(n3878), .B1(n3915), .B2(n3877), .ZN(n3879)
         );
  OAI21_X1 U4741 ( .B1(n3880), .B2(n4180), .A(n3879), .ZN(n3882) );
  NAND3_X1 U4742 ( .A1(n3880), .A2(STATE2_REG_0__SCAN_IN), .A3(n4180), .ZN(
        n3881) );
  OAI211_X1 U4743 ( .C1(n4180), .C2(n3915), .A(n3882), .B(n3881), .ZN(n3897)
         );
  NAND2_X1 U4744 ( .A1(n3884), .A2(n3883), .ZN(n3886) );
  NAND2_X1 U4745 ( .A1(n6461), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4746 ( .A1(n3886), .A2(n3885), .ZN(n3890) );
  XNOR2_X1 U4747 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3889) );
  INV_X1 U4748 ( .A(n3889), .ZN(n3887) );
  XNOR2_X1 U4749 ( .A(n3890), .B(n3887), .ZN(n4179) );
  NAND2_X1 U4750 ( .A1(n3911), .A2(n4179), .ZN(n3893) );
  OAI211_X1 U4751 ( .C1(n4179), .C2(n3888), .A(n3894), .B(n3893), .ZN(n3896)
         );
  XNOR2_X1 U4752 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4753 ( .A1(n3890), .A2(n3889), .ZN(n3892) );
  NAND2_X1 U4754 ( .A1(n4716), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3891) );
  NAND2_X1 U4755 ( .A1(n3892), .A2(n3891), .ZN(n3899) );
  XOR2_X1 U4756 ( .A(n3898), .B(n3899), .Z(n4178) );
  INV_X1 U4757 ( .A(n4122), .ZN(n4062) );
  OAI22_X1 U4758 ( .A1(n3894), .A2(n3893), .B1(n4178), .B2(n4062), .ZN(n3895)
         );
  AOI21_X1 U4759 ( .B1(n3897), .B2(n3896), .A(n3895), .ZN(n3905) );
  NAND2_X1 U4760 ( .A1(n3899), .A2(n3898), .ZN(n3901) );
  NAND2_X1 U4761 ( .A1(n6466), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U4762 ( .A1(n3901), .A2(n3900), .ZN(n3908) );
  NAND2_X1 U4763 ( .A1(n3902), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3909) );
  OR2_X1 U4764 ( .A1(n3908), .A2(n3909), .ZN(n4183) );
  AOI21_X1 U4765 ( .B1(n4178), .B2(n4183), .A(n3903), .ZN(n3904) );
  OAI22_X1 U4766 ( .A1(n3905), .A2(n3904), .B1(n3915), .B2(n4183), .ZN(n3906)
         );
  AOI21_X1 U4767 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6599), .A(n3906), 
        .ZN(n3913) );
  INV_X1 U4768 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6614) );
  AND2_X1 U4769 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6614), .ZN(n3907)
         );
  OR2_X1 U4770 ( .A1(n3908), .A2(n3907), .ZN(n3910) );
  NAND2_X1 U4771 ( .A1(n3911), .A2(n3914), .ZN(n3912) );
  NAND2_X1 U4772 ( .A1(n3913), .A2(n3912), .ZN(n3917) );
  INV_X1 U4773 ( .A(n3914), .ZN(n4182) );
  NAND2_X1 U4774 ( .A1(n3918), .A2(n5072), .ZN(n3919) );
  INV_X1 U4775 ( .A(n6592), .ZN(n4272) );
  MUX2_X1 U4776 ( .A(n3919), .B(n4272), .S(n3187), .Z(n4208) );
  NAND2_X1 U4777 ( .A1(n6452), .A2(n4059), .ZN(n3922) );
  NOR2_X1 U4778 ( .A1(n4202), .A2(n3920), .ZN(n3921) );
  NAND2_X1 U4779 ( .A1(n3922), .A2(n3921), .ZN(n4219) );
  INV_X1 U4780 ( .A(n4219), .ZN(n3923) );
  NAND2_X1 U4781 ( .A1(n4208), .A2(n3923), .ZN(n3925) );
  INV_X1 U4782 ( .A(n4210), .ZN(n5518) );
  NAND2_X1 U4783 ( .A1(n3925), .A2(n5518), .ZN(n4251) );
  OR2_X1 U4784 ( .A1(n4188), .A2(n4348), .ZN(n4201) );
  AND2_X1 U4785 ( .A1(n4251), .A2(n4201), .ZN(n4229) );
  NOR2_X1 U4786 ( .A1(n6452), .A2(n4243), .ZN(n4228) );
  NAND2_X1 U4787 ( .A1(n5524), .A2(n5514), .ZN(n3931) );
  INV_X1 U4788 ( .A(n5279), .ZN(n5454) );
  NAND3_X1 U4789 ( .A1(n5454), .A2(n4257), .A3(n4353), .ZN(n4295) );
  INV_X1 U4790 ( .A(n4295), .ZN(n3929) );
  INV_X4 U4791 ( .A(n3934), .ZN(n4030) );
  NAND3_X1 U4792 ( .A1(n3929), .A2(n3928), .A3(n4030), .ZN(n3930) );
  NAND2_X1 U4793 ( .A1(n3931), .A2(n3930), .ZN(n3933) );
  NAND2_X1 U4794 ( .A1(n3932), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6488) );
  INV_X1 U4795 ( .A(n6488), .ZN(n5528) );
  NOR2_X1 U4796 ( .A1(n5674), .A2(n5454), .ZN(n5672) );
  INV_X2 U4797 ( .A(n5672), .ZN(n5677) );
  NAND2_X1 U4798 ( .A1(n3935), .A2(n5072), .ZN(n3946) );
  NAND2_X1 U4799 ( .A1(n3946), .A2(EBX_REG_0__SCAN_IN), .ZN(n3937) );
  INV_X1 U4800 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U4801 ( .A1(n4262), .A2(n5190), .ZN(n3936) );
  INV_X2 U4802 ( .A(n3938), .ZN(n5307) );
  INV_X1 U4803 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U4804 ( .A1(n3946), .A2(n4215), .ZN(n3941) );
  BUF_X4 U4805 ( .A(n3938), .Z(n4262) );
  INV_X1 U4806 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U4807 ( .A1(n4030), .A2(n3939), .ZN(n3940) );
  NAND3_X1 U4808 ( .A1(n3941), .A2(n4262), .A3(n3940), .ZN(n3942) );
  XNOR2_X1 U4809 ( .A(n4236), .B(n3944), .ZN(n4287) );
  NAND2_X1 U4810 ( .A1(n4290), .A2(n3944), .ZN(n4306) );
  OR2_X1 U4811 ( .A1(n4028), .A2(EBX_REG_2__SCAN_IN), .ZN(n3951) );
  INV_X1 U4812 ( .A(n3946), .ZN(n3954) );
  INV_X1 U4813 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U4814 ( .A1(n4022), .A2(n6346), .ZN(n3949) );
  INV_X1 U4815 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U4816 ( .A1(n4030), .A2(n3947), .ZN(n3948) );
  NAND3_X1 U4817 ( .A1(n3949), .A2(n4262), .A3(n3948), .ZN(n3950) );
  NAND2_X1 U4818 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3955)
         );
  OAI211_X1 U4819 ( .C1(n5530), .C2(EBX_REG_3__SCAN_IN), .A(n4022), .B(n3955), 
        .ZN(n3956) );
  OAI21_X1 U4820 ( .B1(n5272), .B2(EBX_REG_3__SCAN_IN), .A(n3956), .ZN(n4313)
         );
  NOR2_X2 U4821 ( .A1(n4304), .A2(n4313), .ZN(n4311) );
  OR2_X1 U4822 ( .A1(n4028), .A2(EBX_REG_4__SCAN_IN), .ZN(n3960) );
  NAND2_X1 U4823 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3957)
         );
  NAND2_X1 U4824 ( .A1(n4022), .A2(n3957), .ZN(n3958) );
  OAI21_X1 U4825 ( .B1(EBX_REG_4__SCAN_IN), .B2(n5530), .A(n3958), .ZN(n3959)
         );
  NAND2_X1 U4826 ( .A1(n3960), .A2(n3959), .ZN(n4410) );
  NAND2_X1 U4827 ( .A1(n4311), .A2(n4410), .ZN(n4409) );
  NAND2_X1 U4828 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3961)
         );
  OAI211_X1 U4829 ( .C1(n5530), .C2(EBX_REG_5__SCAN_IN), .A(n4022), .B(n3961), 
        .ZN(n3962) );
  OAI21_X1 U4830 ( .B1(n5272), .B2(EBX_REG_5__SCAN_IN), .A(n3962), .ZN(n4415)
         );
  OR2_X1 U4831 ( .A1(n4028), .A2(EBX_REG_6__SCAN_IN), .ZN(n3969) );
  INV_X1 U4832 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U4833 ( .A1(n4022), .A2(n5170), .ZN(n3967) );
  INV_X1 U4834 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U4835 ( .A1(n4030), .A2(n3965), .ZN(n3966) );
  NAND3_X1 U4836 ( .A1(n3967), .A2(n4262), .A3(n3966), .ZN(n3968) );
  NOR2_X2 U4837 ( .A1(n4416), .A2(n4622), .ZN(n4624) );
  MUX2_X1 U4838 ( .A(n5272), .B(n4262), .S(EBX_REG_7__SCAN_IN), .Z(n3970) );
  OAI21_X1 U4839 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5531), .A(n3970), 
        .ZN(n4926) );
  INV_X1 U4840 ( .A(n4926), .ZN(n3971) );
  AND2_X2 U4841 ( .A1(n4624), .A2(n3971), .ZN(n4875) );
  OR2_X1 U4842 ( .A1(n4028), .A2(EBX_REG_8__SCAN_IN), .ZN(n3976) );
  INV_X1 U4843 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U4844 ( .A1(n4022), .A2(n6290), .ZN(n3974) );
  INV_X1 U4845 ( .A(EBX_REG_8__SCAN_IN), .ZN(n3972) );
  NAND2_X1 U4846 ( .A1(n4030), .A2(n3972), .ZN(n3973) );
  NAND3_X1 U4847 ( .A1(n3974), .A2(n4262), .A3(n3973), .ZN(n3975) );
  NAND2_X1 U4848 ( .A1(n3976), .A2(n3975), .ZN(n4876) );
  NAND2_X1 U4849 ( .A1(n4875), .A2(n4876), .ZN(n4874) );
  MUX2_X1 U4850 ( .A(n5272), .B(n4262), .S(EBX_REG_9__SCAN_IN), .Z(n3977) );
  OAI21_X1 U4851 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5531), .A(n3977), 
        .ZN(n5036) );
  OR2_X2 U4852 ( .A1(n4874), .A2(n5036), .ZN(n5184) );
  OR2_X1 U4853 ( .A1(n4028), .A2(EBX_REG_10__SCAN_IN), .ZN(n3981) );
  INV_X1 U4854 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U4855 ( .A1(n4022), .A2(n4133), .ZN(n3979) );
  INV_X1 U4856 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U4857 ( .A1(n4030), .A2(n6077), .ZN(n3978) );
  NAND3_X1 U4858 ( .A1(n3979), .A2(n4262), .A3(n3978), .ZN(n3980) );
  MUX2_X1 U4859 ( .A(n5272), .B(n4262), .S(EBX_REG_11__SCAN_IN), .Z(n3982) );
  OAI21_X1 U4860 ( .B1(n5531), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n3982), 
        .ZN(n3983) );
  INV_X1 U4861 ( .A(n3983), .ZN(n5225) );
  OR2_X1 U4862 ( .A1(n4028), .A2(EBX_REG_12__SCAN_IN), .ZN(n3988) );
  INV_X1 U4863 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U4864 ( .A1(n4022), .A2(n4139), .ZN(n3986) );
  INV_X1 U4865 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3984) );
  NAND2_X1 U4866 ( .A1(n4030), .A2(n3984), .ZN(n3985) );
  NAND3_X1 U4867 ( .A1(n3986), .A2(n4262), .A3(n3985), .ZN(n3987) );
  NAND2_X1 U4868 ( .A1(n3988), .A2(n3987), .ZN(n5233) );
  NAND2_X1 U4869 ( .A1(n5224), .A2(n5233), .ZN(n5232) );
  MUX2_X1 U4870 ( .A(n5272), .B(n4262), .S(EBX_REG_13__SCAN_IN), .Z(n3989) );
  OAI21_X1 U4871 ( .B1(n5531), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n3989), 
        .ZN(n5261) );
  OR2_X2 U4872 ( .A1(n5232), .A2(n5261), .ZN(n5267) );
  OR2_X1 U4873 ( .A1(n4028), .A2(EBX_REG_14__SCAN_IN), .ZN(n3993) );
  NAND2_X1 U4874 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3990) );
  NAND2_X1 U4875 ( .A1(n4022), .A2(n3990), .ZN(n3991) );
  OAI21_X1 U4876 ( .B1(EBX_REG_14__SCAN_IN), .B2(n5530), .A(n3991), .ZN(n3992)
         );
  AND2_X1 U4877 ( .A1(n3993), .A2(n3992), .ZN(n5266) );
  MUX2_X1 U4878 ( .A(n5272), .B(n4262), .S(EBX_REG_15__SCAN_IN), .Z(n3994) );
  OAI21_X1 U4879 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5531), .A(n3994), 
        .ZN(n5594) );
  OR2_X1 U4880 ( .A1(n4028), .A2(EBX_REG_16__SCAN_IN), .ZN(n3998) );
  INV_X1 U4881 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U4882 ( .A1(n4022), .A2(n5964), .ZN(n3996) );
  INV_X1 U4883 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U4884 ( .A1(n4030), .A2(n6029), .ZN(n3995) );
  NAND3_X1 U4885 ( .A1(n3996), .A2(n4262), .A3(n3995), .ZN(n3997) );
  NAND2_X1 U4886 ( .A1(n3998), .A2(n3997), .ZN(n5666) );
  MUX2_X1 U4887 ( .A(n5272), .B(n3938), .S(EBX_REG_17__SCAN_IN), .Z(n3999) );
  OAI21_X1 U4888 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5531), .A(n3999), 
        .ZN(n5581) );
  OR2_X2 U4889 ( .A1(n5580), .A2(n5581), .ZN(n5658) );
  OR2_X1 U4890 ( .A1(n4028), .A2(EBX_REG_19__SCAN_IN), .ZN(n4003) );
  NAND2_X1 U4891 ( .A1(n3938), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U4892 ( .A1(n4022), .A2(n4000), .ZN(n4001) );
  OAI21_X1 U4893 ( .B1(EBX_REG_19__SCAN_IN), .B2(n5530), .A(n4001), .ZN(n4002)
         );
  AND2_X1 U4894 ( .A1(n4003), .A2(n4002), .ZN(n5309) );
  NOR2_X2 U4895 ( .A1(n5658), .A2(n5309), .ZN(n5381) );
  INV_X1 U4896 ( .A(n5531), .ZN(n4238) );
  INV_X1 U4897 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5388) );
  NOR2_X1 U4898 ( .A1(n5530), .A2(EBX_REG_20__SCAN_IN), .ZN(n4004) );
  AOI21_X1 U4899 ( .B1(n4238), .B2(n5388), .A(n4004), .ZN(n5383) );
  OR2_X1 U4900 ( .A1(n5531), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4005)
         );
  INV_X1 U4901 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U4902 ( .A1(n4030), .A2(n5661), .ZN(n5308) );
  NAND2_X1 U4903 ( .A1(n4005), .A2(n5308), .ZN(n5382) );
  NAND2_X1 U4904 ( .A1(n5307), .A2(EBX_REG_20__SCAN_IN), .ZN(n4007) );
  NAND2_X1 U4905 ( .A1(n5382), .A2(n4262), .ZN(n4006) );
  OAI211_X1 U4906 ( .C1(n5383), .C2(n5382), .A(n4007), .B(n4006), .ZN(n4008)
         );
  INV_X1 U4907 ( .A(n4008), .ZN(n4009) );
  AND2_X2 U4908 ( .A1(n5381), .A2(n4009), .ZN(n5648) );
  OR2_X1 U4909 ( .A1(n4028), .A2(EBX_REG_21__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U4910 ( .A1(n3938), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4010) );
  NAND2_X1 U4911 ( .A1(n4022), .A2(n4010), .ZN(n4011) );
  OAI21_X1 U4912 ( .B1(EBX_REG_21__SCAN_IN), .B2(n5530), .A(n4011), .ZN(n4012)
         );
  NAND2_X1 U4913 ( .A1(n4013), .A2(n4012), .ZN(n5647) );
  NAND2_X1 U4914 ( .A1(n5648), .A2(n5647), .ZN(n5640) );
  NAND2_X1 U4915 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4014) );
  OAI211_X1 U4916 ( .C1(n5530), .C2(EBX_REG_22__SCAN_IN), .A(n4022), .B(n4014), 
        .ZN(n4015) );
  OAI21_X1 U4917 ( .B1(n5272), .B2(EBX_REG_22__SCAN_IN), .A(n4015), .ZN(n5641)
         );
  OR2_X1 U4918 ( .A1(n4028), .A2(EBX_REG_23__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U4919 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U4920 ( .A1(n4022), .A2(n4016), .ZN(n4017) );
  OAI21_X1 U4921 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5530), .A(n4017), .ZN(n4018)
         );
  AND2_X1 U4922 ( .A1(n4019), .A2(n4018), .ZN(n5631) );
  MUX2_X1 U4923 ( .A(n5272), .B(n3938), .S(EBX_REG_24__SCAN_IN), .Z(n4021) );
  NAND2_X1 U4924 ( .A1(n4238), .A2(n5417), .ZN(n4020) );
  AND2_X1 U4925 ( .A1(n4021), .A2(n4020), .ZN(n5412) );
  OR2_X1 U4926 ( .A1(n4028), .A2(EBX_REG_25__SCAN_IN), .ZN(n4026) );
  INV_X1 U4927 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U4928 ( .A1(n4022), .A2(n5337), .ZN(n4024) );
  INV_X1 U4929 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U4930 ( .A1(n4030), .A2(n5865), .ZN(n4023) );
  NAND3_X1 U4931 ( .A1(n4024), .A2(n3938), .A3(n4023), .ZN(n4025) );
  NAND2_X1 U4932 ( .A1(n4026), .A2(n4025), .ZN(n5621) );
  NAND2_X1 U4933 ( .A1(n5411), .A2(n5621), .ZN(n5614) );
  MUX2_X1 U4934 ( .A(n5272), .B(n3938), .S(EBX_REG_26__SCAN_IN), .Z(n4027) );
  OAI21_X1 U4935 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5531), .A(n4027), 
        .ZN(n5615) );
  OR2_X1 U4936 ( .A1(n4028), .A2(EBX_REG_27__SCAN_IN), .ZN(n4034) );
  INV_X1 U4937 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U4938 ( .A1(n4022), .A2(n5765), .ZN(n4032) );
  INV_X1 U4939 ( .A(EBX_REG_27__SCAN_IN), .ZN(n4029) );
  NAND2_X1 U4940 ( .A1(n4030), .A2(n4029), .ZN(n4031) );
  NAND3_X1 U4941 ( .A1(n4032), .A2(n4262), .A3(n4031), .ZN(n4033) );
  AND2_X1 U4942 ( .A1(n4034), .A2(n4033), .ZN(n5357) );
  NAND2_X1 U4943 ( .A1(n3938), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4035) );
  OAI211_X1 U4944 ( .C1(n5530), .C2(EBX_REG_28__SCAN_IN), .A(n4022), .B(n4035), 
        .ZN(n4036) );
  OAI21_X1 U4945 ( .B1(n5272), .B2(EBX_REG_28__SCAN_IN), .A(n4036), .ZN(n5550)
         );
  OR2_X1 U4946 ( .A1(n5531), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5273)
         );
  OAI211_X1 U4947 ( .C1(EBX_REG_29__SCAN_IN), .C2(n5530), .A(n5278), .B(n5273), 
        .ZN(n4041) );
  NAND2_X1 U4948 ( .A1(n5531), .A2(EBX_REG_30__SCAN_IN), .ZN(n4038) );
  NAND2_X1 U4949 ( .A1(n5530), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U4950 ( .A1(n4038), .A2(n4037), .ZN(n5534) );
  AOI21_X1 U4951 ( .B1(n4041), .B2(n5278), .A(n5534), .ZN(n4039) );
  NAND2_X1 U4952 ( .A1(n4041), .A2(n3938), .ZN(n5532) );
  INV_X1 U4953 ( .A(n5278), .ZN(n5553) );
  INV_X1 U4954 ( .A(n5534), .ZN(n4040) );
  AOI21_X1 U4955 ( .B1(n5553), .B2(n5307), .A(n4040), .ZN(n4042) );
  NAND2_X1 U4956 ( .A1(n4042), .A2(n4041), .ZN(n4043) );
  INV_X1 U4957 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4045) );
  NAND2_X2 U4958 ( .A1(n5265), .A2(n5264), .ZN(n5636) );
  NOR2_X2 U4959 ( .A1(n5636), .A2(n5593), .ZN(n4051) );
  OR2_X2 U4960 ( .A1(n5654), .A2(n5653), .ZN(n5656) );
  AND2_X1 U4961 ( .A1(n5592), .A2(n4052), .ZN(n5395) );
  OR2_X2 U4962 ( .A1(n4053), .A2(n5395), .ZN(n5322) );
  AND2_X1 U4963 ( .A1(n6599), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U4964 ( .A1(n5056), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6494) );
  NOR2_X2 U4965 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5836) );
  OR2_X1 U4966 ( .A1(n6494), .A2(n5844), .ZN(n5406) );
  NOR2_X1 U4967 ( .A1(n5322), .A2(n5406), .ZN(n4160) );
  NAND2_X1 U4968 ( .A1(n4322), .A2(n4122), .ZN(n4058) );
  XNOR2_X1 U4969 ( .A(n4068), .B(n4067), .ZN(n4055) );
  OAI211_X1 U4970 ( .C1(n4055), .C2(n4272), .A(n4054), .B(n3196), .ZN(n4056)
         );
  INV_X1 U4971 ( .A(n4056), .ZN(n4057) );
  NAND2_X1 U4972 ( .A1(n4058), .A2(n4057), .ZN(n4381) );
  NAND2_X1 U4973 ( .A1(n4059), .A2(n4364), .ZN(n4070) );
  OAI21_X1 U4974 ( .B1(n4272), .B2(n4068), .A(n4070), .ZN(n4060) );
  INV_X1 U4975 ( .A(n4060), .ZN(n4061) );
  OAI21_X2 U4976 ( .B1(n4324), .B2(n4062), .A(n4061), .ZN(n4242) );
  NAND2_X1 U4977 ( .A1(n4242), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4063)
         );
  NAND2_X1 U4978 ( .A1(n4063), .A2(n4215), .ZN(n4064) );
  AND2_X1 U4979 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U4980 ( .A1(n4242), .A2(n6334), .ZN(n4065) );
  AND2_X1 U4981 ( .A1(n4064), .A2(n4065), .ZN(n4382) );
  NAND2_X1 U4982 ( .A1(n4381), .A2(n4382), .ZN(n4066) );
  NAND2_X1 U4983 ( .A1(n4066), .A2(n4065), .ZN(n6245) );
  NAND2_X1 U4984 ( .A1(n6245), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4073)
         );
  NAND2_X1 U4985 ( .A1(n4068), .A2(n4067), .ZN(n4079) );
  XNOR2_X1 U4986 ( .A(n4079), .B(n4069), .ZN(n4071) );
  OAI21_X1 U4987 ( .B1(n4071), .B2(n4272), .A(n4070), .ZN(n4072) );
  AOI21_X1 U4988 ( .B1(n4321), .B2(n4122), .A(n4072), .ZN(n6246) );
  NAND2_X1 U4989 ( .A1(n4073), .A2(n6246), .ZN(n4076) );
  INV_X1 U4990 ( .A(n6245), .ZN(n4074) );
  NAND2_X1 U4991 ( .A1(n4074), .A2(n6346), .ZN(n4075) );
  AND2_X1 U4992 ( .A1(n4076), .A2(n4075), .ZN(n5025) );
  NAND2_X1 U4993 ( .A1(n4077), .A2(n4122), .ZN(n4083) );
  NAND2_X1 U4994 ( .A1(n4079), .A2(n4078), .ZN(n4088) );
  INV_X1 U4995 ( .A(n4087), .ZN(n4080) );
  XNOR2_X1 U4996 ( .A(n4088), .B(n4080), .ZN(n4081) );
  NAND2_X1 U4997 ( .A1(n4081), .A2(n6592), .ZN(n4082) );
  NAND2_X1 U4998 ( .A1(n4083), .A2(n4082), .ZN(n4084) );
  INV_X1 U4999 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6329) );
  XNOR2_X1 U5000 ( .A(n4084), .B(n6329), .ZN(n5024) );
  NAND2_X1 U5001 ( .A1(n5025), .A2(n5024), .ZN(n5022) );
  NAND2_X1 U5002 ( .A1(n4084), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4085)
         );
  NAND2_X1 U5003 ( .A1(n5022), .A2(n4085), .ZN(n6238) );
  NAND2_X1 U5004 ( .A1(n4086), .A2(n4122), .ZN(n4091) );
  NAND2_X1 U5005 ( .A1(n4088), .A2(n4087), .ZN(n4106) );
  XNOR2_X1 U5006 ( .A(n4106), .B(n4104), .ZN(n4089) );
  NAND2_X1 U5007 ( .A1(n4089), .A2(n6592), .ZN(n4090) );
  NAND2_X1 U5008 ( .A1(n4091), .A2(n4090), .ZN(n4092) );
  INV_X1 U5009 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U5010 ( .A(n4092), .B(n6320), .ZN(n6237) );
  NAND2_X1 U5011 ( .A1(n6238), .A2(n6237), .ZN(n6240) );
  NAND2_X1 U5012 ( .A1(n4092), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4093)
         );
  NAND2_X1 U5013 ( .A1(n6240), .A2(n4093), .ZN(n5049) );
  NAND2_X1 U5014 ( .A1(n4094), .A2(n4122), .ZN(n4099) );
  INV_X1 U5015 ( .A(n4104), .ZN(n4095) );
  OR2_X1 U5016 ( .A1(n4106), .A2(n4095), .ZN(n4096) );
  XNOR2_X1 U5017 ( .A(n4096), .B(n4103), .ZN(n4097) );
  NAND2_X1 U5018 ( .A1(n4097), .A2(n6592), .ZN(n4098) );
  NAND2_X1 U5019 ( .A1(n4099), .A2(n4098), .ZN(n4100) );
  INV_X1 U5020 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5168) );
  XNOR2_X1 U5021 ( .A(n4100), .B(n5168), .ZN(n5048) );
  NAND2_X1 U5022 ( .A1(n5049), .A2(n5048), .ZN(n5046) );
  NAND2_X1 U5023 ( .A1(n4100), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4101)
         );
  NAND2_X1 U5024 ( .A1(n5046), .A2(n4101), .ZN(n4676) );
  NAND3_X1 U5025 ( .A1(n4126), .A2(n4102), .A3(n4122), .ZN(n4109) );
  NAND2_X1 U5026 ( .A1(n4104), .A2(n4103), .ZN(n4105) );
  OR2_X1 U5027 ( .A1(n4106), .A2(n4105), .ZN(n4113) );
  XNOR2_X1 U5028 ( .A(n4113), .B(n4114), .ZN(n4107) );
  NAND2_X1 U5029 ( .A1(n4107), .A2(n6592), .ZN(n4108) );
  NAND2_X1 U5030 ( .A1(n4109), .A2(n4108), .ZN(n4110) );
  XNOR2_X1 U5031 ( .A(n4110), .B(n5170), .ZN(n4675) );
  NAND2_X1 U5032 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U5033 ( .A1(n4110), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4111)
         );
  NAND2_X1 U5034 ( .A1(n4674), .A2(n4111), .ZN(n5042) );
  NAND2_X1 U5035 ( .A1(n4112), .A2(n4122), .ZN(n4118) );
  INV_X1 U5036 ( .A(n4113), .ZN(n4115) );
  NAND2_X1 U5037 ( .A1(n4115), .A2(n4114), .ZN(n4128) );
  XNOR2_X1 U5038 ( .A(n4128), .B(n4121), .ZN(n4116) );
  NAND2_X1 U5039 ( .A1(n4116), .A2(n6592), .ZN(n4117) );
  NAND2_X1 U5040 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  INV_X1 U5041 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6285) );
  XNOR2_X1 U5042 ( .A(n4119), .B(n6285), .ZN(n5041) );
  NAND2_X1 U5043 ( .A1(n5042), .A2(n5041), .ZN(n5040) );
  NAND2_X1 U5044 ( .A1(n4119), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4120)
         );
  NAND2_X1 U5045 ( .A1(n5040), .A2(n4120), .ZN(n5403) );
  NAND2_X1 U5046 ( .A1(n4122), .A2(n4121), .ZN(n4124) );
  NOR2_X1 U5047 ( .A1(n4124), .A2(n4123), .ZN(n4125) );
  OR3_X1 U5048 ( .A1(n4128), .A2(n4127), .A3(n4272), .ZN(n4129) );
  NAND2_X1 U5049 ( .A1(n5720), .A2(n4129), .ZN(n4130) );
  XNOR2_X1 U5050 ( .A(n4130), .B(n6290), .ZN(n5402) );
  NAND2_X1 U5051 ( .A1(n5403), .A2(n5402), .ZN(n5401) );
  NAND2_X1 U5052 ( .A1(n4130), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4131)
         );
  INV_X1 U5053 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U5054 ( .A1(n5720), .A2(n5174), .ZN(n5158) );
  NAND2_X1 U5055 ( .A1(n5160), .A2(n5158), .ZN(n4132) );
  NAND2_X1 U5056 ( .A1(n4132), .A2(n5159), .ZN(n5214) );
  NAND2_X1 U5057 ( .A1(n5720), .A2(n4133), .ZN(n5215) );
  INV_X1 U5058 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4134) );
  AND2_X1 U5059 ( .A1(n5720), .A2(n4134), .ZN(n4136) );
  OAI21_X2 U5060 ( .B1(n6220), .B2(n4136), .A(n3019), .ZN(n5246) );
  NOR2_X1 U5061 ( .A1(n5720), .A2(n4139), .ZN(n5941) );
  XNOR2_X1 U5062 ( .A(n5720), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5945)
         );
  INV_X1 U5063 ( .A(n5945), .ZN(n4137) );
  OR2_X1 U5064 ( .A1(n5246), .A2(n4138), .ZN(n4143) );
  NAND2_X1 U5065 ( .A1(n5720), .A2(n4139), .ZN(n5943) );
  INV_X1 U5066 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4140) );
  NAND2_X1 U5067 ( .A1(n5720), .A2(n4140), .ZN(n4141) );
  NAND2_X1 U5068 ( .A1(n4143), .A2(n4142), .ZN(n5297) );
  INV_X1 U5069 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5298) );
  OAI22_X2 U5070 ( .A1(n5297), .A2(n4144), .B1(n5720), .B2(n5298), .ZN(n5745)
         );
  INV_X1 U5071 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5970) );
  NOR2_X1 U5072 ( .A1(n5720), .A2(n5970), .ZN(n4146) );
  NAND2_X1 U5073 ( .A1(n5720), .A2(n5970), .ZN(n4145) );
  OAI21_X1 U5074 ( .B1(n5745), .B2(n4146), .A(n4145), .ZN(n5323) );
  INV_X1 U5075 ( .A(n5323), .ZN(n4148) );
  NAND3_X1 U5076 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n4147) );
  NAND2_X1 U5077 ( .A1(n4148), .A2(n3018), .ZN(n4161) );
  INV_X1 U5078 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5936) );
  INV_X1 U5079 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5832) );
  AND3_X1 U5080 ( .A1(n5964), .A2(n5936), .A3(n5832), .ZN(n4149) );
  NAND2_X1 U5081 ( .A1(n4161), .A2(n4150), .ZN(n5331) );
  INV_X2 U5082 ( .A(n5331), .ZN(n5335) );
  INV_X1 U5083 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U5084 ( .A1(n5335), .A2(n6768), .ZN(n4163) );
  OAI21_X1 U5085 ( .B1(n5335), .B2(n6768), .A(n5378), .ZN(n4151) );
  XNOR2_X1 U5086 ( .A(n4151), .B(n5720), .ZN(n5823) );
  NOR2_X1 U5087 ( .A1(n4219), .A2(n4152), .ZN(n6472) );
  NAND2_X2 U5088 ( .A1(n4373), .A2(n6472), .ZN(n6229) );
  NAND2_X1 U5089 ( .A1(n5844), .A2(n4156), .ZN(n6602) );
  NAND2_X1 U5090 ( .A1(n6602), .A2(n6599), .ZN(n4153) );
  AND2_X2 U5091 ( .A1(n6229), .A2(n4153), .ZN(n6236) );
  NAND2_X1 U5092 ( .A1(n6599), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5093 ( .A1(n6593), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4154) );
  AND2_X1 U5094 ( .A1(n4155), .A2(n4154), .ZN(n4278) );
  INV_X1 U5095 ( .A(n6236), .ZN(n5741) );
  OR2_X1 U5096 ( .A1(n4156), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6281) );
  INV_X2 U5097 ( .A(n6281), .ZN(n6336) );
  NAND2_X1 U5098 ( .A1(n6336), .A2(REIP_REG_19__SCAN_IN), .ZN(n5817) );
  OAI21_X1 U5099 ( .B1(n5741), .B2(n5313), .A(n5817), .ZN(n4157) );
  OR2_X1 U5100 ( .A1(n4160), .A2(n4159), .ZN(U2967) );
  OAI21_X2 U5101 ( .B1(n5723), .B2(n6768), .A(n5720), .ZN(n5377) );
  XNOR2_X1 U5102 ( .A(n5720), .B(n5388), .ZN(n5379) );
  INV_X1 U5103 ( .A(n5379), .ZN(n4162) );
  NAND3_X1 U5104 ( .A1(n4163), .A2(n5377), .A3(n4162), .ZN(n5736) );
  OR2_X1 U5105 ( .A1(n5720), .A2(n5388), .ZN(n5737) );
  INV_X1 U5106 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6785) );
  XNOR2_X1 U5107 ( .A(n5720), .B(n6785), .ZN(n5740) );
  INV_X1 U5108 ( .A(n5740), .ZN(n4164) );
  AND2_X1 U5109 ( .A1(n5737), .A2(n4164), .ZN(n4165) );
  NAND2_X1 U5110 ( .A1(n5736), .A2(n4165), .ZN(n4166) );
  OAI21_X1 U5111 ( .B1(n5824), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n4166), 
        .ZN(n5731) );
  NAND3_X1 U5112 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4167) );
  OAI22_X2 U5113 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5731), .B2(n4167), .ZN(n4168) );
  INV_X1 U5114 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5417) );
  XNOR2_X1 U5115 ( .A(n4168), .B(n5417), .ZN(n5423) );
  INV_X1 U5116 ( .A(n6229), .ZN(n6251) );
  NAND2_X1 U5117 ( .A1(n5423), .A2(n6251), .ZN(n4177) );
  NOR2_X1 U5118 ( .A1(n5636), .A2(n4169), .ZN(n5630) );
  OAI21_X1 U5119 ( .B1(n5630), .B2(n4171), .A(n4170), .ZN(n5686) );
  INV_X1 U5120 ( .A(n5570), .ZN(n4173) );
  NAND2_X1 U5121 ( .A1(n6336), .A2(REIP_REG_24__SCAN_IN), .ZN(n5414) );
  OAI21_X1 U5122 ( .B1(n5741), .B2(n5571), .A(n5414), .ZN(n4172) );
  AOI21_X1 U5123 ( .B1(n4173), .B2(n6224), .A(n4172), .ZN(n4174) );
  NAND2_X1 U5124 ( .A1(n4177), .A2(n4176), .ZN(U2962) );
  INV_X1 U5125 ( .A(n5522), .ZN(n5513) );
  NAND2_X1 U5126 ( .A1(n4373), .A2(n5513), .ZN(n4187) );
  NAND3_X1 U5127 ( .A1(n4180), .A2(n4179), .A3(n4178), .ZN(n4181) );
  NAND2_X1 U5128 ( .A1(n4182), .A2(n4181), .ZN(n4184) );
  AND2_X1 U5129 ( .A1(n4184), .A2(n4183), .ZN(n4220) );
  INV_X1 U5130 ( .A(n4220), .ZN(n5519) );
  AND2_X1 U5131 ( .A1(n4210), .A2(n5519), .ZN(n5520) );
  NAND2_X1 U5132 ( .A1(n5520), .A2(n5528), .ZN(n4186) );
  AND2_X1 U5133 ( .A1(n5836), .A2(n6571), .ZN(n5078) );
  AOI21_X1 U5134 ( .B1(n4186), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5078), .ZN(
        n4185) );
  NAND2_X1 U5135 ( .A1(n4187), .A2(n4185), .ZN(U2788) );
  NOR2_X1 U5136 ( .A1(n5078), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4190) );
  INV_X1 U5137 ( .A(n4188), .ZN(n6597) );
  NOR2_X1 U5138 ( .A1(n6597), .A2(n6592), .ZN(n5526) );
  NAND2_X1 U5139 ( .A1(n6601), .A2(n5526), .ZN(n4189) );
  OAI21_X1 U5140 ( .B1(n6601), .B2(n4190), .A(n4189), .ZN(U3474) );
  INV_X1 U5141 ( .A(n4192), .ZN(n6137) );
  INV_X1 U5142 ( .A(n4296), .ZN(n4198) );
  NOR2_X1 U5143 ( .A1(n4198), .A2(n4197), .ZN(n4199) );
  AND2_X1 U5144 ( .A1(n4196), .A2(n4199), .ZN(n4200) );
  AND2_X1 U5145 ( .A1(n4194), .A2(n4200), .ZN(n4209) );
  NAND2_X1 U5146 ( .A1(n4238), .A2(n4201), .ZN(n4203) );
  AOI22_X1 U5147 ( .A1(n4203), .A2(n3920), .B1(n4202), .B2(n5307), .ZN(n4206)
         );
  NAND2_X1 U5148 ( .A1(n4244), .A2(n4348), .ZN(n4204) );
  AND4_X1 U5149 ( .A1(n4206), .A2(n3185), .A3(n4205), .A4(n4204), .ZN(n4207)
         );
  AND2_X1 U5150 ( .A1(n4208), .A2(n4207), .ZN(n4267) );
  NAND2_X1 U5151 ( .A1(n4209), .A2(n4267), .ZN(n4550) );
  INV_X1 U5152 ( .A(n4550), .ZN(n6453) );
  AND2_X1 U5153 ( .A1(n4210), .A2(n3926), .ZN(n6454) );
  INV_X1 U5154 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4233) );
  NOR3_X1 U5155 ( .A1(n6452), .A2(n5499), .A3(n4212), .ZN(n4213) );
  AOI21_X1 U5156 ( .B1(n6454), .B2(n4233), .A(n4213), .ZN(n4214) );
  OAI21_X1 U5157 ( .B1(n6137), .B2(n6453), .A(n4214), .ZN(n6457) );
  INV_X1 U5158 ( .A(n6579), .ZN(n6574) );
  INV_X1 U5159 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5441) );
  AOI22_X1 U5160 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5441), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4215), .ZN(n5502) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5503) );
  NOR2_X1 U5162 ( .A1(n6571), .A2(n5503), .ZN(n4217) );
  AOI222_X1 U5163 ( .A1(n6457), .A2(n6574), .B1(n5502), .B2(n4217), .C1(n4216), 
        .C2(n5500), .ZN(n4235) );
  INV_X1 U5164 ( .A(n4218), .ZN(n5523) );
  OR2_X1 U5165 ( .A1(n4219), .A2(n5523), .ZN(n4256) );
  OR2_X1 U5166 ( .A1(n5524), .A2(n4256), .ZN(n4223) );
  INV_X1 U5167 ( .A(n4194), .ZN(n4221) );
  NOR2_X1 U5168 ( .A1(n4220), .A2(READY_N), .ZN(n4248) );
  NAND2_X1 U5169 ( .A1(n4221), .A2(n4248), .ZN(n4222) );
  NAND2_X1 U5170 ( .A1(n4223), .A2(n4222), .ZN(n4298) );
  INV_X1 U5171 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U5172 ( .A1(n4224), .A2(n6507), .ZN(n6596) );
  INV_X1 U5173 ( .A(n6596), .ZN(n5525) );
  INV_X1 U5174 ( .A(n4196), .ZN(n4226) );
  NAND2_X1 U5175 ( .A1(n5530), .A2(n6596), .ZN(n4225) );
  AOI22_X1 U5176 ( .A1(n6454), .A2(n5525), .B1(n4226), .B2(n4225), .ZN(n4227)
         );
  OR2_X1 U5177 ( .A1(n4227), .A2(READY_N), .ZN(n4230) );
  NAND2_X1 U5178 ( .A1(n5524), .A2(n4228), .ZN(n4252) );
  OAI211_X1 U5179 ( .C1(n5524), .C2(n4230), .A(n4252), .B(n4229), .ZN(n4231)
         );
  NOR2_X1 U5180 ( .A1(n6571), .A2(n4987), .ZN(n4580) );
  NAND2_X1 U5181 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4580), .ZN(n6568) );
  INV_X1 U5182 ( .A(n6568), .ZN(n4232) );
  AOI22_X1 U5183 ( .A1(n6458), .A2(n5528), .B1(FLUSH_REG_SCAN_IN), .B2(n4232), 
        .ZN(n5990) );
  NAND2_X1 U5184 ( .A1(n6599), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U5185 ( .A1(n5990), .A2(n6569), .ZN(n6576) );
  INV_X1 U5186 ( .A(n6576), .ZN(n5508) );
  NOR2_X1 U5187 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6483), .ZN(n6573)
         );
  INV_X1 U5188 ( .A(n4233), .ZN(n4551) );
  OAI21_X1 U5189 ( .B1(n5508), .B2(n6573), .A(n4551), .ZN(n4234) );
  OAI21_X1 U5190 ( .B1(n4235), .B2(n5508), .A(n4234), .ZN(U3460) );
  INV_X1 U5191 ( .A(n4236), .ZN(n4237) );
  AOI21_X1 U5192 ( .B1(n4238), .B2(n5503), .A(n4237), .ZN(n5193) );
  INV_X1 U5193 ( .A(n5193), .ZN(n4241) );
  XOR2_X1 U5194 ( .A(n4240), .B(n4239), .Z(n5187) );
  INV_X1 U5195 ( .A(n5187), .ZN(n4408) );
  OAI222_X1 U5196 ( .A1(n4241), .A2(n5670), .B1(n5677), .B2(n4408), .C1(n5190), 
        .C2(n5669), .ZN(U2859) );
  XNOR2_X1 U5197 ( .A(n4242), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4283)
         );
  NAND2_X1 U5198 ( .A1(n4243), .A2(n6596), .ZN(n5063) );
  INV_X1 U5199 ( .A(READY_N), .ZN(n6603) );
  NAND2_X1 U5200 ( .A1(n5063), .A2(n6603), .ZN(n4245) );
  OAI211_X1 U5201 ( .C1(n4196), .C2(n4245), .A(n5072), .B(n4244), .ZN(n4247)
         );
  NAND2_X1 U5202 ( .A1(n4247), .A2(n4246), .ZN(n4255) );
  NAND2_X1 U5203 ( .A1(n3926), .A2(n6596), .ZN(n4249) );
  NAND3_X1 U5204 ( .A1(n4249), .A2(n4248), .A3(n4348), .ZN(n4250) );
  NAND3_X1 U5205 ( .A1(n4252), .A2(n4251), .A3(n4250), .ZN(n4253) );
  NAND2_X1 U5206 ( .A1(n4253), .A2(n5528), .ZN(n4254) );
  INV_X1 U5207 ( .A(n4256), .ZN(n4546) );
  OR2_X1 U5208 ( .A1(n4546), .A2(n6472), .ZN(n5512) );
  INV_X1 U5209 ( .A(n5512), .ZN(n4260) );
  OAI22_X1 U5210 ( .A1(n4196), .A2(n5530), .B1(n4257), .B2(n4273), .ZN(n4258)
         );
  INV_X1 U5211 ( .A(n4258), .ZN(n4259) );
  NAND3_X1 U5212 ( .A1(n4260), .A2(n4259), .A3(n4194), .ZN(n4261) );
  NAND2_X1 U5213 ( .A1(n4275), .A2(n4261), .ZN(n6342) );
  NAND2_X1 U5214 ( .A1(n4275), .A2(n5514), .ZN(n5362) );
  INV_X1 U5215 ( .A(n5362), .ZN(n6333) );
  OAI22_X1 U5216 ( .A1(n4296), .A2(n4264), .B1(n4263), .B2(n4262), .ZN(n4265)
         );
  INV_X1 U5217 ( .A(n4265), .ZN(n4266) );
  OR3_X1 U5218 ( .A1(n6452), .A2(n5072), .A3(n4364), .ZN(n4554) );
  NAND3_X1 U5219 ( .A1(n4267), .A2(n4266), .A3(n4554), .ZN(n4268) );
  AND2_X1 U5220 ( .A1(n4275), .A2(n4268), .ZN(n5977) );
  NOR2_X1 U5221 ( .A1(n6333), .A2(n5977), .ZN(n5972) );
  INV_X1 U5222 ( .A(n5972), .ZN(n4271) );
  NAND2_X1 U5223 ( .A1(n5977), .A2(n5503), .ZN(n4270) );
  OR2_X1 U5224 ( .A1(n4275), .A2(n6336), .ZN(n4269) );
  AND2_X1 U5225 ( .A1(n4270), .A2(n4269), .ZN(n5347) );
  OAI21_X1 U5226 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5362), .A(n5347), 
        .ZN(n4384) );
  OAI22_X1 U5227 ( .A1(n4271), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n5975), 
        .B2(n4384), .ZN(n4277) );
  OR2_X1 U5228 ( .A1(n4196), .A2(n4272), .ZN(n6479) );
  OAI21_X1 U5229 ( .B1(n4273), .B2(n3109), .A(n6479), .ZN(n4274) );
  NAND2_X1 U5230 ( .A1(n4275), .A2(n4274), .ZN(n6283) );
  AND2_X1 U5231 ( .A1(n6336), .A2(REIP_REG_0__SCAN_IN), .ZN(n4280) );
  AOI21_X1 U5232 ( .B1(n6338), .B2(n5193), .A(n4280), .ZN(n4276) );
  OAI211_X1 U5233 ( .C1(n4283), .C2(n6342), .A(n4277), .B(n4276), .ZN(U3018)
         );
  INV_X1 U5234 ( .A(n4278), .ZN(n4279) );
  OAI21_X1 U5235 ( .B1(n6236), .B2(n4279), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4282) );
  INV_X2 U5236 ( .A(n5406), .ZN(n6225) );
  AOI21_X1 U5237 ( .B1(n5187), .B2(n6225), .A(n4280), .ZN(n4281) );
  OAI211_X1 U5238 ( .C1(n4283), .C2(n6229), .A(n4282), .B(n4281), .ZN(U2986)
         );
  OAI21_X1 U5239 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n5017) );
  INV_X1 U5240 ( .A(n4287), .ZN(n4288) );
  NAND2_X1 U5241 ( .A1(n4288), .A2(n5530), .ZN(n4289) );
  AND2_X1 U5242 ( .A1(n4290), .A2(n4289), .ZN(n6146) );
  INV_X1 U5243 ( .A(n6146), .ZN(n4291) );
  AOI22_X1 U5244 ( .A1(n5675), .A2(n4291), .B1(EBX_REG_1__SCAN_IN), .B2(n5674), 
        .ZN(n4292) );
  OAI21_X1 U5245 ( .B1(n5677), .B2(n5017), .A(n4292), .ZN(U2858) );
  OR2_X1 U5246 ( .A1(n5522), .A2(READY_N), .ZN(n4293) );
  NOR2_X1 U5247 ( .A1(n4294), .A2(n4293), .ZN(n4316) );
  NAND2_X1 U5248 ( .A1(n4316), .A2(n3926), .ZN(n6196) );
  NOR2_X1 U5249 ( .A1(n4296), .A2(n4295), .ZN(n4297) );
  OAI21_X1 U5250 ( .B1(n4298), .B2(n4297), .A(n5528), .ZN(n4299) );
  NAND2_X1 U5251 ( .A1(n3171), .A2(n5279), .ZN(n4300) );
  INV_X1 U5252 ( .A(n4300), .ZN(n4301) );
  INV_X1 U5253 ( .A(n5689), .ZN(n4672) );
  INV_X1 U5254 ( .A(DATAI_1_), .ZN(n4357) );
  INV_X1 U5255 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6183) );
  OAI222_X1 U5256 ( .A1(n5017), .A2(n5917), .B1(n4672), .B2(n4357), .C1(n5453), 
        .C2(n6183), .ZN(U2890) );
  OAI21_X1 U5257 ( .B1(n4303), .B2(n4302), .A(n4310), .ZN(n6248) );
  CLKBUF_X1 U5258 ( .A(n4304), .Z(n4312) );
  INV_X1 U5259 ( .A(n4312), .ZN(n4305) );
  AOI21_X1 U5260 ( .B1(n4307), .B2(n4306), .A(n4305), .ZN(n6337) );
  AOI22_X1 U5261 ( .A1(n5675), .A2(n6337), .B1(EBX_REG_2__SCAN_IN), .B2(n5674), 
        .ZN(n4308) );
  OAI21_X1 U5262 ( .B1(n6248), .B2(n5677), .A(n4308), .ZN(U2857) );
  INV_X1 U5263 ( .A(DATAI_2_), .ZN(n4349) );
  INV_X1 U5264 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6752) );
  OAI222_X1 U5265 ( .A1(n6248), .A2(n5917), .B1(n4672), .B2(n4349), .C1(n5453), 
        .C2(n6752), .ZN(U2889) );
  XNOR2_X1 U5266 ( .A(n4310), .B(n4309), .ZN(n5157) );
  AOI21_X1 U5267 ( .B1(n4313), .B2(n4312), .A(n4311), .ZN(n6322) );
  AOI22_X1 U5268 ( .A1(n5675), .A2(n6322), .B1(EBX_REG_3__SCAN_IN), .B2(n5674), 
        .ZN(n4314) );
  OAI21_X1 U5269 ( .B1(n5157), .B2(n5677), .A(n4314), .ZN(U2856) );
  INV_X1 U5270 ( .A(n6479), .ZN(n4315) );
  INV_X1 U5271 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4791) );
  NOR2_X2 U5272 ( .A1(n6211), .A2(n4316), .ZN(n6210) );
  NAND2_X1 U5273 ( .A1(n6210), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4317) );
  NAND2_X1 U5274 ( .A1(n6214), .A2(DATAI_6_), .ZN(n4847) );
  OAI211_X1 U5275 ( .C1(n6217), .C2(n4791), .A(n4317), .B(n4847), .ZN(U2930)
         );
  INV_X1 U5276 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4319) );
  NAND2_X1 U5277 ( .A1(n6210), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U5278 ( .A1(n6214), .A2(DATAI_0_), .ZN(n4856) );
  OAI211_X1 U5279 ( .C1(n6217), .C2(n4319), .A(n4318), .B(n4856), .ZN(U2939)
         );
  NAND2_X1 U5280 ( .A1(n6210), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U5281 ( .A1(n6214), .A2(DATAI_1_), .ZN(n4845) );
  OAI211_X1 U5282 ( .C1(n6217), .C2(n6183), .A(n4320), .B(n4845), .ZN(U2940)
         );
  INV_X1 U5283 ( .A(DATAI_3_), .ZN(n4366) );
  INV_X1 U5284 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6180) );
  OAI222_X1 U5285 ( .A1(n5917), .A2(n5157), .B1(n4672), .B2(n4366), .C1(n5453), 
        .C2(n6180), .ZN(U2888) );
  AND2_X1 U5286 ( .A1(n3337), .A2(n5837), .ZN(n4323) );
  AND2_X1 U5287 ( .A1(n5841), .A2(n4323), .ZN(n4333) );
  AND2_X1 U5288 ( .A1(n4333), .A2(n4722), .ZN(n4931) );
  NAND2_X1 U5289 ( .A1(n6225), .A2(DATAI_23_), .ZN(n6399) );
  NAND2_X1 U5290 ( .A1(n6225), .A2(DATAI_31_), .ZN(n6451) );
  INV_X1 U5291 ( .A(n6451), .ZN(n6395) );
  NAND2_X1 U5292 ( .A1(n5837), .A2(n4888), .ZN(n4638) );
  NOR2_X1 U5293 ( .A1(n4638), .A2(n4454), .ZN(n4325) );
  NAND2_X1 U5294 ( .A1(n4325), .A2(n5841), .ZN(n4499) );
  INV_X1 U5295 ( .A(n6569), .ZN(n4326) );
  NOR2_X1 U5296 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5993) );
  NAND2_X1 U5297 ( .A1(n4365), .A2(n5279), .ZN(n5099) );
  INV_X1 U5298 ( .A(n4328), .ZN(n4688) );
  NAND2_X1 U5299 ( .A1(n4632), .A2(n4688), .ZN(n4715) );
  AND2_X1 U5300 ( .A1(n4192), .A2(n5205), .ZN(n4599) );
  INV_X1 U5301 ( .A(n4599), .ZN(n6353) );
  OR2_X1 U5302 ( .A1(n4715), .A2(n6353), .ZN(n4330) );
  NAND2_X1 U5303 ( .A1(n4330), .A2(n4368), .ZN(n4334) );
  AOI22_X1 U5304 ( .A1(n4334), .A2(n5836), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4501), .ZN(n4367) );
  INV_X1 U5305 ( .A(DATAI_7_), .ZN(n4393) );
  NOR2_X1 U5306 ( .A1(n4393), .A2(n4572), .ZN(n6446) );
  INV_X1 U5307 ( .A(n6446), .ZN(n5098) );
  OAI22_X1 U5308 ( .A1(n5099), .A2(n4368), .B1(n4367), .B2(n5098), .ZN(n4332)
         );
  AOI21_X1 U5309 ( .B1(n6395), .B2(n4533), .A(n4332), .ZN(n4339) );
  NAND2_X1 U5310 ( .A1(n5836), .A2(n6593), .ZN(n5088) );
  OAI21_X1 U5311 ( .B1(n4333), .B2(n5406), .A(n5088), .ZN(n4336) );
  INV_X1 U5312 ( .A(n4334), .ZN(n4335) );
  NAND2_X1 U5313 ( .A1(n4336), .A2(n4335), .ZN(n4337) );
  AOI21_X1 U5314 ( .B1(n6455), .B2(STATE2_REG_3__SCAN_IN), .A(n4572), .ZN(
        n4751) );
  OAI211_X1 U5315 ( .C1(n4501), .C2(n5836), .A(n4337), .B(n4751), .ZN(n4370)
         );
  NAND2_X1 U5316 ( .A1(n4370), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4338)
         );
  OAI211_X1 U5317 ( .C1(n4972), .C2(n6399), .A(n4339), .B(n4338), .ZN(U3147)
         );
  NAND2_X1 U5318 ( .A1(n6225), .A2(DATAI_21_), .ZN(n6388) );
  INV_X1 U5319 ( .A(DATAI_29_), .ZN(n4340) );
  NOR2_X1 U5320 ( .A1(n5406), .A2(n4340), .ZN(n6385) );
  NAND2_X1 U5321 ( .A1(n4365), .A2(n3196), .ZN(n5139) );
  INV_X1 U5322 ( .A(DATAI_5_), .ZN(n4418) );
  NOR2_X1 U5323 ( .A1(n4418), .A2(n4572), .ZN(n6383) );
  INV_X1 U5324 ( .A(n6383), .ZN(n5136) );
  OAI22_X1 U5325 ( .A1(n5139), .A2(n4368), .B1(n4367), .B2(n5136), .ZN(n4341)
         );
  AOI21_X1 U5326 ( .B1(n6385), .B2(n4533), .A(n4341), .ZN(n4343) );
  NAND2_X1 U5327 ( .A1(n4370), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4342)
         );
  OAI211_X1 U5328 ( .C1(n4972), .C2(n6388), .A(n4343), .B(n4342), .ZN(U3145)
         );
  NAND2_X1 U5329 ( .A1(n6225), .A2(DATAI_16_), .ZN(n6366) );
  INV_X1 U5330 ( .A(DATAI_24_), .ZN(n4344) );
  NOR2_X1 U5331 ( .A1(n5406), .A2(n4344), .ZN(n6363) );
  NAND2_X1 U5332 ( .A1(n4365), .A2(n5072), .ZN(n5124) );
  INV_X1 U5333 ( .A(DATAI_0_), .ZN(n4407) );
  NOR2_X1 U5334 ( .A1(n4407), .A2(n4572), .ZN(n6355) );
  INV_X1 U5335 ( .A(n6355), .ZN(n5123) );
  OAI22_X1 U5336 ( .A1(n5124), .A2(n4368), .B1(n4367), .B2(n5123), .ZN(n4345)
         );
  AOI21_X1 U5337 ( .B1(n6363), .B2(n4533), .A(n4345), .ZN(n4347) );
  NAND2_X1 U5338 ( .A1(n4370), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4346)
         );
  OAI211_X1 U5339 ( .C1(n4972), .C2(n6366), .A(n4347), .B(n4346), .ZN(U3140)
         );
  NAND2_X1 U5340 ( .A1(n6225), .A2(DATAI_18_), .ZN(n6374) );
  NAND2_X1 U5341 ( .A1(n6225), .A2(DATAI_26_), .ZN(n6422) );
  INV_X1 U5342 ( .A(n6422), .ZN(n6371) );
  NAND2_X1 U5343 ( .A1(n4365), .A2(n4348), .ZN(n5109) );
  NOR2_X1 U5344 ( .A1(n4349), .A2(n4572), .ZN(n6419) );
  INV_X1 U5345 ( .A(n6419), .ZN(n5108) );
  OAI22_X1 U5346 ( .A1(n5109), .A2(n4368), .B1(n4367), .B2(n5108), .ZN(n4350)
         );
  AOI21_X1 U5347 ( .B1(n6371), .B2(n4533), .A(n4350), .ZN(n4352) );
  NAND2_X1 U5348 ( .A1(n4370), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4351)
         );
  OAI211_X1 U5349 ( .C1(n4972), .C2(n6374), .A(n4352), .B(n4351), .ZN(U3142)
         );
  NAND2_X1 U5350 ( .A1(n6225), .A2(DATAI_22_), .ZN(n6392) );
  NAND2_X1 U5351 ( .A1(n6225), .A2(DATAI_30_), .ZN(n6440) );
  INV_X1 U5352 ( .A(n6440), .ZN(n6389) );
  NAND2_X1 U5353 ( .A1(n4365), .A2(n4353), .ZN(n5104) );
  INV_X1 U5354 ( .A(DATAI_6_), .ZN(n4671) );
  NOR2_X1 U5355 ( .A1(n4671), .A2(n4572), .ZN(n6437) );
  INV_X1 U5356 ( .A(n6437), .ZN(n5103) );
  OAI22_X1 U5357 ( .A1(n5104), .A2(n4368), .B1(n4367), .B2(n5103), .ZN(n4354)
         );
  AOI21_X1 U5358 ( .B1(n6389), .B2(n4533), .A(n4354), .ZN(n4356) );
  NAND2_X1 U5359 ( .A1(n4370), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4355)
         );
  OAI211_X1 U5360 ( .C1(n4972), .C2(n6392), .A(n4356), .B(n4355), .ZN(U3146)
         );
  NAND2_X1 U5361 ( .A1(n6225), .A2(DATAI_17_), .ZN(n6370) );
  NAND2_X1 U5362 ( .A1(n6225), .A2(DATAI_25_), .ZN(n6416) );
  INV_X1 U5363 ( .A(n6416), .ZN(n6367) );
  NAND2_X1 U5364 ( .A1(n4365), .A2(n3926), .ZN(n5131) );
  NOR2_X1 U5365 ( .A1(n4357), .A2(n4572), .ZN(n6413) );
  INV_X1 U5366 ( .A(n6413), .ZN(n5130) );
  OAI22_X1 U5367 ( .A1(n5131), .A2(n4368), .B1(n4367), .B2(n5130), .ZN(n4358)
         );
  AOI21_X1 U5368 ( .B1(n6367), .B2(n4533), .A(n4358), .ZN(n4360) );
  NAND2_X1 U5369 ( .A1(n4370), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4359)
         );
  OAI211_X1 U5370 ( .C1(n4972), .C2(n6370), .A(n4360), .B(n4359), .ZN(U3141)
         );
  NAND2_X1 U5371 ( .A1(n6225), .A2(DATAI_20_), .ZN(n6382) );
  NAND2_X1 U5372 ( .A1(n6225), .A2(DATAI_28_), .ZN(n6434) );
  INV_X1 U5373 ( .A(n6434), .ZN(n6379) );
  NAND2_X1 U5374 ( .A1(n4365), .A2(n3109), .ZN(n5114) );
  INV_X1 U5375 ( .A(DATAI_4_), .ZN(n4406) );
  NOR2_X1 U5376 ( .A1(n4406), .A2(n4572), .ZN(n6431) );
  INV_X1 U5377 ( .A(n6431), .ZN(n5113) );
  OAI22_X1 U5378 ( .A1(n5114), .A2(n4368), .B1(n4367), .B2(n5113), .ZN(n4361)
         );
  AOI21_X1 U5379 ( .B1(n6379), .B2(n4533), .A(n4361), .ZN(n4363) );
  NAND2_X1 U5380 ( .A1(n4370), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4362)
         );
  OAI211_X1 U5381 ( .C1(n4972), .C2(n6382), .A(n4363), .B(n4362), .ZN(U3144)
         );
  NAND2_X1 U5382 ( .A1(n6225), .A2(DATAI_19_), .ZN(n6378) );
  NAND2_X1 U5383 ( .A1(n6225), .A2(DATAI_27_), .ZN(n6428) );
  INV_X1 U5384 ( .A(n6428), .ZN(n6375) );
  NAND2_X1 U5385 ( .A1(n4365), .A2(n4364), .ZN(n5119) );
  NOR2_X1 U5386 ( .A1(n4366), .A2(n4572), .ZN(n6425) );
  INV_X1 U5387 ( .A(n6425), .ZN(n5118) );
  OAI22_X1 U5388 ( .A1(n5119), .A2(n4368), .B1(n4367), .B2(n5118), .ZN(n4369)
         );
  AOI21_X1 U5389 ( .B1(n6375), .B2(n4533), .A(n4369), .ZN(n4372) );
  NAND2_X1 U5390 ( .A1(n4370), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4371)
         );
  OAI211_X1 U5391 ( .C1(n4972), .C2(n6378), .A(n4372), .B(n4371), .ZN(U3143)
         );
  INV_X1 U5392 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U5393 ( .A1(n4373), .A2(n6454), .ZN(n4374) );
  NAND2_X1 U5394 ( .A1(n6217), .A2(n4374), .ZN(n4375) );
  NAND2_X1 U5395 ( .A1(n6160), .A2(n5072), .ZN(n4800) );
  NAND2_X1 U5396 ( .A1(n4580), .A2(n6599), .ZN(n6476) );
  AOI22_X1 U5398 ( .A1(n6604), .A2(UWORD_REG_9__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U5399 ( .B1(n4377), .B2(n4800), .A(n4376), .ZN(U2898) );
  INV_X1 U5400 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4379) );
  AOI22_X1 U5401 ( .A1(n6604), .A2(UWORD_REG_13__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4378) );
  OAI21_X1 U5402 ( .B1(n4379), .B2(n4800), .A(n4378), .ZN(U2894) );
  INV_X1 U5403 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6194) );
  AOI22_X1 U5404 ( .A1(n6604), .A2(UWORD_REG_11__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4380) );
  OAI21_X1 U5405 ( .B1(n6194), .B2(n4800), .A(n4380), .ZN(U2896) );
  CLKBUF_X1 U5406 ( .A(n4381), .Z(n4383) );
  XNOR2_X1 U5407 ( .A(n4383), .B(n4382), .ZN(n5021) );
  INV_X1 U5408 ( .A(n5345), .ZN(n4680) );
  NAND2_X1 U5409 ( .A1(n4680), .A2(n5362), .ZN(n5957) );
  INV_X1 U5410 ( .A(n5957), .ZN(n5955) );
  NOR2_X1 U5411 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5975), .ZN(n4677)
         );
  NOR2_X1 U5412 ( .A1(n5955), .A2(n4677), .ZN(n4385) );
  MUX2_X1 U5413 ( .A(n4385), .B(n4384), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4387) );
  NOR2_X1 U5414 ( .A1(n6283), .A2(n6146), .ZN(n4386) );
  AOI211_X1 U5415 ( .C1(n6336), .C2(REIP_REG_1__SCAN_IN), .A(n4387), .B(n4386), 
        .ZN(n4388) );
  OAI21_X1 U5416 ( .B1(n5021), .B2(n6342), .A(n4388), .ZN(U3017) );
  INV_X1 U5417 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U5419 ( .A1(n6604), .A2(UWORD_REG_7__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5420 ( .B1(n4390), .B2(n4800), .A(n4389), .ZN(U2900) );
  INV_X1 U5421 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n4392) );
  INV_X1 U5422 ( .A(DATAI_9_), .ZN(n6615) );
  NOR2_X1 U5423 ( .A1(n6196), .A2(n6615), .ZN(n4396) );
  AOI21_X1 U5424 ( .B1(n6211), .B2(EAX_REG_9__SCAN_IN), .A(n4396), .ZN(n4391)
         );
  OAI21_X1 U5425 ( .B1(n4843), .B2(n4392), .A(n4391), .ZN(U2948) );
  INV_X1 U5426 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4395) );
  NOR2_X1 U5427 ( .A1(n6196), .A2(n4393), .ZN(n4399) );
  AOI21_X1 U5428 ( .B1(n6211), .B2(EAX_REG_23__SCAN_IN), .A(n4399), .ZN(n4394)
         );
  OAI21_X1 U5429 ( .B1(n4843), .B2(n4395), .A(n4394), .ZN(U2931) );
  INV_X1 U5430 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n4398) );
  AOI21_X1 U5431 ( .B1(n6211), .B2(EAX_REG_25__SCAN_IN), .A(n4396), .ZN(n4397)
         );
  OAI21_X1 U5432 ( .B1(n4843), .B2(n4398), .A(n4397), .ZN(U2933) );
  INV_X1 U5433 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4401) );
  AOI21_X1 U5434 ( .B1(n6211), .B2(EAX_REG_7__SCAN_IN), .A(n4399), .ZN(n4400)
         );
  OAI21_X1 U5435 ( .B1(n4843), .B2(n4401), .A(n4400), .ZN(U2946) );
  CLKBUF_X1 U5436 ( .A(n4402), .Z(n4413) );
  OR2_X1 U5437 ( .A1(n4404), .A2(n4403), .ZN(n4405) );
  AND2_X1 U5438 ( .A1(n4413), .A2(n4405), .ZN(n6241) );
  INV_X1 U5439 ( .A(n6241), .ZN(n6126) );
  OAI222_X1 U5440 ( .A1(n6126), .A2(n5917), .B1(n4672), .B2(n4406), .C1(n5453), 
        .C2(n4866), .ZN(U2887) );
  OAI222_X1 U5441 ( .A1(n5917), .A2(n4408), .B1(n4672), .B2(n4407), .C1(n5453), 
        .C2(n4319), .ZN(U2891) );
  OR2_X1 U5442 ( .A1(n4311), .A2(n4410), .ZN(n4411) );
  NAND2_X1 U5443 ( .A1(n4409), .A2(n4411), .ZN(n6313) );
  INV_X1 U5444 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U5445 ( .A1(n6313), .A2(n5670), .B1(n5669), .B2(n6766), .C1(n6126), 
        .C2(n5677), .ZN(U2855) );
  INV_X1 U5446 ( .A(n4620), .ZN(n4412) );
  AOI21_X1 U5447 ( .B1(n4414), .B2(n4413), .A(n4412), .ZN(n5053) );
  INV_X1 U5448 ( .A(n5053), .ZN(n5086) );
  OAI21_X1 U5449 ( .B1(n3964), .B2(n3963), .A(n4623), .ZN(n5082) );
  INV_X1 U5450 ( .A(n5082), .ZN(n6304) );
  AOI22_X1 U5451 ( .A1(n5675), .A2(n6304), .B1(EBX_REG_5__SCAN_IN), .B2(n5674), 
        .ZN(n4417) );
  OAI21_X1 U5452 ( .B1(n5086), .B2(n5677), .A(n4417), .ZN(U2854) );
  OAI222_X1 U5453 ( .A1(n5086), .A2(n5917), .B1(n4672), .B2(n4418), .C1(n5453), 
        .C2(n4861), .ZN(U2886) );
  NAND2_X1 U5454 ( .A1(n5841), .A2(n4454), .ZN(n4607) );
  OAI21_X1 U5455 ( .B1(n4889), .B2(n6593), .A(n5836), .ZN(n4887) );
  NAND2_X1 U5456 ( .A1(n5837), .A2(n4722), .ZN(n4606) );
  NOR2_X1 U5457 ( .A1(n4686), .A2(n4606), .ZN(n4419) );
  NAND2_X1 U5458 ( .A1(n4419), .A2(n4628), .ZN(n4664) );
  INV_X1 U5459 ( .A(n5088), .ZN(n4933) );
  NAND2_X1 U5460 ( .A1(n5205), .A2(n6137), .ZN(n4461) );
  OR2_X1 U5461 ( .A1(n4461), .A2(n4536), .ZN(n4881) );
  OAI21_X1 U5462 ( .B1(n4664), .B2(n4933), .A(n4881), .ZN(n4422) );
  NAND3_X1 U5463 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6466), .A3(n6461), .ZN(n4885) );
  OR2_X1 U5464 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4885), .ZN(n4449)
         );
  NOR2_X1 U5465 ( .A1(n4423), .A2(n4987), .ZN(n6359) );
  INV_X1 U5466 ( .A(n4457), .ZN(n4420) );
  OR2_X1 U5467 ( .A1(n6350), .A2(n4420), .ZN(n4940) );
  INV_X1 U5468 ( .A(n4940), .ZN(n4424) );
  INV_X1 U5469 ( .A(n4572), .ZN(n4500) );
  OAI21_X1 U5470 ( .B1(n4424), .B2(n4987), .A(n4500), .ZN(n4936) );
  AOI211_X1 U5471 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4449), .A(n6359), .B(
        n4936), .ZN(n4421) );
  OAI21_X1 U5472 ( .B1(n4887), .B2(n4422), .A(n4421), .ZN(n4447) );
  NAND2_X1 U5473 ( .A1(n4447), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4428) );
  OR2_X1 U5474 ( .A1(n4632), .A2(n5844), .ZN(n6354) );
  INV_X1 U5475 ( .A(n6354), .ZN(n4425) );
  INV_X1 U5476 ( .A(n4461), .ZN(n4745) );
  AND2_X1 U5477 ( .A1(n4423), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6351) );
  AOI22_X1 U5478 ( .A1(n4425), .A2(n4745), .B1(n4424), .B2(n6351), .ZN(n4448)
         );
  OAI22_X1 U5479 ( .A1(n5109), .A2(n4449), .B1(n4448), .B2(n5108), .ZN(n4426)
         );
  AOI21_X1 U5480 ( .B1(n6371), .B2(n4451), .A(n4426), .ZN(n4427) );
  OAI211_X1 U5481 ( .C1(n4919), .C2(n6374), .A(n4428), .B(n4427), .ZN(U3054)
         );
  NAND2_X1 U5482 ( .A1(n4447), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4431) );
  OAI22_X1 U5483 ( .A1(n5114), .A2(n4449), .B1(n4448), .B2(n5113), .ZN(n4429)
         );
  AOI21_X1 U5484 ( .B1(n6379), .B2(n4451), .A(n4429), .ZN(n4430) );
  OAI211_X1 U5485 ( .C1(n4919), .C2(n6382), .A(n4431), .B(n4430), .ZN(U3056)
         );
  NAND2_X1 U5486 ( .A1(n4447), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4434) );
  OAI22_X1 U5487 ( .A1(n5139), .A2(n4449), .B1(n4448), .B2(n5136), .ZN(n4432)
         );
  AOI21_X1 U5488 ( .B1(n6385), .B2(n4451), .A(n4432), .ZN(n4433) );
  OAI211_X1 U5489 ( .C1(n4919), .C2(n6388), .A(n4434), .B(n4433), .ZN(U3057)
         );
  NAND2_X1 U5490 ( .A1(n4447), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4437) );
  OAI22_X1 U5491 ( .A1(n5131), .A2(n4449), .B1(n4448), .B2(n5130), .ZN(n4435)
         );
  AOI21_X1 U5492 ( .B1(n6367), .B2(n4451), .A(n4435), .ZN(n4436) );
  OAI211_X1 U5493 ( .C1(n4919), .C2(n6370), .A(n4437), .B(n4436), .ZN(U3053)
         );
  NAND2_X1 U5494 ( .A1(n4447), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4440) );
  OAI22_X1 U5495 ( .A1(n5099), .A2(n4449), .B1(n4448), .B2(n5098), .ZN(n4438)
         );
  AOI21_X1 U5496 ( .B1(n6395), .B2(n4451), .A(n4438), .ZN(n4439) );
  OAI211_X1 U5497 ( .C1(n4919), .C2(n6399), .A(n4440), .B(n4439), .ZN(U3059)
         );
  NAND2_X1 U5498 ( .A1(n4447), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4443) );
  OAI22_X1 U5499 ( .A1(n5119), .A2(n4449), .B1(n4448), .B2(n5118), .ZN(n4441)
         );
  AOI21_X1 U5500 ( .B1(n6375), .B2(n4451), .A(n4441), .ZN(n4442) );
  OAI211_X1 U5501 ( .C1(n4919), .C2(n6378), .A(n4443), .B(n4442), .ZN(U3055)
         );
  NAND2_X1 U5502 ( .A1(n4447), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4446) );
  OAI22_X1 U5503 ( .A1(n5104), .A2(n4449), .B1(n4448), .B2(n5103), .ZN(n4444)
         );
  AOI21_X1 U5504 ( .B1(n6389), .B2(n4451), .A(n4444), .ZN(n4445) );
  OAI211_X1 U5505 ( .C1(n4919), .C2(n6392), .A(n4446), .B(n4445), .ZN(U3058)
         );
  NAND2_X1 U5506 ( .A1(n4447), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4453) );
  OAI22_X1 U5507 ( .A1(n5124), .A2(n4449), .B1(n4448), .B2(n5123), .ZN(n4450)
         );
  AOI21_X1 U5508 ( .B1(n6363), .B2(n4451), .A(n4450), .ZN(n4452) );
  OAI211_X1 U5509 ( .C1(n4919), .C2(n6366), .A(n4453), .B(n4452), .ZN(U3052)
         );
  OR2_X1 U5510 ( .A1(n4714), .A2(n4606), .ZN(n4460) );
  NOR2_X1 U5511 ( .A1(n5837), .A2(n4454), .ZN(n4455) );
  NAND2_X1 U5512 ( .A1(n5841), .A2(n4455), .ZN(n4574) );
  AOI21_X1 U5513 ( .B1(n4460), .B2(n4743), .A(n6593), .ZN(n4456) );
  AOI211_X1 U5514 ( .C1(n4745), .C2(n4632), .A(n5844), .B(n4456), .ZN(n4459)
         );
  NOR3_X1 U5515 ( .A1(n4716), .A2(n6466), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4753) );
  INV_X1 U5516 ( .A(n4753), .ZN(n4747) );
  NOR2_X1 U5517 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4747), .ZN(n4492)
         );
  INV_X1 U5518 ( .A(n6359), .ZN(n5095) );
  OR2_X1 U5519 ( .A1(n6350), .A2(n4457), .ZN(n4803) );
  AOI21_X1 U5520 ( .B1(n4803), .B2(STATE2_REG_2__SCAN_IN), .A(n4572), .ZN(
        n4807) );
  OAI211_X1 U5521 ( .C1(n3174), .C2(n4492), .A(n5095), .B(n4807), .ZN(n4458)
         );
  INV_X1 U5522 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4466) );
  INV_X1 U5523 ( .A(n5139), .ZN(n6384) );
  INV_X1 U5524 ( .A(n4632), .ZN(n5153) );
  NOR2_X1 U5525 ( .A1(n5153), .A2(n5844), .ZN(n4805) );
  INV_X1 U5526 ( .A(n4805), .ZN(n4462) );
  INV_X1 U5527 ( .A(n6351), .ZN(n4808) );
  OAI22_X1 U5528 ( .A1(n4462), .A2(n4461), .B1(n4808), .B2(n4803), .ZN(n4491)
         );
  AOI22_X1 U5529 ( .A1(n6384), .A2(n4492), .B1(n6383), .B2(n4491), .ZN(n4463)
         );
  OAI21_X1 U5530 ( .B1(n6388), .B2(n4743), .A(n4463), .ZN(n4464) );
  AOI21_X1 U5531 ( .B1(n6385), .B2(n6441), .A(n4464), .ZN(n4465) );
  OAI21_X1 U5532 ( .B1(n4497), .B2(n4466), .A(n4465), .ZN(U3121) );
  INV_X1 U5533 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4470) );
  INV_X1 U5534 ( .A(n5119), .ZN(n6424) );
  AOI22_X1 U5535 ( .A1(n6424), .A2(n4492), .B1(n6425), .B2(n4491), .ZN(n4467)
         );
  OAI21_X1 U5536 ( .B1(n6378), .B2(n4743), .A(n4467), .ZN(n4468) );
  AOI21_X1 U5537 ( .B1(n6375), .B2(n6441), .A(n4468), .ZN(n4469) );
  OAI21_X1 U5538 ( .B1(n4497), .B2(n4470), .A(n4469), .ZN(U3119) );
  INV_X1 U5539 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4474) );
  INV_X1 U5540 ( .A(n5114), .ZN(n6430) );
  AOI22_X1 U5541 ( .A1(n6430), .A2(n4492), .B1(n6431), .B2(n4491), .ZN(n4471)
         );
  OAI21_X1 U5542 ( .B1(n6382), .B2(n4743), .A(n4471), .ZN(n4472) );
  AOI21_X1 U5543 ( .B1(n6379), .B2(n6441), .A(n4472), .ZN(n4473) );
  OAI21_X1 U5544 ( .B1(n4497), .B2(n4474), .A(n4473), .ZN(U3120) );
  INV_X1 U5545 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4478) );
  INV_X1 U5546 ( .A(n5131), .ZN(n6412) );
  AOI22_X1 U5547 ( .A1(n6412), .A2(n4492), .B1(n6413), .B2(n4491), .ZN(n4475)
         );
  OAI21_X1 U5548 ( .B1(n6370), .B2(n4743), .A(n4475), .ZN(n4476) );
  AOI21_X1 U5549 ( .B1(n6367), .B2(n6441), .A(n4476), .ZN(n4477) );
  OAI21_X1 U5550 ( .B1(n4497), .B2(n4478), .A(n4477), .ZN(U3117) );
  INV_X1 U5551 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4482) );
  INV_X1 U5552 ( .A(n5109), .ZN(n6418) );
  AOI22_X1 U5553 ( .A1(n6418), .A2(n4492), .B1(n6419), .B2(n4491), .ZN(n4479)
         );
  OAI21_X1 U5554 ( .B1(n6374), .B2(n4743), .A(n4479), .ZN(n4480) );
  AOI21_X1 U5555 ( .B1(n6371), .B2(n6441), .A(n4480), .ZN(n4481) );
  OAI21_X1 U5556 ( .B1(n4497), .B2(n4482), .A(n4481), .ZN(U3118) );
  INV_X1 U5557 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4486) );
  INV_X1 U5558 ( .A(n5104), .ZN(n6436) );
  AOI22_X1 U5559 ( .A1(n6436), .A2(n4492), .B1(n6437), .B2(n4491), .ZN(n4483)
         );
  OAI21_X1 U5560 ( .B1(n6392), .B2(n4743), .A(n4483), .ZN(n4484) );
  AOI21_X1 U5561 ( .B1(n6389), .B2(n6441), .A(n4484), .ZN(n4485) );
  OAI21_X1 U5562 ( .B1(n4497), .B2(n4486), .A(n4485), .ZN(U3122) );
  INV_X1 U5563 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4490) );
  INV_X1 U5564 ( .A(n5099), .ZN(n6444) );
  AOI22_X1 U5565 ( .A1(n6444), .A2(n4492), .B1(n6446), .B2(n4491), .ZN(n4487)
         );
  OAI21_X1 U5566 ( .B1(n6399), .B2(n4743), .A(n4487), .ZN(n4488) );
  AOI21_X1 U5567 ( .B1(n6395), .B2(n6441), .A(n4488), .ZN(n4489) );
  OAI21_X1 U5568 ( .B1(n4497), .B2(n4490), .A(n4489), .ZN(U3123) );
  INV_X1 U5569 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4496) );
  INV_X1 U5570 ( .A(n5124), .ZN(n6356) );
  AOI22_X1 U5571 ( .A1(n6356), .A2(n4492), .B1(n6355), .B2(n4491), .ZN(n4493)
         );
  OAI21_X1 U5572 ( .B1(n6366), .B2(n4743), .A(n4493), .ZN(n4494) );
  AOI21_X1 U5573 ( .B1(n6363), .B2(n6441), .A(n4494), .ZN(n4495) );
  OAI21_X1 U5574 ( .B1(n4497), .B2(n4496), .A(n4495), .ZN(U3116) );
  INV_X1 U5575 ( .A(n4574), .ZN(n4498) );
  AOI21_X1 U5576 ( .B1(n4782), .B2(n4499), .A(n6593), .ZN(n4506) );
  NOR2_X1 U5577 ( .A1(n4599), .A2(n5844), .ZN(n6361) );
  INV_X1 U5578 ( .A(n6361), .ZN(n4505) );
  OAI21_X1 U5579 ( .B1(n6350), .B2(n4987), .A(n4500), .ZN(n6358) );
  NOR2_X1 U5580 ( .A1(n6359), .A2(n6358), .ZN(n4504) );
  INV_X1 U5581 ( .A(n4501), .ZN(n4502) );
  OR2_X1 U5582 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4502), .ZN(n4531)
         );
  AOI21_X1 U5583 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4531), .A(n6466), .ZN(
        n4503) );
  OAI211_X1 U5584 ( .C1(n4506), .C2(n4505), .A(n4504), .B(n4503), .ZN(n4529)
         );
  NAND2_X1 U5585 ( .A1(n4529), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4510)
         );
  INV_X1 U5586 ( .A(n6392), .ZN(n6435) );
  NOR2_X1 U5587 ( .A1(n4808), .A2(n6466), .ZN(n4507) );
  AOI22_X1 U5588 ( .A1(n4805), .A2(n4599), .B1(n6350), .B2(n4507), .ZN(n4530)
         );
  OAI22_X1 U5589 ( .A1(n5104), .A2(n4531), .B1(n4530), .B2(n5103), .ZN(n4508)
         );
  AOI21_X1 U5590 ( .B1(n6435), .B2(n4533), .A(n4508), .ZN(n4509) );
  OAI211_X1 U5591 ( .C1(n4782), .C2(n6440), .A(n4510), .B(n4509), .ZN(U3138)
         );
  NAND2_X1 U5592 ( .A1(n4529), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4513)
         );
  INV_X1 U5593 ( .A(n6378), .ZN(n6423) );
  OAI22_X1 U5594 ( .A1(n5119), .A2(n4531), .B1(n4530), .B2(n5118), .ZN(n4511)
         );
  AOI21_X1 U5595 ( .B1(n6423), .B2(n4533), .A(n4511), .ZN(n4512) );
  OAI211_X1 U5596 ( .C1(n4782), .C2(n6428), .A(n4513), .B(n4512), .ZN(U3135)
         );
  NAND2_X1 U5597 ( .A1(n4529), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4516)
         );
  INV_X1 U5598 ( .A(n6382), .ZN(n6429) );
  OAI22_X1 U5599 ( .A1(n5114), .A2(n4531), .B1(n4530), .B2(n5113), .ZN(n4514)
         );
  AOI21_X1 U5600 ( .B1(n6429), .B2(n4533), .A(n4514), .ZN(n4515) );
  OAI211_X1 U5601 ( .C1(n4782), .C2(n6434), .A(n4516), .B(n4515), .ZN(U3136)
         );
  INV_X1 U5602 ( .A(n6385), .ZN(n5145) );
  NAND2_X1 U5603 ( .A1(n4529), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4519)
         );
  INV_X1 U5604 ( .A(n6388), .ZN(n5142) );
  OAI22_X1 U5605 ( .A1(n5139), .A2(n4531), .B1(n4530), .B2(n5136), .ZN(n4517)
         );
  AOI21_X1 U5606 ( .B1(n5142), .B2(n4533), .A(n4517), .ZN(n4518) );
  OAI211_X1 U5607 ( .C1(n4782), .C2(n5145), .A(n4519), .B(n4518), .ZN(U3137)
         );
  INV_X1 U5608 ( .A(n6363), .ZN(n5129) );
  NAND2_X1 U5609 ( .A1(n4529), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4522)
         );
  INV_X1 U5610 ( .A(n6366), .ZN(n5126) );
  OAI22_X1 U5611 ( .A1(n5124), .A2(n4531), .B1(n4530), .B2(n5123), .ZN(n4520)
         );
  AOI21_X1 U5612 ( .B1(n5126), .B2(n4533), .A(n4520), .ZN(n4521) );
  OAI211_X1 U5613 ( .C1(n4782), .C2(n5129), .A(n4522), .B(n4521), .ZN(U3132)
         );
  NAND2_X1 U5614 ( .A1(n4529), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4525)
         );
  INV_X1 U5615 ( .A(n6374), .ZN(n6417) );
  OAI22_X1 U5616 ( .A1(n5109), .A2(n4531), .B1(n4530), .B2(n5108), .ZN(n4523)
         );
  AOI21_X1 U5617 ( .B1(n6417), .B2(n4533), .A(n4523), .ZN(n4524) );
  OAI211_X1 U5618 ( .C1(n4782), .C2(n6422), .A(n4525), .B(n4524), .ZN(U3134)
         );
  NAND2_X1 U5619 ( .A1(n4529), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4528)
         );
  INV_X1 U5620 ( .A(n6370), .ZN(n6411) );
  OAI22_X1 U5621 ( .A1(n5131), .A2(n4531), .B1(n4530), .B2(n5130), .ZN(n4526)
         );
  AOI21_X1 U5622 ( .B1(n6411), .B2(n4533), .A(n4526), .ZN(n4527) );
  OAI211_X1 U5623 ( .C1(n4782), .C2(n6416), .A(n4528), .B(n4527), .ZN(U3133)
         );
  NAND2_X1 U5624 ( .A1(n4529), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4535)
         );
  INV_X1 U5625 ( .A(n6399), .ZN(n6442) );
  OAI22_X1 U5626 ( .A1(n5099), .A2(n4531), .B1(n4530), .B2(n5098), .ZN(n4532)
         );
  AOI21_X1 U5627 ( .B1(n6442), .B2(n4533), .A(n4532), .ZN(n4534) );
  OAI211_X1 U5628 ( .C1(n4782), .C2(n6451), .A(n4535), .B(n4534), .ZN(U3139)
         );
  INV_X1 U5629 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6001) );
  NAND2_X1 U5630 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6001), .ZN(n4569) );
  OAI21_X1 U5631 ( .B1(n6458), .B2(STATE2_REG_1__SCAN_IN), .A(n4569), .ZN(
        n4541) );
  INV_X1 U5632 ( .A(n4536), .ZN(n4537) );
  NOR2_X1 U5633 ( .A1(n4538), .A2(n4537), .ZN(n4539) );
  XOR2_X1 U5634 ( .A(n3902), .B(n4539), .Z(n6115) );
  NOR3_X1 U5635 ( .A1(n6115), .A2(STATE2_REG_1__SCAN_IN), .A3(n4194), .ZN(
        n4540) );
  AOI21_X1 U5636 ( .B1(n4541), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n4540), 
        .ZN(n4571) );
  INV_X1 U5637 ( .A(n4542), .ZN(n4568) );
  INV_X1 U5638 ( .A(n6454), .ZN(n4545) );
  XNOR2_X1 U5639 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4544) );
  XNOR2_X1 U5640 ( .A(n5499), .B(n5510), .ZN(n4547) );
  INV_X1 U5641 ( .A(n4547), .ZN(n4543) );
  OAI22_X1 U5642 ( .A1(n4545), .A2(n4544), .B1(n4554), .B2(n4543), .ZN(n4549)
         );
  NOR2_X1 U5643 ( .A1(n5514), .A2(n4546), .ZN(n4563) );
  NOR2_X1 U5644 ( .A1(n4563), .A2(n4547), .ZN(n4548) );
  AOI211_X1 U5645 ( .C1(n5205), .C2(n4550), .A(n4549), .B(n4548), .ZN(n5501)
         );
  MUX2_X1 U5646 ( .A(n5510), .B(n5501), .S(n6458), .Z(n6464) );
  INV_X1 U5647 ( .A(n6464), .ZN(n4566) );
  NAND2_X1 U5648 ( .A1(n4551), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4552) );
  INV_X1 U5649 ( .A(n4552), .ZN(n4553) );
  MUX2_X1 U5650 ( .A(n4553), .B(n4552), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4560) );
  INV_X1 U5651 ( .A(n4554), .ZN(n4559) );
  INV_X1 U5652 ( .A(n4555), .ZN(n4556) );
  OAI211_X1 U5653 ( .C1(n5499), .C2(n4558), .A(n4557), .B(n4556), .ZN(n5848)
         );
  AOI22_X1 U5654 ( .A1(n6454), .A2(n4560), .B1(n4559), .B2(n5848), .ZN(n4565)
         );
  MUX2_X1 U5655 ( .A(n4561), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5499), 
        .Z(n4562) );
  OR3_X1 U5656 ( .A1(n4563), .A2(n4542), .A3(n4562), .ZN(n4564) );
  OAI211_X1 U5657 ( .C1(n5153), .C2(n6453), .A(n4565), .B(n4564), .ZN(n5847)
         );
  MUX2_X1 U5658 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5847), .S(n6458), 
        .Z(n6467) );
  NAND3_X1 U5659 ( .A1(n4566), .A2(n6467), .A3(n6571), .ZN(n4567) );
  OAI211_X1 U5660 ( .C1(n4569), .C2(n4568), .A(n4567), .B(n4571), .ZN(n6473)
         );
  INV_X1 U5661 ( .A(n6473), .ZN(n4570) );
  AOI21_X1 U5662 ( .B1(n4571), .B2(n4212), .A(n4570), .ZN(n4582) );
  NOR2_X1 U5663 ( .A1(n4582), .A2(FLUSH_REG_SCAN_IN), .ZN(n4573) );
  OAI21_X1 U5664 ( .B1(n4573), .B2(n6568), .A(n4572), .ZN(n6348) );
  OR2_X1 U5665 ( .A1(n4574), .A2(n6593), .ZN(n4748) );
  AND2_X1 U5666 ( .A1(n4748), .A2(n4714), .ZN(n4629) );
  INV_X1 U5667 ( .A(n4607), .ZN(n4575) );
  NAND2_X1 U5668 ( .A1(n4575), .A2(n5840), .ZN(n4598) );
  AOI21_X1 U5669 ( .B1(n4629), .B2(n4598), .A(n5844), .ZN(n4578) );
  INV_X1 U5670 ( .A(n4686), .ZN(n4576) );
  AND2_X1 U5671 ( .A1(n3174), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5842) );
  OAI22_X1 U5672 ( .A1(n4576), .A2(n5088), .B1(n5153), .B2(n5842), .ZN(n4577)
         );
  OAI21_X1 U5673 ( .B1(n4578), .B2(n4577), .A(n6348), .ZN(n4579) );
  OAI21_X1 U5674 ( .B1(n6348), .B2(n6466), .A(n4579), .ZN(U3462) );
  INV_X1 U5675 ( .A(n4580), .ZN(n4581) );
  NOR2_X1 U5676 ( .A1(n4582), .A2(n4581), .ZN(n6482) );
  OAI22_X1 U5677 ( .A1(n4888), .A2(n5844), .B1(n4328), .B2(n5842), .ZN(n4583)
         );
  OAI21_X1 U5678 ( .B1(n6482), .B2(n4583), .A(n6348), .ZN(n4584) );
  OAI21_X1 U5679 ( .B1(n6348), .B2(n6455), .A(n4584), .ZN(U3465) );
  INV_X1 U5680 ( .A(n5840), .ZN(n4585) );
  OAI21_X1 U5681 ( .B1(n4714), .B2(n4585), .A(n5836), .ZN(n4590) );
  OR2_X1 U5682 ( .A1(n5205), .A2(n6137), .ZN(n4631) );
  INV_X1 U5683 ( .A(n4631), .ZN(n4586) );
  AND2_X1 U5684 ( .A1(n4586), .A2(n4632), .ZN(n4981) );
  NOR2_X1 U5685 ( .A1(n4633), .A2(n6466), .ZN(n6443) );
  AOI21_X1 U5686 ( .B1(n4981), .B2(n4688), .A(n6443), .ZN(n4587) );
  NAND3_X1 U5687 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4716), .ZN(n4982) );
  OAI22_X1 U5688 ( .A1(n4590), .A2(n4587), .B1(n4982), .B2(n4987), .ZN(n6445)
         );
  INV_X1 U5689 ( .A(n6445), .ZN(n4597) );
  INV_X1 U5690 ( .A(n4587), .ZN(n4589) );
  AOI21_X1 U5691 ( .B1(n5844), .B2(n4982), .A(n4883), .ZN(n4588) );
  OAI21_X1 U5692 ( .B1(n4590), .B2(n4589), .A(n4588), .ZN(n6447) );
  AOI22_X1 U5693 ( .A1(n6384), .A2(n6443), .B1(n5142), .B2(n6441), .ZN(n4591)
         );
  OAI21_X1 U5694 ( .B1(n6450), .B2(n5145), .A(n4591), .ZN(n4592) );
  AOI21_X1 U5695 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(n6447), .A(n4592), 
        .ZN(n4593) );
  OAI21_X1 U5696 ( .B1(n4597), .B2(n5136), .A(n4593), .ZN(U3113) );
  AOI22_X1 U5697 ( .A1(n6356), .A2(n6443), .B1(n5126), .B2(n6441), .ZN(n4594)
         );
  OAI21_X1 U5698 ( .B1(n6450), .B2(n5129), .A(n4594), .ZN(n4595) );
  AOI21_X1 U5699 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n6447), .A(n4595), 
        .ZN(n4596) );
  OAI21_X1 U5700 ( .B1(n4597), .B2(n5123), .A(n4596), .ZN(U3108) );
  NAND2_X1 U5701 ( .A1(n5836), .A2(n4598), .ZN(n4603) );
  NAND3_X1 U5702 ( .A1(n5153), .A2(n4688), .A3(n4599), .ZN(n4600) );
  AND2_X1 U5703 ( .A1(n4600), .A2(n4605), .ZN(n4604) );
  INV_X1 U5704 ( .A(n4604), .ZN(n4602) );
  AOI21_X1 U5705 ( .B1(n6349), .B2(n5844), .A(n4883), .ZN(n4601) );
  OAI21_X1 U5706 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n6407) );
  OAI22_X1 U5707 ( .A1(n4604), .A2(n4603), .B1(n4987), .B2(n6349), .ZN(n6406)
         );
  AOI22_X1 U5708 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6407), .B1(n6413), 
        .B2(n6406), .ZN(n4609) );
  INV_X1 U5709 ( .A(n4605), .ZN(n6405) );
  NOR2_X2 U5710 ( .A1(n4607), .A2(n4606), .ZN(n6404) );
  AOI22_X1 U5711 ( .A1(n6412), .A2(n6405), .B1(n6411), .B2(n6404), .ZN(n4608)
         );
  OAI211_X1 U5712 ( .C1(n6416), .C2(n6410), .A(n4609), .B(n4608), .ZN(U3077)
         );
  AOI22_X1 U5713 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6407), .B1(n6425), 
        .B2(n6406), .ZN(n4611) );
  AOI22_X1 U5714 ( .A1(n6424), .A2(n6405), .B1(n6423), .B2(n6404), .ZN(n4610)
         );
  OAI211_X1 U5715 ( .C1(n6428), .C2(n6410), .A(n4611), .B(n4610), .ZN(U3079)
         );
  AOI22_X1 U5716 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6407), .B1(n6355), 
        .B2(n6406), .ZN(n4613) );
  AOI22_X1 U5717 ( .A1(n6356), .A2(n6405), .B1(n5126), .B2(n6404), .ZN(n4612)
         );
  OAI211_X1 U5718 ( .C1(n5129), .C2(n6410), .A(n4613), .B(n4612), .ZN(U3076)
         );
  AOI22_X1 U5719 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6407), .B1(n6383), 
        .B2(n6406), .ZN(n4615) );
  AOI22_X1 U5720 ( .A1(n6384), .A2(n6405), .B1(n5142), .B2(n6404), .ZN(n4614)
         );
  OAI211_X1 U5721 ( .C1(n5145), .C2(n6410), .A(n4615), .B(n4614), .ZN(U3081)
         );
  AOI22_X1 U5722 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6407), .B1(n6446), 
        .B2(n6406), .ZN(n4617) );
  AOI22_X1 U5723 ( .A1(n6444), .A2(n6405), .B1(n6442), .B2(n6404), .ZN(n4616)
         );
  OAI211_X1 U5724 ( .C1(n6451), .C2(n6410), .A(n4617), .B(n4616), .ZN(U3083)
         );
  NAND2_X1 U5725 ( .A1(n4620), .A2(n4619), .ZN(n4621) );
  AND2_X1 U5726 ( .A1(n4867), .A2(n4621), .ZN(n6231) );
  INV_X1 U5727 ( .A(n6231), .ZN(n4673) );
  AND2_X1 U5728 ( .A1(n4623), .A2(n4622), .ZN(n4625) );
  OR2_X1 U5729 ( .A1(n4625), .A2(n4624), .ZN(n6109) );
  INV_X1 U5730 ( .A(n6109), .ZN(n4626) );
  AOI22_X1 U5731 ( .A1(n5675), .A2(n4626), .B1(EBX_REG_6__SCAN_IN), .B2(n5674), 
        .ZN(n4627) );
  OAI21_X1 U5732 ( .B1(n4673), .B2(n5677), .A(n4627), .ZN(U2853) );
  NAND3_X1 U5733 ( .A1(n4629), .A2(n4628), .A3(n5840), .ZN(n4630) );
  NAND2_X1 U5734 ( .A1(n4630), .A2(n5836), .ZN(n4643) );
  INV_X1 U5735 ( .A(n4643), .ZN(n4637) );
  NOR2_X1 U5736 ( .A1(n4632), .A2(n4631), .ZN(n5097) );
  NAND2_X1 U5737 ( .A1(n5097), .A2(n4688), .ZN(n4635) );
  INV_X1 U5738 ( .A(n4633), .ZN(n4634) );
  NAND2_X1 U5739 ( .A1(n4634), .A2(n6466), .ZN(n4665) );
  NAND2_X1 U5740 ( .A1(n4635), .A2(n4665), .ZN(n4642) );
  NAND3_X1 U5741 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6466), .A3(n4716), .ZN(n5087) );
  INV_X1 U5742 ( .A(n5087), .ZN(n4636) );
  AOI22_X1 U5743 ( .A1(n4637), .A2(n4642), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4636), .ZN(n4670) );
  NOR3_X1 U5744 ( .A1(n4686), .A2(n5841), .A3(n4638), .ZN(n4639) );
  OAI22_X1 U5745 ( .A1(n5139), .A2(n4665), .B1(n6388), .B2(n4664), .ZN(n4640)
         );
  AOI21_X1 U5746 ( .B1(n6385), .B2(n5141), .A(n4640), .ZN(n4645) );
  AOI21_X1 U5747 ( .B1(n5844), .B2(n5087), .A(n4883), .ZN(n4641) );
  OAI21_X1 U5748 ( .B1(n4643), .B2(n4642), .A(n4641), .ZN(n4667) );
  NAND2_X1 U5749 ( .A1(n4667), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4644) );
  OAI211_X1 U5750 ( .C1(n4670), .C2(n5136), .A(n4645), .B(n4644), .ZN(U3049)
         );
  OAI22_X1 U5751 ( .A1(n5104), .A2(n4665), .B1(n6392), .B2(n4664), .ZN(n4646)
         );
  AOI21_X1 U5752 ( .B1(n6389), .B2(n5141), .A(n4646), .ZN(n4648) );
  NAND2_X1 U5753 ( .A1(n4667), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4647) );
  OAI211_X1 U5754 ( .C1(n4670), .C2(n5103), .A(n4648), .B(n4647), .ZN(U3050)
         );
  OAI22_X1 U5755 ( .A1(n5119), .A2(n4665), .B1(n6378), .B2(n4664), .ZN(n4649)
         );
  AOI21_X1 U5756 ( .B1(n6375), .B2(n5141), .A(n4649), .ZN(n4651) );
  NAND2_X1 U5757 ( .A1(n4667), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4650) );
  OAI211_X1 U5758 ( .C1(n4670), .C2(n5118), .A(n4651), .B(n4650), .ZN(U3047)
         );
  OAI22_X1 U5759 ( .A1(n5131), .A2(n4665), .B1(n6370), .B2(n4664), .ZN(n4652)
         );
  AOI21_X1 U5760 ( .B1(n6367), .B2(n5141), .A(n4652), .ZN(n4654) );
  NAND2_X1 U5761 ( .A1(n4667), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4653) );
  OAI211_X1 U5762 ( .C1(n4670), .C2(n5130), .A(n4654), .B(n4653), .ZN(U3045)
         );
  OAI22_X1 U5763 ( .A1(n5109), .A2(n4665), .B1(n6374), .B2(n4664), .ZN(n4655)
         );
  AOI21_X1 U5764 ( .B1(n6371), .B2(n5141), .A(n4655), .ZN(n4657) );
  NAND2_X1 U5765 ( .A1(n4667), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4656) );
  OAI211_X1 U5766 ( .C1(n4670), .C2(n5108), .A(n4657), .B(n4656), .ZN(U3046)
         );
  OAI22_X1 U5767 ( .A1(n5114), .A2(n4665), .B1(n6382), .B2(n4664), .ZN(n4658)
         );
  AOI21_X1 U5768 ( .B1(n6379), .B2(n5141), .A(n4658), .ZN(n4660) );
  NAND2_X1 U5769 ( .A1(n4667), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4659) );
  OAI211_X1 U5770 ( .C1(n4670), .C2(n5113), .A(n4660), .B(n4659), .ZN(U3048)
         );
  OAI22_X1 U5771 ( .A1(n5124), .A2(n4665), .B1(n6366), .B2(n4664), .ZN(n4661)
         );
  AOI21_X1 U5772 ( .B1(n6363), .B2(n5141), .A(n4661), .ZN(n4663) );
  NAND2_X1 U5773 ( .A1(n4667), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4662) );
  OAI211_X1 U5774 ( .C1(n4670), .C2(n5123), .A(n4663), .B(n4662), .ZN(U3044)
         );
  OAI22_X1 U5775 ( .A1(n5099), .A2(n4665), .B1(n6399), .B2(n4664), .ZN(n4666)
         );
  AOI21_X1 U5776 ( .B1(n6395), .B2(n5141), .A(n4666), .ZN(n4669) );
  NAND2_X1 U5777 ( .A1(n4667), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4668) );
  OAI211_X1 U5778 ( .C1(n4670), .C2(n5098), .A(n4669), .B(n4668), .ZN(U3051)
         );
  OAI222_X1 U5779 ( .A1(n4673), .A2(n5917), .B1(n4672), .B2(n4671), .C1(n5453), 
        .C2(n4849), .ZN(U2885) );
  OAI21_X1 U5780 ( .B1(n4676), .B2(n4675), .A(n4674), .ZN(n6230) );
  NOR2_X1 U5781 ( .A1(n6283), .A2(n6109), .ZN(n4684) );
  INV_X1 U5782 ( .A(n4677), .ZN(n4678) );
  NAND3_X1 U5783 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6331), .ZN(n6305) );
  NAND2_X1 U5784 ( .A1(n5362), .A2(n6305), .ZN(n5173) );
  INV_X1 U5785 ( .A(n5173), .ZN(n6323) );
  AOI21_X1 U5786 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6335) );
  NAND2_X1 U5787 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6316) );
  NOR2_X1 U5788 ( .A1(n6335), .A2(n6316), .ZN(n6301) );
  NAND2_X1 U5789 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6301), .ZN(n5169)
         );
  NOR2_X1 U5790 ( .A1(n6323), .A2(n5169), .ZN(n4682) );
  NAND2_X1 U5791 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5167) );
  INV_X1 U5792 ( .A(n5167), .ZN(n4679) );
  OAI21_X1 U5793 ( .B1(n4680), .B2(n4679), .A(n5347), .ZN(n6332) );
  AOI21_X1 U5794 ( .B1(n5169), .B2(n5957), .A(n6332), .ZN(n6312) );
  INV_X1 U5795 ( .A(n6312), .ZN(n4681) );
  MUX2_X1 U5796 ( .A(n4682), .B(n4681), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4683) );
  AOI211_X1 U5797 ( .C1(n6336), .C2(REIP_REG_6__SCAN_IN), .A(n4684), .B(n4683), 
        .ZN(n4685) );
  OAI21_X1 U5798 ( .B1(n6342), .B2(n6230), .A(n4685), .ZN(U3012) );
  NOR3_X1 U5799 ( .A1(n4686), .A2(n5841), .A3(n5837), .ZN(n4694) );
  NAND2_X1 U5800 ( .A1(n4694), .A2(n4888), .ZN(n4930) );
  INV_X1 U5801 ( .A(n4694), .ZN(n4687) );
  OAI21_X1 U5802 ( .B1(n4687), .B2(n6593), .A(n5836), .ZN(n4692) );
  OR2_X1 U5803 ( .A1(n5205), .A2(n4192), .ZN(n4941) );
  INV_X1 U5804 ( .A(n4941), .ZN(n4811) );
  NAND2_X1 U5805 ( .A1(n5153), .A2(n4811), .ZN(n4932) );
  INV_X1 U5806 ( .A(n4932), .ZN(n4689) );
  NAND3_X1 U5807 ( .A1(n6466), .A2(n4716), .A3(n6461), .ZN(n4935) );
  NOR2_X1 U5808 ( .A1(n6455), .A2(n4935), .ZN(n4711) );
  AOI21_X1 U5809 ( .B1(n4689), .B2(n4688), .A(n4711), .ZN(n4693) );
  INV_X1 U5810 ( .A(n4693), .ZN(n4691) );
  AOI21_X1 U5811 ( .B1(n5844), .B2(n4935), .A(n4883), .ZN(n4690) );
  OAI21_X1 U5812 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n4710) );
  OAI22_X1 U5813 ( .A1(n4693), .A2(n4692), .B1(n4987), .B2(n4935), .ZN(n4709)
         );
  AOI22_X1 U5814 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4710), .B1(n6431), 
        .B2(n4709), .ZN(n4696) );
  NAND2_X1 U5815 ( .A1(n4694), .A2(n4722), .ZN(n5146) );
  AOI22_X1 U5816 ( .A1(n5089), .A2(n6429), .B1(n6430), .B2(n4711), .ZN(n4695)
         );
  OAI211_X1 U5817 ( .C1(n6434), .C2(n4930), .A(n4696), .B(n4695), .ZN(U3032)
         );
  AOI22_X1 U5818 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4710), .B1(n6383), 
        .B2(n4709), .ZN(n4698) );
  AOI22_X1 U5819 ( .A1(n5089), .A2(n5142), .B1(n6384), .B2(n4711), .ZN(n4697)
         );
  OAI211_X1 U5820 ( .C1(n5145), .C2(n4930), .A(n4698), .B(n4697), .ZN(U3033)
         );
  AOI22_X1 U5821 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4710), .B1(n6419), 
        .B2(n4709), .ZN(n4700) );
  AOI22_X1 U5822 ( .A1(n5089), .A2(n6417), .B1(n6418), .B2(n4711), .ZN(n4699)
         );
  OAI211_X1 U5823 ( .C1(n6422), .C2(n4930), .A(n4700), .B(n4699), .ZN(U3030)
         );
  AOI22_X1 U5824 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4710), .B1(n6355), 
        .B2(n4709), .ZN(n4702) );
  AOI22_X1 U5825 ( .A1(n5089), .A2(n5126), .B1(n6356), .B2(n4711), .ZN(n4701)
         );
  OAI211_X1 U5826 ( .C1(n5129), .C2(n4930), .A(n4702), .B(n4701), .ZN(U3028)
         );
  AOI22_X1 U5827 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4710), .B1(n6446), 
        .B2(n4709), .ZN(n4704) );
  AOI22_X1 U5828 ( .A1(n5089), .A2(n6442), .B1(n6444), .B2(n4711), .ZN(n4703)
         );
  OAI211_X1 U5829 ( .C1(n6451), .C2(n4930), .A(n4704), .B(n4703), .ZN(U3035)
         );
  AOI22_X1 U5830 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4710), .B1(n6437), 
        .B2(n4709), .ZN(n4706) );
  AOI22_X1 U5831 ( .A1(n5089), .A2(n6435), .B1(n6436), .B2(n4711), .ZN(n4705)
         );
  OAI211_X1 U5832 ( .C1(n6440), .C2(n4930), .A(n4706), .B(n4705), .ZN(U3034)
         );
  AOI22_X1 U5833 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4710), .B1(n6425), 
        .B2(n4709), .ZN(n4708) );
  AOI22_X1 U5834 ( .A1(n5089), .A2(n6423), .B1(n6424), .B2(n4711), .ZN(n4707)
         );
  OAI211_X1 U5835 ( .C1(n6428), .C2(n4930), .A(n4708), .B(n4707), .ZN(U3031)
         );
  AOI22_X1 U5836 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4710), .B1(n6413), 
        .B2(n4709), .ZN(n4713) );
  AOI22_X1 U5837 ( .A1(n5089), .A2(n6411), .B1(n6412), .B2(n4711), .ZN(n4712)
         );
  OAI211_X1 U5838 ( .C1(n6416), .C2(n4930), .A(n4713), .B(n4712), .ZN(U3029)
         );
  INV_X1 U5839 ( .A(n4715), .ZN(n4746) );
  NAND3_X1 U5840 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4716), .A3(n6461), .ZN(n4802) );
  NOR2_X1 U5841 ( .A1(n6455), .A2(n4802), .ZN(n4740) );
  AOI21_X1 U5842 ( .B1(n4746), .B2(n4811), .A(n4740), .ZN(n4721) );
  INV_X1 U5843 ( .A(n4721), .ZN(n4719) );
  INV_X1 U5844 ( .A(n4723), .ZN(n4717) );
  OAI21_X1 U5845 ( .B1(n4717), .B2(n6593), .A(n5836), .ZN(n4720) );
  AOI21_X1 U5846 ( .B1(n5844), .B2(n4802), .A(n4883), .ZN(n4718) );
  OAI21_X1 U5847 ( .B1(n4719), .B2(n4720), .A(n4718), .ZN(n4739) );
  OAI22_X1 U5848 ( .A1(n4721), .A2(n4720), .B1(n4987), .B2(n4802), .ZN(n4738)
         );
  AOI22_X1 U5849 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4739), .B1(n6413), 
        .B2(n4738), .ZN(n4725) );
  NAND2_X1 U5850 ( .A1(n4723), .A2(n4722), .ZN(n4978) );
  AOI22_X1 U5851 ( .A1(n5013), .A2(n6411), .B1(n6412), .B2(n4740), .ZN(n4724)
         );
  OAI211_X1 U5852 ( .C1(n6416), .C2(n4842), .A(n4725), .B(n4724), .ZN(U3093)
         );
  AOI22_X1 U5853 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4739), .B1(n6446), 
        .B2(n4738), .ZN(n4727) );
  AOI22_X1 U5854 ( .A1(n5013), .A2(n6442), .B1(n6444), .B2(n4740), .ZN(n4726)
         );
  OAI211_X1 U5855 ( .C1(n6451), .C2(n4842), .A(n4727), .B(n4726), .ZN(U3099)
         );
  AOI22_X1 U5856 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4739), .B1(n6419), 
        .B2(n4738), .ZN(n4729) );
  AOI22_X1 U5857 ( .A1(n5013), .A2(n6417), .B1(n6418), .B2(n4740), .ZN(n4728)
         );
  OAI211_X1 U5858 ( .C1(n6422), .C2(n4842), .A(n4729), .B(n4728), .ZN(U3094)
         );
  AOI22_X1 U5859 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4739), .B1(n6355), 
        .B2(n4738), .ZN(n4731) );
  AOI22_X1 U5860 ( .A1(n5013), .A2(n5126), .B1(n6356), .B2(n4740), .ZN(n4730)
         );
  OAI211_X1 U5861 ( .C1(n5129), .C2(n4842), .A(n4731), .B(n4730), .ZN(U3092)
         );
  AOI22_X1 U5862 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4739), .B1(n6431), 
        .B2(n4738), .ZN(n4733) );
  AOI22_X1 U5863 ( .A1(n5013), .A2(n6429), .B1(n6430), .B2(n4740), .ZN(n4732)
         );
  OAI211_X1 U5864 ( .C1(n6434), .C2(n4842), .A(n4733), .B(n4732), .ZN(U3096)
         );
  AOI22_X1 U5865 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4739), .B1(n6425), 
        .B2(n4738), .ZN(n4735) );
  AOI22_X1 U5866 ( .A1(n5013), .A2(n6423), .B1(n6424), .B2(n4740), .ZN(n4734)
         );
  OAI211_X1 U5867 ( .C1(n6428), .C2(n4842), .A(n4735), .B(n4734), .ZN(U3095)
         );
  AOI22_X1 U5868 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4739), .B1(n6383), 
        .B2(n4738), .ZN(n4737) );
  AOI22_X1 U5869 ( .A1(n5013), .A2(n5142), .B1(n6384), .B2(n4740), .ZN(n4736)
         );
  OAI211_X1 U5870 ( .C1(n5145), .C2(n4842), .A(n4737), .B(n4736), .ZN(U3097)
         );
  AOI22_X1 U5871 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4739), .B1(n6437), 
        .B2(n4738), .ZN(n4742) );
  AOI22_X1 U5872 ( .A1(n5013), .A2(n6435), .B1(n6436), .B2(n4740), .ZN(n4741)
         );
  OAI211_X1 U5873 ( .C1(n6440), .C2(n4842), .A(n4742), .B(n4741), .ZN(U3098)
         );
  NOR2_X1 U5874 ( .A1(n6455), .A2(n4747), .ZN(n4744) );
  INV_X1 U5875 ( .A(n4744), .ZN(n4778) );
  AOI21_X1 U5876 ( .B1(n4746), .B2(n4745), .A(n4744), .ZN(n4749) );
  OAI22_X1 U5877 ( .A1(n4749), .A2(n5844), .B1(n4747), .B2(n4987), .ZN(n4776)
         );
  NAND2_X1 U5878 ( .A1(n4749), .A2(n4748), .ZN(n4750) );
  OR2_X1 U5879 ( .A1(n5844), .A2(n4750), .ZN(n4752) );
  OAI211_X1 U5880 ( .C1(n5836), .C2(n4753), .A(n4752), .B(n4751), .ZN(n4775)
         );
  AOI22_X1 U5881 ( .A1(n4776), .A2(n6437), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4775), .ZN(n4754) );
  OAI21_X1 U5882 ( .B1(n5104), .B2(n4778), .A(n4754), .ZN(n4755) );
  AOI21_X1 U5883 ( .B1(n6389), .B2(n4780), .A(n4755), .ZN(n4756) );
  OAI21_X1 U5884 ( .B1(n6392), .B2(n4782), .A(n4756), .ZN(U3130) );
  AOI22_X1 U5885 ( .A1(n4776), .A2(n6425), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4775), .ZN(n4757) );
  OAI21_X1 U5886 ( .B1(n5119), .B2(n4778), .A(n4757), .ZN(n4758) );
  AOI21_X1 U5887 ( .B1(n6375), .B2(n4780), .A(n4758), .ZN(n4759) );
  OAI21_X1 U5888 ( .B1(n6378), .B2(n4782), .A(n4759), .ZN(U3127) );
  AOI22_X1 U5889 ( .A1(n4776), .A2(n6446), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4775), .ZN(n4760) );
  OAI21_X1 U5890 ( .B1(n5099), .B2(n4778), .A(n4760), .ZN(n4761) );
  AOI21_X1 U5891 ( .B1(n6395), .B2(n4780), .A(n4761), .ZN(n4762) );
  OAI21_X1 U5892 ( .B1(n6399), .B2(n4782), .A(n4762), .ZN(U3131) );
  AOI22_X1 U5893 ( .A1(n4776), .A2(n6413), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4775), .ZN(n4763) );
  OAI21_X1 U5894 ( .B1(n5131), .B2(n4778), .A(n4763), .ZN(n4764) );
  AOI21_X1 U5895 ( .B1(n6367), .B2(n4780), .A(n4764), .ZN(n4765) );
  OAI21_X1 U5896 ( .B1(n6370), .B2(n4782), .A(n4765), .ZN(U3125) );
  AOI22_X1 U5897 ( .A1(n4776), .A2(n6419), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4775), .ZN(n4766) );
  OAI21_X1 U5898 ( .B1(n5109), .B2(n4778), .A(n4766), .ZN(n4767) );
  AOI21_X1 U5899 ( .B1(n6371), .B2(n4780), .A(n4767), .ZN(n4768) );
  OAI21_X1 U5900 ( .B1(n6374), .B2(n4782), .A(n4768), .ZN(U3126) );
  AOI22_X1 U5901 ( .A1(n4776), .A2(n6355), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4775), .ZN(n4769) );
  OAI21_X1 U5902 ( .B1(n5124), .B2(n4778), .A(n4769), .ZN(n4770) );
  AOI21_X1 U5903 ( .B1(n6363), .B2(n4780), .A(n4770), .ZN(n4771) );
  OAI21_X1 U5904 ( .B1(n6366), .B2(n4782), .A(n4771), .ZN(U3124) );
  AOI22_X1 U5905 ( .A1(n4776), .A2(n6431), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4775), .ZN(n4772) );
  OAI21_X1 U5906 ( .B1(n5114), .B2(n4778), .A(n4772), .ZN(n4773) );
  AOI21_X1 U5907 ( .B1(n6379), .B2(n4780), .A(n4773), .ZN(n4774) );
  OAI21_X1 U5908 ( .B1(n6382), .B2(n4782), .A(n4774), .ZN(U3128) );
  AOI22_X1 U5909 ( .A1(n4776), .A2(n6383), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4775), .ZN(n4777) );
  OAI21_X1 U5910 ( .B1(n5139), .B2(n4778), .A(n4777), .ZN(n4779) );
  AOI21_X1 U5911 ( .B1(n6385), .B2(n4780), .A(n4779), .ZN(n4781) );
  OAI21_X1 U5912 ( .B1(n6388), .B2(n4782), .A(n4781), .ZN(U3129) );
  INV_X1 U5913 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5914 ( .A1(n6604), .A2(UWORD_REG_14__SCAN_IN), .B1(
        DATAO_REG_30__SCAN_IN), .B2(n6184), .ZN(n4783) );
  OAI21_X1 U5915 ( .B1(n4784), .B2(n4800), .A(n4783), .ZN(U2893) );
  INV_X1 U5916 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4786) );
  AOI22_X1 U5917 ( .A1(n6604), .A2(UWORD_REG_8__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4785) );
  OAI21_X1 U5918 ( .B1(n4786), .B2(n4800), .A(n4785), .ZN(U2899) );
  INV_X1 U5919 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6191) );
  AOI22_X1 U5920 ( .A1(n6604), .A2(UWORD_REG_10__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4787) );
  OAI21_X1 U5921 ( .B1(n6191), .B2(n4800), .A(n4787), .ZN(U2897) );
  INV_X1 U5922 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U5923 ( .A1(n6604), .A2(UWORD_REG_12__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4788) );
  OAI21_X1 U5924 ( .B1(n6626), .B2(n4800), .A(n4788), .ZN(U2895) );
  INV_X1 U5925 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4851) );
  AOI22_X1 U5926 ( .A1(n6604), .A2(UWORD_REG_4__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4789) );
  OAI21_X1 U5927 ( .B1(n4851), .B2(n4800), .A(n4789), .ZN(U2903) );
  AOI22_X1 U5928 ( .A1(n6604), .A2(UWORD_REG_6__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4790) );
  OAI21_X1 U5929 ( .B1(n4791), .B2(n4800), .A(n4790), .ZN(U2901) );
  INV_X1 U5930 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U5931 ( .A1(n6604), .A2(UWORD_REG_0__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4792) );
  OAI21_X1 U5932 ( .B1(n4793), .B2(n4800), .A(n4792), .ZN(U2907) );
  INV_X1 U5933 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5934 ( .A1(n6604), .A2(UWORD_REG_5__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4794) );
  OAI21_X1 U5935 ( .B1(n4795), .B2(n4800), .A(n4794), .ZN(U2902) );
  INV_X1 U5936 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U5937 ( .A1(n6604), .A2(UWORD_REG_3__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4796) );
  OAI21_X1 U5938 ( .B1(n4797), .B2(n4800), .A(n4796), .ZN(U2904) );
  INV_X1 U5939 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U5940 ( .A1(n6604), .A2(UWORD_REG_2__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4798) );
  OAI21_X1 U5941 ( .B1(n4854), .B2(n4800), .A(n4798), .ZN(U2905) );
  INV_X1 U5942 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4801) );
  AOI22_X1 U5943 ( .A1(n6604), .A2(UWORD_REG_1__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4799) );
  OAI21_X1 U5944 ( .B1(n4801), .B2(n4800), .A(n4799), .ZN(U2906) );
  NOR2_X1 U5945 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4802), .ZN(n4809)
         );
  INV_X1 U5946 ( .A(n4809), .ZN(n4837) );
  INV_X1 U5947 ( .A(n4803), .ZN(n4804) );
  AOI22_X1 U5948 ( .A1(n4805), .A2(n4811), .B1(n6359), .B2(n4804), .ZN(n4836)
         );
  OAI22_X1 U5949 ( .A1(n5131), .A2(n4837), .B1(n4836), .B2(n5130), .ZN(n4806)
         );
  AOI21_X1 U5950 ( .B1(n6367), .B2(n6404), .A(n4806), .ZN(n4817) );
  OAI211_X1 U5951 ( .C1(n3174), .C2(n4809), .A(n4808), .B(n4807), .ZN(n4810)
         );
  AOI21_X1 U5952 ( .B1(n4941), .B2(n4933), .A(n4810), .ZN(n4815) );
  INV_X1 U5953 ( .A(n6404), .ZN(n4813) );
  OAI21_X1 U5954 ( .B1(n4811), .B2(n5844), .A(n6354), .ZN(n4812) );
  NAND3_X1 U5955 ( .A1(n4842), .A2(n4813), .A3(n4812), .ZN(n4814) );
  NAND2_X1 U5956 ( .A1(n4815), .A2(n4814), .ZN(n4839) );
  NAND2_X1 U5957 ( .A1(n4839), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4816) );
  OAI211_X1 U5958 ( .C1(n4842), .C2(n6370), .A(n4817), .B(n4816), .ZN(U3085)
         );
  OAI22_X1 U5959 ( .A1(n5124), .A2(n4837), .B1(n4836), .B2(n5123), .ZN(n4818)
         );
  AOI21_X1 U5960 ( .B1(n6363), .B2(n6404), .A(n4818), .ZN(n4820) );
  NAND2_X1 U5961 ( .A1(n4839), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4819) );
  OAI211_X1 U5962 ( .C1(n4842), .C2(n6366), .A(n4820), .B(n4819), .ZN(U3084)
         );
  OAI22_X1 U5963 ( .A1(n5099), .A2(n4837), .B1(n4836), .B2(n5098), .ZN(n4821)
         );
  AOI21_X1 U5964 ( .B1(n6395), .B2(n6404), .A(n4821), .ZN(n4823) );
  NAND2_X1 U5965 ( .A1(n4839), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4822) );
  OAI211_X1 U5966 ( .C1(n4842), .C2(n6399), .A(n4823), .B(n4822), .ZN(U3091)
         );
  OAI22_X1 U5967 ( .A1(n5109), .A2(n4837), .B1(n4836), .B2(n5108), .ZN(n4824)
         );
  AOI21_X1 U5968 ( .B1(n6371), .B2(n6404), .A(n4824), .ZN(n4826) );
  NAND2_X1 U5969 ( .A1(n4839), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4825) );
  OAI211_X1 U5970 ( .C1(n4842), .C2(n6374), .A(n4826), .B(n4825), .ZN(U3086)
         );
  OAI22_X1 U5971 ( .A1(n5119), .A2(n4837), .B1(n4836), .B2(n5118), .ZN(n4827)
         );
  AOI21_X1 U5972 ( .B1(n6375), .B2(n6404), .A(n4827), .ZN(n4829) );
  NAND2_X1 U5973 ( .A1(n4839), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4828) );
  OAI211_X1 U5974 ( .C1(n4842), .C2(n6378), .A(n4829), .B(n4828), .ZN(U3087)
         );
  OAI22_X1 U5975 ( .A1(n5104), .A2(n4837), .B1(n4836), .B2(n5103), .ZN(n4830)
         );
  AOI21_X1 U5976 ( .B1(n6389), .B2(n6404), .A(n4830), .ZN(n4832) );
  NAND2_X1 U5977 ( .A1(n4839), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4831) );
  OAI211_X1 U5978 ( .C1(n4842), .C2(n6392), .A(n4832), .B(n4831), .ZN(U3090)
         );
  OAI22_X1 U5979 ( .A1(n5114), .A2(n4837), .B1(n4836), .B2(n5113), .ZN(n4833)
         );
  AOI21_X1 U5980 ( .B1(n6379), .B2(n6404), .A(n4833), .ZN(n4835) );
  NAND2_X1 U5981 ( .A1(n4839), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4834) );
  OAI211_X1 U5982 ( .C1(n4842), .C2(n6382), .A(n4835), .B(n4834), .ZN(U3088)
         );
  OAI22_X1 U5983 ( .A1(n5139), .A2(n4837), .B1(n4836), .B2(n5136), .ZN(n4838)
         );
  AOI21_X1 U5984 ( .B1(n6385), .B2(n6404), .A(n4838), .ZN(n4841) );
  NAND2_X1 U5985 ( .A1(n4839), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4840) );
  OAI211_X1 U5986 ( .C1(n4842), .C2(n6388), .A(n4841), .B(n4840), .ZN(U3089)
         );
  NAND2_X1 U5987 ( .A1(n6215), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U5988 ( .A1(n6214), .A2(DATAI_2_), .ZN(n4852) );
  OAI211_X1 U5989 ( .C1(n6217), .C2(n6752), .A(n4844), .B(n4852), .ZN(U2941)
         );
  NAND2_X1 U5990 ( .A1(n6215), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4846) );
  OAI211_X1 U5991 ( .C1(n6217), .C2(n4801), .A(n4846), .B(n4845), .ZN(U2925)
         );
  NAND2_X1 U5992 ( .A1(n6215), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4848) );
  OAI211_X1 U5993 ( .C1(n6217), .C2(n4849), .A(n4848), .B(n4847), .ZN(U2945)
         );
  NAND2_X1 U5994 ( .A1(n6215), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U5995 ( .A1(n6214), .A2(DATAI_4_), .ZN(n4864) );
  OAI211_X1 U5996 ( .C1(n6217), .C2(n4851), .A(n4850), .B(n4864), .ZN(U2928)
         );
  NAND2_X1 U5997 ( .A1(n6215), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4853) );
  OAI211_X1 U5998 ( .C1(n6217), .C2(n4854), .A(n4853), .B(n4852), .ZN(U2926)
         );
  NAND2_X1 U5999 ( .A1(n6215), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U6000 ( .A1(n6214), .A2(DATAI_3_), .ZN(n4862) );
  OAI211_X1 U6001 ( .C1(n6217), .C2(n4797), .A(n4855), .B(n4862), .ZN(U2927)
         );
  NAND2_X1 U6002 ( .A1(n6215), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4857) );
  OAI211_X1 U6003 ( .C1(n6217), .C2(n4793), .A(n4857), .B(n4856), .ZN(U2924)
         );
  NAND2_X1 U6004 ( .A1(n6215), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U6005 ( .A1(n6214), .A2(DATAI_5_), .ZN(n4859) );
  OAI211_X1 U6006 ( .C1(n6217), .C2(n4795), .A(n4858), .B(n4859), .ZN(U2929)
         );
  NAND2_X1 U6007 ( .A1(n6215), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4860) );
  OAI211_X1 U6008 ( .C1(n6217), .C2(n4861), .A(n4860), .B(n4859), .ZN(U2944)
         );
  NAND2_X1 U6009 ( .A1(n6215), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4863) );
  OAI211_X1 U6010 ( .C1(n6217), .C2(n6180), .A(n4863), .B(n4862), .ZN(U2942)
         );
  INV_X1 U6011 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4866) );
  NAND2_X1 U6012 ( .A1(n6215), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4865) );
  OAI211_X1 U6013 ( .C1(n6217), .C2(n4866), .A(n4865), .B(n4864), .ZN(U2943)
         );
  XOR2_X1 U6014 ( .A(n4868), .B(n4867), .Z(n5203) );
  INV_X1 U6015 ( .A(n5203), .ZN(n4928) );
  AOI22_X1 U6016 ( .A1(n5689), .A2(DATAI_7_), .B1(n6156), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4869) );
  OAI21_X1 U6017 ( .B1(n4928), .B2(n5917), .A(n4869), .ZN(U2884) );
  OAI21_X1 U6018 ( .B1(n4872), .B2(n4871), .A(n5032), .ZN(n6100) );
  AOI22_X1 U6019 ( .A1(n5689), .A2(DATAI_8_), .B1(n6156), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4873) );
  OAI21_X1 U6020 ( .B1(n6100), .B2(n5917), .A(n4873), .ZN(U2883) );
  OR2_X1 U6021 ( .A1(n4875), .A2(n4876), .ZN(n4877) );
  NAND2_X1 U6022 ( .A1(n5035), .A2(n4877), .ZN(n6282) );
  INV_X1 U6023 ( .A(n6282), .ZN(n4878) );
  AOI22_X1 U6024 ( .A1(n5675), .A2(n4878), .B1(EBX_REG_8__SCAN_IN), .B2(n5674), 
        .ZN(n4879) );
  OAI21_X1 U6025 ( .B1(n6100), .B2(n5677), .A(n4879), .ZN(U2851) );
  NOR2_X1 U6026 ( .A1(n6455), .A2(n4885), .ZN(n4917) );
  INV_X1 U6027 ( .A(n4917), .ZN(n4880) );
  OAI21_X1 U6028 ( .B1(n4881), .B2(n4328), .A(n4880), .ZN(n4884) );
  NOR2_X1 U6029 ( .A1(n4887), .A2(n4884), .ZN(n4882) );
  AOI211_X2 U6030 ( .C1(n4885), .C2(n5844), .A(n4883), .B(n4882), .ZN(n4924)
         );
  INV_X1 U6031 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4893) );
  INV_X1 U6032 ( .A(n4884), .ZN(n4886) );
  OAI22_X1 U6033 ( .A1(n4887), .A2(n4886), .B1(n4885), .B2(n4987), .ZN(n4921)
         );
  AOI22_X1 U6034 ( .A1(n6412), .A2(n4917), .B1(n6411), .B2(n3020), .ZN(n4890)
         );
  OAI21_X1 U6035 ( .B1(n6416), .B2(n4919), .A(n4890), .ZN(n4891) );
  AOI21_X1 U6036 ( .B1(n6413), .B2(n4921), .A(n4891), .ZN(n4892) );
  OAI21_X1 U6037 ( .B1(n4924), .B2(n4893), .A(n4892), .ZN(U3061) );
  INV_X1 U6038 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4897) );
  AOI22_X1 U6039 ( .A1(n6444), .A2(n4917), .B1(n6442), .B2(n3020), .ZN(n4894)
         );
  OAI21_X1 U6040 ( .B1(n6451), .B2(n4919), .A(n4894), .ZN(n4895) );
  AOI21_X1 U6041 ( .B1(n6446), .B2(n4921), .A(n4895), .ZN(n4896) );
  OAI21_X1 U6042 ( .B1(n4924), .B2(n4897), .A(n4896), .ZN(U3067) );
  INV_X1 U6043 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U6044 ( .A1(n6436), .A2(n4917), .B1(n6435), .B2(n3020), .ZN(n4898)
         );
  OAI21_X1 U6045 ( .B1(n6440), .B2(n4919), .A(n4898), .ZN(n4899) );
  AOI21_X1 U6046 ( .B1(n6437), .B2(n4921), .A(n4899), .ZN(n4900) );
  OAI21_X1 U6047 ( .B1(n4924), .B2(n6743), .A(n4900), .ZN(U3066) );
  INV_X1 U6048 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4904) );
  AOI22_X1 U6049 ( .A1(n6418), .A2(n4917), .B1(n6417), .B2(n3020), .ZN(n4901)
         );
  OAI21_X1 U6050 ( .B1(n6422), .B2(n4919), .A(n4901), .ZN(n4902) );
  AOI21_X1 U6051 ( .B1(n6419), .B2(n4921), .A(n4902), .ZN(n4903) );
  OAI21_X1 U6052 ( .B1(n4924), .B2(n4904), .A(n4903), .ZN(U3062) );
  INV_X1 U6053 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4908) );
  AOI22_X1 U6054 ( .A1(n6356), .A2(n4917), .B1(n5126), .B2(n3020), .ZN(n4905)
         );
  OAI21_X1 U6055 ( .B1(n5129), .B2(n4919), .A(n4905), .ZN(n4906) );
  AOI21_X1 U6056 ( .B1(n6355), .B2(n4921), .A(n4906), .ZN(n4907) );
  OAI21_X1 U6057 ( .B1(n4924), .B2(n4908), .A(n4907), .ZN(U3060) );
  INV_X1 U6058 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U6059 ( .A1(n6424), .A2(n4917), .B1(n6423), .B2(n3020), .ZN(n4909)
         );
  OAI21_X1 U6060 ( .B1(n6428), .B2(n4919), .A(n4909), .ZN(n4910) );
  AOI21_X1 U6061 ( .B1(n6425), .B2(n4921), .A(n4910), .ZN(n4911) );
  OAI21_X1 U6062 ( .B1(n4924), .B2(n4912), .A(n4911), .ZN(U3063) );
  INV_X1 U6063 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4916) );
  AOI22_X1 U6064 ( .A1(n6384), .A2(n4917), .B1(n5142), .B2(n3020), .ZN(n4913)
         );
  OAI21_X1 U6065 ( .B1(n5145), .B2(n4919), .A(n4913), .ZN(n4914) );
  AOI21_X1 U6066 ( .B1(n6383), .B2(n4921), .A(n4914), .ZN(n4915) );
  OAI21_X1 U6067 ( .B1(n4924), .B2(n4916), .A(n4915), .ZN(U3065) );
  INV_X1 U6068 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4923) );
  AOI22_X1 U6069 ( .A1(n6430), .A2(n4917), .B1(n6429), .B2(n3020), .ZN(n4918)
         );
  OAI21_X1 U6070 ( .B1(n6434), .B2(n4919), .A(n4918), .ZN(n4920) );
  AOI21_X1 U6071 ( .B1(n6431), .B2(n4921), .A(n4920), .ZN(n4922) );
  OAI21_X1 U6072 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(U3064) );
  INV_X1 U6073 ( .A(n4624), .ZN(n4925) );
  AOI21_X1 U6074 ( .B1(n4926), .B2(n4925), .A(n4875), .ZN(n6293) );
  INV_X1 U6075 ( .A(n6293), .ZN(n4929) );
  INV_X1 U6076 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4927) );
  OAI222_X1 U6077 ( .A1(n4929), .A2(n5670), .B1(n5677), .B2(n4928), .C1(n4927), 
        .C2(n5669), .ZN(U2852) );
  NOR3_X1 U6078 ( .A1(n4974), .A2(n4931), .A3(n5844), .ZN(n4934) );
  OAI21_X1 U6079 ( .B1(n4934), .B2(n4933), .A(n4932), .ZN(n4939) );
  NOR2_X1 U6080 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4935), .ZN(n4970)
         );
  INV_X1 U6081 ( .A(n4970), .ZN(n4937) );
  AOI211_X1 U6082 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4937), .A(n6351), .B(
        n4936), .ZN(n4938) );
  INV_X1 U6083 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4945) );
  OAI22_X1 U6084 ( .A1(n6354), .A2(n4941), .B1(n5095), .B2(n4940), .ZN(n4969)
         );
  AOI22_X1 U6085 ( .A1(n6412), .A2(n4970), .B1(n6413), .B2(n4969), .ZN(n4942)
         );
  OAI21_X1 U6086 ( .B1(n6416), .B2(n4972), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6087 ( .B1(n6411), .B2(n4974), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6088 ( .B1(n4977), .B2(n4945), .A(n4944), .ZN(U3021) );
  INV_X1 U6089 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6090 ( .A1(n6424), .A2(n4970), .B1(n6425), .B2(n4969), .ZN(n4946)
         );
  OAI21_X1 U6091 ( .B1(n6428), .B2(n4972), .A(n4946), .ZN(n4947) );
  AOI21_X1 U6092 ( .B1(n6423), .B2(n4974), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6093 ( .B1(n4977), .B2(n4949), .A(n4948), .ZN(U3023) );
  AOI22_X1 U6094 ( .A1(n6356), .A2(n4970), .B1(n6355), .B2(n4969), .ZN(n4950)
         );
  OAI21_X1 U6095 ( .B1(n5129), .B2(n4972), .A(n4950), .ZN(n4951) );
  AOI21_X1 U6096 ( .B1(n5126), .B2(n4974), .A(n4951), .ZN(n4952) );
  OAI21_X1 U6097 ( .B1(n4977), .B2(n4953), .A(n4952), .ZN(U3020) );
  AOI22_X1 U6098 ( .A1(n6444), .A2(n4970), .B1(n6446), .B2(n4969), .ZN(n4954)
         );
  OAI21_X1 U6099 ( .B1(n6451), .B2(n4972), .A(n4954), .ZN(n4955) );
  AOI21_X1 U6100 ( .B1(n6442), .B2(n4974), .A(n4955), .ZN(n4956) );
  OAI21_X1 U6101 ( .B1(n4977), .B2(n4957), .A(n4956), .ZN(U3027) );
  INV_X1 U6102 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6103 ( .A1(n6436), .A2(n4970), .B1(n6437), .B2(n4969), .ZN(n4958)
         );
  OAI21_X1 U6104 ( .B1(n6440), .B2(n4972), .A(n4958), .ZN(n4959) );
  AOI21_X1 U6105 ( .B1(n6435), .B2(n4974), .A(n4959), .ZN(n4960) );
  OAI21_X1 U6106 ( .B1(n4977), .B2(n4961), .A(n4960), .ZN(U3026) );
  AOI22_X1 U6107 ( .A1(n6384), .A2(n4970), .B1(n6383), .B2(n4969), .ZN(n4962)
         );
  OAI21_X1 U6108 ( .B1(n5145), .B2(n4972), .A(n4962), .ZN(n4963) );
  AOI21_X1 U6109 ( .B1(n5142), .B2(n4974), .A(n4963), .ZN(n4964) );
  OAI21_X1 U6110 ( .B1(n4977), .B2(n3370), .A(n4964), .ZN(U3025) );
  INV_X1 U6111 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U6112 ( .A1(n6418), .A2(n4970), .B1(n6419), .B2(n4969), .ZN(n4965)
         );
  OAI21_X1 U6113 ( .B1(n6422), .B2(n4972), .A(n4965), .ZN(n4966) );
  AOI21_X1 U6114 ( .B1(n6417), .B2(n4974), .A(n4966), .ZN(n4967) );
  OAI21_X1 U6115 ( .B1(n4977), .B2(n4968), .A(n4967), .ZN(U3022) );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U6117 ( .A1(n6430), .A2(n4970), .B1(n6431), .B2(n4969), .ZN(n4971)
         );
  OAI21_X1 U6118 ( .B1(n6434), .B2(n4972), .A(n4971), .ZN(n4973) );
  AOI21_X1 U6119 ( .B1(n6429), .B2(n4974), .A(n4973), .ZN(n4975) );
  OAI21_X1 U6120 ( .B1(n4977), .B2(n4976), .A(n4975), .ZN(U3024) );
  NAND2_X1 U6121 ( .A1(n4978), .A2(n6450), .ZN(n4979) );
  AOI21_X1 U6122 ( .B1(n4979), .B2(STATEBS16_REG_SCAN_IN), .A(n5844), .ZN(
        n4985) );
  NOR2_X1 U6123 ( .A1(n5095), .A2(n6466), .ZN(n4980) );
  AOI22_X1 U6124 ( .A1(n4985), .A2(n4981), .B1(n6350), .B2(n4980), .ZN(n5016)
         );
  NOR2_X1 U6125 ( .A1(n6351), .A2(n6358), .ZN(n5092) );
  INV_X1 U6126 ( .A(n4981), .ZN(n4984) );
  NOR2_X1 U6127 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4982), .ZN(n4988)
         );
  NOR2_X1 U6128 ( .A1(n4988), .A2(n3174), .ZN(n4983) );
  AOI21_X1 U6129 ( .B1(n4985), .B2(n4984), .A(n4983), .ZN(n4986) );
  OAI211_X1 U6130 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4987), .A(n5092), .B(n4986), .ZN(n5010) );
  NAND2_X1 U6131 ( .A1(n5010), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4991)
         );
  INV_X1 U6132 ( .A(n4988), .ZN(n5011) );
  OAI22_X1 U6133 ( .A1(n5139), .A2(n5011), .B1(n6450), .B2(n6388), .ZN(n4989)
         );
  AOI21_X1 U6134 ( .B1(n5013), .B2(n6385), .A(n4989), .ZN(n4990) );
  OAI211_X1 U6135 ( .C1(n5016), .C2(n5136), .A(n4991), .B(n4990), .ZN(U3105)
         );
  NAND2_X1 U6136 ( .A1(n5010), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4994)
         );
  OAI22_X1 U6137 ( .A1(n5099), .A2(n5011), .B1(n6450), .B2(n6399), .ZN(n4992)
         );
  AOI21_X1 U6138 ( .B1(n5013), .B2(n6395), .A(n4992), .ZN(n4993) );
  OAI211_X1 U6139 ( .C1(n5016), .C2(n5098), .A(n4994), .B(n4993), .ZN(U3107)
         );
  NAND2_X1 U6140 ( .A1(n5010), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4997)
         );
  OAI22_X1 U6141 ( .A1(n5131), .A2(n5011), .B1(n6450), .B2(n6370), .ZN(n4995)
         );
  AOI21_X1 U6142 ( .B1(n5013), .B2(n6367), .A(n4995), .ZN(n4996) );
  OAI211_X1 U6143 ( .C1(n5016), .C2(n5130), .A(n4997), .B(n4996), .ZN(U3101)
         );
  NAND2_X1 U6144 ( .A1(n5010), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5000)
         );
  OAI22_X1 U6145 ( .A1(n5114), .A2(n5011), .B1(n6450), .B2(n6382), .ZN(n4998)
         );
  AOI21_X1 U6146 ( .B1(n5013), .B2(n6379), .A(n4998), .ZN(n4999) );
  OAI211_X1 U6147 ( .C1(n5016), .C2(n5113), .A(n5000), .B(n4999), .ZN(U3104)
         );
  NAND2_X1 U6148 ( .A1(n5010), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5003)
         );
  OAI22_X1 U6149 ( .A1(n5124), .A2(n5011), .B1(n6450), .B2(n6366), .ZN(n5001)
         );
  AOI21_X1 U6150 ( .B1(n5013), .B2(n6363), .A(n5001), .ZN(n5002) );
  OAI211_X1 U6151 ( .C1(n5016), .C2(n5123), .A(n5003), .B(n5002), .ZN(U3100)
         );
  NAND2_X1 U6152 ( .A1(n5010), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5006)
         );
  OAI22_X1 U6153 ( .A1(n5104), .A2(n5011), .B1(n6450), .B2(n6392), .ZN(n5004)
         );
  AOI21_X1 U6154 ( .B1(n5013), .B2(n6389), .A(n5004), .ZN(n5005) );
  OAI211_X1 U6155 ( .C1(n5016), .C2(n5103), .A(n5006), .B(n5005), .ZN(U3106)
         );
  NAND2_X1 U6156 ( .A1(n5010), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5009)
         );
  OAI22_X1 U6157 ( .A1(n5109), .A2(n5011), .B1(n6450), .B2(n6374), .ZN(n5007)
         );
  AOI21_X1 U6158 ( .B1(n5013), .B2(n6371), .A(n5007), .ZN(n5008) );
  OAI211_X1 U6159 ( .C1(n5016), .C2(n5108), .A(n5009), .B(n5008), .ZN(U3102)
         );
  NAND2_X1 U6160 ( .A1(n5010), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5015)
         );
  OAI22_X1 U6161 ( .A1(n5119), .A2(n5011), .B1(n6450), .B2(n6378), .ZN(n5012)
         );
  AOI21_X1 U6162 ( .B1(n5013), .B2(n6375), .A(n5012), .ZN(n5014) );
  OAI211_X1 U6163 ( .C1(n5016), .C2(n5118), .A(n5015), .B(n5014), .ZN(U3103)
         );
  INV_X1 U6164 ( .A(n5017), .ZN(n6142) );
  AOI22_X1 U6165 ( .A1(n6236), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6336), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5018) );
  OAI21_X1 U6166 ( .B1(n6255), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5018), 
        .ZN(n5019) );
  AOI21_X1 U6167 ( .B1(n6225), .B2(n6142), .A(n5019), .ZN(n5020) );
  OAI21_X1 U6168 ( .B1(n5021), .B2(n6229), .A(n5020), .ZN(U2985) );
  CLKBUF_X1 U6169 ( .A(n5022), .Z(n5023) );
  OAI21_X1 U6170 ( .B1(n5025), .B2(n5024), .A(n5023), .ZN(n5026) );
  INV_X1 U6171 ( .A(n5026), .ZN(n6325) );
  AND2_X1 U6172 ( .A1(n6336), .A2(REIP_REG_3__SCAN_IN), .ZN(n6321) );
  AOI21_X1 U6173 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6321), 
        .ZN(n5027) );
  OAI21_X1 U6174 ( .B1(n6255), .B2(n5149), .A(n5027), .ZN(n5028) );
  AOI21_X1 U6175 ( .B1(n6325), .B2(n6251), .A(n5028), .ZN(n5029) );
  OAI21_X1 U6176 ( .B1(n5157), .B2(n5406), .A(n5029), .ZN(U2983) );
  AOI21_X1 U6177 ( .B1(n5033), .B2(n5032), .A(n5031), .ZN(n6085) );
  INV_X1 U6178 ( .A(n6085), .ZN(n5039) );
  INV_X1 U6179 ( .A(n5184), .ZN(n5034) );
  AOI21_X1 U6180 ( .B1(n5036), .B2(n5035), .A(n5034), .ZN(n6078) );
  AOI22_X1 U6181 ( .A1(n5675), .A2(n6078), .B1(EBX_REG_9__SCAN_IN), .B2(n5674), 
        .ZN(n5037) );
  OAI21_X1 U6182 ( .B1(n5039), .B2(n5677), .A(n5037), .ZN(U2850) );
  AOI22_X1 U6183 ( .A1(n5689), .A2(DATAI_9_), .B1(n6156), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5038) );
  OAI21_X1 U6184 ( .B1(n5039), .B2(n5917), .A(n5038), .ZN(U2882) );
  OAI21_X1 U6185 ( .B1(n5042), .B2(n5041), .A(n5040), .ZN(n6294) );
  NAND2_X1 U6186 ( .A1(n6336), .A2(REIP_REG_7__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U6187 ( .A1(n6236), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5043)
         );
  OAI211_X1 U6188 ( .C1(n6255), .C2(n5198), .A(n6291), .B(n5043), .ZN(n5044)
         );
  AOI21_X1 U6189 ( .B1(n5203), .B2(n6225), .A(n5044), .ZN(n5045) );
  OAI21_X1 U6190 ( .B1(n6294), .B2(n6229), .A(n5045), .ZN(U2979) );
  CLKBUF_X1 U6191 ( .A(n5046), .Z(n5047) );
  OR2_X1 U6192 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  NAND2_X1 U6193 ( .A1(n5047), .A2(n5050), .ZN(n6306) );
  NAND2_X1 U6194 ( .A1(n6336), .A2(REIP_REG_5__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U6195 ( .A1(n6236), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5051)
         );
  OAI211_X1 U6196 ( .C1(n6255), .C2(n5068), .A(n6302), .B(n5051), .ZN(n5052)
         );
  AOI21_X1 U6197 ( .B1(n5053), .B2(n6225), .A(n5052), .ZN(n5054) );
  OAI21_X1 U6198 ( .B1(n6229), .B2(n6306), .A(n5054), .ZN(U2981) );
  INV_X1 U6199 ( .A(n5993), .ZN(n6598) );
  NOR3_X1 U6200 ( .A1(n6599), .A2(n3174), .A3(n6598), .ZN(n6481) );
  AND2_X1 U6201 ( .A1(n5056), .A2(n5055), .ZN(n6490) );
  OR2_X1 U6202 ( .A1(n6336), .A2(n6490), .ZN(n5057) );
  OR2_X1 U6203 ( .A1(n6481), .A2(n5057), .ZN(n5058) );
  INV_X1 U6204 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5426) );
  INV_X1 U6205 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5060) );
  XNOR2_X1 U6206 ( .A(n5061), .B(n5060), .ZN(n5450) );
  NOR2_X1 U6207 ( .A1(n5450), .A2(n6571), .ZN(n5062) );
  OAI21_X1 U6208 ( .B1(n5075), .B2(n5523), .A(n6099), .ZN(n6141) );
  INV_X1 U6209 ( .A(n6141), .ZN(n6125) );
  NOR2_X1 U6210 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5070) );
  AND3_X1 U6211 ( .A1(n5063), .A2(n5070), .A3(n5072), .ZN(n5064) );
  INV_X1 U6212 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6520) );
  INV_X1 U6213 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6589) );
  INV_X1 U6214 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6517) );
  INV_X1 U6215 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6515) );
  NOR3_X1 U6216 ( .A1(n6589), .A2(n6517), .A3(n6515), .ZN(n6119) );
  NAND2_X1 U6217 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6119), .ZN(n5065) );
  NOR2_X1 U6218 ( .A1(n6520), .A2(n5065), .ZN(n5195) );
  OAI21_X1 U6219 ( .B1(n6083), .B2(n5195), .A(n6066), .ZN(n6111) );
  OAI21_X1 U6220 ( .B1(n6083), .B2(n5065), .A(n6520), .ZN(n5084) );
  INV_X1 U6221 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5605) );
  NOR2_X1 U6222 ( .A1(n5075), .A2(n5605), .ZN(n5539) );
  NOR2_X1 U6223 ( .A1(n5530), .A2(n5070), .ZN(n5066) );
  AND2_X1 U6224 ( .A1(n5450), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5067) );
  INV_X1 U6225 ( .A(n5068), .ZN(n5080) );
  INV_X1 U6226 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5077) );
  INV_X1 U6227 ( .A(n5070), .ZN(n5069) );
  OR2_X1 U6228 ( .A1(n6596), .A2(n5069), .ZN(n6480) );
  AND2_X1 U6229 ( .A1(n6592), .A2(n6480), .ZN(n5538) );
  NOR2_X1 U6230 ( .A1(n5070), .A2(EBX_REG_31__SCAN_IN), .ZN(n5071) );
  AND2_X1 U6231 ( .A1(n5072), .A2(n5071), .ZN(n5073) );
  NOR2_X1 U6232 ( .A1(n5538), .A2(n5073), .ZN(n5074) );
  OAI22_X1 U6233 ( .A1(n5077), .A2(n6138), .B1(n5076), .B2(n6124), .ZN(n5079)
         );
  NAND2_X1 U6234 ( .A1(n6066), .A2(n5078), .ZN(n6122) );
  INV_X1 U6235 ( .A(n6122), .ZN(n6107) );
  AOI211_X1 U6236 ( .C1(n6102), .C2(n5080), .A(n5079), .B(n6107), .ZN(n5081)
         );
  OAI21_X1 U6237 ( .B1(n6145), .B2(n5082), .A(n5081), .ZN(n5083) );
  AOI21_X1 U6238 ( .B1(n6111), .B2(n5084), .A(n5083), .ZN(n5085) );
  OAI21_X1 U6239 ( .B1(n5086), .B2(n6125), .A(n5085), .ZN(U2822) );
  NOR2_X1 U6240 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5087), .ZN(n5094)
         );
  OAI21_X1 U6241 ( .B1(n5089), .B2(n5141), .A(n5088), .ZN(n5091) );
  INV_X1 U6242 ( .A(n5097), .ZN(n5090) );
  NAND2_X1 U6243 ( .A1(n5091), .A2(n5090), .ZN(n5093) );
  OAI221_X1 U6244 ( .B1(n5094), .B2(n3174), .C1(n5094), .C2(n5093), .A(n5092), 
        .ZN(n5135) );
  NAND2_X1 U6245 ( .A1(n5135), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5102) );
  INV_X1 U6246 ( .A(n5094), .ZN(n5138) );
  NOR2_X1 U6247 ( .A1(n5095), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5096)
         );
  AOI22_X1 U6248 ( .A1(n5097), .A2(n5836), .B1(n6350), .B2(n5096), .ZN(n5137)
         );
  OAI22_X1 U6249 ( .A1(n5099), .A2(n5138), .B1(n5137), .B2(n5098), .ZN(n5100)
         );
  AOI21_X1 U6250 ( .B1(n6442), .B2(n5141), .A(n5100), .ZN(n5101) );
  OAI211_X1 U6251 ( .C1(n5146), .C2(n6451), .A(n5102), .B(n5101), .ZN(U3043)
         );
  NAND2_X1 U6252 ( .A1(n5135), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5107) );
  OAI22_X1 U6253 ( .A1(n5104), .A2(n5138), .B1(n5137), .B2(n5103), .ZN(n5105)
         );
  AOI21_X1 U6254 ( .B1(n6435), .B2(n5141), .A(n5105), .ZN(n5106) );
  OAI211_X1 U6255 ( .C1(n5146), .C2(n6440), .A(n5107), .B(n5106), .ZN(U3042)
         );
  NAND2_X1 U6256 ( .A1(n5135), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5112) );
  OAI22_X1 U6257 ( .A1(n5109), .A2(n5138), .B1(n5137), .B2(n5108), .ZN(n5110)
         );
  AOI21_X1 U6258 ( .B1(n6417), .B2(n5141), .A(n5110), .ZN(n5111) );
  OAI211_X1 U6259 ( .C1(n5146), .C2(n6422), .A(n5112), .B(n5111), .ZN(U3038)
         );
  NAND2_X1 U6260 ( .A1(n5135), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U6261 ( .A1(n5114), .A2(n5138), .B1(n5137), .B2(n5113), .ZN(n5115)
         );
  AOI21_X1 U6262 ( .B1(n6429), .B2(n5141), .A(n5115), .ZN(n5116) );
  OAI211_X1 U6263 ( .C1(n5146), .C2(n6434), .A(n5117), .B(n5116), .ZN(U3040)
         );
  NAND2_X1 U6264 ( .A1(n5135), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5122) );
  OAI22_X1 U6265 ( .A1(n5119), .A2(n5138), .B1(n5137), .B2(n5118), .ZN(n5120)
         );
  AOI21_X1 U6266 ( .B1(n6423), .B2(n5141), .A(n5120), .ZN(n5121) );
  OAI211_X1 U6267 ( .C1(n5146), .C2(n6428), .A(n5122), .B(n5121), .ZN(U3039)
         );
  NAND2_X1 U6268 ( .A1(n5135), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5128) );
  OAI22_X1 U6269 ( .A1(n5124), .A2(n5138), .B1(n5137), .B2(n5123), .ZN(n5125)
         );
  AOI21_X1 U6270 ( .B1(n5126), .B2(n5141), .A(n5125), .ZN(n5127) );
  OAI211_X1 U6271 ( .C1(n5146), .C2(n5129), .A(n5128), .B(n5127), .ZN(U3036)
         );
  NAND2_X1 U6272 ( .A1(n5135), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5134) );
  OAI22_X1 U6273 ( .A1(n5131), .A2(n5138), .B1(n5137), .B2(n5130), .ZN(n5132)
         );
  AOI21_X1 U6274 ( .B1(n6411), .B2(n5141), .A(n5132), .ZN(n5133) );
  OAI211_X1 U6275 ( .C1(n6416), .C2(n5146), .A(n5134), .B(n5133), .ZN(U3037)
         );
  NAND2_X1 U6276 ( .A1(n5135), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5144) );
  OAI22_X1 U6277 ( .A1(n5139), .A2(n5138), .B1(n5137), .B2(n5136), .ZN(n5140)
         );
  AOI21_X1 U6278 ( .B1(n5142), .B2(n5141), .A(n5140), .ZN(n5143) );
  OAI211_X1 U6279 ( .C1(n5146), .C2(n5145), .A(n5144), .B(n5143), .ZN(U3041)
         );
  INV_X1 U6280 ( .A(n6083), .ZN(n6120) );
  NAND2_X1 U6281 ( .A1(n6120), .A2(n6589), .ZN(n6143) );
  INV_X1 U6282 ( .A(n6143), .ZN(n5147) );
  INV_X1 U6283 ( .A(n6066), .ZN(n6132) );
  NOR3_X1 U6284 ( .A1(n5147), .A2(n6132), .A3(n6515), .ZN(n5210) );
  OAI21_X1 U6285 ( .B1(n6083), .B2(n6119), .A(n6066), .ZN(n6118) );
  OAI21_X1 U6286 ( .B1(n5210), .B2(REIP_REG_3__SCAN_IN), .A(n6118), .ZN(n5156)
         );
  NAND2_X1 U6287 ( .A1(n5148), .A2(n6597), .ZN(n6136) );
  INV_X1 U6288 ( .A(n5149), .ZN(n5150) );
  AOI22_X1 U6289 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6133), .B1(n6102), 
        .B2(n5150), .ZN(n5152) );
  NAND2_X1 U6290 ( .A1(n2993), .A2(EBX_REG_3__SCAN_IN), .ZN(n5151) );
  OAI211_X1 U6291 ( .C1(n5153), .C2(n6136), .A(n5152), .B(n5151), .ZN(n5154)
         );
  AOI21_X1 U6292 ( .B1(n6079), .B2(n6322), .A(n5154), .ZN(n5155) );
  OAI211_X1 U6293 ( .C1(n5157), .C2(n6125), .A(n5156), .B(n5155), .ZN(U2824)
         );
  NAND2_X1 U6294 ( .A1(n5159), .A2(n5158), .ZN(n5161) );
  XOR2_X1 U6295 ( .A(n5161), .B(n5160), .Z(n5178) );
  INV_X1 U6296 ( .A(n6088), .ZN(n5164) );
  INV_X1 U6297 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5162) );
  NOR2_X1 U6298 ( .A1(n6281), .A2(n5162), .ZN(n5175) );
  AOI21_X1 U6299 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5175), 
        .ZN(n5163) );
  OAI21_X1 U6300 ( .B1(n6255), .B2(n5164), .A(n5163), .ZN(n5165) );
  AOI21_X1 U6301 ( .B1(n6085), .B2(n6225), .A(n5165), .ZN(n5166) );
  OAI21_X1 U6302 ( .B1(n5178), .B2(n6229), .A(n5166), .ZN(U2977) );
  NOR2_X1 U6303 ( .A1(n6285), .A2(n6290), .ZN(n6284) );
  NOR4_X1 U6304 ( .A1(n5168), .A2(n5170), .A3(n5167), .A4(n6316), .ZN(n5343)
         );
  INV_X1 U6305 ( .A(n5343), .ZN(n5172) );
  NOR2_X1 U6306 ( .A1(n5170), .A2(n5169), .ZN(n5341) );
  OAI21_X1 U6307 ( .B1(n5341), .B2(n5362), .A(n5347), .ZN(n5171) );
  AOI21_X1 U6308 ( .B1(n5345), .B2(n5172), .A(n5171), .ZN(n6295) );
  OAI21_X1 U6309 ( .B1(n5955), .B2(n6284), .A(n6295), .ZN(n6273) );
  INV_X1 U6310 ( .A(n6284), .ZN(n5340) );
  NAND2_X1 U6311 ( .A1(n5341), .A2(n5173), .ZN(n6300) );
  NOR2_X1 U6312 ( .A1(n5340), .A2(n6300), .ZN(n6276) );
  AOI22_X1 U6313 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6273), .B1(n6276), 
        .B2(n5174), .ZN(n5177) );
  AOI21_X1 U6314 ( .B1(n6338), .B2(n6078), .A(n5175), .ZN(n5176) );
  OAI211_X1 U6315 ( .C1(n5178), .C2(n6342), .A(n5177), .B(n5176), .ZN(U3009)
         );
  AND2_X1 U6316 ( .A1(n5180), .A2(n5179), .ZN(n5182) );
  OR2_X1 U6317 ( .A1(n5182), .A2(n5181), .ZN(n6072) );
  AOI22_X1 U6318 ( .A1(n5689), .A2(DATAI_10_), .B1(n6156), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5183) );
  OAI21_X1 U6319 ( .B1(n6072), .B2(n5917), .A(n5183), .ZN(U2881) );
  AOI21_X1 U6320 ( .B1(n5185), .B2(n5184), .A(n5226), .ZN(n6272) );
  AOI22_X1 U6321 ( .A1(n5675), .A2(n6272), .B1(EBX_REG_10__SCAN_IN), .B2(n5674), .ZN(n5186) );
  OAI21_X1 U6322 ( .B1(n6072), .B2(n5677), .A(n5186), .ZN(U2849) );
  NAND2_X1 U6323 ( .A1(n6141), .A2(n5187), .ZN(n5189) );
  OAI21_X1 U6324 ( .B1(n6133), .B2(n6102), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5188) );
  OAI211_X1 U6325 ( .C1(n6136), .C2(n4328), .A(n5189), .B(n5188), .ZN(n5192)
         );
  NAND2_X1 U6326 ( .A1(n6083), .A2(n6066), .ZN(n5569) );
  INV_X1 U6327 ( .A(n5569), .ZN(n5883) );
  INV_X1 U6328 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6583) );
  OAI22_X1 U6329 ( .A1(n5883), .A2(n6583), .B1(n5190), .B2(n6138), .ZN(n5191)
         );
  AOI211_X1 U6330 ( .C1(n6079), .C2(n5193), .A(n5192), .B(n5191), .ZN(n5194)
         );
  INV_X1 U6331 ( .A(n5194), .ZN(U2827) );
  INV_X1 U6332 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6522) );
  AND3_X1 U6333 ( .A1(n6120), .A2(n5195), .A3(n6522), .ZN(n6106) );
  OAI21_X1 U6334 ( .B1(n6106), .B2(n6111), .A(REIP_REG_7__SCAN_IN), .ZN(n5197)
         );
  NAND2_X1 U6335 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5195), .ZN(n5235) );
  OR3_X1 U6336 ( .A1(n6083), .A2(REIP_REG_7__SCAN_IN), .A3(n5235), .ZN(n5196)
         );
  OAI211_X1 U6337 ( .C1(n6135), .C2(n5198), .A(n5197), .B(n5196), .ZN(n5202)
         );
  INV_X1 U6338 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5200) );
  AOI22_X1 U6339 ( .A1(EBX_REG_7__SCAN_IN), .A2(n2993), .B1(n6079), .B2(n6293), 
        .ZN(n5199) );
  OAI211_X1 U6340 ( .C1(n6124), .C2(n5200), .A(n5199), .B(n6122), .ZN(n5201)
         );
  AOI211_X1 U6341 ( .C1(n6112), .C2(n5203), .A(n5202), .B(n5201), .ZN(n5204)
         );
  INV_X1 U6342 ( .A(n5204), .ZN(U2820) );
  INV_X1 U6343 ( .A(n5205), .ZN(n5843) );
  INV_X1 U6344 ( .A(n6254), .ZN(n5206) );
  AOI22_X1 U6345 ( .A1(n6133), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6102), 
        .B2(n5206), .ZN(n5208) );
  NAND2_X1 U6346 ( .A1(n2993), .A2(EBX_REG_2__SCAN_IN), .ZN(n5207) );
  OAI211_X1 U6347 ( .C1(n5843), .C2(n6136), .A(n5208), .B(n5207), .ZN(n5212)
         );
  AOI21_X1 U6348 ( .B1(n6120), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5209) );
  NOR2_X1 U6349 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  AOI211_X1 U6350 ( .C1(n6337), .C2(n6079), .A(n5212), .B(n5211), .ZN(n5213)
         );
  OAI21_X1 U6351 ( .B1(n6125), .B2(n6248), .A(n5213), .ZN(U2825) );
  NAND2_X1 U6352 ( .A1(n6219), .A2(n5215), .ZN(n5216) );
  XNOR2_X1 U6353 ( .A(n5214), .B(n5216), .ZN(n6274) );
  NAND2_X1 U6354 ( .A1(n6274), .A2(n6251), .ZN(n5220) );
  NAND2_X1 U6355 ( .A1(n6336), .A2(REIP_REG_10__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U6356 ( .B1(n5741), .B2(n5217), .A(n6270), .ZN(n5218) );
  AOI21_X1 U6357 ( .B1(n6074), .B2(n6224), .A(n5218), .ZN(n5219) );
  OAI211_X1 U6358 ( .C1(n5406), .C2(n6072), .A(n5220), .B(n5219), .ZN(U2976)
         );
  NOR2_X1 U6359 ( .A1(n5181), .A2(n5221), .ZN(n5222) );
  OR2_X1 U6360 ( .A1(n5229), .A2(n5222), .ZN(n6060) );
  AOI22_X1 U6361 ( .A1(n5689), .A2(DATAI_11_), .B1(n6156), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5223) );
  OAI21_X1 U6362 ( .B1(n6060), .B2(n5917), .A(n5223), .ZN(U2880) );
  INV_X1 U6363 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5228) );
  NOR2_X1 U6364 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  OR2_X1 U6365 ( .A1(n5224), .A2(n5227), .ZN(n6057) );
  OAI222_X1 U6366 ( .A1(n6060), .A2(n5677), .B1(n5228), .B2(n5669), .C1(n5670), 
        .C2(n6057), .ZN(U2848) );
  XOR2_X1 U6367 ( .A(n5230), .B(n5229), .Z(n5252) );
  INV_X1 U6368 ( .A(n5252), .ZN(n5245) );
  AOI22_X1 U6369 ( .A1(n5689), .A2(DATAI_12_), .B1(n6156), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5231) );
  OAI21_X1 U6370 ( .B1(n5245), .B2(n5917), .A(n5231), .ZN(U2879) );
  INV_X1 U6371 ( .A(n5250), .ZN(n5241) );
  OR2_X1 U6372 ( .A1(n5224), .A2(n5233), .ZN(n5234) );
  NAND2_X1 U6373 ( .A1(n5232), .A2(n5234), .ZN(n5243) );
  INV_X1 U6374 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6524) );
  NOR2_X1 U6375 ( .A1(n6524), .A2(n5235), .ZN(n6093) );
  NAND2_X1 U6376 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6093), .ZN(n6065) );
  NAND2_X1 U6377 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6067) );
  NOR2_X1 U6378 ( .A1(n6065), .A2(n6067), .ZN(n6058) );
  NAND2_X1 U6379 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6058), .ZN(n5284) );
  INV_X1 U6380 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U6381 ( .A1(n6120), .A2(n6531), .ZN(n5236) );
  OAI22_X1 U6382 ( .A1(n6145), .A2(n5243), .B1(n5284), .B2(n5236), .ZN(n5240)
         );
  INV_X1 U6383 ( .A(n5284), .ZN(n5237) );
  NOR2_X1 U6384 ( .A1(n6083), .A2(n5237), .ZN(n6059) );
  NOR2_X1 U6385 ( .A1(n6059), .A2(n6132), .ZN(n6047) );
  AOI22_X1 U6386 ( .A1(EBX_REG_12__SCAN_IN), .A2(n2993), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6133), .ZN(n5238) );
  OAI211_X1 U6387 ( .C1(n6047), .C2(n6531), .A(n5238), .B(n6122), .ZN(n5239)
         );
  AOI211_X1 U6388 ( .C1(n6102), .C2(n5241), .A(n5240), .B(n5239), .ZN(n5242)
         );
  OAI21_X1 U6389 ( .B1(n5245), .B2(n6099), .A(n5242), .ZN(U2815) );
  INV_X1 U6390 ( .A(n5243), .ZN(n6258) );
  AOI22_X1 U6391 ( .A1(n6258), .A2(n5675), .B1(EBX_REG_12__SCAN_IN), .B2(n5674), .ZN(n5244) );
  OAI21_X1 U6392 ( .B1(n5245), .B2(n5677), .A(n5244), .ZN(U2847) );
  INV_X1 U6393 ( .A(n5941), .ZN(n5247) );
  NAND2_X1 U6394 ( .A1(n5247), .A2(n5943), .ZN(n5248) );
  XNOR2_X1 U6395 ( .A(n5942), .B(n5248), .ZN(n6259) );
  INV_X1 U6396 ( .A(n6259), .ZN(n5254) );
  AOI22_X1 U6397 ( .A1(n6236), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6336), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5249) );
  OAI21_X1 U6398 ( .B1(n6255), .B2(n5250), .A(n5249), .ZN(n5251) );
  AOI21_X1 U6399 ( .B1(n5252), .B2(n6225), .A(n5251), .ZN(n5253) );
  OAI21_X1 U6400 ( .B1(n5254), .B2(n6229), .A(n5253), .ZN(U2974) );
  NAND2_X1 U6401 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  AND2_X1 U6402 ( .A1(n5258), .A2(n5257), .ZN(n6053) );
  INV_X1 U6403 ( .A(n6053), .ZN(n5263) );
  AOI22_X1 U6404 ( .A1(n5689), .A2(DATAI_13_), .B1(n6156), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5259) );
  OAI21_X1 U6405 ( .B1(n5263), .B2(n5917), .A(n5259), .ZN(U2878) );
  INV_X1 U6406 ( .A(n5267), .ZN(n5260) );
  AOI21_X1 U6407 ( .B1(n5261), .B2(n5232), .A(n5260), .ZN(n6048) );
  AOI22_X1 U6408 ( .A1(n6048), .A2(n5675), .B1(EBX_REG_13__SCAN_IN), .B2(n5674), .ZN(n5262) );
  OAI21_X1 U6409 ( .B1(n5263), .B2(n5677), .A(n5262), .ZN(U2846) );
  OAI21_X1 U6410 ( .B1(n5265), .B2(n5264), .A(n5636), .ZN(n6040) );
  INV_X1 U6411 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6412 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  NAND2_X1 U6413 ( .A1(n5595), .A2(n5268), .ZN(n6037) );
  OAI222_X1 U6414 ( .A1(n6040), .A2(n5677), .B1(n5269), .B2(n5669), .C1(n5670), 
        .C2(n6037), .ZN(U2845) );
  INV_X1 U6415 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5291) );
  INV_X1 U6416 ( .A(n5272), .ZN(n5276) );
  INV_X1 U6417 ( .A(n5273), .ZN(n5274) );
  MUX2_X1 U6418 ( .A(EBX_REG_29__SCAN_IN), .B(n5274), .S(n3938), .Z(n5275) );
  AOI21_X1 U6419 ( .B1(n5276), .B2(n5291), .A(n5275), .ZN(n5277) );
  NAND2_X1 U6420 ( .A1(n5278), .A2(n5277), .ZN(n5533) );
  OAI21_X1 U6421 ( .B1(n5278), .B2(n5277), .A(n5533), .ZN(n5283) );
  OAI222_X1 U6422 ( .A1(n5677), .A2(n5470), .B1(n5291), .B2(n5669), .C1(n5283), 
        .C2(n5670), .ZN(U2830) );
  AND2_X1 U6423 ( .A1(n5453), .A2(n3198), .ZN(n6153) );
  AOI22_X1 U6424 ( .A1(n6153), .A2(DATAI_29_), .B1(n6156), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5282) );
  AND2_X1 U6425 ( .A1(n3161), .A2(n5279), .ZN(n5280) );
  NAND2_X1 U6426 ( .A1(n6157), .A2(DATAI_13_), .ZN(n5281) );
  OAI211_X1 U6427 ( .C1(n5470), .C2(n5917), .A(n5282), .B(n5281), .ZN(U2862)
         );
  INV_X1 U6428 ( .A(n5283), .ZN(n5468) );
  NAND2_X1 U6429 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5868) );
  INV_X1 U6430 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U6431 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5293) );
  NOR2_X1 U6432 ( .A1(n6531), .A2(n5284), .ZN(n6035) );
  NAND3_X1 U6433 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n6035), .ZN(n5292) );
  NOR2_X1 U6434 ( .A1(n6132), .A2(n5292), .ZN(n5599) );
  NAND4_X1 U6435 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5599), .ZN(n5311) );
  NOR3_X1 U6436 ( .A1(n6542), .A2(n5293), .A3(n5311), .ZN(n5882) );
  NAND4_X1 U6437 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5882), .ZN(n5568) );
  NOR2_X1 U6438 ( .A1(n5868), .A2(n5568), .ZN(n5285) );
  NAND2_X1 U6439 ( .A1(n5285), .A2(REIP_REG_26__SCAN_IN), .ZN(n5286) );
  AND2_X1 U6440 ( .A1(n5286), .A2(n5569), .ZN(n5856) );
  AND2_X1 U6441 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5287) );
  NOR2_X1 U6442 ( .A1(n6083), .A2(n5287), .ZN(n5288) );
  OR2_X1 U6443 ( .A1(n5856), .A2(n5288), .ZN(n5556) );
  NAND2_X1 U6444 ( .A1(n5556), .A2(REIP_REG_29__SCAN_IN), .ZN(n5290) );
  AOI22_X1 U6445 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6133), .B1(n6102), 
        .B2(n5471), .ZN(n5289) );
  OAI211_X1 U6446 ( .C1(n5291), .C2(n6138), .A(n5290), .B(n5289), .ZN(n5295)
         );
  NOR2_X1 U6447 ( .A1(n6083), .A2(n5292), .ZN(n5585) );
  NAND4_X1 U6448 ( .A1(n5585), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5314) );
  NOR2_X1 U6449 ( .A1(n5314), .A2(n5293), .ZN(n5906) );
  NAND2_X1 U6450 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5906), .ZN(n5884) );
  INV_X1 U6451 ( .A(n5884), .ZN(n5897) );
  INV_X1 U6452 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6547) );
  INV_X1 U6453 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6545) );
  NOR2_X1 U6454 ( .A1(n6547), .A2(n6545), .ZN(n5885) );
  AND2_X1 U6455 ( .A1(n5897), .A2(n5885), .ZN(n5877) );
  NAND2_X1 U6456 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5877), .ZN(n5867) );
  NOR2_X1 U6457 ( .A1(n5867), .A2(n5868), .ZN(n5857) );
  NAND3_X1 U6458 ( .A1(n5857), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .ZN(n5549) );
  INV_X1 U6459 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6555) );
  NOR3_X1 U6460 ( .A1(n5549), .A2(REIP_REG_29__SCAN_IN), .A3(n6555), .ZN(n5294) );
  AOI211_X1 U6461 ( .C1(n5468), .C2(n6079), .A(n5295), .B(n5294), .ZN(n5296)
         );
  OAI21_X1 U6462 ( .B1(n5470), .B2(n6099), .A(n5296), .ZN(U2798) );
  XNOR2_X1 U6463 ( .A(n5720), .B(n5298), .ZN(n5299) );
  XNOR2_X1 U6464 ( .A(n5300), .B(n5299), .ZN(n5979) );
  INV_X1 U6465 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5301) );
  OAI22_X1 U6466 ( .A1(n5741), .A2(n6038), .B1(n6281), .B2(n5301), .ZN(n5303)
         );
  NOR2_X1 U6467 ( .A1(n6040), .A2(n5406), .ZN(n5302) );
  AOI211_X1 U6468 ( .C1(n6224), .C2(n6041), .A(n5303), .B(n5302), .ZN(n5304)
         );
  OAI21_X1 U6469 ( .B1(n6229), .B2(n5979), .A(n5304), .ZN(U2972) );
  AOI22_X1 U6470 ( .A1(n6153), .A2(DATAI_19_), .B1(n6156), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6471 ( .A1(n6157), .A2(DATAI_3_), .ZN(n5305) );
  OAI211_X1 U6472 ( .C1(n5322), .C2(n5917), .A(n5306), .B(n5305), .ZN(U2872)
         );
  MUX2_X1 U6473 ( .A(n5382), .B(n5308), .S(n5307), .Z(n5657) );
  NOR2_X1 U6474 ( .A1(n5658), .A2(n5657), .ZN(n5660) );
  XNOR2_X1 U6475 ( .A(n5660), .B(n5309), .ZN(n5816) );
  AOI22_X1 U6476 ( .A1(n5816), .A2(n5675), .B1(EBX_REG_19__SCAN_IN), .B2(n5674), .ZN(n5310) );
  OAI21_X1 U6477 ( .B1(n5322), .B2(n5677), .A(n5310), .ZN(U2840) );
  NAND2_X1 U6478 ( .A1(n5569), .A2(n5311), .ZN(n5587) );
  INV_X1 U6479 ( .A(n5587), .ZN(n6017) );
  NOR2_X1 U6480 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5314), .ZN(n6016) );
  OAI21_X1 U6481 ( .B1(n6017), .B2(n6016), .A(REIP_REG_19__SCAN_IN), .ZN(n5312) );
  OAI211_X1 U6482 ( .C1(n6124), .C2(n5313), .A(n5312), .B(n6122), .ZN(n5320)
         );
  INV_X1 U6483 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6540) );
  NOR3_X1 U6484 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5314), .A3(n6540), .ZN(n5319) );
  INV_X1 U6485 ( .A(n5816), .ZN(n5317) );
  AOI22_X1 U6486 ( .A1(n2993), .A2(EBX_REG_19__SCAN_IN), .B1(n5315), .B2(n6102), .ZN(n5316) );
  OAI21_X1 U6487 ( .B1(n5317), .B2(n6145), .A(n5316), .ZN(n5318) );
  NOR3_X1 U6488 ( .A1(n5320), .A2(n5319), .A3(n5318), .ZN(n5321) );
  OAI21_X1 U6489 ( .B1(n5322), .B2(n6099), .A(n5321), .ZN(U2808) );
  XNOR2_X1 U6490 ( .A(n5720), .B(n5964), .ZN(n5324) );
  XNOR2_X1 U6491 ( .A(n5825), .B(n5324), .ZN(n5960) );
  INV_X1 U6492 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5326) );
  INV_X1 U6493 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5325) );
  OAI22_X1 U6494 ( .A1(n5741), .A2(n5326), .B1(n6281), .B2(n5325), .ZN(n5329)
         );
  NOR2_X1 U6495 ( .A1(n5665), .A2(n5406), .ZN(n5328) );
  AOI211_X1 U6496 ( .C1(n6224), .C2(n6031), .A(n5329), .B(n5328), .ZN(n5330)
         );
  OAI21_X1 U6497 ( .B1(n6229), .B2(n5960), .A(n5330), .ZN(U2970) );
  AND2_X1 U6498 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5797) );
  AND2_X1 U6499 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5719) );
  AND2_X1 U6500 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5353) );
  AND3_X1 U6501 ( .A1(n5797), .A2(n5719), .A3(n5353), .ZN(n5366) );
  NAND2_X1 U6502 ( .A1(n5331), .A2(n5366), .ZN(n5332) );
  NAND2_X1 U6503 ( .A1(n5332), .A2(n5720), .ZN(n5336) );
  NAND2_X1 U6504 ( .A1(n5720), .A2(n5337), .ZN(n5459) );
  INV_X1 U6505 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5693) );
  NOR2_X1 U6506 ( .A1(n5824), .A2(n5693), .ZN(n5705) );
  NOR2_X1 U6507 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5803) );
  INV_X1 U6508 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5796) );
  NAND4_X1 U6509 ( .A1(n5803), .A2(n5417), .A3(n5388), .A4(n5796), .ZN(n5333)
         );
  NOR2_X1 U6510 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5333), .ZN(n5334)
         );
  NAND2_X1 U6511 ( .A1(n5457), .A2(n5336), .ZN(n5713) );
  NOR2_X1 U6512 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5704)
         );
  AND2_X1 U6513 ( .A1(n5704), .A2(n5337), .ZN(n5338) );
  NAND2_X1 U6514 ( .A1(n5713), .A2(n5338), .ZN(n5695) );
  NAND2_X1 U6515 ( .A1(n5438), .A2(n5695), .ZN(n5339) );
  XNOR2_X1 U6516 ( .A(n5339), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5376)
         );
  NAND2_X1 U6517 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6275) );
  NOR2_X1 U6518 ( .A1(n5340), .A2(n6275), .ZN(n5956) );
  NAND2_X1 U6519 ( .A1(n5956), .A2(n5341), .ZN(n5361) );
  INV_X1 U6520 ( .A(n5361), .ZN(n5342) );
  NAND2_X1 U6521 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6257) );
  INV_X1 U6522 ( .A(n6257), .ZN(n5973) );
  NAND2_X1 U6523 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5973), .ZN(n5978) );
  OR2_X1 U6524 ( .A1(n5298), .A2(n5978), .ZN(n5958) );
  NOR3_X1 U6525 ( .A1(n5970), .A2(n5964), .A3(n5958), .ZN(n5363) );
  AND2_X1 U6526 ( .A1(n5342), .A2(n5363), .ZN(n5348) );
  AND2_X1 U6527 ( .A1(n5343), .A2(n5956), .ZN(n5360) );
  NAND2_X1 U6528 ( .A1(n5363), .A2(n5360), .ZN(n5344) );
  NAND2_X1 U6529 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  OAI211_X1 U6530 ( .C1(n5348), .C2(n5362), .A(n5347), .B(n5346), .ZN(n5949)
         );
  INV_X1 U6531 ( .A(n5949), .ZN(n5351) );
  NAND2_X1 U6532 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5365) );
  INV_X1 U6533 ( .A(n5365), .ZN(n5349) );
  NAND2_X1 U6534 ( .A1(n5719), .A2(n5349), .ZN(n5416) );
  NAND2_X1 U6535 ( .A1(n5957), .A2(n5416), .ZN(n5350) );
  NAND2_X1 U6536 ( .A1(n5351), .A2(n5350), .ZN(n5810) );
  INV_X1 U6537 ( .A(n5797), .ZN(n5804) );
  AND2_X1 U6538 ( .A1(n5957), .A2(n5804), .ZN(n5352) );
  OR2_X1 U6539 ( .A1(n5810), .A2(n5352), .ZN(n5795) );
  NOR2_X1 U6540 ( .A1(n6331), .A2(n6333), .ZN(n5385) );
  NOR2_X1 U6541 ( .A1(n5385), .A2(n5353), .ZN(n5354) );
  NOR2_X1 U6542 ( .A1(n5795), .A2(n5354), .ZN(n5776) );
  NAND2_X1 U6543 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U6544 ( .A1(n5957), .A2(n5778), .ZN(n5355) );
  NAND2_X1 U6545 ( .A1(n5776), .A2(n5355), .ZN(n5771) );
  AND2_X1 U6546 ( .A1(n6336), .A2(REIP_REG_27__SCAN_IN), .ZN(n5370) );
  INV_X1 U6547 ( .A(n5551), .ZN(n5356) );
  AOI21_X1 U6548 ( .B1(n5357), .B2(n5617), .A(n5356), .ZN(n5608) );
  INV_X1 U6549 ( .A(n5608), .ZN(n5358) );
  NOR2_X1 U6550 ( .A1(n5358), .A2(n6283), .ZN(n5359) );
  AOI211_X1 U6551 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5771), .A(n5370), .B(n5359), .ZN(n5367) );
  NOR2_X1 U6552 ( .A1(n5362), .A2(n5361), .ZN(n5976) );
  INV_X1 U6553 ( .A(n5363), .ZN(n5364) );
  NOR2_X1 U6554 ( .A1(n5831), .A2(n5365), .ZN(n5821) );
  NAND2_X1 U6555 ( .A1(n5821), .A2(n5366), .ZN(n5785) );
  NOR2_X1 U6556 ( .A1(n5785), .A2(n5778), .ZN(n5764) );
  NAND2_X1 U6557 ( .A1(n5764), .A2(n5765), .ZN(n5770) );
  OAI211_X1 U6558 ( .C1(n5376), .C2(n6342), .A(n5367), .B(n5770), .ZN(U2991)
         );
  OAI21_X1 U6559 ( .B1(n5612), .B2(n5369), .A(n5368), .ZN(n5683) );
  INV_X1 U6560 ( .A(n5683), .ZN(n5374) );
  INV_X1 U6561 ( .A(n5562), .ZN(n5372) );
  AOI21_X1 U6562 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5370), 
        .ZN(n5371) );
  OAI21_X1 U6563 ( .B1(n6255), .B2(n5372), .A(n5371), .ZN(n5373) );
  AOI21_X1 U6564 ( .B1(n5374), .B2(n6225), .A(n5373), .ZN(n5375) );
  OAI21_X1 U6565 ( .B1(n5376), .B2(n6229), .A(n5375), .ZN(U2959) );
  NAND2_X1 U6566 ( .A1(n5378), .A2(n5377), .ZN(n5380) );
  XNOR2_X1 U6567 ( .A(n5380), .B(n5379), .ZN(n5400) );
  MUX2_X1 U6568 ( .A(n3938), .B(n5382), .S(n5381), .Z(n5384) );
  XNOR2_X1 U6569 ( .A(n5384), .B(n5383), .ZN(n5904) );
  INV_X1 U6570 ( .A(n5385), .ZN(n5386) );
  AOI21_X1 U6571 ( .B1(n5386), .B2(n5936), .A(n5949), .ZN(n5828) );
  INV_X1 U6572 ( .A(n5828), .ZN(n5387) );
  AOI21_X1 U6573 ( .B1(n5832), .B2(n5957), .A(n5387), .ZN(n5819) );
  NAND2_X1 U6574 ( .A1(n6336), .A2(REIP_REG_20__SCAN_IN), .ZN(n5397) );
  OAI21_X1 U6575 ( .B1(n5819), .B2(n5388), .A(n5397), .ZN(n5389) );
  AOI21_X1 U6576 ( .B1(n6338), .B2(n5904), .A(n5389), .ZN(n5392) );
  INV_X1 U6577 ( .A(n5719), .ZN(n5390) );
  OAI211_X1 U6578 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5821), .B(n5390), .ZN(n5391) );
  OAI211_X1 U6579 ( .C1(n5400), .C2(n6342), .A(n5392), .B(n5391), .ZN(U2998)
         );
  NAND2_X1 U6580 ( .A1(n5592), .A2(n5393), .ZN(n5645) );
  INV_X1 U6581 ( .A(n5652), .ZN(n5927) );
  NAND2_X1 U6582 ( .A1(n6236), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5396)
         );
  OAI211_X1 U6583 ( .C1(n6255), .C2(n5902), .A(n5397), .B(n5396), .ZN(n5398)
         );
  AOI21_X1 U6584 ( .B1(n5927), .B2(n6225), .A(n5398), .ZN(n5399) );
  OAI21_X1 U6585 ( .B1(n5400), .B2(n6229), .A(n5399), .ZN(U2966) );
  OAI21_X1 U6586 ( .B1(n5403), .B2(n5402), .A(n5401), .ZN(n6280) );
  INV_X1 U6587 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5404) );
  OAI22_X1 U6588 ( .A1(n5741), .A2(n5405), .B1(n6281), .B2(n5404), .ZN(n5408)
         );
  NOR2_X1 U6589 ( .A1(n6100), .A2(n5406), .ZN(n5407) );
  AOI211_X1 U6590 ( .C1(n6224), .C2(n6103), .A(n5408), .B(n5407), .ZN(n5409)
         );
  OAI21_X1 U6591 ( .B1(n6229), .B2(n6280), .A(n5409), .ZN(U2978) );
  AOI22_X1 U6592 ( .A1(n5689), .A2(DATAI_14_), .B1(n6156), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5410) );
  OAI21_X1 U6593 ( .B1(n6040), .B2(n5917), .A(n5410), .ZN(U2877) );
  NOR2_X1 U6594 ( .A1(n5633), .A2(n5412), .ZN(n5413) );
  OR2_X1 U6595 ( .A1(n5411), .A2(n5413), .ZN(n5625) );
  OAI21_X1 U6596 ( .B1(n5625), .B2(n6283), .A(n5414), .ZN(n5415) );
  NOR2_X1 U6597 ( .A1(n5831), .A2(n5416), .ZN(n5813) );
  NAND3_X1 U6598 ( .A1(n5813), .A2(n5797), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5418) );
  AOI21_X1 U6599 ( .B1(n5418), .B2(n5417), .A(n5776), .ZN(n5419) );
  AOI21_X1 U6600 ( .B1(n5423), .B2(n6324), .A(n5422), .ZN(n5424) );
  INV_X1 U6601 ( .A(n5424), .ZN(U2994) );
  INV_X1 U6602 ( .A(n5425), .ZN(n5494) );
  OAI22_X1 U6603 ( .A1(n5426), .A2(n6124), .B1(n6135), .B2(n5494), .ZN(n5428)
         );
  INV_X1 U6604 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6560) );
  NOR3_X1 U6605 ( .A1(n5549), .A2(n6560), .A3(n6555), .ZN(n5537) );
  OAI21_X1 U6606 ( .B1(n6083), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n5431) );
  NOR2_X1 U6607 ( .A1(n5556), .A2(n5431), .ZN(n5543) );
  INV_X1 U6608 ( .A(n5543), .ZN(n5432) );
  OAI21_X1 U6609 ( .B1(n5537), .B2(REIP_REG_30__SCAN_IN), .A(n5432), .ZN(n5433) );
  OAI211_X1 U6610 ( .C1(n5437), .C2(n6099), .A(n5434), .B(n5433), .ZN(U2797)
         );
  AOI22_X1 U6611 ( .A1(n6153), .A2(DATAI_30_), .B1(n6156), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6612 ( .A1(n6157), .A2(DATAI_14_), .ZN(n5435) );
  OAI211_X1 U6613 ( .C1(n5437), .C2(n5917), .A(n5436), .B(n5435), .ZN(U2861)
         );
  NAND2_X1 U6614 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5466) );
  AND2_X1 U6615 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U6616 ( .A(n5720), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5712)
         );
  NAND2_X1 U6617 ( .A1(n5713), .A2(n5712), .ZN(n5711) );
  NOR2_X1 U6618 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6619 ( .A1(n5704), .A2(n5439), .ZN(n5463) );
  NOR4_X1 U6620 ( .A1(n5711), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5463), .ZN(n5440) );
  AOI21_X1 U6621 ( .B1(n5481), .B2(n5754), .A(n5440), .ZN(n5442) );
  XNOR2_X1 U6622 ( .A(n5442), .B(n5441), .ZN(n5762) );
  AOI22_X1 U6623 ( .A1(n5446), .A2(EAX_REG_31__SCAN_IN), .B1(n5445), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5447) );
  AND2_X1 U6624 ( .A1(n6336), .A2(REIP_REG_31__SCAN_IN), .ZN(n5758) );
  AOI21_X1 U6625 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5758), 
        .ZN(n5449) );
  OAI21_X1 U6626 ( .B1(n6255), .B2(n5450), .A(n5449), .ZN(n5451) );
  OAI21_X1 U6627 ( .B1(n5762), .B2(n6229), .A(n5452), .ZN(U2955) );
  NAND3_X1 U6628 ( .A1(n5529), .A2(n5454), .A3(n5453), .ZN(n5456) );
  AOI22_X1 U6629 ( .A1(n6153), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6156), .ZN(n5455) );
  NAND2_X1 U6630 ( .A1(n5456), .A2(n5455), .ZN(U2860) );
  NAND2_X1 U6631 ( .A1(n5458), .A2(n5457), .ZN(n5462) );
  INV_X1 U6632 ( .A(n5459), .ZN(n5460) );
  OR2_X1 U6633 ( .A1(n5460), .A2(n5712), .ZN(n5461) );
  AND2_X1 U6634 ( .A1(n6336), .A2(REIP_REG_29__SCAN_IN), .ZN(n5472) );
  INV_X1 U6635 ( .A(n5466), .ZN(n5465) );
  NAND2_X1 U6636 ( .A1(n5764), .A2(n5465), .ZN(n5756) );
  AOI21_X1 U6637 ( .B1(n5466), .B2(n5957), .A(n5771), .ZN(n5753) );
  AND2_X1 U6638 ( .A1(n5753), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5486)
         );
  AOI21_X1 U6639 ( .B1(n5756), .B2(n5479), .A(n5486), .ZN(n5467) );
  AOI211_X1 U6640 ( .C1(n5468), .C2(n6338), .A(n5472), .B(n5467), .ZN(n5469)
         );
  OAI21_X1 U6641 ( .B1(n5478), .B2(n6342), .A(n5469), .ZN(U2989) );
  INV_X1 U6642 ( .A(n5470), .ZN(n5476) );
  INV_X1 U6643 ( .A(n5471), .ZN(n5474) );
  AOI21_X1 U6644 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5472), 
        .ZN(n5473) );
  OAI21_X1 U6645 ( .B1(n6255), .B2(n5474), .A(n5473), .ZN(n5475) );
  AOI21_X1 U6646 ( .B1(n5476), .B2(n6225), .A(n5475), .ZN(n5477) );
  OAI21_X1 U6647 ( .B1(n5478), .B2(n6229), .A(n5477), .ZN(U2957) );
  NAND2_X1 U6648 ( .A1(n5480), .A2(n5479), .ZN(n5483) );
  NAND2_X1 U6649 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  XNOR2_X1 U6650 ( .A(n5484), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5498)
         );
  NOR2_X1 U6651 ( .A1(n5485), .A2(n6283), .ZN(n5490) );
  NOR3_X1 U6652 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5479), 
        .ZN(n5489) );
  AND2_X1 U6653 ( .A1(n6336), .A2(REIP_REG_30__SCAN_IN), .ZN(n5492) );
  INV_X1 U6654 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5487) );
  AOI211_X1 U6655 ( .C1(n5955), .C2(n5776), .A(n5487), .B(n5486), .ZN(n5488)
         );
  NOR4_X1 U6656 ( .A1(n5490), .A2(n5489), .A3(n5492), .A4(n5488), .ZN(n5491)
         );
  OAI21_X1 U6657 ( .B1(n5498), .B2(n6342), .A(n5491), .ZN(U2988) );
  AOI21_X1 U6658 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5492), 
        .ZN(n5493) );
  OAI21_X1 U6659 ( .B1(n6255), .B2(n5494), .A(n5493), .ZN(n5495) );
  AOI21_X1 U6660 ( .B1(n5496), .B2(n6225), .A(n5495), .ZN(n5497) );
  OAI21_X1 U6661 ( .B1(n5498), .B2(n6229), .A(n5497), .ZN(U2956) );
  INV_X1 U6662 ( .A(n5499), .ZN(n5504) );
  AOI21_X1 U6663 ( .B1(n5500), .B2(n5504), .A(n5508), .ZN(n5511) );
  INV_X1 U6664 ( .A(n5501), .ZN(n5507) );
  NOR3_X1 U6665 ( .A1(n6571), .A2(n5503), .A3(n5502), .ZN(n5506) );
  NOR3_X1 U6666 ( .A1(n5504), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6483), 
        .ZN(n5505) );
  AOI211_X1 U6667 ( .C1(n5507), .C2(n6574), .A(n5506), .B(n5505), .ZN(n5509)
         );
  OAI22_X1 U6668 ( .A1(n5511), .A2(n5510), .B1(n5509), .B2(n5508), .ZN(U3459)
         );
  OAI21_X1 U6669 ( .B1(n5513), .B2(n5512), .A(n5524), .ZN(n5517) );
  INV_X1 U6670 ( .A(n5514), .ZN(n5515) );
  OR2_X1 U6671 ( .A1(n5524), .A2(n5515), .ZN(n5516) );
  OAI211_X1 U6672 ( .C1(n5519), .C2(n5518), .A(n5517), .B(n5516), .ZN(n6470)
         );
  INV_X1 U6673 ( .A(n5520), .ZN(n5521) );
  AOI22_X1 U6674 ( .A1(n5524), .A2(n5523), .B1(n5522), .B2(n5521), .ZN(n5994)
         );
  OAI21_X1 U6675 ( .B1(n5526), .B2(n5525), .A(n6603), .ZN(n5527) );
  NAND2_X1 U6676 ( .A1(n5994), .A2(n5527), .ZN(n6469) );
  AND2_X1 U6677 ( .A1(n6469), .A2(n5528), .ZN(n6002) );
  MUX2_X1 U6678 ( .A(MORE_REG_SCAN_IN), .B(n6470), .S(n6002), .Z(U3471) );
  INV_X1 U6679 ( .A(n5529), .ZN(n5546) );
  OAI22_X1 U6680 ( .A1(n5531), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5530), .ZN(n5536) );
  OAI21_X1 U6681 ( .B1(n5534), .B2(n5533), .A(n5532), .ZN(n5535) );
  NAND2_X1 U6682 ( .A1(n5569), .A2(REIP_REG_31__SCAN_IN), .ZN(n5542) );
  INV_X1 U6683 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6564) );
  NAND3_X1 U6684 ( .A1(n5537), .A2(REIP_REG_30__SCAN_IN), .A3(n6564), .ZN(
        n5541) );
  AOI22_X1 U6685 ( .A1(n5539), .A2(n5538), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n6133), .ZN(n5540) );
  OAI211_X1 U6686 ( .C1(n5543), .C2(n5542), .A(n5541), .B(n5540), .ZN(n5544)
         );
  AOI21_X1 U6687 ( .B1(n3023), .B2(n6079), .A(n5544), .ZN(n5545) );
  OAI21_X1 U6688 ( .B1(n5546), .B2(n6099), .A(n5545), .ZN(U2796) );
  INV_X1 U6689 ( .A(n5701), .ZN(n5680) );
  INV_X1 U6690 ( .A(n5549), .ZN(n5560) );
  NAND2_X1 U6691 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  NAND2_X1 U6692 ( .A1(n5553), .A2(n5552), .ZN(n5763) );
  OAI22_X1 U6693 ( .A1(n5554), .A2(n6124), .B1(n6135), .B2(n5699), .ZN(n5555)
         );
  AOI21_X1 U6694 ( .B1(n2993), .B2(EBX_REG_28__SCAN_IN), .A(n5555), .ZN(n5558)
         );
  NAND2_X1 U6695 ( .A1(n5556), .A2(REIP_REG_28__SCAN_IN), .ZN(n5557) );
  OAI211_X1 U6696 ( .C1(n5763), .C2(n6145), .A(n5558), .B(n5557), .ZN(n5559)
         );
  AOI21_X1 U6697 ( .B1(n5560), .B2(n6555), .A(n5559), .ZN(n5561) );
  OAI21_X1 U6698 ( .B1(n5680), .B2(n6099), .A(n5561), .ZN(U2799) );
  NAND2_X1 U6699 ( .A1(n5856), .A2(REIP_REG_27__SCAN_IN), .ZN(n5564) );
  AOI22_X1 U6700 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6133), .B1(n6102), 
        .B2(n5562), .ZN(n5563) );
  OAI211_X1 U6701 ( .C1(n6138), .C2(n4029), .A(n5564), .B(n5563), .ZN(n5565)
         );
  AOI21_X1 U6702 ( .B1(n5608), .B2(n6079), .A(n5565), .ZN(n5567) );
  INV_X1 U6703 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6553) );
  NAND3_X1 U6704 ( .A1(n5857), .A2(REIP_REG_26__SCAN_IN), .A3(n6553), .ZN(
        n5566) );
  OAI211_X1 U6705 ( .C1(n5683), .C2(n6099), .A(n5567), .B(n5566), .ZN(U2800)
         );
  INV_X1 U6706 ( .A(n5625), .ZN(n5575) );
  INV_X1 U6707 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U6708 ( .A1(n5569), .A2(n5568), .ZN(n5861) );
  OAI22_X1 U6709 ( .A1(n5571), .A2(n6124), .B1(n5570), .B2(n6135), .ZN(n5572)
         );
  AOI21_X1 U6710 ( .B1(EBX_REG_24__SCAN_IN), .B2(n2993), .A(n5572), .ZN(n5573)
         );
  OAI221_X1 U6711 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5867), .C1(n6549), .C2(
        n5861), .A(n5573), .ZN(n5574) );
  AOI21_X1 U6712 ( .B1(n6079), .B2(n5575), .A(n5574), .ZN(n5576) );
  OAI21_X1 U6713 ( .B1(n5686), .B2(n6099), .A(n5576), .ZN(U2803) );
  INV_X1 U6714 ( .A(n5654), .ZN(n5577) );
  AOI21_X1 U6715 ( .B1(n5579), .B2(n5578), .A(n5577), .ZN(n6150) );
  INV_X1 U6716 ( .A(n6150), .ZN(n5664) );
  NAND2_X1 U6717 ( .A1(n5580), .A2(n5581), .ZN(n5582) );
  AND2_X1 U6718 ( .A1(n5658), .A2(n5582), .ZN(n5950) );
  INV_X1 U6719 ( .A(n5938), .ZN(n5584) );
  NAND2_X1 U6720 ( .A1(n2993), .A2(EBX_REG_17__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U6721 ( .C1(n5584), .C2(n6135), .A(n5583), .B(n6122), .ZN(n5590)
         );
  INV_X1 U6722 ( .A(n5585), .ZN(n5597) );
  INV_X1 U6723 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6536) );
  NOR2_X1 U6724 ( .A1(n5597), .A2(n6536), .ZN(n6024) );
  AOI21_X1 U6725 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6024), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5588) );
  OAI22_X1 U6726 ( .A1(n5588), .A2(n5587), .B1(n5586), .B2(n6124), .ZN(n5589)
         );
  AOI211_X1 U6727 ( .C1(n6079), .C2(n5950), .A(n5590), .B(n5589), .ZN(n5591)
         );
  OAI21_X1 U6728 ( .B1(n5664), .B2(n6099), .A(n5591), .ZN(U2810) );
  AOI21_X1 U6729 ( .B1(n5593), .B2(n5636), .A(n5592), .ZN(n5750) );
  INV_X1 U6730 ( .A(n5750), .ZN(n5691) );
  AND2_X1 U6731 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  NOR2_X1 U6732 ( .A1(n5667), .A2(n5596), .ZN(n5966) );
  NOR2_X1 U6733 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5597), .ZN(n6025) );
  INV_X1 U6734 ( .A(n6025), .ZN(n5598) );
  OAI21_X1 U6735 ( .B1(n6135), .B2(n5748), .A(n5598), .ZN(n5603) );
  NOR2_X1 U6736 ( .A1(n5883), .A2(n5599), .ZN(n6036) );
  AOI22_X1 U6737 ( .A1(EBX_REG_15__SCAN_IN), .A2(n2993), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6036), .ZN(n5600) );
  OAI211_X1 U6738 ( .C1(n6124), .C2(n5601), .A(n5600), .B(n6122), .ZN(n5602)
         );
  AOI211_X1 U6739 ( .C1(n5966), .C2(n6079), .A(n5603), .B(n5602), .ZN(n5604)
         );
  OAI21_X1 U6740 ( .B1(n5691), .B2(n6099), .A(n5604), .ZN(U2812) );
  INV_X1 U6741 ( .A(n3023), .ZN(n5606) );
  OAI22_X1 U6742 ( .A1(n5606), .A2(n5670), .B1(n5669), .B2(n5605), .ZN(U2828)
         );
  INV_X1 U6743 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5607) );
  OAI222_X1 U6744 ( .A1(n5677), .A2(n5680), .B1(n5607), .B2(n5669), .C1(n5763), 
        .C2(n5670), .ZN(U2831) );
  AOI22_X1 U6745 ( .A1(n5608), .A2(n5675), .B1(EBX_REG_27__SCAN_IN), .B2(n5674), .ZN(n5609) );
  OAI21_X1 U6746 ( .B1(n5683), .B2(n5677), .A(n5609), .ZN(U2832) );
  AND2_X1 U6747 ( .A1(n5610), .A2(n5611), .ZN(n5613) );
  OR2_X1 U6748 ( .A1(n5613), .A2(n5612), .ZN(n5913) );
  INV_X1 U6749 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6750 ( .A1(n5614), .A2(n5615), .ZN(n5616) );
  NAND2_X1 U6751 ( .A1(n5617), .A2(n5616), .ZN(n5854) );
  OAI222_X1 U6752 ( .A1(n5677), .A2(n5913), .B1(n5618), .B2(n5669), .C1(n5854), 
        .C2(n5670), .ZN(U2833) );
  NAND2_X1 U6753 ( .A1(n4170), .A2(n5619), .ZN(n5620) );
  AND2_X1 U6754 ( .A1(n5610), .A2(n5620), .ZN(n5918) );
  OR2_X1 U6755 ( .A1(n5411), .A2(n5621), .ZN(n5622) );
  NAND2_X1 U6756 ( .A1(n5614), .A2(n5622), .ZN(n5872) );
  OAI22_X1 U6757 ( .A1(n5872), .A2(n5670), .B1(n5865), .B2(n5669), .ZN(n5623)
         );
  AOI21_X1 U6758 ( .B1(n5918), .B2(n5672), .A(n5623), .ZN(n5624) );
  INV_X1 U6759 ( .A(n5624), .ZN(U2834) );
  INV_X1 U6760 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5626) );
  OAI222_X1 U6761 ( .A1(n5677), .A2(n5686), .B1(n5626), .B2(n5669), .C1(n5625), 
        .C2(n5670), .ZN(U2835) );
  NOR2_X1 U6762 ( .A1(n5636), .A2(n5627), .ZN(n5638) );
  NOR2_X1 U6763 ( .A1(n5638), .A2(n5628), .ZN(n5629) );
  INV_X1 U6764 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6755) );
  AND2_X1 U6765 ( .A1(n5632), .A2(n5631), .ZN(n5634) );
  OR2_X1 U6766 ( .A1(n5634), .A2(n5633), .ZN(n5874) );
  OAI222_X1 U6767 ( .A1(n5677), .A2(n5875), .B1(n5669), .B2(n6755), .C1(n5874), 
        .C2(n5670), .ZN(U2836) );
  OR2_X1 U6768 ( .A1(n5636), .A2(n5635), .ZN(n5643) );
  AND2_X1 U6769 ( .A1(n5643), .A2(n5637), .ZN(n5639) );
  INV_X1 U6770 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5642) );
  XNOR2_X1 U6771 ( .A(n5640), .B(n5641), .ZN(n5889) );
  OAI222_X1 U6772 ( .A1(n5677), .A2(n5732), .B1(n5642), .B2(n5669), .C1(n5889), 
        .C2(n5670), .ZN(U2837) );
  INV_X1 U6773 ( .A(n5643), .ZN(n5644) );
  INV_X1 U6774 ( .A(n5924), .ZN(n5650) );
  INV_X1 U6775 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5895) );
  OR2_X1 U6776 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  NAND2_X1 U6777 ( .A1(n5640), .A2(n5649), .ZN(n5901) );
  OAI222_X1 U6778 ( .A1(n5650), .A2(n5677), .B1(n5669), .B2(n5895), .C1(n5901), 
        .C2(n5670), .ZN(U2838) );
  AOI22_X1 U6779 ( .A1(n5904), .A2(n5675), .B1(EBX_REG_20__SCAN_IN), .B2(n5674), .ZN(n5651) );
  OAI21_X1 U6780 ( .B1(n5652), .B2(n5677), .A(n5651), .ZN(U2839) );
  NAND2_X1 U6781 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  INV_X1 U6782 ( .A(n6147), .ZN(n5662) );
  AND2_X1 U6783 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  NOR2_X1 U6784 ( .A1(n5660), .A2(n5659), .ZN(n5830) );
  INV_X1 U6785 ( .A(n5830), .ZN(n6020) );
  OAI222_X1 U6786 ( .A1(n5662), .A2(n5677), .B1(n5661), .B2(n5669), .C1(n5670), 
        .C2(n6020), .ZN(U2841) );
  AOI22_X1 U6787 ( .A1(n5950), .A2(n5675), .B1(EBX_REG_17__SCAN_IN), .B2(n5674), .ZN(n5663) );
  OAI21_X1 U6788 ( .B1(n5664), .B2(n5677), .A(n5663), .ZN(U2842) );
  INV_X1 U6789 ( .A(n5665), .ZN(n6155) );
  OR2_X1 U6790 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  NAND2_X1 U6791 ( .A1(n5580), .A2(n5668), .ZN(n6034) );
  OAI22_X1 U6792 ( .A1(n6034), .A2(n5670), .B1(n6029), .B2(n5669), .ZN(n5671)
         );
  AOI21_X1 U6793 ( .B1(n6155), .B2(n5672), .A(n5671), .ZN(n5673) );
  INV_X1 U6794 ( .A(n5673), .ZN(U2843) );
  AOI22_X1 U6795 ( .A1(n5966), .A2(n5675), .B1(EBX_REG_15__SCAN_IN), .B2(n5674), .ZN(n5676) );
  OAI21_X1 U6796 ( .B1(n5691), .B2(n5677), .A(n5676), .ZN(U2844) );
  AOI22_X1 U6797 ( .A1(n6153), .A2(DATAI_28_), .B1(n6156), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6798 ( .A1(n6157), .A2(DATAI_12_), .ZN(n5678) );
  OAI211_X1 U6799 ( .C1(n5680), .C2(n5917), .A(n5679), .B(n5678), .ZN(U2863)
         );
  AOI22_X1 U6800 ( .A1(n6153), .A2(DATAI_27_), .B1(n6156), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6801 ( .A1(n6157), .A2(DATAI_11_), .ZN(n5681) );
  OAI211_X1 U6802 ( .C1(n5683), .C2(n5917), .A(n5682), .B(n5681), .ZN(U2864)
         );
  AOI22_X1 U6803 ( .A1(n6153), .A2(DATAI_24_), .B1(n6156), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U6804 ( .A1(n6157), .A2(DATAI_8_), .ZN(n5684) );
  OAI211_X1 U6805 ( .C1(n5686), .C2(n5917), .A(n5685), .B(n5684), .ZN(U2867)
         );
  AOI22_X1 U6806 ( .A1(n6157), .A2(DATAI_7_), .B1(n6156), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U6807 ( .A1(n6153), .A2(DATAI_23_), .ZN(n5687) );
  OAI211_X1 U6808 ( .C1(n5875), .C2(n5917), .A(n5688), .B(n5687), .ZN(U2868)
         );
  AOI22_X1 U6809 ( .A1(n5689), .A2(DATAI_15_), .B1(n6156), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5690) );
  OAI21_X1 U6810 ( .B1(n5691), .B2(n5917), .A(n5690), .ZN(U2876) );
  AND2_X1 U6811 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5692)
         );
  AND2_X1 U6812 ( .A1(n5693), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5694)
         );
  XNOR2_X1 U6813 ( .A(n5697), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5775)
         );
  AND2_X1 U6814 ( .A1(n6336), .A2(REIP_REG_28__SCAN_IN), .ZN(n5768) );
  AOI21_X1 U6815 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5768), 
        .ZN(n5698) );
  OAI21_X1 U6816 ( .B1(n6255), .B2(n5699), .A(n5698), .ZN(n5700) );
  AOI21_X1 U6817 ( .B1(n5701), .B2(n6225), .A(n5700), .ZN(n5702) );
  OAI21_X1 U6818 ( .B1(n6229), .B2(n5775), .A(n5702), .ZN(U2958) );
  NOR2_X1 U6819 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  XOR2_X1 U6820 ( .A(n5703), .B(n5706), .Z(n5784) );
  INV_X1 U6821 ( .A(n5913), .ZN(n5709) );
  AND2_X1 U6822 ( .A1(n6336), .A2(REIP_REG_26__SCAN_IN), .ZN(n5777) );
  AOI21_X1 U6823 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5777), 
        .ZN(n5707) );
  OAI21_X1 U6824 ( .B1(n6255), .B2(n5852), .A(n5707), .ZN(n5708) );
  AOI21_X1 U6825 ( .B1(n5709), .B2(n6225), .A(n5708), .ZN(n5710) );
  OAI21_X1 U6826 ( .B1(n5784), .B2(n6229), .A(n5710), .ZN(U2960) );
  OAI21_X1 U6827 ( .B1(n5713), .B2(n5712), .A(n5711), .ZN(n5791) );
  INV_X1 U6828 ( .A(n5791), .ZN(n5718) );
  INV_X1 U6829 ( .A(n5862), .ZN(n5715) );
  AND2_X1 U6830 ( .A1(n6336), .A2(REIP_REG_25__SCAN_IN), .ZN(n5786) );
  AOI21_X1 U6831 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5786), 
        .ZN(n5714) );
  OAI21_X1 U6832 ( .B1(n6255), .B2(n5715), .A(n5714), .ZN(n5716) );
  AOI21_X1 U6833 ( .B1(n5918), .B2(n6225), .A(n5716), .ZN(n5717) );
  OAI21_X1 U6834 ( .B1(n5718), .B2(n6229), .A(n5717), .ZN(U2961) );
  NAND3_X1 U6835 ( .A1(n5720), .A2(n5797), .A3(n5719), .ZN(n5722) );
  OAI21_X1 U6836 ( .B1(n2996), .B2(n5722), .A(n5721), .ZN(n5724) );
  XNOR2_X1 U6837 ( .A(n5724), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5800)
         );
  AND2_X1 U6838 ( .A1(n6336), .A2(REIP_REG_23__SCAN_IN), .ZN(n5794) );
  NOR2_X1 U6839 ( .A1(n5741), .A2(n5881), .ZN(n5725) );
  AOI211_X1 U6840 ( .C1(n6224), .C2(n5873), .A(n5794), .B(n5725), .ZN(n5728)
         );
  INV_X1 U6841 ( .A(n5875), .ZN(n5726) );
  NAND2_X1 U6842 ( .A1(n5726), .A2(n6225), .ZN(n5727) );
  OAI211_X1 U6843 ( .C1(n5800), .C2(n6229), .A(n5728), .B(n5727), .ZN(U2963)
         );
  AOI21_X1 U6844 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5720), .A(n5729), 
        .ZN(n5730) );
  XNOR2_X1 U6845 ( .A(n5731), .B(n5730), .ZN(n5808) );
  NOR2_X1 U6846 ( .A1(n6281), .A2(n6547), .ZN(n5802) );
  AOI21_X1 U6847 ( .B1(n6236), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5802), 
        .ZN(n5733) );
  OAI21_X1 U6848 ( .B1(n6255), .B2(n5893), .A(n5733), .ZN(n5734) );
  AOI21_X1 U6849 ( .B1(n5921), .B2(n6225), .A(n5734), .ZN(n5735) );
  OAI21_X1 U6850 ( .B1(n5808), .B2(n6229), .A(n5735), .ZN(U2964) );
  NAND2_X1 U6851 ( .A1(n5736), .A2(n5737), .ZN(n5739) );
  AOI21_X1 U6852 ( .B1(n5740), .B2(n5739), .A(n5738), .ZN(n5815) );
  NOR2_X1 U6853 ( .A1(n6281), .A2(n6545), .ZN(n5809) );
  NOR2_X1 U6854 ( .A1(n5741), .A2(n5894), .ZN(n5742) );
  AOI211_X1 U6855 ( .C1(n6224), .C2(n5898), .A(n5809), .B(n5742), .ZN(n5744)
         );
  NAND2_X1 U6856 ( .A1(n5924), .A2(n6225), .ZN(n5743) );
  OAI211_X1 U6857 ( .C1(n5815), .C2(n6229), .A(n5744), .B(n5743), .ZN(U2965)
         );
  XNOR2_X1 U6858 ( .A(n5720), .B(n5970), .ZN(n5746) );
  XNOR2_X1 U6859 ( .A(n5745), .B(n5746), .ZN(n5967) );
  INV_X1 U6860 ( .A(n5967), .ZN(n5752) );
  AOI22_X1 U6861 ( .A1(n6236), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6336), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5747) );
  OAI21_X1 U6862 ( .B1(n6255), .B2(n5748), .A(n5747), .ZN(n5749) );
  AOI21_X1 U6863 ( .B1(n5750), .B2(n6225), .A(n5749), .ZN(n5751) );
  OAI21_X1 U6864 ( .B1(n5752), .B2(n6229), .A(n5751), .ZN(U2971) );
  OAI21_X1 U6865 ( .B1(n5955), .B2(n5754), .A(n5753), .ZN(n5759) );
  INV_X1 U6866 ( .A(n5754), .ZN(n5755) );
  NOR3_X1 U6867 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5755), 
        .ZN(n5757) );
  AOI211_X1 U6868 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n5759), .A(n5758), .B(n5757), .ZN(n5761) );
  NAND2_X1 U6869 ( .A1(n3023), .A2(n6338), .ZN(n5760) );
  OAI211_X1 U6870 ( .C1(n5762), .C2(n6342), .A(n5761), .B(n5760), .ZN(U2987)
         );
  INV_X1 U6871 ( .A(n5763), .ZN(n5769) );
  INV_X1 U6872 ( .A(n5764), .ZN(n5766) );
  NOR3_X1 U6873 ( .A1(n5766), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5765), 
        .ZN(n5767) );
  AOI211_X1 U6874 ( .C1(n5769), .C2(n6338), .A(n5768), .B(n5767), .ZN(n5774)
         );
  INV_X1 U6875 ( .A(n5770), .ZN(n5772) );
  OAI21_X1 U6876 ( .B1(n5772), .B2(n5771), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n5773) );
  OAI211_X1 U6877 ( .C1(n5775), .C2(n6342), .A(n5774), .B(n5773), .ZN(U2990)
         );
  INV_X1 U6878 ( .A(n5776), .ZN(n5787) );
  AOI21_X1 U6879 ( .B1(n5787), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5777), 
        .ZN(n5781) );
  OAI21_X1 U6880 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5778), .ZN(n5779) );
  OR2_X1 U6881 ( .A1(n5785), .A2(n5779), .ZN(n5780) );
  OAI211_X1 U6882 ( .C1(n5854), .C2(n6283), .A(n5781), .B(n5780), .ZN(n5782)
         );
  INV_X1 U6883 ( .A(n5782), .ZN(n5783) );
  OAI21_X1 U6884 ( .B1(n5784), .B2(n6342), .A(n5783), .ZN(U2992) );
  NOR2_X1 U6885 ( .A1(n5785), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5790)
         );
  AOI21_X1 U6886 ( .B1(n5787), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5786), 
        .ZN(n5788) );
  OAI21_X1 U6887 ( .B1(n5872), .B2(n6283), .A(n5788), .ZN(n5789) );
  AOI211_X1 U6888 ( .C1(n5791), .C2(n6324), .A(n5790), .B(n5789), .ZN(n5792)
         );
  INV_X1 U6889 ( .A(n5792), .ZN(U2993) );
  NOR2_X1 U6890 ( .A1(n5874), .A2(n6283), .ZN(n5793) );
  AOI211_X1 U6891 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5795), .A(n5794), .B(n5793), .ZN(n5799) );
  NAND3_X1 U6892 ( .A1(n5813), .A2(n5797), .A3(n5796), .ZN(n5798) );
  OAI211_X1 U6893 ( .C1(n5800), .C2(n6342), .A(n5799), .B(n5798), .ZN(U2995)
         );
  NOR2_X1 U6894 ( .A1(n5889), .A2(n6283), .ZN(n5801) );
  AOI211_X1 U6895 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5810), .A(n5802), .B(n5801), .ZN(n5807) );
  INV_X1 U6896 ( .A(n5803), .ZN(n5805) );
  NAND3_X1 U6897 ( .A1(n5813), .A2(n5805), .A3(n5804), .ZN(n5806) );
  OAI211_X1 U6898 ( .C1(n5808), .C2(n6342), .A(n5807), .B(n5806), .ZN(U2996)
         );
  AOI21_X1 U6899 ( .B1(n5810), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5809), 
        .ZN(n5811) );
  OAI21_X1 U6900 ( .B1(n5901), .B2(n6283), .A(n5811), .ZN(n5812) );
  AOI21_X1 U6901 ( .B1(n5813), .B2(n6785), .A(n5812), .ZN(n5814) );
  OAI21_X1 U6902 ( .B1(n5815), .B2(n6342), .A(n5814), .ZN(U2997) );
  NAND2_X1 U6903 ( .A1(n5816), .A2(n6338), .ZN(n5818) );
  OAI211_X1 U6904 ( .C1(n5819), .C2(n6768), .A(n5818), .B(n5817), .ZN(n5820)
         );
  AOI21_X1 U6905 ( .B1(n5821), .B2(n6768), .A(n5820), .ZN(n5822) );
  OAI21_X1 U6906 ( .B1(n5823), .B2(n6342), .A(n5822), .ZN(U2999) );
  NAND3_X1 U6907 ( .A1(n5825), .A2(n5824), .A3(n5964), .ZN(n5933) );
  NOR3_X1 U6908 ( .A1(n5825), .A2(n5824), .A3(n5964), .ZN(n5935) );
  NAND2_X1 U6909 ( .A1(n5935), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5826) );
  OAI21_X1 U6910 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5933), .A(n5826), 
        .ZN(n5827) );
  XNOR2_X1 U6911 ( .A(n5827), .B(n5832), .ZN(n5930) );
  INV_X1 U6912 ( .A(n5930), .ZN(n5835) );
  OAI22_X1 U6913 ( .A1(n5828), .A2(n5832), .B1(n6281), .B2(n6540), .ZN(n5829)
         );
  AOI21_X1 U6914 ( .B1(n6338), .B2(n5830), .A(n5829), .ZN(n5834) );
  INV_X1 U6915 ( .A(n5831), .ZN(n5951) );
  NAND3_X1 U6916 ( .A1(n5951), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5832), .ZN(n5833) );
  OAI211_X1 U6917 ( .C1(n5835), .C2(n6342), .A(n5834), .B(n5833), .ZN(U3000)
         );
  OAI21_X1 U6918 ( .B1(n5837), .B2(STATEBS16_REG_SCAN_IN), .A(n5836), .ZN(
        n5838) );
  OAI22_X1 U6919 ( .A1(n5838), .A2(n5840), .B1(n6137), .B2(n5842), .ZN(n5839)
         );
  MUX2_X1 U6920 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5839), .S(n6348), 
        .Z(U3464) );
  XNOR2_X1 U6921 ( .A(n5841), .B(n5840), .ZN(n5845) );
  OAI22_X1 U6922 ( .A1(n5845), .A2(n5844), .B1(n5843), .B2(n5842), .ZN(n5846)
         );
  MUX2_X1 U6923 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5846), .S(n6348), 
        .Z(U3463) );
  INV_X1 U6924 ( .A(n5847), .ZN(n5850) );
  INV_X1 U6925 ( .A(n5848), .ZN(n5849) );
  OAI22_X1 U6926 ( .A1(n5850), .A2(n6579), .B1(n5849), .B2(n6483), .ZN(n5851)
         );
  MUX2_X1 U6927 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5851), .S(n6576), 
        .Z(U3456) );
  AND2_X1 U6928 ( .A1(n6175), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI22_X1 U6929 ( .A1(n6737), .A2(n6124), .B1(n5852), .B2(n6135), .ZN(n5853)
         );
  AOI21_X1 U6930 ( .B1(EBX_REG_26__SCAN_IN), .B2(n2993), .A(n5853), .ZN(n5860)
         );
  OAI22_X1 U6931 ( .A1(n5913), .A2(n6099), .B1(n6145), .B2(n5854), .ZN(n5855)
         );
  INV_X1 U6932 ( .A(n5855), .ZN(n5859) );
  OAI21_X1 U6933 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5857), .A(n5856), .ZN(n5858) );
  NAND3_X1 U6934 ( .A1(n5860), .A2(n5859), .A3(n5858), .ZN(U2801) );
  INV_X1 U6935 ( .A(n5861), .ZN(n5878) );
  NAND2_X1 U6936 ( .A1(n5878), .A2(REIP_REG_25__SCAN_IN), .ZN(n5864) );
  AOI22_X1 U6937 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6133), .B1(n6102), 
        .B2(n5862), .ZN(n5863) );
  OAI211_X1 U6938 ( .C1(n5865), .C2(n6138), .A(n5864), .B(n5863), .ZN(n5866)
         );
  AOI21_X1 U6939 ( .B1(n5918), .B2(n6112), .A(n5866), .ZN(n5871) );
  INV_X1 U6940 ( .A(n5867), .ZN(n5869) );
  OAI211_X1 U6941 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5869), .B(n5868), .ZN(n5870) );
  OAI211_X1 U6942 ( .C1(n5872), .C2(n6145), .A(n5871), .B(n5870), .ZN(U2802)
         );
  AOI22_X1 U6943 ( .A1(EBX_REG_23__SCAN_IN), .A2(n2993), .B1(n5873), .B2(n6102), .ZN(n5880) );
  OAI22_X1 U6944 ( .A1(n5875), .A2(n6099), .B1(n5874), .B2(n6145), .ZN(n5876)
         );
  AOI221_X1 U6945 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5878), .C1(n5877), .C2(
        n5878), .A(n5876), .ZN(n5879) );
  OAI211_X1 U6946 ( .C1(n5881), .C2(n6124), .A(n5880), .B(n5879), .ZN(U2804)
         );
  NOR2_X1 U6947 ( .A1(n5883), .A2(n5882), .ZN(n5905) );
  AOI211_X1 U6948 ( .C1(n6547), .C2(n6545), .A(n5885), .B(n5884), .ZN(n5888)
         );
  AOI22_X1 U6949 ( .A1(EBX_REG_22__SCAN_IN), .A2(n2993), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6133), .ZN(n5886) );
  INV_X1 U6950 ( .A(n5886), .ZN(n5887) );
  AOI211_X1 U6951 ( .C1(REIP_REG_22__SCAN_IN), .C2(n5905), .A(n5888), .B(n5887), .ZN(n5892) );
  INV_X1 U6952 ( .A(n5889), .ZN(n5890) );
  AOI22_X1 U6953 ( .A1(n5921), .A2(n6112), .B1(n5890), .B2(n6079), .ZN(n5891)
         );
  OAI211_X1 U6954 ( .C1(n5893), .C2(n6135), .A(n5892), .B(n5891), .ZN(U2805)
         );
  OAI22_X1 U6955 ( .A1(n5895), .A2(n6138), .B1(n5894), .B2(n6124), .ZN(n5896)
         );
  AOI221_X1 U6956 ( .B1(n5905), .B2(REIP_REG_21__SCAN_IN), .C1(n5897), .C2(
        n6545), .A(n5896), .ZN(n5900) );
  AOI22_X1 U6957 ( .A1(n5924), .A2(n6112), .B1(n6102), .B2(n5898), .ZN(n5899)
         );
  OAI211_X1 U6958 ( .C1(n5901), .C2(n6145), .A(n5900), .B(n5899), .ZN(U2806)
         );
  AOI22_X1 U6959 ( .A1(EBX_REG_20__SCAN_IN), .A2(n2993), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6133), .ZN(n5910) );
  INV_X1 U6960 ( .A(n5902), .ZN(n5903) );
  AOI22_X1 U6961 ( .A1(n5927), .A2(n6112), .B1(n5903), .B2(n6102), .ZN(n5909)
         );
  NAND2_X1 U6962 ( .A1(n6079), .A2(n5904), .ZN(n5908) );
  OAI21_X1 U6963 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5906), .A(n5905), .ZN(n5907) );
  NAND4_X1 U6964 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(U2807)
         );
  INV_X1 U6965 ( .A(n6153), .ZN(n5912) );
  INV_X1 U6966 ( .A(DATAI_26_), .ZN(n5911) );
  OAI22_X1 U6967 ( .A1(n5913), .A2(n5917), .B1(n5912), .B2(n5911), .ZN(n5914)
         );
  INV_X1 U6968 ( .A(n5914), .ZN(n5916) );
  AOI22_X1 U6969 ( .A1(n6157), .A2(DATAI_10_), .B1(n6156), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U6970 ( .A1(n5916), .A2(n5915), .ZN(U2865) );
  INV_X1 U6971 ( .A(n5917), .ZN(n6154) );
  AOI22_X1 U6972 ( .A1(n5918), .A2(n6154), .B1(n6153), .B2(DATAI_25_), .ZN(
        n5920) );
  AOI22_X1 U6973 ( .A1(n6157), .A2(DATAI_9_), .B1(n6156), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U6974 ( .A1(n5920), .A2(n5919), .ZN(U2866) );
  AOI22_X1 U6975 ( .A1(n5921), .A2(n6154), .B1(n6153), .B2(DATAI_22_), .ZN(
        n5923) );
  AOI22_X1 U6976 ( .A1(n6157), .A2(DATAI_6_), .B1(n6156), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U6977 ( .A1(n5923), .A2(n5922), .ZN(U2869) );
  AOI22_X1 U6978 ( .A1(n5924), .A2(n6154), .B1(n6153), .B2(DATAI_21_), .ZN(
        n5926) );
  AOI22_X1 U6979 ( .A1(n6157), .A2(DATAI_5_), .B1(n6156), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U6980 ( .A1(n5926), .A2(n5925), .ZN(U2870) );
  AOI22_X1 U6981 ( .A1(n5927), .A2(n6154), .B1(n6153), .B2(DATAI_20_), .ZN(
        n5929) );
  AOI22_X1 U6982 ( .A1(n6157), .A2(DATAI_4_), .B1(n6156), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U6983 ( .A1(n5929), .A2(n5928), .ZN(U2871) );
  AOI22_X1 U6984 ( .A1(n6336), .A2(REIP_REG_18__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5932) );
  AOI22_X1 U6985 ( .A1(n5930), .A2(n6251), .B1(n6225), .B2(n6147), .ZN(n5931)
         );
  OAI211_X1 U6986 ( .C1(n6255), .C2(n6023), .A(n5932), .B(n5931), .ZN(U2968)
         );
  INV_X1 U6987 ( .A(n5933), .ZN(n5934) );
  NOR2_X1 U6988 ( .A1(n5935), .A2(n5934), .ZN(n5937) );
  XNOR2_X1 U6989 ( .A(n5937), .B(n5936), .ZN(n5954) );
  AOI22_X1 U6990 ( .A1(n6336), .A2(REIP_REG_17__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5940) );
  AOI22_X1 U6991 ( .A1(n6150), .A2(n6225), .B1(n6224), .B2(n5938), .ZN(n5939)
         );
  OAI211_X1 U6992 ( .C1(n5954), .C2(n6229), .A(n5940), .B(n5939), .ZN(U2969)
         );
  AOI22_X1 U6993 ( .A1(n6336), .A2(REIP_REG_13__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5948) );
  OR2_X1 U6994 ( .A1(n5942), .A2(n5941), .ZN(n5944) );
  NAND2_X1 U6995 ( .A1(n5944), .A2(n5943), .ZN(n5946) );
  XNOR2_X1 U6996 ( .A(n5946), .B(n5945), .ZN(n5986) );
  AOI22_X1 U6997 ( .A1(n5986), .A2(n6251), .B1(n6225), .B2(n6053), .ZN(n5947)
         );
  OAI211_X1 U6998 ( .C1(n6255), .C2(n6056), .A(n5948), .B(n5947), .ZN(U2973)
         );
  AOI22_X1 U6999 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5949), .B1(n6336), .B2(REIP_REG_17__SCAN_IN), .ZN(n5953) );
  AOI22_X1 U7000 ( .A1(n5951), .A2(n5936), .B1(n6338), .B2(n5950), .ZN(n5952)
         );
  OAI211_X1 U7001 ( .C1(n5954), .C2(n6342), .A(n5953), .B(n5952), .ZN(U3001)
         );
  OAI21_X1 U7002 ( .B1(n5956), .B2(n5955), .A(n6295), .ZN(n6266) );
  AOI21_X1 U7003 ( .B1(n5958), .B2(n5957), .A(n6266), .ZN(n5971) );
  NOR2_X1 U7004 ( .A1(n5958), .A2(n5984), .ZN(n5965) );
  OAI221_X1 U7005 ( .B1(n5970), .B2(n5964), .C1(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C2(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .A(n5965), .ZN(n5959) );
  INV_X1 U7006 ( .A(n5959), .ZN(n5962) );
  OAI22_X1 U7007 ( .A1(n5960), .A2(n6342), .B1(n6283), .B2(n6034), .ZN(n5961)
         );
  AOI211_X1 U7008 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6336), .A(n5962), .B(n5961), .ZN(n5963) );
  OAI21_X1 U7009 ( .B1(n5971), .B2(n5964), .A(n5963), .ZN(U3002) );
  AOI22_X1 U7010 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6336), .B1(n5965), .B2(
        n5970), .ZN(n5969) );
  AOI22_X1 U7011 ( .A1(n5967), .A2(n6324), .B1(n6338), .B2(n5966), .ZN(n5968)
         );
  OAI211_X1 U7012 ( .C1(n5971), .C2(n5970), .A(n5969), .B(n5968), .ZN(U3003)
         );
  NOR2_X1 U7013 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  AOI211_X1 U7014 ( .C1(n5975), .C2(n5978), .A(n5974), .B(n6266), .ZN(n5989)
         );
  OAI21_X1 U7015 ( .B1(n5977), .B2(n5976), .A(n4140), .ZN(n5983) );
  NOR3_X1 U7016 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5984), .A3(n5978), 
        .ZN(n5981) );
  OAI22_X1 U7017 ( .A1(n5979), .A2(n6342), .B1(n6283), .B2(n6037), .ZN(n5980)
         );
  AOI211_X1 U7018 ( .C1(REIP_REG_14__SCAN_IN), .C2(n6336), .A(n5981), .B(n5980), .ZN(n5982) );
  OAI221_X1 U7019 ( .B1(n5298), .B2(n5989), .C1(n5298), .C2(n5983), .A(n5982), 
        .ZN(U3004) );
  AOI22_X1 U7020 ( .A1(n6048), .A2(n6338), .B1(n6336), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5988) );
  INV_X1 U7021 ( .A(n5984), .ZN(n6265) );
  NOR2_X1 U7022 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6257), .ZN(n5985)
         );
  AOI22_X1 U7023 ( .A1(n5986), .A2(n6324), .B1(n6265), .B2(n5985), .ZN(n5987)
         );
  OAI211_X1 U7024 ( .C1(n5989), .C2(n4140), .A(n5988), .B(n5987), .ZN(U3005)
         );
  OR4_X1 U7025 ( .A1(n5990), .A2(n6115), .A3(n4194), .A4(n6579), .ZN(n5991) );
  OAI21_X1 U7026 ( .B1(n6576), .B2(n3902), .A(n5991), .ZN(U3455) );
  INV_X1 U7027 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6503) );
  NOR2_X1 U7028 ( .A1(n6503), .A2(STATE_REG_0__SCAN_IN), .ZN(n6535) );
  OAI21_X1 U7029 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6503), .A(
        STATE_REG_0__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U7030 ( .A1(ADS_N_REG_SCAN_IN), .A2(n5999), .ZN(n5992) );
  NOR2_X1 U7031 ( .A1(n6535), .A2(n5992), .ZN(U2789) );
  NAND2_X1 U7032 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5993), .ZN(n5997) );
  INV_X1 U7033 ( .A(n5994), .ZN(n5995) );
  OAI21_X1 U7034 ( .B1(n5995), .B2(n6488), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5996) );
  OAI21_X1 U7035 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5997), .A(n5996), .ZN(
        U2790) );
  NOR2_X1 U7036 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6000) );
  OAI21_X1 U7037 ( .B1(n6000), .B2(D_C_N_REG_SCAN_IN), .A(n6607), .ZN(n5998)
         );
  OAI21_X1 U7038 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6607), .A(n5998), .ZN(
        U2791) );
  NAND2_X1 U7039 ( .A1(n6607), .A2(n5999), .ZN(n6608) );
  INV_X1 U7040 ( .A(n6608), .ZN(n6567) );
  OAI21_X1 U7041 ( .B1(n6000), .B2(BS16_N), .A(n6567), .ZN(n6566) );
  OAI21_X1 U7042 ( .B1(n6567), .B2(n6593), .A(n6566), .ZN(U2792) );
  OAI21_X1 U7043 ( .B1(n6002), .B2(n6001), .A(n6229), .ZN(U2793) );
  NOR4_X1 U7044 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6012) );
  NOR4_X1 U7045 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6011) );
  AOI211_X1 U7046 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_18__SCAN_IN), .B(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6003) );
  INV_X1 U7047 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6736) );
  INV_X1 U7048 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6629) );
  NAND3_X1 U7049 ( .A1(n6003), .A2(n6736), .A3(n6629), .ZN(n6009) );
  NOR4_X1 U7050 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6007) );
  NOR4_X1 U7051 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6006) );
  NOR4_X1 U7052 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6005) );
  NOR4_X1 U7053 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6004) );
  NAND4_X1 U7054 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n6008)
         );
  NOR4_X1 U7055 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(n6009), .A4(n6008), .ZN(n6010) );
  NAND3_X1 U7056 ( .A1(n6012), .A2(n6011), .A3(n6010), .ZN(n6590) );
  INV_X1 U7057 ( .A(n6590), .ZN(n6587) );
  NAND2_X1 U7058 ( .A1(n6587), .A2(n6583), .ZN(n6586) );
  NOR3_X1 U7059 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6586), .ZN(n6014) );
  AOI21_X1 U7060 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6590), .A(n6014), .ZN(
        n6013) );
  OAI21_X1 U7061 ( .B1(n6589), .B2(n6590), .A(n6013), .ZN(U2794) );
  NAND2_X1 U7062 ( .A1(n6587), .A2(n6589), .ZN(n6581) );
  AOI21_X1 U7063 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n6590), .A(n6014), .ZN(
        n6015) );
  OAI21_X1 U7064 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6581), .A(n6015), .ZN(
        U2795) );
  AOI211_X1 U7065 ( .C1(n6133), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6016), 
        .B(n6107), .ZN(n6019) );
  AOI22_X1 U7066 ( .A1(EBX_REG_18__SCAN_IN), .A2(n2993), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6017), .ZN(n6018) );
  OAI211_X1 U7067 ( .C1(n6145), .C2(n6020), .A(n6019), .B(n6018), .ZN(n6021)
         );
  AOI21_X1 U7068 ( .B1(n6147), .B2(n6112), .A(n6021), .ZN(n6022) );
  OAI21_X1 U7069 ( .B1(n6023), .B2(n6135), .A(n6022), .ZN(U2809) );
  INV_X1 U7070 ( .A(n6024), .ZN(n6027) );
  NOR2_X1 U7071 ( .A1(n6036), .A2(n6025), .ZN(n6026) );
  MUX2_X1 U7072 ( .A(n6027), .B(n6026), .S(REIP_REG_16__SCAN_IN), .Z(n6028) );
  OAI21_X1 U7073 ( .B1(n6029), .B2(n6138), .A(n6028), .ZN(n6030) );
  AOI211_X1 U7074 ( .C1(n6133), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6107), 
        .B(n6030), .ZN(n6033) );
  AOI22_X1 U7075 ( .A1(n6155), .A2(n6112), .B1(n6102), .B2(n6031), .ZN(n6032)
         );
  OAI211_X1 U7076 ( .C1(n6145), .C2(n6034), .A(n6033), .B(n6032), .ZN(U2811)
         );
  AND2_X1 U7077 ( .A1(n6120), .A2(n6035), .ZN(n6052) );
  AOI21_X1 U7078 ( .B1(REIP_REG_13__SCAN_IN), .B2(n6052), .A(
        REIP_REG_14__SCAN_IN), .ZN(n6046) );
  INV_X1 U7079 ( .A(n6036), .ZN(n6045) );
  OAI22_X1 U7080 ( .A1(n6038), .A2(n6124), .B1(n6145), .B2(n6037), .ZN(n6039)
         );
  AOI211_X1 U7081 ( .C1(n2993), .C2(EBX_REG_14__SCAN_IN), .A(n6107), .B(n6039), 
        .ZN(n6044) );
  INV_X1 U7082 ( .A(n6040), .ZN(n6042) );
  AOI22_X1 U7083 ( .A1(n6042), .A2(n6112), .B1(n6102), .B2(n6041), .ZN(n6043)
         );
  OAI211_X1 U7084 ( .C1(n6046), .C2(n6045), .A(n6044), .B(n6043), .ZN(U2813)
         );
  INV_X1 U7085 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U7086 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6083), .A(n6047), .ZN(n6051) );
  AOI22_X1 U7087 ( .A1(EBX_REG_13__SCAN_IN), .A2(n2993), .B1(n6079), .B2(n6048), .ZN(n6049) );
  OAI211_X1 U7088 ( .C1(n6124), .C2(n3500), .A(n6049), .B(n6122), .ZN(n6050)
         );
  AOI221_X1 U7089 ( .B1(n6052), .B2(n6533), .C1(n6051), .C2(
        REIP_REG_13__SCAN_IN), .A(n6050), .ZN(n6055) );
  NAND2_X1 U7090 ( .A1(n6053), .A2(n6112), .ZN(n6054) );
  OAI211_X1 U7091 ( .C1(n6135), .C2(n6056), .A(n6055), .B(n6054), .ZN(U2814)
         );
  INV_X1 U7092 ( .A(n6057), .ZN(n6264) );
  AOI22_X1 U7093 ( .A1(EBX_REG_11__SCAN_IN), .A2(n2993), .B1(n6079), .B2(n6264), .ZN(n6064) );
  AOI22_X1 U7094 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6133), .B1(n6132), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6063) );
  AOI221_X1 U7095 ( .B1(REIP_REG_11__SCAN_IN), .B2(n6059), .C1(n6058), .C2(
        n6059), .A(n6107), .ZN(n6062) );
  INV_X1 U7096 ( .A(n6060), .ZN(n6226) );
  AOI22_X1 U7097 ( .A1(n6226), .A2(n6112), .B1(n6102), .B2(n6223), .ZN(n6061)
         );
  NAND4_X1 U7098 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(U2816)
         );
  INV_X1 U7099 ( .A(n6065), .ZN(n6080) );
  OR2_X1 U7100 ( .A1(n6083), .A2(n6080), .ZN(n6096) );
  NAND2_X1 U7101 ( .A1(n6066), .A2(n6096), .ZN(n6092) );
  AOI22_X1 U7102 ( .A1(n6079), .A2(n6272), .B1(REIP_REG_10__SCAN_IN), .B2(
        n6092), .ZN(n6076) );
  OAI211_X1 U7103 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n6067), .B(n6080), .ZN(n6069) );
  NAND2_X1 U7104 ( .A1(n6133), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6068)
         );
  OAI211_X1 U7105 ( .C1(n6083), .C2(n6069), .A(n6122), .B(n6068), .ZN(n6070)
         );
  INV_X1 U7106 ( .A(n6070), .ZN(n6071) );
  OAI21_X1 U7107 ( .B1(n6072), .B2(n6099), .A(n6071), .ZN(n6073) );
  AOI21_X1 U7108 ( .B1(n6074), .B2(n6102), .A(n6073), .ZN(n6075) );
  OAI211_X1 U7109 ( .C1(n6077), .C2(n6138), .A(n6076), .B(n6075), .ZN(U2817)
         );
  INV_X1 U7110 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6091) );
  AOI22_X1 U7111 ( .A1(n6079), .A2(n6078), .B1(REIP_REG_9__SCAN_IN), .B2(n6092), .ZN(n6090) );
  NAND2_X1 U7112 ( .A1(n6080), .A2(n5162), .ZN(n6082) );
  NAND2_X1 U7113 ( .A1(n6133), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6081)
         );
  OAI211_X1 U7114 ( .C1(n6083), .C2(n6082), .A(n6122), .B(n6081), .ZN(n6084)
         );
  AOI21_X1 U7115 ( .B1(n6085), .B2(n6112), .A(n6084), .ZN(n6086) );
  INV_X1 U7116 ( .A(n6086), .ZN(n6087) );
  AOI21_X1 U7117 ( .B1(n6088), .B2(n6102), .A(n6087), .ZN(n6089) );
  OAI211_X1 U7118 ( .C1(n6091), .C2(n6138), .A(n6090), .B(n6089), .ZN(U2818)
         );
  AOI22_X1 U7119 ( .A1(EBX_REG_8__SCAN_IN), .A2(n2993), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6092), .ZN(n6105) );
  INV_X1 U7120 ( .A(n6093), .ZN(n6095) );
  NAND2_X1 U7121 ( .A1(n6133), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6094)
         );
  OAI211_X1 U7122 ( .C1(n6096), .C2(n6095), .A(n6122), .B(n6094), .ZN(n6097)
         );
  INV_X1 U7123 ( .A(n6097), .ZN(n6098) );
  OAI21_X1 U7124 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n6101) );
  AOI21_X1 U7125 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(n6104) );
  OAI211_X1 U7126 ( .C1(n6145), .C2(n6282), .A(n6105), .B(n6104), .ZN(U2819)
         );
  AOI211_X1 U7127 ( .C1(n6133), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6107), 
        .B(n6106), .ZN(n6108) );
  OAI21_X1 U7128 ( .B1(n6145), .B2(n6109), .A(n6108), .ZN(n6110) );
  AOI21_X1 U7129 ( .B1(EBX_REG_6__SCAN_IN), .B2(n2993), .A(n6110), .ZN(n6114)
         );
  AOI22_X1 U7130 ( .A1(n6231), .A2(n6112), .B1(REIP_REG_6__SCAN_IN), .B2(n6111), .ZN(n6113) );
  OAI211_X1 U7131 ( .C1(n6235), .C2(n6135), .A(n6114), .B(n6113), .ZN(U2821)
         );
  INV_X1 U7132 ( .A(n6136), .ZN(n6117) );
  INV_X1 U7133 ( .A(n6115), .ZN(n6116) );
  AOI22_X1 U7134 ( .A1(n6118), .A2(REIP_REG_4__SCAN_IN), .B1(n6117), .B2(n6116), .ZN(n6131) );
  INV_X1 U7135 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6123) );
  INV_X1 U7136 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6519) );
  NAND3_X1 U7137 ( .A1(n6120), .A2(n6119), .A3(n6519), .ZN(n6121) );
  OAI211_X1 U7138 ( .C1(n6124), .C2(n6123), .A(n6122), .B(n6121), .ZN(n6128)
         );
  OAI22_X1 U7139 ( .A1(n6126), .A2(n6125), .B1(n6244), .B2(n6135), .ZN(n6127)
         );
  AOI211_X1 U7140 ( .C1(EBX_REG_4__SCAN_IN), .C2(n2993), .A(n6128), .B(n6127), 
        .ZN(n6130) );
  OAI211_X1 U7141 ( .C1(n6145), .C2(n6313), .A(n6131), .B(n6130), .ZN(U2823)
         );
  AOI22_X1 U7142 ( .A1(n6133), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6132), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6134) );
  OAI21_X1 U7143 ( .B1(n6135), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6134), 
        .ZN(n6140) );
  OAI22_X1 U7144 ( .A1(n6138), .A2(n3939), .B1(n6137), .B2(n6136), .ZN(n6139)
         );
  AOI211_X1 U7145 ( .C1(n6142), .C2(n6141), .A(n6140), .B(n6139), .ZN(n6144)
         );
  OAI211_X1 U7146 ( .C1(n6146), .C2(n6145), .A(n6144), .B(n6143), .ZN(U2826)
         );
  AOI22_X1 U7147 ( .A1(n6147), .A2(n6154), .B1(n6153), .B2(DATAI_18_), .ZN(
        n6149) );
  AOI22_X1 U7148 ( .A1(n6157), .A2(DATAI_2_), .B1(n6156), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7149 ( .A1(n6149), .A2(n6148), .ZN(U2873) );
  AOI22_X1 U7150 ( .A1(n6150), .A2(n6154), .B1(n6153), .B2(DATAI_17_), .ZN(
        n6152) );
  AOI22_X1 U7151 ( .A1(n6157), .A2(DATAI_1_), .B1(n6156), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7152 ( .A1(n6152), .A2(n6151), .ZN(U2874) );
  AOI22_X1 U7153 ( .A1(n6155), .A2(n6154), .B1(n6153), .B2(DATAI_16_), .ZN(
        n6159) );
  AOI22_X1 U7154 ( .A1(n6157), .A2(DATAI_0_), .B1(n6156), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7155 ( .A1(n6159), .A2(n6158), .ZN(U2875) );
  INV_X1 U7156 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6218) );
  AOI22_X1 U7157 ( .A1(n6604), .A2(LWORD_REG_15__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6161) );
  OAI21_X1 U7158 ( .B1(n6218), .B2(n6187), .A(n6161), .ZN(U2908) );
  INV_X1 U7159 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6163) );
  AOI22_X1 U7160 ( .A1(n6604), .A2(LWORD_REG_14__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U7161 ( .B1(n6163), .B2(n6187), .A(n6162), .ZN(U2909) );
  INV_X1 U7162 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6165) );
  AOI22_X1 U7163 ( .A1(n6604), .A2(LWORD_REG_13__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6164) );
  OAI21_X1 U7164 ( .B1(n6165), .B2(n6187), .A(n6164), .ZN(U2910) );
  INV_X1 U7165 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7166 ( .A1(n6604), .A2(LWORD_REG_12__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6166) );
  OAI21_X1 U7167 ( .B1(n6612), .B2(n6187), .A(n6166), .ZN(U2911) );
  INV_X1 U7168 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6168) );
  AOI22_X1 U7169 ( .A1(n6604), .A2(LWORD_REG_11__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6167) );
  OAI21_X1 U7170 ( .B1(n6168), .B2(n6187), .A(n6167), .ZN(U2912) );
  INV_X1 U7171 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U7172 ( .A1(n6604), .A2(LWORD_REG_10__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6169) );
  OAI21_X1 U7173 ( .B1(n6746), .B2(n6187), .A(n6169), .ZN(U2913) );
  INV_X1 U7174 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6171) );
  AOI22_X1 U7175 ( .A1(n6604), .A2(LWORD_REG_9__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6170) );
  OAI21_X1 U7176 ( .B1(n6171), .B2(n6187), .A(n6170), .ZN(U2914) );
  INV_X1 U7177 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6173) );
  AOI22_X1 U7178 ( .A1(n6604), .A2(LWORD_REG_8__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6172) );
  OAI21_X1 U7179 ( .B1(n6173), .B2(n6187), .A(n6172), .ZN(U2915) );
  AOI22_X1 U7180 ( .A1(n6604), .A2(LWORD_REG_7__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U7181 ( .B1(n3416), .B2(n6187), .A(n6174), .ZN(U2916) );
  AOI22_X1 U7182 ( .A1(n6604), .A2(LWORD_REG_6__SCAN_IN), .B1(n6175), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7183 ( .B1(n4849), .B2(n6187), .A(n6176), .ZN(U2917) );
  AOI22_X1 U7184 ( .A1(n6604), .A2(LWORD_REG_5__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6177) );
  OAI21_X1 U7185 ( .B1(n4861), .B2(n6187), .A(n6177), .ZN(U2918) );
  AOI22_X1 U7186 ( .A1(n6604), .A2(LWORD_REG_4__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6178) );
  OAI21_X1 U7187 ( .B1(n4866), .B2(n6187), .A(n6178), .ZN(U2919) );
  AOI22_X1 U7188 ( .A1(n6604), .A2(LWORD_REG_3__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6179) );
  OAI21_X1 U7189 ( .B1(n6180), .B2(n6187), .A(n6179), .ZN(U2920) );
  AOI22_X1 U7190 ( .A1(n6604), .A2(LWORD_REG_2__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6181) );
  OAI21_X1 U7191 ( .B1(n6752), .B2(n6187), .A(n6181), .ZN(U2921) );
  AOI22_X1 U7192 ( .A1(n6604), .A2(LWORD_REG_1__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6182) );
  OAI21_X1 U7193 ( .B1(n6183), .B2(n6187), .A(n6182), .ZN(U2922) );
  AOI22_X1 U7194 ( .A1(n6604), .A2(LWORD_REG_0__SCAN_IN), .B1(n6184), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U7195 ( .B1(n4319), .B2(n6187), .A(n6186), .ZN(U2923) );
  AOI22_X1 U7196 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6211), .B1(n6210), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7197 ( .A1(n6214), .A2(DATAI_8_), .ZN(n6200) );
  NAND2_X1 U7198 ( .A1(n6188), .A2(n6200), .ZN(U2932) );
  INV_X1 U7199 ( .A(DATAI_10_), .ZN(n6189) );
  NOR2_X1 U7200 ( .A1(n6196), .A2(n6189), .ZN(n6202) );
  AOI21_X1 U7201 ( .B1(n6210), .B2(UWORD_REG_10__SCAN_IN), .A(n6202), .ZN(
        n6190) );
  OAI21_X1 U7202 ( .B1(n6191), .B2(n6217), .A(n6190), .ZN(U2934) );
  NAND2_X1 U7203 ( .A1(n6214), .A2(DATAI_11_), .ZN(n6204) );
  INV_X1 U7204 ( .A(n6204), .ZN(n6192) );
  AOI21_X1 U7205 ( .B1(n6210), .B2(UWORD_REG_11__SCAN_IN), .A(n6192), .ZN(
        n6193) );
  OAI21_X1 U7206 ( .B1(n6194), .B2(n6217), .A(n6193), .ZN(U2935) );
  INV_X1 U7207 ( .A(DATAI_12_), .ZN(n6195) );
  NOR2_X1 U7208 ( .A1(n6196), .A2(n6195), .ZN(n6206) );
  AOI21_X1 U7209 ( .B1(n6210), .B2(UWORD_REG_12__SCAN_IN), .A(n6206), .ZN(
        n6197) );
  OAI21_X1 U7210 ( .B1(n6626), .B2(n6217), .A(n6197), .ZN(U2936) );
  AOI22_X1 U7211 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6211), .B1(n6215), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7212 ( .A1(n6214), .A2(DATAI_13_), .ZN(n6208) );
  NAND2_X1 U7213 ( .A1(n6198), .A2(n6208), .ZN(U2937) );
  AOI22_X1 U7214 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6211), .B1(n6210), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7215 ( .A1(n6214), .A2(DATAI_14_), .ZN(n6212) );
  NAND2_X1 U7216 ( .A1(n6199), .A2(n6212), .ZN(U2938) );
  AOI22_X1 U7217 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6211), .B1(n6210), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7218 ( .A1(n6201), .A2(n6200), .ZN(U2947) );
  AOI21_X1 U7219 ( .B1(n6210), .B2(LWORD_REG_10__SCAN_IN), .A(n6202), .ZN(
        n6203) );
  OAI21_X1 U7220 ( .B1(n6746), .B2(n6217), .A(n6203), .ZN(U2949) );
  AOI22_X1 U7221 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6211), .B1(n6210), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7222 ( .A1(n6205), .A2(n6204), .ZN(U2950) );
  AOI21_X1 U7223 ( .B1(n6210), .B2(LWORD_REG_12__SCAN_IN), .A(n6206), .ZN(
        n6207) );
  OAI21_X1 U7224 ( .B1(n6612), .B2(n6217), .A(n6207), .ZN(U2951) );
  AOI22_X1 U7225 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6211), .B1(n6210), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7226 ( .A1(n6209), .A2(n6208), .ZN(U2952) );
  AOI22_X1 U7227 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6211), .B1(n6210), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7228 ( .A1(n6213), .A2(n6212), .ZN(U2953) );
  AOI22_X1 U7229 ( .A1(n6215), .A2(LWORD_REG_15__SCAN_IN), .B1(n6214), .B2(
        DATAI_15_), .ZN(n6216) );
  OAI21_X1 U7230 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(U2954) );
  NAND2_X1 U7231 ( .A1(n6220), .A2(n6219), .ZN(n6222) );
  XNOR2_X1 U7232 ( .A(n5720), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6221)
         );
  XNOR2_X1 U7233 ( .A(n6222), .B(n6221), .ZN(n6269) );
  AOI22_X1 U7234 ( .A1(n6336), .A2(REIP_REG_11__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6228) );
  AOI22_X1 U7235 ( .A1(n6226), .A2(n6225), .B1(n6224), .B2(n6223), .ZN(n6227)
         );
  OAI211_X1 U7236 ( .C1(n6269), .C2(n6229), .A(n6228), .B(n6227), .ZN(U2975)
         );
  AOI22_X1 U7237 ( .A1(n6336), .A2(REIP_REG_6__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6234) );
  INV_X1 U7238 ( .A(n6230), .ZN(n6232) );
  AOI22_X1 U7239 ( .A1(n6232), .A2(n6251), .B1(n6225), .B2(n6231), .ZN(n6233)
         );
  OAI211_X1 U7240 ( .C1(n6255), .C2(n6235), .A(n6234), .B(n6233), .ZN(U2980)
         );
  AOI22_X1 U7241 ( .A1(n6336), .A2(REIP_REG_4__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6243) );
  OR2_X1 U7242 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  AND2_X1 U7243 ( .A1(n6240), .A2(n6239), .ZN(n6315) );
  AOI22_X1 U7244 ( .A1(n6315), .A2(n6251), .B1(n6241), .B2(n6225), .ZN(n6242)
         );
  OAI211_X1 U7245 ( .C1(n6255), .C2(n6244), .A(n6243), .B(n6242), .ZN(U2982)
         );
  AOI22_X1 U7246 ( .A1(n6336), .A2(REIP_REG_2__SCAN_IN), .B1(n6236), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6253) );
  XNOR2_X1 U7247 ( .A(n6245), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6247)
         );
  XNOR2_X1 U7248 ( .A(n6247), .B(n6246), .ZN(n6341) );
  INV_X1 U7249 ( .A(n6341), .ZN(n6250) );
  INV_X1 U7250 ( .A(n6248), .ZN(n6249) );
  AOI22_X1 U7251 ( .A1(n6251), .A2(n6250), .B1(n6249), .B2(n6225), .ZN(n6252)
         );
  OAI211_X1 U7252 ( .C1(n6255), .C2(n6254), .A(n6253), .B(n6252), .ZN(U2984)
         );
  AOI221_X1 U7253 ( .B1(n6333), .B2(n6257), .C1(n6256), .C2(n6257), .A(n6266), 
        .ZN(n6263) );
  AOI21_X1 U7254 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6265), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6262) );
  AOI22_X1 U7255 ( .A1(n6259), .A2(n6324), .B1(n6338), .B2(n6258), .ZN(n6261)
         );
  NAND2_X1 U7256 ( .A1(n6336), .A2(REIP_REG_12__SCAN_IN), .ZN(n6260) );
  OAI211_X1 U7257 ( .C1(n6263), .C2(n6262), .A(n6261), .B(n6260), .ZN(U3006)
         );
  AOI22_X1 U7258 ( .A1(n6338), .A2(n6264), .B1(n6336), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6268) );
  AOI22_X1 U7259 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6266), .B1(n6265), .B2(n4134), .ZN(n6267) );
  OAI211_X1 U7260 ( .C1(n6269), .C2(n6342), .A(n6268), .B(n6267), .ZN(U3007)
         );
  INV_X1 U7261 ( .A(n6270), .ZN(n6271) );
  AOI21_X1 U7262 ( .B1(n6338), .B2(n6272), .A(n6271), .ZN(n6279) );
  AOI22_X1 U7263 ( .A1(n6274), .A2(n6324), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6273), .ZN(n6278) );
  OAI211_X1 U7264 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6276), .B(n6275), .ZN(n6277) );
  NAND3_X1 U7265 ( .A1(n6279), .A2(n6278), .A3(n6277), .ZN(U3008) );
  INV_X1 U7266 ( .A(n6280), .ZN(n6288) );
  OAI22_X1 U7267 ( .A1(n6283), .A2(n6282), .B1(n5404), .B2(n6281), .ZN(n6287)
         );
  AOI211_X1 U7268 ( .C1(n6285), .C2(n6290), .A(n6284), .B(n6300), .ZN(n6286)
         );
  AOI211_X1 U7269 ( .C1(n6288), .C2(n6324), .A(n6287), .B(n6286), .ZN(n6289)
         );
  OAI21_X1 U7270 ( .B1(n6295), .B2(n6290), .A(n6289), .ZN(U3010) );
  INV_X1 U7271 ( .A(n6291), .ZN(n6292) );
  AOI21_X1 U7272 ( .B1(n6338), .B2(n6293), .A(n6292), .ZN(n6299) );
  INV_X1 U7273 ( .A(n6294), .ZN(n6297) );
  INV_X1 U7274 ( .A(n6295), .ZN(n6296) );
  AOI22_X1 U7275 ( .A1(n6297), .A2(n6324), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6296), .ZN(n6298) );
  OAI211_X1 U7276 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6300), .A(n6299), 
        .B(n6298), .ZN(U3011) );
  AOI21_X1 U7277 ( .B1(n6333), .B2(n6301), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6311) );
  INV_X1 U7278 ( .A(n6302), .ZN(n6303) );
  AOI21_X1 U7279 ( .B1(n6338), .B2(n6304), .A(n6303), .ZN(n6310) );
  NOR3_X1 U7280 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6316), .A3(n6305), 
        .ZN(n6308) );
  NOR2_X1 U7281 ( .A1(n6306), .A2(n6342), .ZN(n6307) );
  NOR2_X1 U7282 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  OAI211_X1 U7283 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n6309), .ZN(U3013)
         );
  AOI21_X1 U7284 ( .B1(n6333), .B2(n6335), .A(n6332), .ZN(n6330) );
  INV_X1 U7285 ( .A(n6313), .ZN(n6314) );
  AOI22_X1 U7286 ( .A1(n6338), .A2(n6314), .B1(n6336), .B2(REIP_REG_4__SCAN_IN), .ZN(n6319) );
  AOI211_X1 U7287 ( .C1(n6329), .C2(n6320), .A(n6323), .B(n6335), .ZN(n6317)
         );
  AOI22_X1 U7288 ( .A1(n6317), .A2(n6316), .B1(n6324), .B2(n6315), .ZN(n6318)
         );
  OAI211_X1 U7289 ( .C1(n6330), .C2(n6320), .A(n6319), .B(n6318), .ZN(U3014)
         );
  AOI21_X1 U7290 ( .B1(n6338), .B2(n6322), .A(n6321), .ZN(n6328) );
  NOR2_X1 U7291 ( .A1(n6335), .A2(n6323), .ZN(n6326) );
  AOI22_X1 U7292 ( .A1(n6326), .A2(n6329), .B1(n6325), .B2(n6324), .ZN(n6327)
         );
  OAI211_X1 U7293 ( .C1(n6330), .C2(n6329), .A(n6328), .B(n6327), .ZN(U3015)
         );
  NAND2_X1 U7294 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6331), .ZN(n6347)
         );
  INV_X1 U7295 ( .A(n6332), .ZN(n6345) );
  OAI221_X1 U7296 ( .B1(n6335), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .C1(n6335), .C2(n6334), .A(n6333), .ZN(n6340) );
  AOI22_X1 U7297 ( .A1(n6338), .A2(n6337), .B1(n6336), .B2(REIP_REG_2__SCAN_IN), .ZN(n6339) );
  OAI211_X1 U7298 ( .C1(n6342), .C2(n6341), .A(n6340), .B(n6339), .ZN(n6343)
         );
  INV_X1 U7299 ( .A(n6343), .ZN(n6344) );
  OAI221_X1 U7300 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6347), .C1(n6346), .C2(n6345), .A(n6344), .ZN(U3016) );
  NOR2_X1 U7301 ( .A1(n6614), .A2(n6348), .ZN(U3019) );
  NOR2_X1 U7302 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6349), .ZN(n6394)
         );
  NAND3_X1 U7303 ( .A1(n6351), .A2(n6350), .A3(n6466), .ZN(n6352) );
  OAI21_X1 U7304 ( .B1(n6354), .B2(n6353), .A(n6352), .ZN(n6393) );
  AOI22_X1 U7305 ( .A1(n6356), .A2(n6394), .B1(n6355), .B2(n6393), .ZN(n6365)
         );
  INV_X1 U7306 ( .A(n6410), .ZN(n6357) );
  OAI21_X1 U7307 ( .B1(n3020), .B2(n6357), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6360) );
  AOI211_X1 U7308 ( .C1(n6361), .C2(n6360), .A(n6359), .B(n6358), .ZN(n6362)
         );
  OAI211_X1 U7309 ( .C1(n6394), .C2(n3174), .A(n6362), .B(n6466), .ZN(n6396)
         );
  AOI22_X1 U7310 ( .A1(n6396), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6363), 
        .B2(n3020), .ZN(n6364) );
  OAI211_X1 U7311 ( .C1(n6366), .C2(n6410), .A(n6365), .B(n6364), .ZN(U3068)
         );
  AOI22_X1 U7312 ( .A1(n6412), .A2(n6394), .B1(n6413), .B2(n6393), .ZN(n6369)
         );
  AOI22_X1 U7313 ( .A1(n6396), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6367), 
        .B2(n3020), .ZN(n6368) );
  OAI211_X1 U7314 ( .C1(n6370), .C2(n6410), .A(n6369), .B(n6368), .ZN(U3069)
         );
  AOI22_X1 U7315 ( .A1(n6418), .A2(n6394), .B1(n6419), .B2(n6393), .ZN(n6373)
         );
  AOI22_X1 U7316 ( .A1(n6396), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6371), 
        .B2(n3020), .ZN(n6372) );
  OAI211_X1 U7317 ( .C1(n6374), .C2(n6410), .A(n6373), .B(n6372), .ZN(U3070)
         );
  AOI22_X1 U7318 ( .A1(n6424), .A2(n6394), .B1(n6425), .B2(n6393), .ZN(n6377)
         );
  AOI22_X1 U7319 ( .A1(n6396), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6375), 
        .B2(n3020), .ZN(n6376) );
  OAI211_X1 U7320 ( .C1(n6378), .C2(n6410), .A(n6377), .B(n6376), .ZN(U3071)
         );
  AOI22_X1 U7321 ( .A1(n6430), .A2(n6394), .B1(n6431), .B2(n6393), .ZN(n6381)
         );
  AOI22_X1 U7322 ( .A1(n6396), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6379), 
        .B2(n3020), .ZN(n6380) );
  OAI211_X1 U7323 ( .C1(n6382), .C2(n6410), .A(n6381), .B(n6380), .ZN(U3072)
         );
  AOI22_X1 U7324 ( .A1(n6384), .A2(n6394), .B1(n6383), .B2(n6393), .ZN(n6387)
         );
  AOI22_X1 U7325 ( .A1(n6396), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6385), 
        .B2(n3020), .ZN(n6386) );
  OAI211_X1 U7326 ( .C1(n6388), .C2(n6410), .A(n6387), .B(n6386), .ZN(U3073)
         );
  AOI22_X1 U7327 ( .A1(n6436), .A2(n6394), .B1(n6437), .B2(n6393), .ZN(n6391)
         );
  AOI22_X1 U7328 ( .A1(n6396), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6389), 
        .B2(n3020), .ZN(n6390) );
  OAI211_X1 U7329 ( .C1(n6392), .C2(n6410), .A(n6391), .B(n6390), .ZN(U3074)
         );
  AOI22_X1 U7330 ( .A1(n6444), .A2(n6394), .B1(n6446), .B2(n6393), .ZN(n6398)
         );
  AOI22_X1 U7331 ( .A1(n6396), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6395), 
        .B2(n3020), .ZN(n6397) );
  OAI211_X1 U7332 ( .C1(n6399), .C2(n6410), .A(n6398), .B(n6397), .ZN(U3075)
         );
  AOI22_X1 U7333 ( .A1(n6418), .A2(n6405), .B1(n6417), .B2(n6404), .ZN(n6401)
         );
  AOI22_X1 U7334 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6407), .B1(n6419), 
        .B2(n6406), .ZN(n6400) );
  OAI211_X1 U7335 ( .C1(n6422), .C2(n6410), .A(n6401), .B(n6400), .ZN(U3078)
         );
  AOI22_X1 U7336 ( .A1(n6430), .A2(n6405), .B1(n6429), .B2(n6404), .ZN(n6403)
         );
  AOI22_X1 U7337 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6407), .B1(n6431), 
        .B2(n6406), .ZN(n6402) );
  OAI211_X1 U7338 ( .C1(n6434), .C2(n6410), .A(n6403), .B(n6402), .ZN(U3080)
         );
  AOI22_X1 U7339 ( .A1(n6436), .A2(n6405), .B1(n6435), .B2(n6404), .ZN(n6409)
         );
  AOI22_X1 U7340 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6407), .B1(n6437), 
        .B2(n6406), .ZN(n6408) );
  OAI211_X1 U7341 ( .C1(n6440), .C2(n6410), .A(n6409), .B(n6408), .ZN(U3082)
         );
  AOI22_X1 U7342 ( .A1(n6412), .A2(n6443), .B1(n6411), .B2(n6441), .ZN(n6415)
         );
  AOI22_X1 U7343 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6447), .B1(n6413), 
        .B2(n6445), .ZN(n6414) );
  OAI211_X1 U7344 ( .C1(n6416), .C2(n6450), .A(n6415), .B(n6414), .ZN(U3109)
         );
  AOI22_X1 U7345 ( .A1(n6418), .A2(n6443), .B1(n6417), .B2(n6441), .ZN(n6421)
         );
  AOI22_X1 U7346 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6447), .B1(n6419), 
        .B2(n6445), .ZN(n6420) );
  OAI211_X1 U7347 ( .C1(n6422), .C2(n6450), .A(n6421), .B(n6420), .ZN(U3110)
         );
  AOI22_X1 U7348 ( .A1(n6424), .A2(n6443), .B1(n6423), .B2(n6441), .ZN(n6427)
         );
  AOI22_X1 U7349 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6447), .B1(n6425), 
        .B2(n6445), .ZN(n6426) );
  OAI211_X1 U7350 ( .C1(n6428), .C2(n6450), .A(n6427), .B(n6426), .ZN(U3111)
         );
  AOI22_X1 U7351 ( .A1(n6430), .A2(n6443), .B1(n6429), .B2(n6441), .ZN(n6433)
         );
  AOI22_X1 U7352 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6447), .B1(n6431), 
        .B2(n6445), .ZN(n6432) );
  OAI211_X1 U7353 ( .C1(n6434), .C2(n6450), .A(n6433), .B(n6432), .ZN(U3112)
         );
  AOI22_X1 U7354 ( .A1(n6436), .A2(n6443), .B1(n6435), .B2(n6441), .ZN(n6439)
         );
  AOI22_X1 U7355 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6447), .B1(n6437), 
        .B2(n6445), .ZN(n6438) );
  OAI211_X1 U7356 ( .C1(n6440), .C2(n6450), .A(n6439), .B(n6438), .ZN(U3114)
         );
  AOI22_X1 U7357 ( .A1(n6444), .A2(n6443), .B1(n6442), .B2(n6441), .ZN(n6449)
         );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6447), .B1(n6446), 
        .B2(n6445), .ZN(n6448) );
  OAI211_X1 U7359 ( .C1(n6451), .C2(n6450), .A(n6449), .B(n6448), .ZN(U3115)
         );
  OAI22_X1 U7360 ( .A1(n4328), .A2(n6453), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6452), .ZN(n6575) );
  NAND2_X1 U7361 ( .A1(n6454), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6580) );
  INV_X1 U7362 ( .A(n6580), .ZN(n6456) );
  OR3_X1 U7363 ( .A1(n6575), .A2(n6456), .A3(n6455), .ZN(n6462) );
  AOI22_X1 U7364 ( .A1(n6458), .A2(n6457), .B1(n6461), .B2(n6462), .ZN(n6459)
         );
  INV_X1 U7365 ( .A(n6459), .ZN(n6460) );
  OAI21_X1 U7366 ( .B1(n6462), .B2(n6461), .A(n6460), .ZN(n6463) );
  AOI222_X1 U7367 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6464), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6463), .C1(n6464), .C2(n6463), 
        .ZN(n6465) );
  AOI222_X1 U7368 ( .A1(n6467), .A2(n6466), .B1(n6467), .B2(n6465), .C1(n6466), 
        .C2(n6465), .ZN(n6475) );
  NOR2_X1 U7369 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6468) );
  NOR2_X1 U7370 ( .A1(n6469), .A2(n6468), .ZN(n6471) );
  NOR4_X1 U7371 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6474)
         );
  OAI21_X1 U7372 ( .B1(n6475), .B2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6474), 
        .ZN(n6477) );
  INV_X1 U7373 ( .A(n6477), .ZN(n6486) );
  OAI22_X1 U7374 ( .A1(n6477), .A2(n6488), .B1(n6603), .B2(n6476), .ZN(n6478)
         );
  OAI21_X1 U7375 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n6570) );
  OAI21_X1 U7376 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6603), .A(n6570), .ZN(
        n6487) );
  AOI221_X1 U7377 ( .B1(n6482), .B2(STATE2_REG_0__SCAN_IN), .C1(n6487), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6481), .ZN(n6485) );
  OAI211_X1 U7378 ( .C1(n6598), .C2(n6483), .A(n6599), .B(n6570), .ZN(n6484)
         );
  OAI211_X1 U7379 ( .C1(n6486), .C2(n6488), .A(n6485), .B(n6484), .ZN(U3148)
         );
  NOR2_X1 U7380 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6496) );
  NAND2_X1 U7381 ( .A1(n6487), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6493) );
  OAI21_X1 U7382 ( .B1(READY_N), .B2(n6489), .A(n6488), .ZN(n6491) );
  AOI21_X1 U7383 ( .B1(n6570), .B2(n6491), .A(n6490), .ZN(n6492) );
  OAI21_X1 U7384 ( .B1(n6496), .B2(n6493), .A(n6492), .ZN(U3149) );
  OAI211_X1 U7385 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6603), .A(n6568), .B(
        n6598), .ZN(n6495) );
  OAI21_X1 U7386 ( .B1(n6496), .B2(n6495), .A(n6494), .ZN(U3150) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6608), .ZN(U3151) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6608), .ZN(U3152) );
  NOR2_X1 U7389 ( .A1(n6567), .A2(n6629), .ZN(U3153) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6608), .ZN(U3154) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6608), .ZN(U3155) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6608), .ZN(U3156) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6608), .ZN(U3157) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6608), .ZN(U3158) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6608), .ZN(U3159) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6608), .ZN(U3160) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6608), .ZN(U3161) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6608), .ZN(U3162) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6608), .ZN(U3163) );
  INV_X1 U7400 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6742) );
  NOR2_X1 U7401 ( .A1(n6567), .A2(n6742), .ZN(U3164) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6608), .ZN(U3166) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6608), .ZN(U3167) );
  NOR2_X1 U7404 ( .A1(n6567), .A2(n6736), .ZN(U3168) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6608), .ZN(U3169) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6608), .ZN(U3170) );
  AND2_X1 U7407 ( .A1(n6608), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6608), .ZN(U3172) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6608), .ZN(U3173) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6608), .ZN(U3174) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6608), .ZN(U3175) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6608), .ZN(U3176) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6608), .ZN(U3177) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6608), .ZN(U3178) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6608), .ZN(U3179) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6608), .ZN(U3180) );
  NOR2_X1 U7417 ( .A1(n6497), .A2(n6503), .ZN(n6504) );
  AOI22_X1 U7418 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6512) );
  AND2_X1 U7419 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6501) );
  INV_X1 U7420 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6499) );
  INV_X1 U7421 ( .A(NA_N), .ZN(n6505) );
  AOI221_X1 U7422 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6505), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6509) );
  AOI221_X1 U7423 ( .B1(n6501), .B2(n6607), .C1(n6499), .C2(n6607), .A(n6509), 
        .ZN(n6498) );
  OAI21_X1 U7424 ( .B1(n6504), .B2(n6512), .A(n6498), .ZN(U3181) );
  NOR2_X1 U7425 ( .A1(n6507), .A2(n6499), .ZN(n6506) );
  NAND2_X1 U7426 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6500) );
  OAI21_X1 U7427 ( .B1(n6506), .B2(n6501), .A(n6500), .ZN(n6502) );
  OAI211_X1 U7428 ( .C1(n6503), .C2(n6603), .A(n6596), .B(n6502), .ZN(U3182)
         );
  AOI21_X1 U7429 ( .B1(n6506), .B2(n6505), .A(n6504), .ZN(n6511) );
  AOI221_X1 U7430 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6603), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6508) );
  AOI221_X1 U7431 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6508), .C2(HOLD), .A(n6507), .ZN(n6510) );
  OAI22_X1 U7432 ( .A1(n6512), .A2(n6511), .B1(n6510), .B2(n6509), .ZN(U3183)
         );
  NAND2_X1 U7433 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6535), .ZN(n6559) );
  NOR2_X2 U7434 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6607), .ZN(n6557) );
  AOI22_X1 U7435 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6607), .ZN(n6513) );
  OAI21_X1 U7436 ( .B1(n6589), .B2(n6559), .A(n6513), .ZN(U3184) );
  AOI22_X1 U7437 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6607), .ZN(n6514) );
  OAI21_X1 U7438 ( .B1(n6515), .B2(n6559), .A(n6514), .ZN(U3185) );
  AOI22_X1 U7439 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6607), .ZN(n6516) );
  OAI21_X1 U7440 ( .B1(n6517), .B2(n6559), .A(n6516), .ZN(U3186) );
  AOI22_X1 U7441 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6607), .ZN(n6518) );
  OAI21_X1 U7442 ( .B1(n6519), .B2(n6559), .A(n6518), .ZN(U3187) );
  INV_X1 U7443 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6745) );
  INV_X1 U7444 ( .A(n6557), .ZN(n6563) );
  OAI222_X1 U7445 ( .A1(n6559), .A2(n6520), .B1(n6745), .B2(n6535), .C1(n6522), 
        .C2(n6563), .ZN(U3188) );
  AOI22_X1 U7446 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6607), .ZN(n6521) );
  OAI21_X1 U7447 ( .B1(n6522), .B2(n6559), .A(n6521), .ZN(U3189) );
  AOI22_X1 U7448 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6607), .ZN(n6523) );
  OAI21_X1 U7449 ( .B1(n6524), .B2(n6559), .A(n6523), .ZN(U3190) );
  AOI22_X1 U7450 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6607), .ZN(n6525) );
  OAI21_X1 U7451 ( .B1(n5404), .B2(n6559), .A(n6525), .ZN(U3191) );
  AOI22_X1 U7452 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6607), .ZN(n6526) );
  OAI21_X1 U7453 ( .B1(n5162), .B2(n6559), .A(n6526), .ZN(U3192) );
  INV_X1 U7454 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7455 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6607), .ZN(n6527) );
  OAI21_X1 U7456 ( .B1(n6528), .B2(n6559), .A(n6527), .ZN(U3193) );
  INV_X1 U7457 ( .A(n6559), .ZN(n6561) );
  AOI22_X1 U7458 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6607), .ZN(n6529) );
  OAI21_X1 U7459 ( .B1(n6531), .B2(n6563), .A(n6529), .ZN(U3194) );
  AOI22_X1 U7460 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6607), .ZN(n6530) );
  OAI21_X1 U7461 ( .B1(n6531), .B2(n6559), .A(n6530), .ZN(U3195) );
  AOI22_X1 U7462 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6607), .ZN(n6532) );
  OAI21_X1 U7463 ( .B1(n6533), .B2(n6559), .A(n6532), .ZN(U3196) );
  AOI22_X1 U7464 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6607), .ZN(n6534) );
  OAI21_X1 U7465 ( .B1(n6536), .B2(n6563), .A(n6534), .ZN(U3197) );
  INV_X1 U7466 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6740) );
  OAI222_X1 U7467 ( .A1(n6559), .A2(n6536), .B1(n6740), .B2(n6535), .C1(n5325), 
        .C2(n6563), .ZN(U3198) );
  AOI22_X1 U7468 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6607), .ZN(n6537) );
  OAI21_X1 U7469 ( .B1(n5325), .B2(n6559), .A(n6537), .ZN(U3199) );
  AOI22_X1 U7470 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6607), .ZN(n6538) );
  OAI21_X1 U7471 ( .B1(n6540), .B2(n6563), .A(n6538), .ZN(U3200) );
  AOI22_X1 U7472 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6607), .ZN(n6539) );
  OAI21_X1 U7473 ( .B1(n6540), .B2(n6559), .A(n6539), .ZN(U3201) );
  AOI22_X1 U7474 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6607), .ZN(n6541) );
  OAI21_X1 U7475 ( .B1(n6542), .B2(n6563), .A(n6541), .ZN(U3202) );
  AOI22_X1 U7476 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6607), .ZN(n6543) );
  OAI21_X1 U7477 ( .B1(n6545), .B2(n6563), .A(n6543), .ZN(U3203) );
  AOI22_X1 U7478 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6607), .ZN(n6544) );
  OAI21_X1 U7479 ( .B1(n6545), .B2(n6559), .A(n6544), .ZN(U3204) );
  AOI22_X1 U7480 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6607), .ZN(n6546) );
  OAI21_X1 U7481 ( .B1(n6547), .B2(n6559), .A(n6546), .ZN(U3205) );
  AOI22_X1 U7482 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6607), .ZN(n6548) );
  OAI21_X1 U7483 ( .B1(n6549), .B2(n6563), .A(n6548), .ZN(U3206) );
  AOI222_X1 U7484 ( .A1(n6557), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6607), .C1(REIP_REG_24__SCAN_IN), .C2(
        n6561), .ZN(n6550) );
  INV_X1 U7485 ( .A(n6550), .ZN(U3207) );
  INV_X1 U7486 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6773) );
  AOI22_X1 U7487 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6607), .ZN(n6551) );
  OAI21_X1 U7488 ( .B1(n6773), .B2(n6559), .A(n6551), .ZN(U3208) );
  AOI22_X1 U7489 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6607), .ZN(n6552) );
  OAI21_X1 U7490 ( .B1(n6553), .B2(n6563), .A(n6552), .ZN(U3209) );
  AOI22_X1 U7491 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6607), .ZN(n6554) );
  OAI21_X1 U7492 ( .B1(n6555), .B2(n6563), .A(n6554), .ZN(U3210) );
  AOI22_X1 U7493 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6607), .ZN(n6556) );
  OAI21_X1 U7494 ( .B1(n6560), .B2(n6563), .A(n6556), .ZN(U3211) );
  AOI22_X1 U7495 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6557), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6607), .ZN(n6558) );
  OAI21_X1 U7496 ( .B1(n6560), .B2(n6559), .A(n6558), .ZN(U3212) );
  AOI22_X1 U7497 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6607), .ZN(n6562) );
  OAI21_X1 U7498 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(U3213) );
  MUX2_X1 U7499 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6607), .Z(U3445) );
  MUX2_X1 U7500 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6607), .Z(U3446) );
  MUX2_X1 U7501 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6607), .Z(U3447) );
  MUX2_X1 U7502 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6607), .Z(U3448) );
  OAI21_X1 U7503 ( .B1(n6567), .B2(DATAWIDTH_REG_0__SCAN_IN), .A(n6566), .ZN(
        n6565) );
  INV_X1 U7504 ( .A(n6565), .ZN(U3451) );
  INV_X1 U7505 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6582) );
  OAI21_X1 U7506 ( .B1(n6567), .B2(n6582), .A(n6566), .ZN(U3452) );
  OAI211_X1 U7507 ( .C1(n6570), .C2(n3174), .A(n6569), .B(n6568), .ZN(U3453)
         );
  NOR2_X1 U7508 ( .A1(n6571), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6572)
         );
  AOI211_X1 U7509 ( .C1(n6575), .C2(n6574), .A(n6573), .B(n6572), .ZN(n6577)
         );
  MUX2_X1 U7510 ( .A(n3304), .B(n6577), .S(n6576), .Z(n6578) );
  OAI21_X1 U7511 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(U3461) );
  INV_X1 U7512 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6783) );
  AOI221_X1 U7513 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6583), .C1(n6783), 
        .C2(n6582), .A(n6581), .ZN(n6585) );
  OAI22_X1 U7514 ( .A1(n6587), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(n6589), 
        .B2(n6586), .ZN(n6584) );
  NOR2_X1 U7515 ( .A1(n6585), .A2(n6584), .ZN(U3468) );
  OAI21_X1 U7516 ( .B1(n6587), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6586), .ZN(
        n6588) );
  OAI21_X1 U7517 ( .B1(n6590), .B2(n6589), .A(n6588), .ZN(U3469) );
  NAND2_X1 U7518 ( .A1(n6607), .A2(W_R_N_REG_SCAN_IN), .ZN(n6591) );
  OAI21_X1 U7519 ( .B1(n6607), .B2(READREQUEST_REG_SCAN_IN), .A(n6591), .ZN(
        U3470) );
  OAI21_X1 U7520 ( .B1(n6596), .B2(n6593), .A(n6592), .ZN(n6594) );
  NAND3_X1 U7521 ( .A1(n6594), .A2(STATE2_REG_2__SCAN_IN), .A3(n6603), .ZN(
        n6595) );
  AOI21_X1 U7522 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(n6600) );
  OAI21_X1 U7523 ( .B1(n6600), .B2(n6599), .A(n6598), .ZN(n6606) );
  AOI211_X1 U7524 ( .C1(n6604), .C2(n6603), .A(n6602), .B(n6601), .ZN(n6605)
         );
  MUX2_X1 U7525 ( .A(n6606), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6605), .Z(
        U3472) );
  MUX2_X1 U7526 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6607), .Z(U3473) );
  NAND2_X1 U7527 ( .A1(n6608), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6802) );
  INV_X1 U7528 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6610) );
  INV_X1 U7529 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6770) );
  AOI22_X1 U7530 ( .A1(n6610), .A2(keyinput80), .B1(keyinput97), .B2(n6770), 
        .ZN(n6609) );
  OAI221_X1 U7531 ( .B1(n6610), .B2(keyinput80), .C1(n6770), .C2(keyinput97), 
        .A(n6609), .ZN(n6622) );
  AOI22_X1 U7532 ( .A1(n6746), .A2(keyinput94), .B1(keyinput84), .B2(n6612), 
        .ZN(n6611) );
  OAI221_X1 U7533 ( .B1(n6746), .B2(keyinput94), .C1(n6612), .C2(keyinput84), 
        .A(n6611), .ZN(n6621) );
  AOI22_X1 U7534 ( .A1(n6615), .A2(keyinput71), .B1(n6614), .B2(keyinput127), 
        .ZN(n6613) );
  OAI221_X1 U7535 ( .B1(n6615), .B2(keyinput71), .C1(n6614), .C2(keyinput127), 
        .A(n6613), .ZN(n6620) );
  INV_X1 U7536 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6616) );
  XOR2_X1 U7537 ( .A(keyinput90), .B(n6616), .Z(n6618) );
  XNOR2_X1 U7538 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput72), .ZN(n6617)
         );
  NAND2_X1 U7539 ( .A1(n6618), .A2(n6617), .ZN(n6619) );
  NOR4_X1 U7540 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6662)
         );
  AOI22_X1 U7541 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput102), 
        .B1(INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput96), .ZN(n6623) );
  OAI221_X1 U7542 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput102), 
        .C1(INSTQUEUE_REG_4__6__SCAN_IN), .C2(keyinput96), .A(n6623), .ZN(
        n6633) );
  AOI22_X1 U7543 ( .A1(EBX_REG_4__SCAN_IN), .A2(keyinput113), .B1(
        INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput88), .ZN(n6624) );
  OAI221_X1 U7544 ( .B1(EBX_REG_4__SCAN_IN), .B2(keyinput113), .C1(
        INSTQUEUE_REG_6__4__SCAN_IN), .C2(keyinput88), .A(n6624), .ZN(n6632)
         );
  AOI22_X1 U7545 ( .A1(n6768), .A2(keyinput76), .B1(keyinput99), .B2(n6626), 
        .ZN(n6625) );
  OAI221_X1 U7546 ( .B1(n6768), .B2(keyinput76), .C1(n6626), .C2(keyinput99), 
        .A(n6625), .ZN(n6631) );
  INV_X1 U7547 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6628) );
  AOI22_X1 U7548 ( .A1(n6629), .A2(keyinput70), .B1(n6628), .B2(keyinput114), 
        .ZN(n6627) );
  OAI221_X1 U7549 ( .B1(n6629), .B2(keyinput70), .C1(n6628), .C2(keyinput114), 
        .A(n6627), .ZN(n6630) );
  NOR4_X1 U7550 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6661)
         );
  AOI22_X1 U7551 ( .A1(n5911), .A2(keyinput73), .B1(n3174), .B2(keyinput107), 
        .ZN(n6634) );
  OAI221_X1 U7552 ( .B1(n5911), .B2(keyinput73), .C1(n3174), .C2(keyinput107), 
        .A(n6634), .ZN(n6635) );
  INV_X1 U7553 ( .A(n6635), .ZN(n6647) );
  INV_X1 U7554 ( .A(DATAI_22_), .ZN(n6638) );
  INV_X1 U7555 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6637) );
  AOI22_X1 U7556 ( .A1(n6638), .A2(keyinput86), .B1(n6637), .B2(keyinput126), 
        .ZN(n6636) );
  OAI221_X1 U7557 ( .B1(n6638), .B2(keyinput86), .C1(n6637), .C2(keyinput126), 
        .A(n6636), .ZN(n6641) );
  INV_X1 U7558 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n6639) );
  XNOR2_X1 U7559 ( .A(n6639), .B(keyinput124), .ZN(n6640) );
  NOR2_X1 U7560 ( .A1(n6641), .A2(n6640), .ZN(n6646) );
  AOI22_X1 U7561 ( .A1(n4923), .A2(keyinput64), .B1(keyinput110), .B2(n6737), 
        .ZN(n6642) );
  OAI221_X1 U7562 ( .B1(n4923), .B2(keyinput64), .C1(n6737), .C2(keyinput110), 
        .A(n6642), .ZN(n6643) );
  INV_X1 U7563 ( .A(n6643), .ZN(n6645) );
  XNOR2_X1 U7564 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput111), .ZN(n6644) );
  AND4_X1 U7565 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6660)
         );
  INV_X1 U7566 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7567 ( .A1(n3630), .A2(keyinput82), .B1(keyinput104), .B2(n6649), 
        .ZN(n6648) );
  OAI221_X1 U7568 ( .B1(n3630), .B2(keyinput82), .C1(n6649), .C2(keyinput104), 
        .A(n6648), .ZN(n6658) );
  INV_X1 U7569 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6652) );
  INV_X1 U7570 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U7571 ( .A1(n6652), .A2(keyinput100), .B1(keyinput93), .B2(n6651), 
        .ZN(n6650) );
  OAI221_X1 U7572 ( .B1(n6652), .B2(keyinput100), .C1(n6651), .C2(keyinput93), 
        .A(n6650), .ZN(n6657) );
  AOI22_X1 U7573 ( .A1(n6752), .A2(keyinput125), .B1(n6771), .B2(keyinput83), 
        .ZN(n6653) );
  OAI221_X1 U7574 ( .B1(n6752), .B2(keyinput125), .C1(n6771), .C2(keyinput83), 
        .A(n6653), .ZN(n6656) );
  AOI22_X1 U7575 ( .A1(n6757), .A2(keyinput103), .B1(keyinput123), .B2(n6745), 
        .ZN(n6654) );
  OAI221_X1 U7576 ( .B1(n6757), .B2(keyinput103), .C1(n6745), .C2(keyinput123), 
        .A(n6654), .ZN(n6655) );
  NOR4_X1 U7577 ( .A1(n6658), .A2(n6657), .A3(n6656), .A4(n6655), .ZN(n6659)
         );
  AND4_X1 U7578 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6800)
         );
  OAI22_X1 U7579 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput79), .B1(
        keyinput119), .B2(DATAO_REG_17__SCAN_IN), .ZN(n6663) );
  AOI221_X1 U7580 ( .B1(INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput79), .C1(
        DATAO_REG_17__SCAN_IN), .C2(keyinput119), .A(n6663), .ZN(n6670) );
  OAI22_X1 U7581 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput105), .B1(
        keyinput109), .B2(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6664) );
  AOI221_X1 U7582 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput105), .C1(
        DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput109), .A(n6664), .ZN(n6669) );
  OAI22_X1 U7583 ( .A1(LWORD_REG_5__SCAN_IN), .A2(keyinput77), .B1(keyinput108), .B2(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6665) );
  AOI221_X1 U7584 ( .B1(LWORD_REG_5__SCAN_IN), .B2(keyinput77), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(keyinput108), .A(n6665), .ZN(n6668) );
  OAI22_X1 U7585 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput117), .B1(
        keyinput98), .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6666) );
  AOI221_X1 U7586 ( .B1(INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput117), .C1(
        INSTQUEUE_REG_14__6__SCAN_IN), .C2(keyinput98), .A(n6666), .ZN(n6667)
         );
  NAND4_X1 U7587 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6698)
         );
  OAI22_X1 U7588 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput121), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput101), .ZN(n6671) );
  AOI221_X1 U7589 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput121), .C1(
        keyinput101), .C2(DATAWIDTH_REG_0__SCAN_IN), .A(n6671), .ZN(n6678) );
  OAI22_X1 U7590 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(keyinput116), .B1(
        keyinput89), .B2(REIP_REG_24__SCAN_IN), .ZN(n6672) );
  AOI221_X1 U7591 ( .B1(INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput116), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput89), .A(n6672), .ZN(n6677) );
  OAI22_X1 U7592 ( .A1(EBX_REG_7__SCAN_IN), .A2(keyinput75), .B1(keyinput81), 
        .B2(EAX_REG_6__SCAN_IN), .ZN(n6673) );
  AOI221_X1 U7593 ( .B1(EBX_REG_7__SCAN_IN), .B2(keyinput75), .C1(
        EAX_REG_6__SCAN_IN), .C2(keyinput81), .A(n6673), .ZN(n6676) );
  OAI22_X1 U7594 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(keyinput65), .B1(
        keyinput91), .B2(DATAO_REG_9__SCAN_IN), .ZN(n6674) );
  AOI221_X1 U7595 ( .B1(INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput65), .C1(
        DATAO_REG_9__SCAN_IN), .C2(keyinput91), .A(n6674), .ZN(n6675) );
  NAND4_X1 U7596 ( .A1(n6678), .A2(n6677), .A3(n6676), .A4(n6675), .ZN(n6697)
         );
  OAI22_X1 U7597 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput120), .B1(
        DATAI_0_), .B2(keyinput67), .ZN(n6679) );
  AOI221_X1 U7598 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput120), .C1(
        keyinput67), .C2(DATAI_0_), .A(n6679), .ZN(n6686) );
  OAI22_X1 U7599 ( .A1(EBX_REG_25__SCAN_IN), .A2(keyinput122), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput66), .ZN(n6680) );
  AOI221_X1 U7600 ( .B1(EBX_REG_25__SCAN_IN), .B2(keyinput122), .C1(keyinput66), .C2(DATAO_REG_0__SCAN_IN), .A(n6680), .ZN(n6685) );
  OAI22_X1 U7601 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput118), .B1(
        keyinput92), .B2(ADDRESS_REG_14__SCAN_IN), .ZN(n6681) );
  AOI221_X1 U7602 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput118), 
        .C1(ADDRESS_REG_14__SCAN_IN), .C2(keyinput92), .A(n6681), .ZN(n6684)
         );
  OAI22_X1 U7603 ( .A1(EAX_REG_27__SCAN_IN), .A2(keyinput69), .B1(keyinput87), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n6682) );
  AOI221_X1 U7604 ( .B1(EAX_REG_27__SCAN_IN), .B2(keyinput69), .C1(
        REIP_REG_8__SCAN_IN), .C2(keyinput87), .A(n6682), .ZN(n6683) );
  NAND4_X1 U7605 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n6696)
         );
  OAI22_X1 U7606 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(keyinput68), .B1(
        keyinput115), .B2(EBX_REG_23__SCAN_IN), .ZN(n6687) );
  AOI221_X1 U7607 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(keyinput68), 
        .C1(EBX_REG_23__SCAN_IN), .C2(keyinput115), .A(n6687), .ZN(n6694) );
  OAI22_X1 U7608 ( .A1(DATAI_28_), .A2(keyinput106), .B1(keyinput85), .B2(
        ADDRESS_REG_23__SCAN_IN), .ZN(n6688) );
  AOI221_X1 U7609 ( .B1(DATAI_28_), .B2(keyinput106), .C1(
        ADDRESS_REG_23__SCAN_IN), .C2(keyinput85), .A(n6688), .ZN(n6693) );
  OAI22_X1 U7610 ( .A1(EAX_REG_31__SCAN_IN), .A2(keyinput95), .B1(keyinput74), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n6689) );
  AOI221_X1 U7611 ( .B1(EAX_REG_31__SCAN_IN), .B2(keyinput95), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput74), .A(n6689), .ZN(n6692) );
  OAI22_X1 U7612 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput78), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput112), .ZN(n6690) );
  AOI221_X1 U7613 ( .B1(INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput78), .C1(
        keyinput112), .C2(DATAWIDTH_REG_18__SCAN_IN), .A(n6690), .ZN(n6691) );
  NAND4_X1 U7614 ( .A1(n6694), .A2(n6693), .A3(n6692), .A4(n6691), .ZN(n6695)
         );
  NOR4_X1 U7615 ( .A1(n6698), .A2(n6697), .A3(n6696), .A4(n6695), .ZN(n6799)
         );
  AOI22_X1 U7616 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput56), .B1(
        INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput53), .ZN(n6699) );
  OAI221_X1 U7617 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput56), .C1(
        INSTQUEUE_REG_9__0__SCAN_IN), .C2(keyinput53), .A(n6699), .ZN(n6706)
         );
  AOI22_X1 U7618 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput44), .B1(
        DATAI_28_), .B2(keyinput42), .ZN(n6700) );
  OAI221_X1 U7619 ( .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput44), .C1(
        DATAI_28_), .C2(keyinput42), .A(n6700), .ZN(n6705) );
  AOI22_X1 U7620 ( .A1(EBX_REG_25__SCAN_IN), .A2(keyinput58), .B1(
        INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput50), .ZN(n6701) );
  OAI221_X1 U7621 ( .B1(EBX_REG_25__SCAN_IN), .B2(keyinput58), .C1(
        INSTQUEUE_REG_14__0__SCAN_IN), .C2(keyinput50), .A(n6701), .ZN(n6704)
         );
  AOI22_X1 U7622 ( .A1(EAX_REG_6__SCAN_IN), .A2(keyinput17), .B1(
        INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput32), .ZN(n6702) );
  OAI221_X1 U7623 ( .B1(EAX_REG_6__SCAN_IN), .B2(keyinput17), .C1(
        INSTQUEUE_REG_4__6__SCAN_IN), .C2(keyinput32), .A(n6702), .ZN(n6703)
         );
  NOR4_X1 U7624 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n6734)
         );
  AOI22_X1 U7625 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(keyinput6), .B1(
        INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput16), .ZN(n6707) );
  OAI221_X1 U7626 ( .B1(DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput6), .C1(
        INSTQUEUE_REG_13__2__SCAN_IN), .C2(keyinput16), .A(n6707), .ZN(n6714)
         );
  AOI22_X1 U7627 ( .A1(UWORD_REG_13__SCAN_IN), .A2(keyinput29), .B1(
        EAX_REG_12__SCAN_IN), .B2(keyinput20), .ZN(n6708) );
  OAI221_X1 U7628 ( .B1(UWORD_REG_13__SCAN_IN), .B2(keyinput29), .C1(
        EAX_REG_12__SCAN_IN), .C2(keyinput20), .A(n6708), .ZN(n6713) );
  AOI22_X1 U7629 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput25), .B1(
        INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput0), .ZN(n6709) );
  OAI221_X1 U7630 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput25), .C1(
        INSTQUEUE_REG_5__4__SCAN_IN), .C2(keyinput0), .A(n6709), .ZN(n6712) );
  AOI22_X1 U7631 ( .A1(DATAO_REG_16__SCAN_IN), .A2(keyinput60), .B1(
        EAX_REG_28__SCAN_IN), .B2(keyinput35), .ZN(n6710) );
  OAI221_X1 U7632 ( .B1(DATAO_REG_16__SCAN_IN), .B2(keyinput60), .C1(
        EAX_REG_28__SCAN_IN), .C2(keyinput35), .A(n6710), .ZN(n6711) );
  NOR4_X1 U7633 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6733)
         );
  AOI22_X1 U7634 ( .A1(DATAI_22_), .A2(keyinput22), .B1(DATAI_9_), .B2(
        keyinput7), .ZN(n6715) );
  OAI221_X1 U7635 ( .B1(DATAI_22_), .B2(keyinput22), .C1(DATAI_9_), .C2(
        keyinput7), .A(n6715), .ZN(n6722) );
  AOI22_X1 U7636 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput27), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput18), .ZN(n6716) );
  OAI221_X1 U7637 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput27), .C1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput18), .A(n6716), .ZN(n6721) );
  AOI22_X1 U7638 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(keyinput4), .B1(
        INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput24), .ZN(n6717) );
  OAI221_X1 U7639 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(keyinput4), .C1(
        INSTQUEUE_REG_6__4__SCAN_IN), .C2(keyinput24), .A(n6717), .ZN(n6720)
         );
  AOI22_X1 U7640 ( .A1(DATAO_REG_8__SCAN_IN), .A2(keyinput26), .B1(DATAI_26_), 
        .B2(keyinput9), .ZN(n6718) );
  OAI221_X1 U7641 ( .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput26), .C1(DATAI_26_), 
        .C2(keyinput9), .A(n6718), .ZN(n6719) );
  NOR4_X1 U7642 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n6732)
         );
  AOI22_X1 U7643 ( .A1(UWORD_REG_8__SCAN_IN), .A2(keyinput36), .B1(
        EAX_REG_27__SCAN_IN), .B2(keyinput5), .ZN(n6723) );
  OAI221_X1 U7644 ( .B1(UWORD_REG_8__SCAN_IN), .B2(keyinput36), .C1(
        EAX_REG_27__SCAN_IN), .C2(keyinput5), .A(n6723), .ZN(n6730) );
  AOI22_X1 U7645 ( .A1(LWORD_REG_10__SCAN_IN), .A2(keyinput40), .B1(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput63), .ZN(n6724) );
  OAI221_X1 U7646 ( .B1(LWORD_REG_10__SCAN_IN), .B2(keyinput40), .C1(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(keyinput63), .A(n6724), .ZN(
        n6729) );
  AOI22_X1 U7647 ( .A1(REIP_REG_8__SCAN_IN), .A2(keyinput23), .B1(
        INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput62), .ZN(n6725) );
  OAI221_X1 U7648 ( .B1(REIP_REG_8__SCAN_IN), .B2(keyinput23), .C1(
        INSTQUEUE_REG_8__7__SCAN_IN), .C2(keyinput62), .A(n6725), .ZN(n6728)
         );
  AOI22_X1 U7649 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput21), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput2), .ZN(n6726) );
  OAI221_X1 U7650 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput21), .C1(
        DATAO_REG_0__SCAN_IN), .C2(keyinput2), .A(n6726), .ZN(n6727) );
  NOR4_X1 U7651 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6731)
         );
  NAND4_X1 U7652 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n6798)
         );
  AOI22_X1 U7653 ( .A1(n6737), .A2(keyinput46), .B1(keyinput45), .B2(n6736), 
        .ZN(n6735) );
  OAI221_X1 U7654 ( .B1(n6737), .B2(keyinput46), .C1(n6736), .C2(keyinput45), 
        .A(n6735), .ZN(n6750) );
  INV_X1 U7655 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U7656 ( .A1(n6740), .A2(keyinput28), .B1(n6739), .B2(keyinput57), 
        .ZN(n6738) );
  OAI221_X1 U7657 ( .B1(n6740), .B2(keyinput28), .C1(n6739), .C2(keyinput57), 
        .A(n6738), .ZN(n6749) );
  AOI22_X1 U7658 ( .A1(n6743), .A2(keyinput1), .B1(keyinput48), .B2(n6742), 
        .ZN(n6741) );
  OAI221_X1 U7659 ( .B1(n6743), .B2(keyinput1), .C1(n6742), .C2(keyinput48), 
        .A(n6741), .ZN(n6748) );
  AOI22_X1 U7660 ( .A1(n6746), .A2(keyinput30), .B1(keyinput59), .B2(n6745), 
        .ZN(n6744) );
  OAI221_X1 U7661 ( .B1(n6746), .B2(keyinput30), .C1(n6745), .C2(keyinput59), 
        .A(n6744), .ZN(n6747) );
  NOR4_X1 U7662 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6796)
         );
  INV_X1 U7663 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6753) );
  AOI22_X1 U7664 ( .A1(n6753), .A2(keyinput34), .B1(keyinput61), .B2(n6752), 
        .ZN(n6751) );
  OAI221_X1 U7665 ( .B1(n6753), .B2(keyinput34), .C1(n6752), .C2(keyinput61), 
        .A(n6751), .ZN(n6763) );
  AOI22_X1 U7666 ( .A1(EAX_REG_31__SCAN_IN), .A2(keyinput31), .B1(n6755), .B2(
        keyinput51), .ZN(n6754) );
  OAI221_X1 U7667 ( .B1(EAX_REG_31__SCAN_IN), .B2(keyinput31), .C1(n6755), 
        .C2(keyinput51), .A(n6754), .ZN(n6762) );
  AOI22_X1 U7668 ( .A1(DATAI_0_), .A2(keyinput3), .B1(STATE2_REG_3__SCAN_IN), 
        .B2(keyinput43), .ZN(n6756) );
  OAI221_X1 U7669 ( .B1(DATAI_0_), .B2(keyinput3), .C1(STATE2_REG_3__SCAN_IN), 
        .C2(keyinput43), .A(n6756), .ZN(n6761) );
  XOR2_X1 U7670 ( .A(n6757), .B(keyinput39), .Z(n6759) );
  XNOR2_X1 U7671 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput47), .ZN(n6758)
         );
  NAND2_X1 U7672 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NOR4_X1 U7673 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6795)
         );
  INV_X1 U7674 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U7675 ( .A1(n6766), .A2(keyinput49), .B1(keyinput13), .B2(n6765), 
        .ZN(n6764) );
  OAI221_X1 U7676 ( .B1(n6766), .B2(keyinput49), .C1(n6765), .C2(keyinput13), 
        .A(n6764), .ZN(n6778) );
  AOI22_X1 U7677 ( .A1(n4927), .A2(keyinput11), .B1(keyinput12), .B2(n6768), 
        .ZN(n6767) );
  OAI221_X1 U7678 ( .B1(n4927), .B2(keyinput11), .C1(n6768), .C2(keyinput12), 
        .A(n6767), .ZN(n6777) );
  AOI22_X1 U7679 ( .A1(n6771), .A2(keyinput19), .B1(keyinput33), .B2(n6770), 
        .ZN(n6769) );
  OAI221_X1 U7680 ( .B1(n6771), .B2(keyinput19), .C1(n6770), .C2(keyinput33), 
        .A(n6769), .ZN(n6776) );
  INV_X1 U7681 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U7682 ( .A1(n6774), .A2(keyinput52), .B1(keyinput10), .B2(n6773), 
        .ZN(n6772) );
  OAI221_X1 U7683 ( .B1(n6774), .B2(keyinput52), .C1(n6773), .C2(keyinput10), 
        .A(n6772), .ZN(n6775) );
  NOR4_X1 U7684 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6794)
         );
  INV_X1 U7685 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6780) );
  AOI22_X1 U7686 ( .A1(n4470), .A2(keyinput14), .B1(keyinput41), .B2(n6780), 
        .ZN(n6779) );
  OAI221_X1 U7687 ( .B1(n4470), .B2(keyinput14), .C1(n6780), .C2(keyinput41), 
        .A(n6779), .ZN(n6792) );
  AOI22_X1 U7688 ( .A1(n6783), .A2(keyinput37), .B1(n6782), .B2(keyinput54), 
        .ZN(n6781) );
  OAI221_X1 U7689 ( .B1(n6783), .B2(keyinput37), .C1(n6782), .C2(keyinput54), 
        .A(n6781), .ZN(n6791) );
  INV_X1 U7690 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6786) );
  AOI22_X1 U7691 ( .A1(n6786), .A2(keyinput55), .B1(n6785), .B2(keyinput38), 
        .ZN(n6784) );
  OAI221_X1 U7692 ( .B1(n6786), .B2(keyinput55), .C1(n6785), .C2(keyinput38), 
        .A(n6784), .ZN(n6790) );
  XNOR2_X1 U7693 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput8), .ZN(n6788)
         );
  XNOR2_X1 U7694 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .B(keyinput15), .ZN(n6787)
         );
  NAND2_X1 U7695 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  NOR4_X1 U7696 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6793)
         );
  NAND4_X1 U7697 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n6797)
         );
  AOI211_X1 U7698 ( .C1(n6800), .C2(n6799), .A(n6798), .B(n6797), .ZN(n6801)
         );
  XNOR2_X1 U7699 ( .A(n6802), .B(n6801), .ZN(U3165) );
  CLKBUF_X1 U3442 ( .A(n3780), .Z(n3006) );
  CLKBUF_X1 U34620 ( .A(n3089), .Z(n3759) );
  AND2_X1 U34690 ( .A1(n3168), .A2(n3167), .ZN(n3918) );
  CLKBUF_X1 U3480 ( .A(n3074), .Z(n3754) );
  CLKBUF_X1 U3484 ( .A(n3118), .Z(n3781) );
  AND2_X1 U3491 ( .A1(n5229), .A2(n5230), .ZN(n3503) );
  CLKBUF_X1 U3520 ( .A(n3934), .Z(n5530) );
  CLKBUF_X1 U3566 ( .A(n4051), .Z(n5592) );
  CLKBUF_X1 U3585 ( .A(n5723), .Z(n2996) );
  CLKBUF_X2 U3586 ( .A(n3927), .Z(n5072) );
  CLKBUF_X1 U3587 ( .A(n6175), .Z(n6184) );
  INV_X2 U3594 ( .A(n6476), .ZN(n6604) );
endmodule

