

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4718;

  INV_X2 U2249 ( .A(n4510), .ZN(n4299) );
  INV_X1 U2250 ( .A(n4094), .ZN(n3700) );
  INV_X1 U2251 ( .A(n2357), .ZN(n2697) );
  CLKBUF_X2 U2252 ( .A(n2328), .Z(n3739) );
  NAND2_X1 U2253 ( .A1(n3029), .A2(n2759), .ZN(n3508) );
  NAND2_X1 U2254 ( .A1(n2717), .A2(IR_REG_31__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U2255 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2385) );
  NAND2_X1 U2256 ( .A1(n2695), .A2(n3874), .ZN(n2760) );
  INV_X2 U2257 ( .A(n3506), .ZN(n2934) );
  CLKBUF_X3 U2258 ( .A(n3012), .Z(n3372) );
  INV_X1 U2259 ( .A(n4132), .ZN(n4092) );
  NAND2_X1 U2261 ( .A1(n3735), .A2(n3865), .ZN(n4076) );
  NAND4_X2 U2262 ( .A1(n2332), .A2(n2331), .A3(n2330), .A4(n2329), .ZN(n3594)
         );
  AND2_X1 U2263 ( .A1(n2751), .A2(n3874), .ZN(n4544) );
  INV_X2 U2264 ( .A(n4515), .ZN(n4313) );
  INV_X1 U2265 ( .A(n3899), .ZN(U4043) );
  XNOR2_X2 U2266 ( .A(n2715), .B(IR_REG_26__SCAN_IN), .ZN(n2738) );
  NOR2_X1 U2267 ( .A1(n4496), .A2(n4497), .ZN(n4495) );
  NAND2_X2 U2268 ( .A1(n2954), .A2(n2953), .ZN(n2952) );
  NAND2_X2 U2269 ( .A1(n3807), .A2(n3810), .ZN(n2953) );
  MUX2_X2 U2270 ( .A(REG0_REG_28__SCAN_IN), .B(n2754), .S(n4553), .Z(n2755) );
  MUX2_X2 U2271 ( .A(REG1_REG_28__SCAN_IN), .B(n2754), .S(n4561), .Z(n2744) );
  NAND2_X2 U2272 ( .A1(n2302), .A2(IR_REG_31__SCAN_IN), .ZN(n2303) );
  XNOR2_X2 U2273 ( .A(n2785), .B(n2827), .ZN(n2821) );
  NAND2_X2 U2274 ( .A1(n3915), .A2(n2784), .ZN(n2785) );
  OAI211_X4 U2275 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_1__SCAN_IN), .A(n2101), 
        .B(n2100), .ZN(n2792) );
  OAI21_X2 U2276 ( .B1(n3145), .B2(n3816), .A(n3830), .ZN(n2998) );
  NAND2_X2 U2277 ( .A1(n2170), .A2(n3815), .ZN(n3145) );
  BUF_X4 U2278 ( .A(n3012), .Z(n2007) );
  INV_X1 U2279 ( .A(n3508), .ZN(n3012) );
  XNOR2_X2 U2280 ( .A(n2832), .B(n2828), .ZN(n2831) );
  NAND2_X2 U2281 ( .A1(n2132), .A2(n2786), .ZN(n2832) );
  XNOR2_X2 U2282 ( .A(n2719), .B(n2718), .ZN(n2736) );
  XNOR2_X2 U2283 ( .A(n3996), .B(n4009), .ZN(n3989) );
  NOR2_X1 U2284 ( .A1(n4495), .A2(n2148), .ZN(n2147) );
  OAI21_X1 U2285 ( .B1(n2206), .B2(n2212), .A(n2620), .ZN(n2063) );
  NAND2_X1 U2286 ( .A1(n4002), .A2(n4003), .ZN(n4024) );
  NOR2_X2 U2287 ( .A1(n4118), .A2(n2748), .ZN(n4097) );
  AOI21_X1 U2288 ( .B1(n3944), .B2(n3223), .A(n2143), .ZN(n2140) );
  NAND2_X1 U2289 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  INV_X2 U2290 ( .A(n2011), .ZN(n3509) );
  NAND2_X1 U2291 ( .A1(n2928), .A2(n2341), .ZN(n3807) );
  INV_X1 U2292 ( .A(n3594), .ZN(n2928) );
  INV_X2 U2293 ( .A(n4456), .ZN(n2305) );
  NOR2_X1 U2294 ( .A1(n2333), .A2(n2281), .ZN(n2339) );
  AOI21_X1 U2295 ( .B1(n4332), .B2(n4547), .A(n2172), .ZN(n2171) );
  XNOR2_X1 U2296 ( .A(n2063), .B(n2062), .ZN(n4336) );
  NAND2_X1 U2297 ( .A1(n4024), .A2(n2149), .ZN(n4496) );
  NAND2_X1 U2298 ( .A1(n3562), .A2(n3447), .ZN(n3565) );
  AOI21_X1 U2299 ( .B1(n2609), .B2(n2204), .A(n2202), .ZN(n2201) );
  NAND2_X1 U2300 ( .A1(n4482), .A2(n4285), .ZN(n4481) );
  AOI21_X1 U2301 ( .B1(n4184), .B2(n2582), .A(n2284), .ZN(n4165) );
  OAI21_X1 U2302 ( .B1(n2205), .B2(n2203), .A(n2638), .ZN(n2202) );
  OR2_X1 U2303 ( .A1(n3363), .A2(n2079), .ZN(n2074) );
  NOR2_X1 U2304 ( .A1(n4334), .A2(n4528), .ZN(n2172) );
  NAND2_X1 U2305 ( .A1(n4282), .A2(n4281), .ZN(n4280) );
  OAI21_X1 U2306 ( .B1(n4100), .B2(n4099), .A(n4098), .ZN(n4409) );
  NAND2_X1 U2307 ( .A1(n3303), .A2(n2258), .ZN(n2256) );
  OAI21_X1 U2308 ( .B1(n3941), .B2(n2141), .A(n2140), .ZN(n3953) );
  NOR2_X1 U2309 ( .A1(n2077), .A2(n3617), .ZN(n2071) );
  AOI21_X1 U2310 ( .B1(n2252), .B2(n2250), .A(n2288), .ZN(n2249) );
  NOR2_X1 U2311 ( .A1(n2255), .A2(n3645), .ZN(n2250) );
  AOI21_X1 U2312 ( .B1(n2258), .B2(n2261), .A(n2035), .ZN(n2257) );
  OAI21_X1 U2313 ( .B1(n2028), .B2(n2254), .A(n3408), .ZN(n2253) );
  INV_X1 U2314 ( .A(n2028), .ZN(n2255) );
  OR2_X1 U2315 ( .A1(n3407), .A2(n3629), .ZN(n3408) );
  OAI22_X1 U2316 ( .A1(n2098), .A2(n2096), .B1(n3112), .B2(n2099), .ZN(n2095)
         );
  NAND2_X1 U2317 ( .A1(n3162), .A2(n2019), .ZN(n3336) );
  AND2_X1 U2318 ( .A1(n4249), .A2(n2031), .ZN(n2225) );
  OAI211_X1 U2319 ( .C1(n2125), .C2(n2180), .A(n2123), .B(n2280), .ZN(n3934)
         );
  AND2_X1 U2320 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  XNOR2_X1 U2321 ( .A(n2181), .B(n3124), .ZN(n2987) );
  NAND2_X1 U2322 ( .A1(n2549), .A2(REG3_REG_19__SCAN_IN), .ZN(n2564) );
  AOI22_X1 U2323 ( .A1(n2846), .A2(REG1_REG_6__SCAN_IN), .B1(n4463), .B2(n2845), .ZN(n2984) );
  NOR2_X2 U2324 ( .A1(n2932), .A2(n4544), .ZN(n2971) );
  INV_X2 U2325 ( .A(n2932), .ZN(n3456) );
  AND2_X1 U2326 ( .A1(n3812), .A2(n3809), .ZN(n3781) );
  AND2_X1 U2327 ( .A1(n3813), .A2(n3815), .ZN(n3778) );
  OR2_X1 U2328 ( .A1(n3100), .A2(n3898), .ZN(n3812) );
  NAND2_X1 U2329 ( .A1(n2675), .A2(n3825), .ZN(n3820) );
  INV_X1 U2330 ( .A(n2760), .ZN(n3029) );
  XNOR2_X1 U2331 ( .A(n2844), .B(n4463), .ZN(n2846) );
  NAND2_X1 U2332 ( .A1(n3205), .A2(n3245), .ZN(n3825) );
  NAND4_X1 U2333 ( .A1(n2364), .A2(n2363), .A3(n2362), .A4(n2361), .ZN(n3897)
         );
  NAND2_X1 U2334 ( .A1(n2317), .A2(n2318), .ZN(n2745) );
  NAND3_X2 U2335 ( .A1(n2738), .A2(n4458), .A3(n2737), .ZN(n2759) );
  CLKBUF_X3 U2336 ( .A(n2360), .Z(n3742) );
  OAI21_X1 U2337 ( .B1(n2661), .B2(n2282), .A(n2660), .ZN(n3800) );
  CLKBUF_X3 U2338 ( .A(n2344), .Z(n2642) );
  XNOR2_X1 U2339 ( .A(n2721), .B(n4688), .ZN(n2735) );
  NAND2_X1 U2340 ( .A1(n2720), .A2(IR_REG_31__SCAN_IN), .ZN(n2721) );
  AOI21_X1 U2341 ( .B1(n2026), .B2(n2664), .A(n2663), .ZN(n2666) );
  OAI21_X1 U2342 ( .B1(n2720), .B2(IR_REG_25__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2715) );
  XNOR2_X1 U2343 ( .A(n2668), .B(IR_REG_22__SCAN_IN), .ZN(n3884) );
  INV_X1 U2344 ( .A(n2306), .ZN(n4455) );
  OR2_X1 U2345 ( .A1(n2704), .A2(IR_REG_27__SCAN_IN), .ZN(n2314) );
  OAI21_X1 U2346 ( .B1(n2794), .B2(REG2_REG_2__SCAN_IN), .A(n2066), .ZN(n3917)
         );
  NAND2_X1 U2347 ( .A1(n2312), .A2(IR_REG_31__SCAN_IN), .ZN(n2704) );
  NAND2_X2 U2348 ( .A1(n2339), .A2(n2338), .ZN(n2794) );
  AND2_X1 U2349 ( .A1(n2367), .A2(n2300), .ZN(n2237) );
  INV_X1 U2350 ( .A(n2334), .ZN(n2367) );
  AND2_X1 U2351 ( .A1(n2530), .A2(n2294), .ZN(n2656) );
  NOR2_X1 U2352 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2291)
         );
  INV_X1 U2353 ( .A(IR_REG_22__SCAN_IN), .ZN(n2711) );
  NOR2_X1 U2354 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2530)
         );
  NOR2_X1 U2355 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2290)
         );
  NOR2_X1 U2356 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2289)
         );
  INV_X1 U2357 ( .A(IR_REG_25__SCAN_IN), .ZN(n4688) );
  AND2_X1 U2358 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2664)
         );
  NOR2_X1 U2359 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2300)
         );
  NOR2_X1 U2360 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2296)
         );
  NOR2_X1 U2361 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2297)
         );
  INV_X1 U2362 ( .A(IR_REG_13__SCAN_IN), .ZN(n2527) );
  AND2_X1 U2363 ( .A1(n2658), .A2(n2657), .ZN(n2712) );
  AND2_X2 U2364 ( .A1(n4718), .A2(n2367), .ZN(n2658) );
  OAI21_X2 U2365 ( .B1(n4109), .B2(n2692), .A(n3867), .ZN(n4077) );
  NAND2_X2 U2366 ( .A1(n4128), .A2(n3861), .ZN(n4109) );
  INV_X1 U2367 ( .A(IR_REG_31__SCAN_IN), .ZN(n2008) );
  NOR2_X2 U2368 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2713)
         );
  NAND2_X1 U2369 ( .A1(n4163), .A2(n2591), .ZN(n4144) );
  AOI22_X2 U2370 ( .A1(n3323), .A2(n2481), .B1(n3378), .B2(n3890), .ZN(n3295)
         );
  XNOR2_X2 U2371 ( .A(n2850), .B(n2839), .ZN(n2849) );
  NAND2_X2 U2372 ( .A1(n2892), .A2(n2837), .ZN(n2850) );
  AOI22_X2 U2373 ( .A1(n4201), .A2(n2572), .B1(n4214), .B2(n4231), .ZN(n4184)
         );
  AOI21_X2 U2374 ( .B1(n4144), .B2(n2600), .A(n2599), .ZN(n4126) );
  BUF_X4 U2375 ( .A(n3743), .Z(n2009) );
  BUF_X4 U2376 ( .A(n3743), .Z(n2010) );
  NAND2_X2 U2377 ( .A1(n2313), .A2(n2314), .ZN(n3743) );
  NAND4_X4 U2378 ( .A1(n2310), .A2(n2153), .A3(n2308), .A4(n2309), .ZN(n2325)
         );
  NOR2_X4 U2379 ( .A1(n3086), .A2(n3310), .ZN(n3162) );
  OR2_X2 U2380 ( .A1(n3244), .A2(n3196), .ZN(n3086) );
  CLKBUF_X3 U2381 ( .A(n2971), .Z(n2011) );
  NAND2_X1 U2382 ( .A1(n4455), .A2(n4456), .ZN(n2344) );
  NAND2_X1 U2383 ( .A1(n2233), .A2(n2231), .ZN(n2230) );
  NOR2_X1 U2384 ( .A1(n2232), .A2(n2443), .ZN(n2231) );
  INV_X1 U2385 ( .A(n2234), .ZN(n2232) );
  NOR2_X1 U2386 ( .A1(n2222), .A2(n2027), .ZN(n2221) );
  INV_X1 U2387 ( .A(n2253), .ZN(n2252) );
  AND2_X1 U2388 ( .A1(n2695), .A2(n3884), .ZN(n2908) );
  NAND2_X1 U2389 ( .A1(n2238), .A2(n2018), .ZN(n2665) );
  INV_X1 U2390 ( .A(n2558), .ZN(n2238) );
  INV_X1 U2391 ( .A(IR_REG_18__SCAN_IN), .ZN(n2239) );
  XNOR2_X1 U2392 ( .A(n2082), .B(n2934), .ZN(n3009) );
  NAND2_X1 U2393 ( .A1(n2084), .A2(n2083), .ZN(n2082) );
  NAND2_X1 U2394 ( .A1(n3456), .A2(n3094), .ZN(n2083) );
  NAND2_X1 U2395 ( .A1(n3898), .A2(n2007), .ZN(n2084) );
  NAND2_X1 U2396 ( .A1(n2236), .A2(n3453), .ZN(n3471) );
  NAND2_X1 U2397 ( .A1(n3565), .A2(n3452), .ZN(n2236) );
  OR2_X2 U2398 ( .A1(n2564), .A2(n3658), .ZN(n2575) );
  NAND2_X1 U2399 ( .A1(n2080), .A2(n3367), .ZN(n2079) );
  INV_X1 U2400 ( .A(n2642), .ZN(n2702) );
  NAND2_X1 U2401 ( .A1(n2608), .A2(n2034), .ZN(n2212) );
  INV_X1 U2402 ( .A(n2510), .ZN(n2509) );
  NOR2_X1 U2403 ( .A1(n3779), .A2(n2229), .ZN(n2228) );
  INV_X1 U2404 ( .A(n2442), .ZN(n2229) );
  AND2_X1 U2405 ( .A1(n3800), .A2(n2707), .ZN(n2751) );
  NAND2_X1 U2406 ( .A1(n3467), .A2(IR_REG_31__SCAN_IN), .ZN(n2067) );
  NAND2_X1 U2407 ( .A1(n2152), .A2(n2151), .ZN(n2150) );
  NOR2_X1 U2408 ( .A1(n3784), .A2(n2670), .ZN(n2151) );
  INV_X1 U2409 ( .A(n3783), .ZN(n2152) );
  INV_X1 U2410 ( .A(n3858), .ZN(n2162) );
  INV_X1 U2411 ( .A(n3856), .ZN(n2168) );
  INV_X1 U2412 ( .A(n2259), .ZN(n2258) );
  OAI21_X1 U2413 ( .B1(n2261), .B2(n3302), .A(n2260), .ZN(n2259) );
  INV_X1 U2414 ( .A(n3343), .ZN(n2260) );
  INV_X1 U2415 ( .A(n2890), .ZN(n2116) );
  INV_X1 U2416 ( .A(n3923), .ZN(n2125) );
  INV_X1 U2417 ( .A(n2190), .ZN(n2189) );
  OAI21_X1 U2418 ( .B1(n3935), .B2(n2191), .A(n3956), .ZN(n2190) );
  INV_X1 U2419 ( .A(n2111), .ZN(n2108) );
  OR2_X1 U2420 ( .A1(n2111), .A2(n2106), .ZN(n2105) );
  INV_X1 U2421 ( .A(n4469), .ZN(n2106) );
  NAND2_X1 U2422 ( .A1(n4013), .A2(REG2_REG_15__SCAN_IN), .ZN(n2137) );
  NAND2_X1 U2423 ( .A1(n2164), .A2(n2168), .ZN(n2163) );
  INV_X1 U2424 ( .A(n3853), .ZN(n2164) );
  AND2_X1 U2425 ( .A1(n2169), .A2(n3851), .ZN(n2167) );
  INV_X1 U2426 ( .A(n3854), .ZN(n2169) );
  NAND2_X1 U2427 ( .A1(n3648), .A2(n4290), .ZN(n2521) );
  INV_X1 U2428 ( .A(n2216), .ZN(n2215) );
  OAI21_X1 U2429 ( .B1(n3294), .B2(n2217), .A(n2508), .ZN(n2216) );
  AND2_X1 U2430 ( .A1(n4077), .A2(n4076), .ZN(n2175) );
  NOR2_X1 U2431 ( .A1(n2590), .A2(n2277), .ZN(n2276) );
  INV_X1 U2432 ( .A(n4156), .ZN(n2277) );
  AND2_X1 U2433 ( .A1(n2273), .A2(n4271), .ZN(n2272) );
  NOR2_X1 U2434 ( .A1(n4290), .A2(n4305), .ZN(n2273) );
  AND2_X1 U2435 ( .A1(n2671), .A2(n2923), .ZN(n2864) );
  INV_X1 U2436 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U2437 ( .A1(n2446), .A2(REG3_REG_11__SCAN_IN), .ZN(n2455) );
  INV_X1 U2438 ( .A(n2447), .ZN(n2446) );
  OR2_X2 U2439 ( .A1(n2455), .A2(n2454), .ZN(n2469) );
  INV_X1 U2440 ( .A(n2052), .ZN(n2261) );
  NOR2_X1 U2441 ( .A1(n3677), .A2(n2087), .ZN(n2086) );
  INV_X1 U2442 ( .A(n2262), .ZN(n2087) );
  INV_X1 U2443 ( .A(n2079), .ZN(n2076) );
  INV_X1 U2444 ( .A(n2249), .ZN(n2077) );
  NAND2_X1 U2445 ( .A1(n2252), .A2(n3415), .ZN(n2251) );
  INV_X1 U2446 ( .A(n3366), .ZN(n2073) );
  OR2_X1 U2447 ( .A1(n2344), .A2(n2881), .ZN(n2321) );
  NAND2_X1 U2448 ( .A1(n2179), .A2(n2178), .ZN(n2829) );
  NAND2_X1 U2449 ( .A1(n2779), .A2(n4465), .ZN(n2178) );
  NAND2_X1 U2450 ( .A1(n2822), .A2(REG1_REG_3__SCAN_IN), .ZN(n2179) );
  XNOR2_X1 U2451 ( .A(n2829), .B(n2828), .ZN(n2830) );
  AND2_X1 U2452 ( .A1(n2118), .A2(n2117), .ZN(n2844) );
  NAND2_X1 U2453 ( .A1(n2836), .A2(REG1_REG_5__SCAN_IN), .ZN(n2117) );
  OR2_X1 U2454 ( .A1(n2181), .A2(n3130), .ZN(n2180) );
  XNOR2_X1 U2455 ( .A(n3934), .B(n3132), .ZN(n3133) );
  NAND2_X1 U2456 ( .A1(n3133), .A2(REG1_REG_10__SCAN_IN), .ZN(n3936) );
  XNOR2_X1 U2457 ( .A(n3970), .B(n3972), .ZN(n3958) );
  NAND2_X1 U2458 ( .A1(n3970), .A2(n4460), .ZN(n2177) );
  NAND2_X1 U2459 ( .A1(n4484), .A2(n4483), .ZN(n2176) );
  AOI21_X1 U2460 ( .B1(n2128), .B2(n2127), .A(n2053), .ZN(n2126) );
  INV_X1 U2461 ( .A(n4017), .ZN(n2127) );
  INV_X1 U2462 ( .A(n2188), .ZN(n2130) );
  NOR2_X1 U2463 ( .A1(n2268), .A2(n4062), .ZN(n2267) );
  INV_X1 U2464 ( .A(n2269), .ZN(n2268) );
  NAND2_X1 U2465 ( .A1(n2611), .A2(n2610), .ZN(n2622) );
  INV_X1 U2466 ( .A(n2612), .ZN(n2611) );
  INV_X1 U2467 ( .A(n4153), .ZN(n4117) );
  OR2_X2 U2468 ( .A1(n2592), .A2(n3567), .ZN(n2612) );
  INV_X1 U2469 ( .A(n2551), .ZN(n2549) );
  AOI21_X1 U2470 ( .B1(n2225), .B2(n2223), .A(n2012), .ZN(n2222) );
  INV_X1 U2471 ( .A(n2538), .ZN(n2223) );
  INV_X1 U2472 ( .A(n2225), .ZN(n2224) );
  AND2_X1 U2474 ( .A1(n2526), .A2(n2525), .ZN(n4294) );
  OR2_X2 U2475 ( .A1(n2494), .A2(n2493), .ZN(n2510) );
  NAND2_X1 U2476 ( .A1(n3295), .A2(n3294), .ZN(n3293) );
  AND2_X1 U2477 ( .A1(n3274), .A2(n3275), .ZN(n3779) );
  OAI21_X1 U2478 ( .B1(n3081), .B2(n3079), .A(n3827), .ZN(n3158) );
  AOI21_X1 U2479 ( .B1(n2015), .B2(n2030), .A(n2235), .ZN(n2234) );
  NOR2_X1 U2480 ( .A1(n3894), .A2(n3310), .ZN(n2235) );
  NAND2_X1 U2481 ( .A1(n3053), .A2(n2227), .ZN(n2233) );
  AND2_X1 U2482 ( .A1(n2422), .A2(n2030), .ZN(n2227) );
  OR2_X2 U2483 ( .A1(n2424), .A2(n3306), .ZN(n2435) );
  OR2_X1 U2484 ( .A1(n3094), .A2(n3898), .ZN(n2350) );
  NAND2_X1 U2485 ( .A1(n3743), .A2(n2315), .ZN(n2318) );
  NAND2_X1 U2486 ( .A1(n2316), .A2(n2792), .ZN(n2317) );
  XNOR2_X1 U2487 ( .A(n2057), .B(n4323), .ZN(n2056) );
  NAND2_X1 U2488 ( .A1(n4097), .A2(n2269), .ZN(n4058) );
  OAI21_X1 U2489 ( .B1(n2670), .B2(n2864), .A(n2863), .ZN(n3031) );
  NOR2_X1 U2490 ( .A1(n4508), .A2(n3884), .ZN(n4537) );
  NAND2_X1 U2491 ( .A1(n2738), .A2(n2723), .ZN(n2815) );
  AND2_X1 U2492 ( .A1(n2759), .A2(n4517), .ZN(n3026) );
  NOR2_X1 U2493 ( .A1(n2654), .A2(n2293), .ZN(n2295) );
  AND2_X1 U2494 ( .A1(n2295), .A2(n2656), .ZN(n2311) );
  NAND2_X1 U2495 ( .A1(n2716), .A2(IR_REG_31__SCAN_IN), .ZN(n2740) );
  OR2_X1 U2496 ( .A1(n2653), .A2(n2652), .ZN(n2282) );
  INV_X1 U2497 ( .A(n2665), .ZN(n2661) );
  INV_X1 U2498 ( .A(IR_REG_6__SCAN_IN), .ZN(n2392) );
  NOR2_X1 U2499 ( .A1(n2378), .A2(IR_REG_5__SCAN_IN), .ZN(n2393) );
  INV_X1 U2500 ( .A(n3009), .ZN(n2081) );
  INV_X1 U2501 ( .A(n2091), .ZN(n3303) );
  OAI211_X1 U2502 ( .C1(n3113), .C2(n2040), .A(n2092), .B(n2020), .ZN(n2091)
         );
  NAND2_X1 U2503 ( .A1(n2095), .A2(n3214), .ZN(n2092) );
  INV_X1 U2504 ( .A(n2248), .ZN(n3647) );
  AOI21_X1 U2505 ( .B1(n3551), .B2(n2255), .A(n2253), .ZN(n2248) );
  INV_X1 U2506 ( .A(n4171), .ZN(n4208) );
  INV_X1 U2507 ( .A(n4294), .ZN(n3889) );
  NAND4_X1 U2508 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .ZN(n3893)
         );
  NAND4_X1 U2509 ( .A1(n2418), .A2(n2417), .A3(n2416), .A4(n2415), .ZN(n3216)
         );
  NAND2_X1 U2510 ( .A1(n2305), .A2(n2017), .ZN(n2153) );
  OAI211_X1 U2511 ( .C1(n2792), .C2(n2781), .A(n3903), .B(n2145), .ZN(n3901)
         );
  NAND2_X1 U2512 ( .A1(n2792), .A2(n2781), .ZN(n2145) );
  INV_X1 U2513 ( .A(n3929), .ZN(n2136) );
  XNOR2_X1 U2514 ( .A(n3943), .B(n3132), .ZN(n3941) );
  NAND2_X1 U2515 ( .A1(n3968), .A2(n3967), .ZN(n3985) );
  XNOR2_X1 U2516 ( .A(n2483), .B(n2482), .ZN(n4009) );
  NAND2_X1 U2517 ( .A1(n4006), .A2(n4275), .ZN(n2149) );
  OR2_X1 U2518 ( .A1(n2185), .A2(n4491), .ZN(n2184) );
  AND2_X1 U2519 ( .A1(n4027), .A2(n2128), .ZN(n4491) );
  NAND2_X1 U2520 ( .A1(n2186), .A2(n4486), .ZN(n2185) );
  NAND2_X1 U2521 ( .A1(n2187), .A2(n4492), .ZN(n2186) );
  AOI21_X1 U2522 ( .B1(n4494), .B2(ADDR_REG_18__SCAN_IN), .A(n4493), .ZN(n2183) );
  INV_X1 U2523 ( .A(n4495), .ZN(n2058) );
  NAND2_X2 U2524 ( .A1(n2563), .A2(n2562), .ZN(n4034) );
  INV_X1 U2525 ( .A(n4090), .ZN(n2062) );
  INV_X1 U2526 ( .A(n2609), .ZN(n2206) );
  INV_X2 U2527 ( .A(n4559), .ZN(n4561) );
  NAND2_X1 U2528 ( .A1(n3937), .A2(n3942), .ZN(n2191) );
  OR2_X1 U2529 ( .A1(n3955), .A2(n3954), .ZN(n3956) );
  NOR2_X1 U2530 ( .A1(n2194), .A2(n2433), .ZN(n2193) );
  OR2_X1 U2531 ( .A1(n4521), .A2(n4014), .ZN(n2111) );
  NAND2_X1 U2532 ( .A1(n3778), .A2(n2365), .ZN(n2198) );
  NOR2_X1 U2533 ( .A1(n2385), .A2(n2384), .ZN(n2401) );
  NAND2_X1 U2534 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2384) );
  INV_X1 U2535 ( .A(IR_REG_28__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U2536 ( .A1(n3785), .A2(n2150), .ZN(n3786) );
  NAND2_X1 U2537 ( .A1(n2986), .A2(n2182), .ZN(n2181) );
  NAND2_X1 U2538 ( .A1(n2985), .A2(n2399), .ZN(n2182) );
  NOR2_X1 U2539 ( .A1(n2125), .A2(n2411), .ZN(n2124) );
  NAND2_X1 U2540 ( .A1(n4006), .A2(n4373), .ZN(n2188) );
  AND2_X1 U2541 ( .A1(n4013), .A2(REG1_REG_15__SCAN_IN), .ZN(n4014) );
  INV_X1 U2542 ( .A(n2210), .ZN(n2203) );
  AND2_X1 U2543 ( .A1(n4114), .A2(n4099), .ZN(n3758) );
  NAND2_X1 U2544 ( .A1(n2162), .A2(n2163), .ZN(n2161) );
  AND2_X1 U2545 ( .A1(n3732), .A2(n2160), .ZN(n2159) );
  NOR2_X1 U2546 ( .A1(n2221), .A2(n2283), .ZN(n2220) );
  OR2_X1 U2547 ( .A1(n3557), .A2(n4307), .ZN(n3723) );
  INV_X1 U2548 ( .A(n2815), .ZN(n2903) );
  NOR2_X1 U2549 ( .A1(n3543), .A2(n4055), .ZN(n2269) );
  NOR2_X1 U2550 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2659)
         );
  INV_X1 U2551 ( .A(IR_REG_21__SCAN_IN), .ZN(n2653) );
  INV_X1 U2552 ( .A(IR_REG_17__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U2553 ( .A1(n2336), .A2(n2335), .ZN(n2334) );
  OR2_X2 U2554 ( .A1(n2435), .A2(n2434), .ZN(n2447) );
  INV_X1 U2555 ( .A(n3588), .ZN(n3427) );
  INV_X1 U2556 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2412) );
  INV_X1 U2557 ( .A(n3214), .ZN(n2093) );
  NAND2_X1 U2558 ( .A1(n2940), .A2(n2939), .ZN(n3598) );
  INV_X1 U2559 ( .A(n3401), .ZN(n2254) );
  NAND2_X1 U2560 ( .A1(n3607), .A2(n3654), .ZN(n3653) );
  AOI21_X1 U2561 ( .B1(n2265), .B2(n2264), .A(n2263), .ZN(n2262) );
  INV_X1 U2562 ( .A(n3654), .ZN(n2264) );
  INV_X1 U2563 ( .A(n3605), .ZN(n2263) );
  NAND2_X1 U2564 ( .A1(n3585), .A2(n2089), .ZN(n2088) );
  NOR2_X1 U2565 ( .A1(n2266), .A2(n2090), .ZN(n2089) );
  INV_X1 U2566 ( .A(n3429), .ZN(n2090) );
  XNOR2_X1 U2567 ( .A(n2935), .B(n2934), .ZN(n2943) );
  OR2_X1 U2568 ( .A1(n2357), .A2(n2327), .ZN(n2331) );
  NAND2_X1 U2569 ( .A1(n2328), .A2(REG1_REG_1__SCAN_IN), .ZN(n2308) );
  OR2_X1 U2570 ( .A1(n2369), .A2(n2763), .ZN(n2320) );
  AND2_X1 U2571 ( .A1(n2116), .A2(REG1_REG_4__SCAN_IN), .ZN(n2114) );
  AND2_X1 U2572 ( .A1(n2829), .A2(n2113), .ZN(n2112) );
  AND2_X1 U2573 ( .A1(n2116), .A2(n4464), .ZN(n2113) );
  NAND2_X1 U2574 ( .A1(n2983), .A2(n2982), .ZN(n3125) );
  NAND2_X1 U2575 ( .A1(n2987), .A2(REG1_REG_8__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U2576 ( .A1(n3958), .A2(REG1_REG_12__SCAN_IN), .ZN(n3971) );
  OAI211_X1 U2577 ( .C1(n2177), .C2(n2122), .A(n2119), .B(n3981), .ZN(n4007)
         );
  NOR2_X1 U2578 ( .A1(n2122), .A2(n2121), .ZN(n2120) );
  AND2_X1 U2579 ( .A1(n2105), .A2(n2110), .ZN(n2104) );
  NAND2_X1 U2580 ( .A1(n4481), .A2(n4001), .ZN(n4002) );
  NAND2_X1 U2581 ( .A1(n4027), .A2(n2188), .ZN(n2187) );
  NAND2_X1 U2582 ( .A1(n2026), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U2583 ( .A1(n2211), .A2(n2620), .ZN(n2210) );
  INV_X1 U2584 ( .A(n2630), .ZN(n2211) );
  INV_X1 U2585 ( .A(n2208), .ZN(n2207) );
  OAI21_X1 U2586 ( .B1(n2630), .B2(n2209), .A(n2629), .ZN(n2208) );
  NAND2_X1 U2587 ( .A1(n2212), .A2(n2620), .ZN(n2209) );
  OR2_X1 U2588 ( .A1(n2583), .A2(n3678), .ZN(n2592) );
  AND2_X1 U2589 ( .A1(n2571), .A2(n2570), .ZN(n4187) );
  NAND2_X1 U2590 ( .A1(n2158), .A2(n2163), .ZN(n4186) );
  NAND2_X1 U2591 ( .A1(n4287), .A2(n2165), .ZN(n2158) );
  NAND2_X1 U2592 ( .A1(n4287), .A2(n2167), .ZN(n4204) );
  OR2_X1 U2593 ( .A1(n2541), .A2(n2540), .ZN(n2551) );
  NAND2_X1 U2594 ( .A1(n4287), .A2(n3851), .ZN(n4261) );
  NAND2_X1 U2595 ( .A1(n2218), .A2(n2490), .ZN(n2214) );
  OR2_X1 U2596 ( .A1(n2215), .A2(n2507), .ZN(n2213) );
  NAND2_X1 U2597 ( .A1(n2467), .A2(REG3_REG_13__SCAN_IN), .ZN(n2494) );
  AOI21_X1 U2598 ( .B1(n2157), .B2(n3780), .A(n2156), .ZN(n2155) );
  INV_X1 U2599 ( .A(n3723), .ZN(n2156) );
  NAND2_X1 U2600 ( .A1(n2684), .A2(n3843), .ZN(n3727) );
  OR2_X1 U2601 ( .A1(n2413), .A2(n2412), .ZN(n2424) );
  CLKBUF_X1 U2602 ( .A(n2996), .Z(n2997) );
  INV_X1 U2603 ( .A(n3778), .ZN(n2199) );
  INV_X1 U2604 ( .A(n3064), .ZN(n2200) );
  INV_X1 U2605 ( .A(n3094), .ZN(n3100) );
  NAND2_X1 U2606 ( .A1(n2955), .A2(n3807), .ZN(n3093) );
  INV_X1 U2607 ( .A(n4262), .ZN(n4306) );
  AND2_X1 U2608 ( .A1(n2174), .A2(n2173), .ZN(n4333) );
  AOI21_X1 U2609 ( .B1(n4079), .B2(n4266), .A(n4078), .ZN(n2173) );
  OAI21_X1 U2610 ( .B1(n4075), .B2(n2175), .A(n4304), .ZN(n2174) );
  NAND2_X1 U2611 ( .A1(n4192), .A2(n2051), .ZN(n4118) );
  NAND2_X1 U2612 ( .A1(n4192), .A2(n2024), .ZN(n4136) );
  AND2_X1 U2613 ( .A1(n4192), .A2(n4179), .ZN(n4352) );
  INV_X1 U2614 ( .A(n3659), .ZN(n4214) );
  AND2_X1 U2615 ( .A1(n4298), .A2(n2050), .ZN(n4236) );
  INV_X1 U2616 ( .A(n3420), .ZN(n4235) );
  NAND2_X1 U2617 ( .A1(n3162), .A2(n2014), .ZN(n3334) );
  NAND2_X1 U2618 ( .A1(n3162), .A2(n2013), .ZN(n3283) );
  AND2_X1 U2619 ( .A1(n3162), .A2(n3576), .ZN(n3177) );
  NOR2_X1 U2620 ( .A1(n2025), .A2(n3151), .ZN(n3150) );
  AND2_X1 U2621 ( .A1(n3150), .A2(n3250), .ZN(n3246) );
  INV_X1 U2622 ( .A(n3120), .ZN(n3250) );
  AND2_X1 U2623 ( .A1(n4212), .A2(n4529), .ZN(n4539) );
  NOR2_X1 U2624 ( .A1(n2962), .A2(n2341), .ZN(n3101) );
  INV_X1 U2625 ( .A(IR_REG_11__SCAN_IN), .ZN(n2476) );
  INV_X1 U2626 ( .A(IR_REG_7__SCAN_IN), .ZN(n2394) );
  XNOR2_X1 U2627 ( .A(n2368), .B(IR_REG_5__SCAN_IN), .ZN(n2836) );
  NOR2_X2 U2628 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2336)
         );
  AND2_X1 U2629 ( .A1(n2008), .A2(n2335), .ZN(n2281) );
  INV_X1 U2630 ( .A(n2334), .ZN(n2333) );
  OAI21_X1 U2631 ( .B1(n3113), .B2(n2097), .A(n2094), .ZN(n3213) );
  INV_X1 U2632 ( .A(n2095), .ZN(n2094) );
  AND2_X1 U2633 ( .A1(n2650), .A2(n2649), .ZN(n4066) );
  AOI21_X1 U2634 ( .B1(n3694), .B2(n3540), .A(n3539), .ZN(n3542) );
  INV_X1 U2635 ( .A(n3695), .ZN(n3539) );
  AND2_X1 U2636 ( .A1(n2640), .A2(n2632), .ZN(n4081) );
  NAND2_X1 U2637 ( .A1(n2256), .A2(n2257), .ZN(n3579) );
  INV_X1 U2638 ( .A(n2745), .ZN(n3596) );
  AND4_X1 U2639 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), .ZN(n3621)
         );
  NOR2_X1 U2640 ( .A1(n2048), .A2(n3366), .ZN(n3619) );
  NAND2_X1 U2641 ( .A1(n3044), .A2(n3043), .ZN(n3047) );
  NAND2_X1 U2642 ( .A1(n2246), .A2(n2244), .ZN(n3044) );
  AND2_X1 U2643 ( .A1(n2246), .A2(n2247), .ZN(n3017) );
  AOI21_X1 U2644 ( .B1(n3303), .B2(n3302), .A(n2261), .ZN(n3344) );
  INV_X1 U2645 ( .A(n4244), .ZN(n3688) );
  NAND2_X1 U2646 ( .A1(n2072), .A2(n2080), .ZN(n2078) );
  NAND2_X1 U2647 ( .A1(n2073), .A2(n2016), .ZN(n2072) );
  INV_X1 U2648 ( .A(n3719), .ZN(n3699) );
  INV_X1 U2649 ( .A(n3715), .ZN(n3668) );
  AOI21_X1 U2650 ( .B1(n2071), .B2(n2069), .A(n2037), .ZN(n2068) );
  INV_X1 U2651 ( .A(n2071), .ZN(n2070) );
  NAND2_X1 U2652 ( .A1(n3368), .A2(n2032), .ZN(n2075) );
  AND3_X1 U2653 ( .A1(n2516), .A2(n2515), .A3(n2514), .ZN(n4312) );
  INV_X1 U2654 ( .A(n3706), .ZN(n3713) );
  AOI21_X1 U2655 ( .B1(n2703), .B2(n2702), .A(n2701), .ZN(n3799) );
  INV_X1 U2656 ( .A(n4066), .ZN(n4079) );
  NAND2_X1 U2657 ( .A1(n2619), .A2(n2618), .ZN(n4132) );
  NAND2_X1 U2658 ( .A1(n2606), .A2(n2605), .ZN(n4153) );
  NAND2_X1 U2659 ( .A1(n2581), .A2(n2580), .ZN(n4171) );
  INV_X1 U2660 ( .A(n4187), .ZN(n4231) );
  OR2_X1 U2661 ( .A1(n2500), .A2(n2499), .ZN(n4291) );
  INV_X1 U2662 ( .A(n3621), .ZN(n3890) );
  NAND4_X1 U2663 ( .A1(n2429), .A2(n2428), .A3(n2427), .A4(n2426), .ZN(n3894)
         );
  AND2_X1 U2664 ( .A1(n2346), .A2(n2347), .ZN(n2085) );
  OR2_X1 U2665 ( .A1(n3742), .A2(n3102), .ZN(n2345) );
  OAI21_X1 U2666 ( .B1(n2792), .B2(REG2_REG_1__SCAN_IN), .A(n2144), .ZN(n3902)
         );
  NAND2_X1 U2667 ( .A1(n2792), .A2(REG2_REG_1__SCAN_IN), .ZN(n2144) );
  NAND2_X1 U2668 ( .A1(n2794), .A2(REG2_REG_2__SCAN_IN), .ZN(n2066) );
  AND2_X1 U2669 ( .A1(n2115), .A2(n2054), .ZN(n2891) );
  NAND2_X1 U2670 ( .A1(n2830), .A2(REG1_REG_4__SCAN_IN), .ZN(n2115) );
  NAND2_X1 U2671 ( .A1(n3129), .A2(n2180), .ZN(n3924) );
  NAND2_X1 U2672 ( .A1(n3924), .A2(n3923), .ZN(n3922) );
  NAND2_X1 U2673 ( .A1(n3126), .A2(n2135), .ZN(n3930) );
  NAND2_X1 U2674 ( .A1(n3123), .A2(REG2_REG_8__SCAN_IN), .ZN(n2135) );
  INV_X1 U2675 ( .A(n3945), .ZN(n2143) );
  NAND2_X1 U2676 ( .A1(n3938), .A2(n3937), .ZN(n3957) );
  NAND2_X1 U2677 ( .A1(n3936), .A2(n2195), .ZN(n3938) );
  NAND2_X1 U2678 ( .A1(n3934), .A2(n3942), .ZN(n2195) );
  NAND2_X1 U2679 ( .A1(n3971), .A2(n2177), .ZN(n3974) );
  NAND2_X1 U2680 ( .A1(n3974), .A2(n3973), .ZN(n3982) );
  XNOR2_X1 U2681 ( .A(n4007), .B(n4009), .ZN(n3983) );
  AND2_X1 U2682 ( .A1(n3999), .A2(n3998), .ZN(n2139) );
  INV_X1 U2683 ( .A(n2138), .ZN(n4473) );
  NOR2_X1 U2684 ( .A1(n4519), .A2(n2545), .ZN(n2148) );
  INV_X1 U2685 ( .A(n4025), .ZN(n2146) );
  OAI21_X1 U2686 ( .B1(n4016), .B2(n2129), .A(n2126), .ZN(n2131) );
  AND2_X1 U2687 ( .A1(n2271), .A2(n2270), .ZN(n4322) );
  OAI21_X1 U2688 ( .B1(n2064), .B2(n2224), .A(n2222), .ZN(n4222) );
  NAND2_X1 U2689 ( .A1(n2226), .A2(n2225), .ZN(n4248) );
  AND2_X1 U2690 ( .A1(n2226), .A2(n2031), .ZN(n4250) );
  NAND2_X1 U2691 ( .A1(n2064), .A2(n2538), .ZN(n2226) );
  NAND2_X1 U2692 ( .A1(n4298), .A2(n2746), .ZN(n4283) );
  NAND2_X1 U2693 ( .A1(n3293), .A2(n2490), .ZN(n4297) );
  NAND2_X1 U2694 ( .A1(n2230), .A2(n2442), .ZN(n3170) );
  NAND2_X1 U2695 ( .A1(n2233), .A2(n2234), .ZN(n3156) );
  AOI21_X1 U2696 ( .B1(n3053), .B2(n2422), .A(n2015), .ZN(n3080) );
  INV_X1 U2697 ( .A(n4316), .ZN(n4257) );
  AND2_X1 U2698 ( .A1(n4252), .A2(n4544), .ZN(n4503) );
  XNOR2_X1 U2699 ( .A(n2670), .B(n3802), .ZN(n2868) );
  AND2_X1 U2700 ( .A1(n3026), .A2(n2921), .ZN(n4510) );
  INV_X2 U2701 ( .A(n4552), .ZN(n4553) );
  INV_X1 U2702 ( .A(IR_REG_29__SCAN_IN), .ZN(n2196) );
  INV_X1 U2703 ( .A(IR_REG_30__SCAN_IN), .ZN(n3468) );
  AND2_X1 U2704 ( .A1(n2237), .A2(n4718), .ZN(n2301) );
  AND2_X1 U2705 ( .A1(n2973), .A2(STATE_REG_SCAN_IN), .ZN(n4517) );
  XNOR2_X1 U2706 ( .A(n2432), .B(IR_REG_9__SCAN_IN), .ZN(n4461) );
  OR3_X1 U2707 ( .A1(n2430), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2431) );
  NAND2_X1 U2708 ( .A1(n2103), .A2(n2102), .ZN(n2101) );
  INV_X1 U2709 ( .A(IR_REG_1__SCAN_IN), .ZN(n2103) );
  NAND2_X1 U2710 ( .A1(n3111), .A2(n3110), .ZN(n3112) );
  NAND2_X1 U2711 ( .A1(n2059), .A2(n2058), .ZN(n4499) );
  OR2_X1 U2712 ( .A1(n4409), .A2(n4395), .ZN(n2060) );
  OR2_X1 U2713 ( .A1(n4409), .A2(n4453), .ZN(n2061) );
  AND2_X1 U2714 ( .A1(n2548), .A2(n3362), .ZN(n2012) );
  INV_X1 U2715 ( .A(IR_REG_31__SCAN_IN), .ZN(n2652) );
  NAND4_X1 U2716 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n4307)
         );
  AND2_X1 U2717 ( .A1(n3576), .A2(n3357), .ZN(n2013) );
  AND2_X1 U2718 ( .A1(n2013), .A2(n3278), .ZN(n2014) );
  NOR2_X1 U2719 ( .A1(n3196), .A2(n3216), .ZN(n2015) );
  NAND2_X1 U2720 ( .A1(n2207), .A2(n2033), .ZN(n2205) );
  NAND2_X1 U2721 ( .A1(n3374), .A2(n3373), .ZN(n2016) );
  AND2_X1 U2722 ( .A1(n2306), .A2(REG0_REG_1__SCAN_IN), .ZN(n2017) );
  AND2_X1 U2723 ( .A1(n2651), .A2(n2239), .ZN(n2018) );
  AND2_X1 U2724 ( .A1(n2014), .A2(n3670), .ZN(n2019) );
  OR2_X1 U2725 ( .A1(n3195), .A2(n3194), .ZN(n2020) );
  NAND2_X1 U2726 ( .A1(n2192), .A2(n2189), .ZN(n3970) );
  AND2_X1 U2727 ( .A1(n2155), .A2(n2049), .ZN(n2021) );
  AND2_X1 U2728 ( .A1(n2656), .A2(n2196), .ZN(n2022) );
  AND2_X1 U2729 ( .A1(n4298), .A2(n2273), .ZN(n2023) );
  INV_X1 U2730 ( .A(n3362), .ZN(n2274) );
  AND2_X1 U2731 ( .A1(n2276), .A2(n4137), .ZN(n2024) );
  OR2_X1 U2732 ( .A1(n3099), .A2(n3067), .ZN(n2025) );
  NAND2_X1 U2733 ( .A1(n2074), .A2(n2078), .ZN(n3551) );
  OR2_X1 U2734 ( .A1(n2558), .A2(IR_REG_18__SCAN_IN), .ZN(n2026) );
  NAND2_X1 U2735 ( .A1(n4192), .A2(n2276), .ZN(n4135) );
  NAND2_X1 U2736 ( .A1(n4097), .A2(n4080), .ZN(n2749) );
  NAND2_X1 U2737 ( .A1(n3585), .A2(n3429), .ZN(n3607) );
  AND2_X1 U2738 ( .A1(n4244), .A2(n3420), .ZN(n2027) );
  NAND2_X1 U2739 ( .A1(n3400), .A2(n3399), .ZN(n2028) );
  OR2_X1 U2740 ( .A1(n2357), .A2(n2322), .ZN(n2029) );
  NAND2_X1 U2741 ( .A1(n3894), .A2(n3310), .ZN(n2030) );
  INV_X1 U2742 ( .A(n2369), .ZN(n2328) );
  NAND2_X1 U2743 ( .A1(n2088), .A2(n2262), .ZN(n3675) );
  NOR2_X1 U2744 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2366)
         );
  NAND2_X1 U2745 ( .A1(n3889), .A2(n3410), .ZN(n2031) );
  AND2_X1 U2746 ( .A1(n2249), .A2(n2076), .ZN(n2032) );
  OR2_X1 U2747 ( .A1(n4094), .A2(n3543), .ZN(n2033) );
  OR2_X1 U2748 ( .A1(n4132), .A2(n4113), .ZN(n2034) );
  AND2_X1 U2749 ( .A1(n3342), .A2(n3341), .ZN(n2035) );
  OR2_X1 U2750 ( .A1(n2745), .A2(n2932), .ZN(n2036) );
  AND2_X1 U2751 ( .A1(n2249), .A2(n2251), .ZN(n2037) );
  NOR2_X1 U2752 ( .A1(n4468), .A2(n4014), .ZN(n2038) );
  INV_X1 U2753 ( .A(n2205), .ZN(n2204) );
  INV_X1 U2754 ( .A(n2490), .ZN(n2217) );
  NAND2_X1 U2755 ( .A1(n3716), .A2(n3557), .ZN(n2490) );
  AND2_X1 U2756 ( .A1(n2154), .A2(n2155), .ZN(n2039) );
  INV_X1 U2757 ( .A(n3617), .ZN(n2080) );
  OR2_X1 U2758 ( .A1(n2097), .A2(n2093), .ZN(n2040) );
  OR2_X1 U2759 ( .A1(n2708), .A2(n2709), .ZN(n2041) );
  INV_X1 U2760 ( .A(n3645), .ZN(n3415) );
  INV_X1 U2761 ( .A(n2266), .ZN(n2265) );
  NAND2_X1 U2762 ( .A1(n3606), .A2(n3656), .ZN(n2266) );
  NAND2_X1 U2763 ( .A1(n3653), .A2(n3656), .ZN(n2042) );
  OR2_X1 U2764 ( .A1(n2609), .A2(n2210), .ZN(n2043) );
  INV_X1 U2765 ( .A(n3185), .ZN(n2099) );
  NAND2_X1 U2766 ( .A1(n2535), .A2(n2534), .ZN(n2558) );
  AND2_X1 U2767 ( .A1(n2257), .A2(n3349), .ZN(n2044) );
  AND2_X1 U2768 ( .A1(n4675), .A2(IR_REG_27__SCAN_IN), .ZN(n2045) );
  AND2_X1 U2769 ( .A1(n2184), .A2(n2183), .ZN(n2046) );
  INV_X1 U2770 ( .A(n2507), .ZN(n2218) );
  AND2_X1 U2771 ( .A1(n2685), .A2(n2746), .ZN(n2507) );
  INV_X1 U2772 ( .A(n2166), .ZN(n2165) );
  NAND2_X1 U2773 ( .A1(n2167), .A2(n2168), .ZN(n2166) );
  OR2_X1 U2774 ( .A1(n2224), .A2(n2027), .ZN(n2047) );
  INV_X1 U2775 ( .A(n3800), .ZN(n2695) );
  INV_X1 U2776 ( .A(n3973), .ZN(n2122) );
  NAND2_X1 U2777 ( .A1(n3169), .A2(n2453), .ZN(n3282) );
  NAND2_X1 U2778 ( .A1(n3113), .A2(n3112), .ZN(n3186) );
  INV_X1 U2779 ( .A(n3937), .ZN(n2194) );
  AND2_X1 U2780 ( .A1(n3368), .A2(n3367), .ZN(n2048) );
  INV_X1 U2781 ( .A(n3670), .ZN(n3378) );
  AND2_X1 U2782 ( .A1(n3726), .A2(n3725), .ZN(n2049) );
  NAND2_X1 U2783 ( .A1(n2230), .A2(n2228), .ZN(n3169) );
  NOR2_X1 U2784 ( .A1(n4234), .A2(n4214), .ZN(n2747) );
  AND2_X1 U2785 ( .A1(n2683), .A2(n3322), .ZN(n3843) );
  INV_X1 U2786 ( .A(n3843), .ZN(n2157) );
  NAND2_X1 U2787 ( .A1(n4298), .A2(n2272), .ZN(n2275) );
  INV_X1 U2788 ( .A(n4312), .ZN(n3648) );
  INV_X1 U2789 ( .A(n4271), .ZN(n3410) );
  AND2_X1 U2790 ( .A1(n2272), .A2(n3362), .ZN(n2050) );
  AND2_X1 U2791 ( .A1(n2878), .A2(n3881), .ZN(n4498) );
  AND2_X1 U2792 ( .A1(n2878), .A2(n2780), .ZN(n4486) );
  INV_X1 U2793 ( .A(n2016), .ZN(n2069) );
  INV_X1 U2794 ( .A(n3543), .ZN(n4080) );
  INV_X1 U2795 ( .A(n3455), .ZN(n4137) );
  AND2_X1 U2796 ( .A1(n2024), .A2(n4119), .ZN(n2051) );
  NAND2_X1 U2797 ( .A1(n3201), .A2(n3200), .ZN(n2052) );
  INV_X1 U2798 ( .A(n2129), .ZN(n2128) );
  OR2_X1 U2799 ( .A1(n4492), .A2(n2130), .ZN(n2129) );
  INV_X1 U2800 ( .A(n2285), .ZN(n2247) );
  OR2_X1 U2801 ( .A1(n4469), .A2(n2520), .ZN(n2109) );
  INV_X1 U2802 ( .A(n4029), .ZN(n4519) );
  AND2_X1 U2803 ( .A1(n4029), .A2(REG1_REG_18__SCAN_IN), .ZN(n2053) );
  NAND2_X1 U2804 ( .A1(n2829), .A2(n4464), .ZN(n2054) );
  INV_X1 U2805 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2121) );
  NAND2_X1 U2806 ( .A1(n3917), .A2(n3916), .ZN(n3915) );
  NAND2_X1 U2807 ( .A1(n2893), .A2(n2894), .ZN(n2892) );
  XNOR2_X1 U2808 ( .A(n2147), .B(n2146), .ZN(n4039) );
  INV_X1 U2809 ( .A(n2201), .ZN(n4054) );
  NAND2_X2 U2810 ( .A1(n3806), .A2(n3803), .ZN(n2670) );
  NAND2_X2 U2811 ( .A1(n2319), .A2(n3596), .ZN(n3806) );
  OAI21_X1 U2812 ( .B1(n3538), .B2(n4539), .A(n3533), .ZN(n2754) );
  INV_X1 U2813 ( .A(n2219), .ZN(n4201) );
  OAI21_X1 U2814 ( .B1(n4259), .B2(n2047), .A(n2220), .ZN(n2219) );
  NAND2_X2 U2815 ( .A1(n4126), .A2(n2607), .ZN(n2609) );
  OAI21_X1 U2816 ( .B1(n3802), .B2(n2670), .A(n3806), .ZN(n2956) );
  OAI21_X1 U2817 ( .B1(n3239), .B2(n2676), .A(n3825), .ZN(n3055) );
  INV_X1 U2818 ( .A(n3066), .ZN(n2055) );
  NOR2_X1 U2819 ( .A1(n4075), .A2(n2693), .ZN(n2694) );
  NAND4_X1 U2820 ( .A1(n4330), .A2(n4329), .A3(n4328), .A4(n4331), .ZN(n4405)
         );
  AOI21_X2 U2821 ( .B1(n2056), .B2(n4304), .A(n4067), .ZN(n4330) );
  NAND3_X2 U2822 ( .A1(n2348), .A2(n2085), .A3(n2345), .ZN(n3898) );
  INV_X1 U2823 ( .A(n4061), .ZN(n2057) );
  NAND2_X1 U2824 ( .A1(n2055), .A2(n3813), .ZN(n2170) );
  NAND2_X1 U2825 ( .A1(n2672), .A2(n3812), .ZN(n3066) );
  NAND2_X1 U2826 ( .A1(n2678), .A2(n3838), .ZN(n3277) );
  NAND2_X1 U2827 ( .A1(n2154), .A2(n2021), .ZN(n4303) );
  AOI21_X1 U2828 ( .B1(n2704), .B2(IR_REG_28__SCAN_IN), .A(n2045), .ZN(n2313)
         );
  AOI21_X2 U2829 ( .B1(n2710), .B2(n4304), .A(n2041), .ZN(n3533) );
  NAND2_X1 U2830 ( .A1(n2065), .A2(n3780), .ZN(n2154) );
  NOR2_X2 U2831 ( .A1(n3989), .A2(n2485), .ZN(n3997) );
  AOI21_X1 U2832 ( .B1(n4496), .B2(n4497), .A(n4038), .ZN(n2059) );
  NOR2_X1 U2833 ( .A1(n2336), .A2(n2008), .ZN(n2337) );
  XNOR2_X2 U2834 ( .A(n4054), .B(n4053), .ZN(n3538) );
  NAND2_X1 U2835 ( .A1(n4280), .A2(n2521), .ZN(n4259) );
  NAND2_X1 U2836 ( .A1(n4165), .A2(n4164), .ZN(n4163) );
  NAND2_X1 U2837 ( .A1(n4338), .A2(n2060), .ZN(U3544) );
  NAND2_X1 U2838 ( .A1(n4408), .A2(n2061), .ZN(U3512) );
  INV_X1 U2839 ( .A(n2684), .ZN(n2065) );
  NAND2_X2 U2840 ( .A1(n2996), .A2(n2409), .ZN(n3053) );
  NAND2_X2 U2841 ( .A1(n4289), .A2(n4288), .ZN(n4287) );
  NAND2_X1 U2842 ( .A1(n2677), .A2(n3824), .ZN(n3081) );
  NAND2_X1 U2843 ( .A1(n3158), .A2(n3839), .ZN(n2678) );
  XNOR2_X2 U2844 ( .A(n3966), .B(n3972), .ZN(n3965) );
  NOR2_X1 U2845 ( .A1(n3997), .A2(n2139), .ZN(n4474) );
  AOI21_X2 U2846 ( .B1(n3282), .B2(n2466), .A(n2465), .ZN(n3323) );
  NAND2_X1 U2847 ( .A1(n2043), .A2(n2207), .ZN(n4073) );
  NAND2_X1 U2848 ( .A1(n4333), .A2(n2171), .ZN(n4406) );
  XNOR2_X2 U2849 ( .A(n2067), .B(n3468), .ZN(n2306) );
  NAND4_X1 U2850 ( .A1(n2237), .A2(n2295), .A3(n4718), .A4(n2022), .ZN(n3467)
         );
  OAI211_X2 U2851 ( .C1(n2073), .C2(n2070), .A(n2075), .B(n2068), .ZN(n3684)
         );
  XNOR2_X1 U2852 ( .A(n3008), .B(n2081), .ZN(n3010) );
  NAND2_X1 U2853 ( .A1(n2088), .A2(n2086), .ZN(n3562) );
  INV_X1 U2854 ( .A(n3184), .ZN(n2096) );
  NOR2_X1 U2855 ( .A1(n3185), .A2(n3184), .ZN(n2097) );
  AND2_X1 U2856 ( .A1(n3112), .A2(n2099), .ZN(n2098) );
  INV_X1 U2857 ( .A(IR_REG_0__SCAN_IN), .ZN(n2102) );
  NAND3_X1 U2858 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2100) );
  NOR2_X1 U2859 ( .A1(n4470), .A2(n4469), .ZN(n4468) );
  NAND2_X1 U2860 ( .A1(n4470), .A2(n2108), .ZN(n2107) );
  OAI211_X1 U2861 ( .C1(n4470), .C2(n2109), .A(n2107), .B(n2104), .ZN(n4484)
         );
  NAND2_X1 U2862 ( .A1(n4521), .A2(n4014), .ZN(n2110) );
  AOI21_X1 U2863 ( .B1(n2830), .B2(n2114), .A(n2112), .ZN(n2118) );
  INV_X1 U2864 ( .A(n2118), .ZN(n2889) );
  NAND2_X1 U2865 ( .A1(n3958), .A2(n2120), .ZN(n2119) );
  NAND2_X1 U2866 ( .A1(n2987), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2867 ( .A1(n4016), .A2(n4017), .ZN(n4027) );
  INV_X1 U2868 ( .A(n2131), .ZN(n4031) );
  NAND2_X1 U2869 ( .A1(n2831), .A2(REG2_REG_4__SCAN_IN), .ZN(n2834) );
  NAND2_X1 U2870 ( .A1(n2821), .A2(REG2_REG_3__SCAN_IN), .ZN(n2132) );
  OAI21_X2 U2871 ( .B1(n3123), .B2(n2134), .A(n2133), .ZN(n3928) );
  AOI21_X2 U2872 ( .B1(n3126), .B2(n3232), .A(n2136), .ZN(n2133) );
  INV_X1 U2873 ( .A(n3126), .ZN(n2134) );
  NAND2_X2 U2874 ( .A1(n3928), .A2(n3128), .ZN(n3943) );
  XNOR2_X2 U2875 ( .A(n4000), .B(n2520), .ZN(n4482) );
  AND2_X2 U2876 ( .A1(n2138), .A2(n2137), .ZN(n4000) );
  OR2_X2 U2877 ( .A1(n4474), .A2(n4475), .ZN(n2138) );
  INV_X1 U2878 ( .A(n3944), .ZN(n2141) );
  NAND2_X1 U2879 ( .A1(n2142), .A2(n3944), .ZN(n3946) );
  NAND2_X1 U2880 ( .A1(n3941), .A2(REG2_REG_10__SCAN_IN), .ZN(n2142) );
  NAND2_X2 U2881 ( .A1(n3953), .A2(n3952), .ZN(n3966) );
  OAI21_X2 U2882 ( .B1(n3985), .B2(n3984), .A(n3988), .ZN(n3996) );
  NAND2_X2 U2883 ( .A1(n2306), .A2(n2305), .ZN(n2357) );
  OAI21_X2 U2884 ( .B1(n4287), .B2(n2161), .A(n2159), .ZN(n4128) );
  NAND3_X1 U2885 ( .A1(n2162), .A2(n2163), .A3(n2166), .ZN(n2160) );
  NOR2_X2 U2886 ( .A1(n4077), .A2(n4076), .ZN(n4075) );
  NAND2_X1 U2888 ( .A1(n2337), .A2(IR_REG_2__SCAN_IN), .ZN(n2338) );
  NAND2_X1 U2889 ( .A1(n2176), .A2(n4015), .ZN(n4016) );
  OAI21_X1 U2890 ( .B1(n4484), .B2(n4483), .A(n2176), .ZN(n4485) );
  NAND2_X1 U2891 ( .A1(n3133), .A2(n2193), .ZN(n2192) );
  AND2_X2 U2892 ( .A1(n2863), .A2(n2326), .ZN(n2954) );
  NAND2_X1 U2893 ( .A1(n2670), .A2(n2864), .ZN(n2863) );
  NAND2_X1 U2894 ( .A1(n2325), .A2(n2745), .ZN(n3803) );
  NAND2_X1 U2895 ( .A1(n2301), .A2(n2311), .ZN(n2302) );
  NAND2_X1 U2896 ( .A1(n3064), .A2(n2365), .ZN(n2197) );
  NAND3_X1 U2897 ( .A1(n2197), .A2(n2198), .A3(n2375), .ZN(n2377) );
  NAND2_X1 U2898 ( .A1(n3063), .A2(n2365), .ZN(n3143) );
  NAND2_X1 U2899 ( .A1(n2200), .A2(n2199), .ZN(n3063) );
  NAND2_X1 U2900 ( .A1(n2609), .A2(n2608), .ZN(n4107) );
  OAI21_X2 U2901 ( .B1(n3295), .B2(n2214), .A(n2213), .ZN(n4282) );
  INV_X1 U2902 ( .A(n3597), .ZN(n2941) );
  XNOR2_X1 U2903 ( .A(n2943), .B(n2942), .ZN(n3597) );
  OAI21_X2 U2904 ( .B1(n3472), .B2(n3489), .A(n3471), .ZN(n3477) );
  AND2_X2 U2905 ( .A1(n3565), .A2(n3451), .ZN(n3472) );
  NAND2_X1 U2906 ( .A1(n3011), .A2(n3010), .ZN(n2246) );
  NAND3_X2 U2907 ( .A1(n2242), .A2(n3046), .A3(n2240), .ZN(n3113) );
  NAND2_X1 U2908 ( .A1(n2241), .A2(n3043), .ZN(n2240) );
  INV_X1 U2909 ( .A(n2244), .ZN(n2241) );
  NAND2_X1 U2910 ( .A1(n3011), .A2(n2243), .ZN(n2242) );
  AND2_X1 U2911 ( .A1(n3010), .A2(n3043), .ZN(n2243) );
  INV_X1 U2912 ( .A(n3016), .ZN(n2245) );
  NOR2_X2 U2913 ( .A1(n2285), .A2(n2245), .ZN(n2244) );
  NAND2_X1 U2914 ( .A1(n2256), .A2(n2044), .ZN(n3577) );
  NAND2_X1 U2915 ( .A1(n4097), .A2(n2267), .ZN(n2271) );
  INV_X1 U2916 ( .A(n2271), .ZN(n4057) );
  NAND2_X1 U2917 ( .A1(n4058), .A2(n4062), .ZN(n2270) );
  INV_X1 U2918 ( .A(n2275), .ZN(n4270) );
  INV_X1 U2919 ( .A(n3011), .ZN(n2972) );
  OR2_X1 U2920 ( .A1(n4034), .A2(n2812), .ZN(n4508) );
  INV_X1 U2921 ( .A(n4034), .ZN(n4459) );
  NAND2_X1 U2922 ( .A1(n2666), .A2(n2665), .ZN(n3874) );
  NOR2_X1 U2923 ( .A1(n2712), .A2(n2659), .ZN(n2660) );
  AND2_X1 U2924 ( .A1(n2967), .A2(n2968), .ZN(n2969) );
  NAND2_X1 U2925 ( .A1(n4236), .A2(n4235), .ZN(n4234) );
  OAI22_X1 U2926 ( .A1(n3508), .A2(n2928), .B1(n2932), .B2(n2927), .ZN(n2929)
         );
  NAND2_X1 U2927 ( .A1(n3246), .A2(n3245), .ZN(n3244) );
  NAND2_X1 U2928 ( .A1(n2306), .A2(n4456), .ZN(n2369) );
  NAND2_X1 U2929 ( .A1(n2871), .A2(n2745), .ZN(n2962) );
  OAI21_X1 U2930 ( .B1(n3684), .B2(n3417), .A(n3686), .ZN(n3418) );
  NAND2_X1 U2931 ( .A1(n4054), .A2(n4053), .ZN(n4327) );
  OR2_X1 U2932 ( .A1(n2759), .A2(n2763), .ZN(n2278) );
  OR2_X1 U2933 ( .A1(n3352), .A2(n3351), .ZN(n2279) );
  AND2_X1 U2934 ( .A1(n2589), .A2(n2588), .ZN(n4151) );
  INV_X1 U2935 ( .A(n4151), .ZN(n4189) );
  OR2_X1 U2936 ( .A1(n3925), .A2(n3131), .ZN(n2280) );
  AND2_X1 U2937 ( .A1(n3688), .A2(n4235), .ZN(n2283) );
  AND2_X1 U2938 ( .A1(n4208), .A2(n4194), .ZN(n2284) );
  AND2_X1 U2939 ( .A1(n3009), .A2(n3008), .ZN(n2285) );
  INV_X1 U2940 ( .A(n4099), .ZN(n2748) );
  AND2_X2 U2941 ( .A1(n3028), .A2(n4299), .ZN(n4515) );
  INV_X1 U2942 ( .A(IR_REG_2__SCAN_IN), .ZN(n2335) );
  INV_X1 U2943 ( .A(n2590), .ZN(n4179) );
  OR2_X1 U2944 ( .A1(n3530), .A2(n4453), .ZN(n2286) );
  OR2_X1 U2945 ( .A1(n3530), .A2(n4395), .ZN(n2287) );
  AND2_X1 U2946 ( .A1(n3414), .A2(n3413), .ZN(n2288) );
  INV_X1 U2947 ( .A(IR_REG_9__SCAN_IN), .ZN(n4689) );
  INV_X1 U2948 ( .A(IR_REG_26__SCAN_IN), .ZN(n2292) );
  NAND2_X1 U2949 ( .A1(n2671), .A2(n2007), .ZN(n2762) );
  AND2_X1 U2950 ( .A1(n3759), .A2(n4087), .ZN(n3862) );
  OR2_X1 U2951 ( .A1(n2686), .A2(n4224), .ZN(n3854) );
  NOR2_X1 U2952 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2294)
         );
  INV_X1 U2953 ( .A(n3580), .ZN(n3349) );
  NAND2_X1 U2954 ( .A1(n2938), .A2(n2934), .ZN(n2939) );
  INV_X1 U2955 ( .A(n3742), .ZN(n2643) );
  INV_X1 U2956 ( .A(n2575), .ZN(n2573) );
  INV_X1 U2957 ( .A(n3942), .ZN(n3132) );
  INV_X1 U2958 ( .A(n2622), .ZN(n2621) );
  INV_X1 U2959 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2434) );
  INV_X1 U2960 ( .A(n2927), .ZN(n2341) );
  OR2_X1 U2961 ( .A1(n2501), .A2(IR_REG_14__SCAN_IN), .ZN(n2502) );
  AND2_X1 U2962 ( .A1(n3386), .A2(n3385), .ZN(n3396) );
  AND2_X1 U2963 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  INV_X1 U2964 ( .A(n3041), .ZN(n3042) );
  INV_X1 U2965 ( .A(n2469), .ZN(n2467) );
  NAND2_X1 U2966 ( .A1(n2573), .A2(REG3_REG_21__SCAN_IN), .ZN(n2583) );
  OR2_X1 U2967 ( .A1(n3987), .A2(n4390), .ZN(n3981) );
  NAND2_X1 U2968 ( .A1(n4074), .A2(n4099), .ZN(n2629) );
  NAND2_X1 U2969 ( .A1(n2621), .A2(REG3_REG_26__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U2970 ( .A1(n4189), .A2(n2590), .ZN(n2591) );
  INV_X1 U2971 ( .A(n4305), .ZN(n2746) );
  NAND2_X1 U2972 ( .A1(n2751), .A2(n2812), .ZN(n4262) );
  INV_X1 U2973 ( .A(n3557), .ZN(n3384) );
  INV_X1 U2974 ( .A(n4263), .ZN(n4308) );
  INV_X1 U2975 ( .A(IR_REG_24__SCAN_IN), .ZN(n2718) );
  OR2_X1 U2976 ( .A1(n2631), .A2(n3545), .ZN(n2640) );
  INV_X1 U2977 ( .A(n3348), .ZN(n3576) );
  INV_X1 U2978 ( .A(n4290), .ZN(n3640) );
  NAND2_X1 U2979 ( .A1(n2509), .A2(REG3_REG_16__SCAN_IN), .ZN(n2541) );
  AND2_X1 U2980 ( .A1(n3380), .A2(n3379), .ZN(n3664) );
  INV_X1 U2981 ( .A(n3667), .ZN(n3717) );
  OR2_X1 U2982 ( .A1(n4102), .A2(n2642), .ZN(n2628) );
  OR2_X1 U2983 ( .A1(n2360), .A2(n2398), .ZN(n2407) );
  INV_X1 U2984 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3306) );
  INV_X1 U2985 ( .A(n4311), .ZN(n4266) );
  INV_X1 U2986 ( .A(n4304), .ZN(n4268) );
  INV_X1 U2987 ( .A(IR_REG_23__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U2988 ( .A1(n2401), .A2(REG3_REG_7__SCAN_IN), .ZN(n2413) );
  INV_X1 U2989 ( .A(n4158), .ZN(n3570) );
  OAI21_X1 U2990 ( .B1(n3685), .B2(n3419), .A(n3418), .ZN(n3587) );
  AND2_X1 U2991 ( .A1(n2622), .A2(n2613), .ZN(n4121) );
  INV_X1 U2992 ( .A(n3073), .ZN(n3067) );
  NAND2_X1 U2993 ( .A1(n2922), .A2(n4299), .ZN(n3719) );
  NAND2_X1 U2994 ( .A1(n2977), .A2(n2976), .ZN(n3703) );
  NAND2_X1 U2995 ( .A1(n2637), .A2(n2636), .ZN(n4094) );
  OAI211_X1 U2996 ( .C1(n3742), .C2(n2545), .A(n2544), .B(n2543), .ZN(n4265)
         );
  OR2_X1 U2997 ( .A1(n2646), .A2(n2433), .ZN(n2439) );
  OR2_X1 U2998 ( .A1(n2642), .A2(REG3_REG_3__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U2999 ( .A1(n3983), .A2(REG1_REG_14__SCAN_IN), .ZN(n4008) );
  AND2_X1 U3000 ( .A1(n2773), .A2(n2772), .ZN(n2878) );
  AND2_X1 U3001 ( .A1(n4313), .A2(n4034), .ZN(n4252) );
  NAND2_X1 U3002 ( .A1(n3878), .A2(n2696), .ZN(n4304) );
  AND2_X1 U3003 ( .A1(n4313), .A2(n3030), .ZN(n4512) );
  NAND2_X1 U3004 ( .A1(n2724), .A2(n2816), .ZN(n3025) );
  INV_X1 U3005 ( .A(n4539), .ZN(n4547) );
  INV_X1 U3006 ( .A(n3025), .ZN(n2904) );
  AND2_X1 U3007 ( .A1(n2506), .A2(n2517), .ZN(n4013) );
  NAND2_X1 U3008 ( .A1(n2419), .A2(n2396), .ZN(n2985) );
  AND2_X1 U3009 ( .A1(n2774), .A2(n2773), .ZN(n4494) );
  NAND2_X1 U3010 ( .A1(n2907), .A2(n4467), .ZN(n3715) );
  OR2_X1 U3011 ( .A1(n2919), .A2(n2917), .ZN(n3706) );
  INV_X1 U3012 ( .A(n3703), .ZN(n3722) );
  INV_X1 U3013 ( .A(n4074), .ZN(n4114) );
  NAND2_X1 U3014 ( .A1(n2557), .A2(n2556), .ZN(n4244) );
  INV_X1 U3015 ( .A(n4486), .ZN(n4490) );
  NAND2_X1 U3016 ( .A1(n4313), .A2(n3141), .ZN(n4316) );
  INV_X1 U3017 ( .A(n4503), .ZN(n4272) );
  NAND2_X1 U3018 ( .A1(n4561), .A2(n4544), .ZN(n4395) );
  OR2_X1 U3019 ( .A1(n3025), .A2(n2753), .ZN(n4559) );
  NAND2_X1 U3020 ( .A1(n4553), .A2(n4544), .ZN(n4453) );
  OR2_X1 U3021 ( .A1(n2904), .A2(n2753), .ZN(n4552) );
  INV_X1 U3022 ( .A(n4562), .ZN(n4516) );
  NAND2_X1 U3023 ( .A1(n2815), .A2(n3026), .ZN(n4562) );
  INV_X1 U3024 ( .A(n2735), .ZN(n4458) );
  XNOR2_X1 U3025 ( .A(n2519), .B(n2518), .ZN(n4521) );
  NOR2_X2 U3026 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2529)
         );
  NAND4_X1 U3027 ( .A1(n2529), .A2(n2291), .A3(n2290), .A4(n2289), .ZN(n2654)
         );
  NAND4_X1 U3028 ( .A1(n2713), .A2(n2711), .A3(n2292), .A4(n4688), .ZN(n2293)
         );
  XNOR2_X2 U3031 ( .A(n2303), .B(IR_REG_29__SCAN_IN), .ZN(n4456) );
  NAND2_X2 U3032 ( .A1(n4455), .A2(n2305), .ZN(n2360) );
  INV_X1 U3033 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2781) );
  OR2_X1 U3034 ( .A1(n2360), .A2(n2781), .ZN(n2310) );
  INV_X1 U3035 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2304) );
  OR2_X1 U3036 ( .A1(n2344), .A2(n2304), .ZN(n2309) );
  INV_X1 U3037 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2307) );
  INV_X1 U3038 ( .A(n2325), .ZN(n2319) );
  NAND2_X1 U3039 ( .A1(n2311), .A2(n2658), .ZN(n2312) );
  INV_X1 U3040 ( .A(DATAI_1_), .ZN(n2315) );
  INV_X1 U3041 ( .A(n3743), .ZN(n2316) );
  INV_X1 U3042 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2881) );
  INV_X1 U3043 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2763) );
  AND2_X1 U3044 ( .A1(n2321), .A2(n2320), .ZN(n2324) );
  INV_X1 U3045 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2322) );
  INV_X1 U3046 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2758) );
  OR2_X1 U3047 ( .A1(n2360), .A2(n2758), .ZN(n2323) );
  NAND3_X2 U3048 ( .A1(n2324), .A2(n2029), .A3(n2323), .ZN(n2671) );
  MUX2_X1 U3049 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2009), .Z(n2923) );
  NAND2_X1 U3050 ( .A1(n2325), .A2(n3596), .ZN(n2326) );
  INV_X1 U3051 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4674) );
  OR2_X1 U3052 ( .A1(n2344), .A2(n4674), .ZN(n2332) );
  INV_X1 U3053 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2327) );
  NAND2_X1 U3054 ( .A1(n2328), .A2(REG1_REG_2__SCAN_IN), .ZN(n2330) );
  INV_X1 U3055 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2783) );
  OR2_X1 U3056 ( .A1(n2360), .A2(n2783), .ZN(n2329) );
  INV_X1 U3057 ( .A(DATAI_2_), .ZN(n2340) );
  MUX2_X1 U3058 ( .A(n2794), .B(n2340), .S(n2010), .Z(n2927) );
  NAND2_X1 U3059 ( .A1(n3594), .A2(n2927), .ZN(n3810) );
  OR2_X1 U3060 ( .A1(n2341), .A2(n3594), .ZN(n2342) );
  NAND2_X1 U3061 ( .A1(n2952), .A2(n2342), .ZN(n3092) );
  NAND2_X1 U3062 ( .A1(n3739), .A2(REG1_REG_3__SCAN_IN), .ZN(n2348) );
  INV_X1 U3063 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2343) );
  OR2_X1 U3064 ( .A1(n2357), .A2(n2343), .ZN(n2347) );
  INV_X1 U3065 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3102) );
  OR2_X1 U3066 ( .A1(n2367), .A2(n2652), .ZN(n2353) );
  XNOR2_X2 U3067 ( .A(n2353), .B(IR_REG_3__SCAN_IN), .ZN(n4465) );
  MUX2_X1 U3068 ( .A(n4465), .B(DATAI_3_), .S(n2010), .Z(n3094) );
  NAND2_X1 U3069 ( .A1(n3898), .A2(n3094), .ZN(n2349) );
  NAND2_X1 U3070 ( .A1(n3092), .A2(n2349), .ZN(n2351) );
  NAND2_X1 U3071 ( .A1(n2351), .A2(n2350), .ZN(n3064) );
  INV_X1 U3072 ( .A(IR_REG_3__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3073 ( .A1(n2353), .A2(n2352), .ZN(n2354) );
  NAND2_X1 U3074 ( .A1(n2354), .A2(IR_REG_31__SCAN_IN), .ZN(n2355) );
  INV_X1 U3075 ( .A(IR_REG_4__SCAN_IN), .ZN(n4710) );
  XNOR2_X1 U3076 ( .A(n2355), .B(n4710), .ZN(n2828) );
  INV_X1 U3077 ( .A(DATAI_4_), .ZN(n2356) );
  MUX2_X1 U3078 ( .A(n2828), .B(n2356), .S(n2009), .Z(n3073) );
  NAND2_X1 U3079 ( .A1(n3739), .A2(REG1_REG_4__SCAN_IN), .ZN(n2364) );
  INV_X1 U3080 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2358) );
  OR2_X1 U3081 ( .A1(n2357), .A2(n2358), .ZN(n2363) );
  OAI21_X1 U3082 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2385), .ZN(n3075) );
  OR2_X1 U3083 ( .A1(n2642), .A2(n3075), .ZN(n2362) );
  INV_X1 U3084 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2359) );
  OR2_X1 U3085 ( .A1(n3742), .A2(n2359), .ZN(n2361) );
  OR2_X1 U3086 ( .A1(n3073), .A2(n3897), .ZN(n3813) );
  NAND2_X1 U3087 ( .A1(n3897), .A2(n3073), .ZN(n3815) );
  NAND2_X1 U3088 ( .A1(n3897), .A2(n3067), .ZN(n2365) );
  NAND2_X1 U3089 ( .A1(n2367), .A2(n2366), .ZN(n2378) );
  NAND2_X1 U3090 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2368) );
  MUX2_X1 U3091 ( .A(n2836), .B(DATAI_5_), .S(n2010), .Z(n3151) );
  NAND2_X1 U3092 ( .A1(n2697), .A2(REG0_REG_5__SCAN_IN), .ZN(n2374) );
  INV_X1 U3093 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2370) );
  OR2_X1 U3094 ( .A1(n2646), .A2(n2370), .ZN(n2373) );
  INV_X1 U3095 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2383) );
  XNOR2_X1 U3096 ( .A(n2385), .B(n2383), .ZN(n3152) );
  OR2_X1 U3097 ( .A1(n2642), .A2(n3152), .ZN(n2372) );
  INV_X1 U3098 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2835) );
  OR2_X1 U3099 ( .A1(n3742), .A2(n2835), .ZN(n2371) );
  NAND4_X1 U3100 ( .A1(n2374), .A2(n2373), .A3(n2372), .A4(n2371), .ZN(n3896)
         );
  OR2_X1 U3101 ( .A1(n3151), .A2(n3896), .ZN(n2375) );
  NAND2_X1 U3102 ( .A1(n3896), .A2(n3151), .ZN(n2376) );
  NAND2_X1 U3103 ( .A1(n2377), .A2(n2376), .ZN(n2996) );
  INV_X1 U3104 ( .A(n2393), .ZN(n2379) );
  NAND2_X1 U3105 ( .A1(n2379), .A2(IR_REG_31__SCAN_IN), .ZN(n2380) );
  XNOR2_X1 U3106 ( .A(n2380), .B(IR_REG_6__SCAN_IN), .ZN(n4463) );
  MUX2_X1 U3107 ( .A(n4463), .B(DATAI_6_), .S(n2010), .Z(n3120) );
  NAND2_X1 U3108 ( .A1(n3739), .A2(REG1_REG_6__SCAN_IN), .ZN(n2391) );
  INV_X1 U3109 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2381) );
  OR2_X1 U3110 ( .A1(n2357), .A2(n2381), .ZN(n2390) );
  INV_X1 U3111 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2382) );
  OAI21_X1 U3112 ( .B1(n2385), .B2(n2383), .A(n2382), .ZN(n2386) );
  INV_X1 U3113 ( .A(n2401), .ZN(n2402) );
  NAND2_X1 U3114 ( .A1(n2386), .A2(n2402), .ZN(n3266) );
  OR2_X1 U3115 ( .A1(n2642), .A2(n3266), .ZN(n2389) );
  INV_X1 U3116 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2387) );
  OR2_X1 U3117 ( .A1(n3742), .A2(n2387), .ZN(n2388) );
  NAND4_X1 U3118 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n3895)
         );
  NAND2_X1 U3119 ( .A1(n2393), .A2(n2392), .ZN(n2430) );
  NAND2_X1 U3120 ( .A1(n2430), .A2(IR_REG_31__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3121 ( .A1(n2395), .A2(n2394), .ZN(n2419) );
  OR2_X1 U3122 ( .A1(n2395), .A2(n2394), .ZN(n2396) );
  INV_X1 U3123 ( .A(DATAI_7_), .ZN(n2397) );
  MUX2_X1 U3124 ( .A(n2985), .B(n2397), .S(n2009), .Z(n3245) );
  INV_X1 U3125 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2398) );
  INV_X1 U3126 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2399) );
  OR2_X1 U3127 ( .A1(n2646), .A2(n2399), .ZN(n2406) );
  INV_X1 U3128 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2400) );
  OR2_X1 U3129 ( .A1(n2357), .A2(n2400), .ZN(n2405) );
  INV_X1 U3130 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U3131 ( .A1(n2402), .A2(n4563), .ZN(n2403) );
  NAND2_X1 U3132 ( .A1(n2413), .A2(n2403), .ZN(n3247) );
  OR2_X1 U3133 ( .A1(n2642), .A2(n3247), .ZN(n2404) );
  NAND4_X1 U3134 ( .A1(n2407), .A2(n2406), .A3(n2405), .A4(n2404), .ZN(n3205)
         );
  OR2_X1 U3135 ( .A1(n3245), .A2(n3205), .ZN(n2675) );
  OAI21_X1 U3136 ( .B1(n3120), .B2(n3895), .A(n3820), .ZN(n2408) );
  INV_X1 U3137 ( .A(n2408), .ZN(n2409) );
  AND2_X1 U3138 ( .A1(n3895), .A2(n3120), .ZN(n2410) );
  INV_X1 U3139 ( .A(n3245), .ZN(n3240) );
  AOI22_X1 U3140 ( .A1(n3820), .A2(n2410), .B1(n3240), .B2(n3205), .ZN(n3052)
         );
  NAND2_X1 U3141 ( .A1(n2697), .A2(REG0_REG_8__SCAN_IN), .ZN(n2418) );
  INV_X1 U3142 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2411) );
  OR2_X1 U3143 ( .A1(n2646), .A2(n2411), .ZN(n2417) );
  NAND2_X1 U3144 ( .A1(n2413), .A2(n2412), .ZN(n2414) );
  NAND2_X1 U3145 ( .A1(n2424), .A2(n2414), .ZN(n3231) );
  OR2_X1 U3146 ( .A1(n2642), .A2(n3231), .ZN(n2416) );
  INV_X1 U3147 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3232) );
  OR2_X1 U31480 ( .A1(n3742), .A2(n3232), .ZN(n2415) );
  NAND2_X1 U31490 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2420) );
  XNOR2_X1 U3150 ( .A(n2420), .B(IR_REG_8__SCAN_IN), .ZN(n3124) );
  MUX2_X1 U3151 ( .A(n3124), .B(DATAI_8_), .S(n2009), .Z(n3196) );
  NAND2_X1 U3152 ( .A1(n3216), .A2(n3196), .ZN(n2421) );
  AND2_X1 U3153 ( .A1(n3052), .A2(n2421), .ZN(n2422) );
  NAND2_X1 U3154 ( .A1(n3739), .A2(REG1_REG_9__SCAN_IN), .ZN(n2429) );
  INV_X1 U3155 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2423) );
  OR2_X1 U3156 ( .A1(n2357), .A2(n2423), .ZN(n2428) );
  NAND2_X1 U3157 ( .A1(n2424), .A2(n3306), .ZN(n2425) );
  NAND2_X1 U3158 ( .A1(n2435), .A2(n2425), .ZN(n3313) );
  OR2_X1 U3159 ( .A1(n2642), .A2(n3313), .ZN(n2427) );
  INV_X1 U3160 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3127) );
  OR2_X1 U3161 ( .A1(n3742), .A2(n3127), .ZN(n2426) );
  NAND2_X1 U3162 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  MUX2_X1 U3163 ( .A(n4461), .B(DATAI_9_), .S(n2009), .Z(n3310) );
  NAND2_X1 U3164 ( .A1(n2697), .A2(REG0_REG_10__SCAN_IN), .ZN(n2440) );
  INV_X1 U3165 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3166 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  NAND2_X1 U3167 ( .A1(n2447), .A2(n2436), .ZN(n3573) );
  OR2_X1 U3168 ( .A1(n2642), .A2(n3573), .ZN(n2438) );
  INV_X1 U3169 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3223) );
  OR2_X1 U3170 ( .A1(n3742), .A2(n3223), .ZN(n2437) );
  OR2_X1 U3171 ( .A1(n2658), .A2(n2652), .ZN(n2441) );
  XNOR2_X1 U3172 ( .A(n2441), .B(IR_REG_10__SCAN_IN), .ZN(n3942) );
  MUX2_X1 U3173 ( .A(n3942), .B(DATAI_10_), .S(n2010), .Z(n3348) );
  NOR2_X1 U3174 ( .A1(n3893), .A2(n3348), .ZN(n2443) );
  NAND2_X1 U3175 ( .A1(n3893), .A2(n3348), .ZN(n2442) );
  INV_X1 U3176 ( .A(IR_REG_10__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3177 ( .A1(n2658), .A2(n2444), .ZN(n2478) );
  NAND2_X1 U3178 ( .A1(n2478), .A2(IR_REG_31__SCAN_IN), .ZN(n2462) );
  XNOR2_X1 U3179 ( .A(n2462), .B(n2476), .ZN(n3955) );
  INV_X1 U3180 ( .A(DATAI_11_), .ZN(n2445) );
  MUX2_X1 U3181 ( .A(n3955), .B(n2445), .S(n2009), .Z(n3357) );
  NAND2_X1 U3182 ( .A1(n2697), .A2(REG0_REG_11__SCAN_IN), .ZN(n2452) );
  INV_X1 U3183 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3954) );
  OR2_X1 U3184 ( .A1(n2646), .A2(n3954), .ZN(n2451) );
  INV_X1 U3185 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U3186 ( .A1(n2447), .A2(n4564), .ZN(n2448) );
  NAND2_X1 U3187 ( .A1(n2455), .A2(n2448), .ZN(n3179) );
  OR2_X1 U3188 ( .A1(n2642), .A2(n3179), .ZN(n2450) );
  INV_X1 U3189 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3951) );
  OR2_X1 U3190 ( .A1(n3742), .A2(n3951), .ZN(n2449) );
  NAND4_X1 U3191 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n3892)
         );
  OR2_X1 U3192 ( .A1(n3357), .A2(n3892), .ZN(n3274) );
  NAND2_X1 U3193 ( .A1(n3892), .A2(n3357), .ZN(n3275) );
  INV_X1 U3194 ( .A(n3357), .ZN(n3353) );
  OR2_X1 U3195 ( .A1(n3353), .A2(n3892), .ZN(n2453) );
  NAND2_X1 U3196 ( .A1(n3739), .A2(REG1_REG_12__SCAN_IN), .ZN(n2461) );
  INV_X1 U3197 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4451) );
  OR2_X1 U3198 ( .A1(n2357), .A2(n4451), .ZN(n2460) );
  NAND2_X1 U3199 ( .A1(n2455), .A2(n2454), .ZN(n2456) );
  NAND2_X1 U3200 ( .A1(n2469), .A2(n2456), .ZN(n3627) );
  OR2_X1 U3201 ( .A1(n2642), .A2(n3627), .ZN(n2459) );
  INV_X1 U3202 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2457) );
  OR2_X1 U3203 ( .A1(n3742), .A2(n2457), .ZN(n2458) );
  NAND4_X1 U3204 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3891)
         );
  NAND2_X1 U3205 ( .A1(n2462), .A2(n2476), .ZN(n2463) );
  NAND2_X1 U3206 ( .A1(n2463), .A2(IR_REG_31__SCAN_IN), .ZN(n2464) );
  XNOR2_X1 U3207 ( .A(n2464), .B(IR_REG_12__SCAN_IN), .ZN(n4460) );
  MUX2_X1 U3208 ( .A(n4460), .B(DATAI_12_), .S(n2010), .Z(n3624) );
  NAND2_X1 U3209 ( .A1(n3891), .A2(n3624), .ZN(n2466) );
  NOR2_X1 U32100 ( .A1(n3891), .A2(n3624), .ZN(n2465) );
  NAND2_X1 U32110 ( .A1(n3739), .A2(REG1_REG_13__SCAN_IN), .ZN(n2474) );
  INV_X1 U32120 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4447) );
  OR2_X1 U32130 ( .A1(n2357), .A2(n4447), .ZN(n2473) );
  INV_X1 U32140 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U32150 ( .A1(n2469), .A2(n2468), .ZN(n2470) );
  NAND2_X1 U32160 ( .A1(n2494), .A2(n2470), .ZN(n3337) );
  OR2_X1 U32170 ( .A1(n2642), .A2(n3337), .ZN(n2472) );
  INV_X1 U32180 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3986) );
  OR2_X1 U32190 ( .A1(n3742), .A2(n3986), .ZN(n2471) );
  INV_X1 U32200 ( .A(IR_REG_12__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U32210 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  OAI21_X1 U32220 ( .B1(n2478), .B2(n2477), .A(IR_REG_31__SCAN_IN), .ZN(n2479)
         );
  XNOR2_X1 U32230 ( .A(n2479), .B(n2527), .ZN(n3987) );
  INV_X1 U32240 ( .A(DATAI_13_), .ZN(n2480) );
  MUX2_X1 U32250 ( .A(n3987), .B(n2480), .S(n2010), .Z(n3670) );
  NAND2_X1 U32260 ( .A1(n3621), .A2(n3670), .ZN(n2481) );
  NAND2_X1 U32270 ( .A1(n2658), .A2(n2656), .ZN(n2501) );
  NAND2_X1 U32280 ( .A1(n2501), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  INV_X1 U32290 ( .A(IR_REG_14__SCAN_IN), .ZN(n2482) );
  INV_X1 U32300 ( .A(DATAI_14_), .ZN(n2484) );
  MUX2_X1 U32310 ( .A(n4009), .B(n2484), .S(n2009), .Z(n3557) );
  XNOR2_X1 U32320 ( .A(n2494), .B(REG3_REG_14__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U32330 ( .A1(n2702), .A2(n3559), .ZN(n2489) );
  INV_X1 U32340 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4443) );
  OR2_X1 U32350 ( .A1(n2357), .A2(n4443), .ZN(n2488) );
  INV_X1 U32360 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4385) );
  OR2_X1 U32370 ( .A1(n2646), .A2(n4385), .ZN(n2487) );
  INV_X1 U32380 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2485) );
  OR2_X1 U32390 ( .A1(n3742), .A2(n2485), .ZN(n2486) );
  NAND2_X1 U32400 ( .A1(n4307), .A2(n3557), .ZN(n3724) );
  NAND2_X1 U32410 ( .A1(n3723), .A2(n3724), .ZN(n3294) );
  INV_X1 U32420 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2492) );
  INV_X1 U32430 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2491) );
  OAI21_X1 U32440 ( .B1(n2494), .B2(n2492), .A(n2491), .ZN(n2495) );
  NAND2_X1 U32450 ( .A1(REG3_REG_15__SCAN_IN), .A2(REG3_REG_14__SCAN_IN), .ZN(
        n2493) );
  NAND2_X1 U32460 ( .A1(n2495), .A2(n2510), .ZN(n4300) );
  INV_X1 U32470 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4301) );
  OR2_X1 U32480 ( .A1(n3742), .A2(n4301), .ZN(n2496) );
  OAI21_X1 U32490 ( .B1(n4300), .B2(n2642), .A(n2496), .ZN(n2500) );
  NAND2_X1 U32500 ( .A1(n2697), .A2(REG0_REG_15__SCAN_IN), .ZN(n2498) );
  INV_X1 U32510 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4012) );
  OR2_X1 U32520 ( .A1(n2646), .A2(n4012), .ZN(n2497) );
  NAND2_X1 U32530 ( .A1(n2498), .A2(n2497), .ZN(n2499) );
  NAND2_X1 U32540 ( .A1(n2502), .A2(IR_REG_31__SCAN_IN), .ZN(n2505) );
  INV_X1 U32550 ( .A(n2505), .ZN(n2503) );
  NAND2_X1 U32560 ( .A1(n2503), .A2(IR_REG_15__SCAN_IN), .ZN(n2506) );
  INV_X1 U32570 ( .A(IR_REG_15__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U32580 ( .A1(n2505), .A2(n2504), .ZN(n2517) );
  MUX2_X1 U32590 ( .A(n4013), .B(DATAI_15_), .S(n2010), .Z(n4305) );
  NAND2_X1 U32600 ( .A1(n4291), .A2(n4305), .ZN(n2508) );
  INV_X1 U32610 ( .A(n4291), .ZN(n2685) );
  INV_X1 U32620 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U32630 ( .A1(n2510), .A2(n4578), .ZN(n2511) );
  NAND2_X1 U32640 ( .A1(n2541), .A2(n2511), .ZN(n4284) );
  OR2_X1 U32650 ( .A1(n4284), .A2(n2642), .ZN(n2516) );
  INV_X1 U32660 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4483) );
  OR2_X1 U32670 ( .A1(n2646), .A2(n4483), .ZN(n2513) );
  INV_X1 U32680 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4667) );
  OR2_X1 U32690 ( .A1(n2357), .A2(n4667), .ZN(n2512) );
  AND2_X1 U32700 ( .A1(n2513), .A2(n2512), .ZN(n2515) );
  INV_X1 U32710 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4285) );
  OR2_X1 U32720 ( .A1(n3742), .A2(n4285), .ZN(n2514) );
  NAND2_X1 U32730 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2519) );
  INV_X1 U32740 ( .A(IR_REG_16__SCAN_IN), .ZN(n2518) );
  INV_X1 U32750 ( .A(n4521), .ZN(n2520) );
  MUX2_X1 U32760 ( .A(n2520), .B(DATAI_16_), .S(n2010), .Z(n4290) );
  NAND2_X1 U32770 ( .A1(n4312), .A2(n4290), .ZN(n3849) );
  NAND2_X1 U32780 ( .A1(n3648), .A2(n3640), .ZN(n3851) );
  NAND2_X1 U32790 ( .A1(n3849), .A2(n3851), .ZN(n4281) );
  XNOR2_X1 U32800 ( .A(n2541), .B(REG3_REG_17__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U32810 ( .A1(n4273), .A2(n2702), .ZN(n2526) );
  INV_X1 U32820 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U32830 ( .A1(n2697), .A2(REG0_REG_17__SCAN_IN), .ZN(n2523) );
  INV_X1 U32840 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4373) );
  OR2_X1 U32850 ( .A1(n2646), .A2(n4373), .ZN(n2522) );
  OAI211_X1 U32860 ( .C1(n4275), .C2(n3742), .A(n2523), .B(n2522), .ZN(n2524)
         );
  INV_X1 U32870 ( .A(n2524), .ZN(n2525) );
  NOR2_X1 U32880 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2528) );
  AND4_X1 U32890 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n2531)
         );
  NAND2_X1 U32900 ( .A1(n2658), .A2(n2531), .ZN(n2533) );
  NAND2_X1 U32910 ( .A1(n2533), .A2(IR_REG_31__SCAN_IN), .ZN(n2532) );
  MUX2_X1 U32920 ( .A(IR_REG_31__SCAN_IN), .B(n2532), .S(IR_REG_17__SCAN_IN), 
        .Z(n2536) );
  INV_X1 U32930 ( .A(n2533), .ZN(n2535) );
  NAND2_X1 U32940 ( .A1(n2536), .A2(n2558), .ZN(n4006) );
  INV_X1 U32950 ( .A(DATAI_17_), .ZN(n2537) );
  MUX2_X1 U32960 ( .A(n4006), .B(n2537), .S(n2009), .Z(n4271) );
  NAND2_X1 U32970 ( .A1(n4294), .A2(n4271), .ZN(n2538) );
  INV_X1 U32980 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2545) );
  INV_X1 U32990 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4668) );
  INV_X1 U33000 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2539) );
  OAI21_X1 U33010 ( .B1(n2541), .B2(n4668), .A(n2539), .ZN(n2542) );
  NAND2_X1 U33020 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2540) );
  AND2_X1 U33030 ( .A1(n2542), .A2(n2551), .ZN(n4253) );
  NAND2_X1 U33040 ( .A1(n4253), .A2(n2702), .ZN(n2544) );
  AOI22_X1 U33050 ( .A1(n3739), .A2(REG1_REG_18__SCAN_IN), .B1(n2697), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U33060 ( .A1(n2558), .A2(IR_REG_31__SCAN_IN), .ZN(n2546) );
  XNOR2_X1 U33070 ( .A(n2546), .B(IR_REG_18__SCAN_IN), .ZN(n4029) );
  INV_X1 U33080 ( .A(DATAI_18_), .ZN(n2547) );
  MUX2_X1 U33090 ( .A(n4519), .B(n2547), .S(n2009), .Z(n3362) );
  OR2_X1 U33100 ( .A1(n4265), .A2(n3362), .ZN(n4225) );
  NAND2_X1 U33110 ( .A1(n4265), .A2(n3362), .ZN(n4226) );
  NAND2_X1 U33120 ( .A1(n4225), .A2(n4226), .ZN(n4249) );
  INV_X1 U33130 ( .A(n4265), .ZN(n2548) );
  INV_X1 U33140 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U33150 ( .A1(n2551), .A2(n2550), .ZN(n2552) );
  NAND2_X1 U33160 ( .A1(n2564), .A2(n2552), .ZN(n4237) );
  OR2_X1 U33170 ( .A1(n4237), .A2(n2642), .ZN(n2557) );
  INV_X1 U33180 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U33190 ( .A1(n3739), .A2(REG1_REG_19__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U33200 ( .A1(n2697), .A2(REG0_REG_19__SCAN_IN), .ZN(n2553) );
  OAI211_X1 U33210 ( .C1(n4238), .C2(n3742), .A(n2554), .B(n2553), .ZN(n2555)
         );
  INV_X1 U33220 ( .A(n2555), .ZN(n2556) );
  INV_X1 U33230 ( .A(IR_REG_19__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U33240 ( .A1(n2560), .A2(n2559), .ZN(n2563) );
  INV_X1 U33250 ( .A(n2560), .ZN(n2561) );
  NAND2_X1 U33260 ( .A1(n2561), .A2(IR_REG_19__SCAN_IN), .ZN(n2562) );
  MUX2_X1 U33270 ( .A(n4459), .B(DATAI_19_), .S(n2010), .Z(n3420) );
  INV_X1 U33280 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3658) );
  NAND2_X1 U33290 ( .A1(n2564), .A2(n3658), .ZN(n2565) );
  AND2_X1 U33300 ( .A1(n2575), .A2(n2565), .ZN(n4217) );
  NAND2_X1 U33310 ( .A1(n4217), .A2(n2702), .ZN(n2571) );
  INV_X1 U33320 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U33330 ( .A1(n3739), .A2(REG1_REG_20__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U33340 ( .A1(n2697), .A2(REG0_REG_20__SCAN_IN), .ZN(n2566) );
  OAI211_X1 U33350 ( .C1(n2568), .C2(n3742), .A(n2567), .B(n2566), .ZN(n2569)
         );
  INV_X1 U33360 ( .A(n2569), .ZN(n2570) );
  NAND2_X1 U33370 ( .A1(n2009), .A2(DATAI_20_), .ZN(n3659) );
  NAND2_X1 U33380 ( .A1(n4187), .A2(n3659), .ZN(n2572) );
  INV_X1 U33390 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33400 ( .A1(n2575), .A2(n2574), .ZN(n2576) );
  NAND2_X1 U33410 ( .A1(n2583), .A2(n2576), .ZN(n3612) );
  OR2_X1 U33420 ( .A1(n3612), .A2(n2642), .ZN(n2581) );
  INV_X1 U33430 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U33440 ( .A1(n2643), .A2(REG2_REG_21__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U33450 ( .A1(n2697), .A2(REG0_REG_21__SCAN_IN), .ZN(n2577) );
  OAI211_X1 U33460 ( .C1(n2646), .C2(n4680), .A(n2578), .B(n2577), .ZN(n2579)
         );
  INV_X1 U33470 ( .A(n2579), .ZN(n2580) );
  AND2_X1 U33480 ( .A1(n2010), .A2(DATAI_21_), .ZN(n3611) );
  NAND2_X1 U33490 ( .A1(n4171), .A2(n3611), .ZN(n2582) );
  INV_X1 U33500 ( .A(n3611), .ZN(n4194) );
  INV_X1 U33510 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U33520 ( .A1(n2583), .A2(n3678), .ZN(n2584) );
  NAND2_X1 U3353 ( .A1(n2592), .A2(n2584), .ZN(n4177) );
  OR2_X1 U33540 ( .A1(n4177), .A2(n2642), .ZN(n2589) );
  INV_X1 U3355 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4176) );
  NAND2_X1 U3356 ( .A1(n2697), .A2(REG0_REG_22__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U3357 ( .A1(n3739), .A2(REG1_REG_22__SCAN_IN), .ZN(n2585) );
  OAI211_X1 U3358 ( .C1(n4176), .C2(n3742), .A(n2586), .B(n2585), .ZN(n2587)
         );
  INV_X1 U3359 ( .A(n2587), .ZN(n2588) );
  AND2_X1 U3360 ( .A1(n2009), .A2(DATAI_22_), .ZN(n2590) );
  NAND2_X1 U3361 ( .A1(n4151), .A2(n2590), .ZN(n4148) );
  NAND2_X1 U3362 ( .A1(n4189), .A2(n4179), .ZN(n2691) );
  NAND2_X1 U3363 ( .A1(n4148), .A2(n2691), .ZN(n4164) );
  INV_X1 U3364 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U3365 ( .A1(n2592), .A2(n3567), .ZN(n2593) );
  NAND2_X1 U3366 ( .A1(n2612), .A2(n2593), .ZN(n4158) );
  NAND2_X1 U3367 ( .A1(n3570), .A2(n2702), .ZN(n2598) );
  INV_X1 U3368 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4157) );
  NAND2_X1 U3369 ( .A1(n3739), .A2(REG1_REG_23__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U3370 ( .A1(n2697), .A2(REG0_REG_23__SCAN_IN), .ZN(n2594) );
  OAI211_X1 U3371 ( .C1(n4157), .C2(n3742), .A(n2595), .B(n2594), .ZN(n2596)
         );
  INV_X1 U3372 ( .A(n2596), .ZN(n2597) );
  AND2_X2 U3373 ( .A1(n2598), .A2(n2597), .ZN(n4173) );
  NAND2_X1 U3374 ( .A1(n2010), .A2(DATAI_23_), .ZN(n4156) );
  NAND2_X1 U3375 ( .A1(n4173), .A2(n4156), .ZN(n2600) );
  NOR2_X1 U3376 ( .A1(n4173), .A2(n4156), .ZN(n2599) );
  XNOR2_X1 U3377 ( .A(n2612), .B(REG3_REG_24__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U3378 ( .A1(n4139), .A2(n2702), .ZN(n2606) );
  INV_X1 U3379 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3380 ( .A1(n3739), .A2(REG1_REG_24__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3381 ( .A1(n2697), .A2(REG0_REG_24__SCAN_IN), .ZN(n2601) );
  OAI211_X1 U3382 ( .C1(n2603), .C2(n3742), .A(n2602), .B(n2601), .ZN(n2604)
         );
  INV_X1 U3383 ( .A(n2604), .ZN(n2605) );
  AND2_X1 U3384 ( .A1(n2010), .A2(DATAI_24_), .ZN(n3455) );
  NAND2_X1 U3385 ( .A1(n4153), .A2(n3455), .ZN(n2607) );
  NAND2_X1 U3386 ( .A1(n4117), .A2(n4137), .ZN(n2608) );
  AND2_X1 U3387 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .ZN(
        n2610) );
  INV_X1 U3388 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3462) );
  INV_X1 U3389 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3479) );
  OAI21_X1 U3390 ( .B1(n2612), .B2(n3462), .A(n3479), .ZN(n2613) );
  NAND2_X1 U3391 ( .A1(n4121), .A2(n2702), .ZN(n2619) );
  INV_X1 U3392 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U3393 ( .A1(n3739), .A2(REG1_REG_25__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U3394 ( .A1(n2697), .A2(REG0_REG_25__SCAN_IN), .ZN(n2614) );
  OAI211_X1 U3395 ( .C1(n2616), .C2(n3742), .A(n2615), .B(n2614), .ZN(n2617)
         );
  INV_X1 U3396 ( .A(n2617), .ZN(n2618) );
  AND2_X1 U3397 ( .A1(n2009), .A2(DATAI_25_), .ZN(n4113) );
  NAND2_X1 U3398 ( .A1(n4132), .A2(n4113), .ZN(n2620) );
  INV_X1 U3399 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U3400 ( .A1(n2622), .A2(n4705), .ZN(n2623) );
  NAND2_X1 U3401 ( .A1(n2631), .A2(n2623), .ZN(n4102) );
  INV_X1 U3402 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U3403 ( .A1(n3739), .A2(REG1_REG_26__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3404 ( .A1(n2643), .A2(REG2_REG_26__SCAN_IN), .ZN(n2624) );
  OAI211_X1 U3405 ( .C1(n2357), .C2(n4679), .A(n2625), .B(n2624), .ZN(n2626)
         );
  INV_X1 U3406 ( .A(n2626), .ZN(n2627) );
  AND2_X2 U3407 ( .A1(n2628), .A2(n2627), .ZN(n4074) );
  NAND2_X1 U3408 ( .A1(n2009), .A2(DATAI_26_), .ZN(n4099) );
  NOR2_X1 U3409 ( .A1(n4074), .A2(n4099), .ZN(n2630) );
  INV_X1 U3410 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3545) );
  NAND2_X1 U3411 ( .A1(n2631), .A2(n3545), .ZN(n2632) );
  NAND2_X1 U3412 ( .A1(n4081), .A2(n2702), .ZN(n2637) );
  INV_X1 U3413 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U3414 ( .A1(n2643), .A2(REG2_REG_27__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3415 ( .A1(n2697), .A2(REG0_REG_27__SCAN_IN), .ZN(n2633) );
  OAI211_X1 U3416 ( .C1(n2646), .C2(n4575), .A(n2634), .B(n2633), .ZN(n2635)
         );
  INV_X1 U3417 ( .A(n2635), .ZN(n2636) );
  AND2_X1 U3418 ( .A1(n2010), .A2(DATAI_27_), .ZN(n3543) );
  NAND2_X1 U3419 ( .A1(n4094), .A2(n3543), .ZN(n2638) );
  INV_X1 U3420 ( .A(n2640), .ZN(n2639) );
  NAND2_X1 U3421 ( .A1(n2639), .A2(REG3_REG_28__SCAN_IN), .ZN(n4068) );
  INV_X1 U3422 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U3423 ( .A1(n2640), .A2(n3518), .ZN(n2641) );
  NAND2_X1 U3424 ( .A1(n4068), .A2(n2641), .ZN(n3532) );
  OR2_X1 U3425 ( .A1(n3532), .A2(n2642), .ZN(n2650) );
  INV_X1 U3426 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3427 ( .A1(n2643), .A2(REG2_REG_28__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3428 ( .A1(n2697), .A2(REG0_REG_28__SCAN_IN), .ZN(n2644) );
  OAI211_X1 U3429 ( .C1(n2647), .C2(n2646), .A(n2645), .B(n2644), .ZN(n2648)
         );
  INV_X1 U3430 ( .A(n2648), .ZN(n2649) );
  AND2_X1 U3431 ( .A1(n2010), .A2(DATAI_28_), .ZN(n4055) );
  NAND2_X1 U3432 ( .A1(n4066), .A2(n4055), .ZN(n3736) );
  INV_X1 U3433 ( .A(n4055), .ZN(n3519) );
  NAND2_X1 U3434 ( .A1(n4079), .A2(n3519), .ZN(n4059) );
  NAND2_X1 U3435 ( .A1(n3736), .A2(n4059), .ZN(n4053) );
  NOR2_X1 U3436 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2651)
         );
  INV_X1 U3437 ( .A(n2654), .ZN(n2655) );
  AND2_X1 U3438 ( .A1(n2656), .A2(n2655), .ZN(n2657) );
  INV_X1 U3439 ( .A(n2712), .ZN(n2667) );
  NAND2_X1 U3440 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2662) );
  AOI22_X1 U3441 ( .A1(IR_REG_20__SCAN_IN), .A2(n2652), .B1(n2662), .B2(
        IR_REG_31__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3442 ( .A1(n2667), .A2(IR_REG_31__SCAN_IN), .ZN(n2668) );
  XNOR2_X1 U3443 ( .A(n2760), .B(n3884), .ZN(n2669) );
  NAND2_X1 U3444 ( .A1(n2669), .A2(n4034), .ZN(n4212) );
  INV_X1 U3445 ( .A(n3874), .ZN(n2812) );
  INV_X1 U3446 ( .A(n4537), .ZN(n4529) );
  INV_X2 U3447 ( .A(n2923), .ZN(n2871) );
  INV_X1 U3448 ( .A(n2953), .ZN(n3782) );
  NAND2_X1 U3449 ( .A1(n2956), .A2(n3782), .ZN(n2955) );
  NAND2_X1 U3450 ( .A1(n3898), .A2(n3100), .ZN(n3809) );
  NAND2_X1 U3451 ( .A1(n3093), .A2(n3781), .ZN(n2672) );
  INV_X1 U3452 ( .A(n3151), .ZN(n2673) );
  AND2_X1 U3453 ( .A1(n3896), .A2(n2673), .ZN(n3816) );
  OR2_X1 U3454 ( .A1(n2673), .A2(n3896), .ZN(n3830) );
  NAND2_X1 U3455 ( .A1(n3895), .A2(n3250), .ZN(n3831) );
  NAND2_X1 U3456 ( .A1(n2998), .A2(n3831), .ZN(n2674) );
  OR2_X1 U3457 ( .A1(n3250), .A2(n3895), .ZN(n3819) );
  NAND2_X1 U34580 ( .A1(n2674), .A2(n3819), .ZN(n3239) );
  INV_X1 U34590 ( .A(n2675), .ZN(n2676) );
  INV_X1 U3460 ( .A(n3196), .ZN(n3208) );
  OR2_X1 U3461 ( .A1(n3208), .A2(n3216), .ZN(n3826) );
  NAND2_X1 U3462 ( .A1(n3055), .A2(n3826), .ZN(n2677) );
  NAND2_X1 U3463 ( .A1(n3216), .A2(n3208), .ZN(n3824) );
  INV_X1 U3464 ( .A(n3310), .ZN(n3082) );
  AND2_X1 U3465 ( .A1(n3894), .A2(n3082), .ZN(n3079) );
  OR2_X1 U3466 ( .A1(n3082), .A2(n3894), .ZN(n3827) );
  NAND2_X1 U34670 ( .A1(n3893), .A2(n3576), .ZN(n3839) );
  OR2_X1 U3468 ( .A1(n3576), .A2(n3893), .ZN(n3838) );
  INV_X1 U34690 ( .A(n3624), .ZN(n3278) );
  NAND2_X1 U3470 ( .A1(n3891), .A2(n3278), .ZN(n3324) );
  NAND2_X1 U34710 ( .A1(n3890), .A2(n3670), .ZN(n3321) );
  NAND2_X1 U3472 ( .A1(n3324), .A2(n3321), .ZN(n2680) );
  INV_X1 U34730 ( .A(n3275), .ZN(n2679) );
  NOR2_X1 U3474 ( .A1(n2680), .A2(n2679), .ZN(n3840) );
  NAND2_X1 U34750 ( .A1(n3277), .A2(n3840), .ZN(n2684) );
  INV_X1 U3476 ( .A(n2680), .ZN(n2682) );
  OR2_X1 U34770 ( .A1(n3278), .A2(n3891), .ZN(n3326) );
  NAND2_X1 U3478 ( .A1(n3326), .A2(n3274), .ZN(n2681) );
  NAND2_X1 U34790 ( .A1(n2682), .A2(n2681), .ZN(n2683) );
  NAND2_X1 U3480 ( .A1(n3621), .A2(n3378), .ZN(n3322) );
  INV_X1 U34810 ( .A(n3294), .ZN(n3780) );
  NAND2_X1 U3482 ( .A1(n2685), .A2(n4305), .ZN(n3726) );
  NAND2_X1 U34830 ( .A1(n4291), .A2(n2746), .ZN(n3725) );
  NAND2_X1 U3484 ( .A1(n4303), .A2(n3725), .ZN(n4289) );
  INV_X1 U34850 ( .A(n4281), .ZN(n4288) );
  NAND2_X1 U3486 ( .A1(n4244), .A2(n4235), .ZN(n3769) );
  NAND2_X1 U34870 ( .A1(n3769), .A2(n4226), .ZN(n2686) );
  AND2_X1 U3488 ( .A1(n3889), .A2(n4271), .ZN(n4224) );
  INV_X1 U34890 ( .A(n2686), .ZN(n2688) );
  OR2_X1 U3490 ( .A1(n3889), .A2(n4271), .ZN(n4223) );
  NAND2_X1 U34910 ( .A1(n4225), .A2(n4223), .ZN(n2687) );
  NAND2_X1 U3492 ( .A1(n2688), .A2(n2687), .ZN(n2689) );
  NAND2_X1 U34930 ( .A1(n3688), .A2(n3420), .ZN(n3770) );
  NAND2_X1 U3494 ( .A1(n2689), .A2(n3770), .ZN(n4202) );
  NOR2_X1 U34950 ( .A1(n4231), .A2(n3659), .ZN(n2690) );
  NOR2_X1 U3496 ( .A1(n4202), .A2(n2690), .ZN(n3853) );
  AND2_X1 U34970 ( .A1(n4231), .A2(n3659), .ZN(n3856) );
  NAND2_X1 U3498 ( .A1(n4208), .A2(n3611), .ZN(n4146) );
  NAND2_X1 U34990 ( .A1(n4148), .A2(n4146), .ZN(n3858) );
  AND2_X1 U3500 ( .A1(n4171), .A2(n4194), .ZN(n3857) );
  INV_X1 U35010 ( .A(n4173), .ZN(n3888) );
  NAND2_X1 U3502 ( .A1(n3888), .A2(n4156), .ZN(n3791) );
  NAND2_X1 U35030 ( .A1(n3791), .A2(n2691), .ZN(n3863) );
  AOI21_X1 U3504 ( .B1(n3857), .B2(n4148), .A(n3863), .ZN(n3732) );
  NOR2_X1 U35050 ( .A1(n4153), .A2(n4137), .ZN(n3794) );
  NOR2_X1 U35060 ( .A1(n3888), .A2(n4156), .ZN(n3790) );
  NOR2_X1 U35070 ( .A1(n3794), .A2(n3790), .ZN(n3861) );
  NAND2_X1 U35080 ( .A1(n4074), .A2(n2748), .ZN(n3759) );
  NAND2_X1 U35090 ( .A1(n4092), .A2(n4113), .ZN(n4087) );
  INV_X1 U35100 ( .A(n3862), .ZN(n2692) );
  INV_X1 U35110 ( .A(n4113), .ZN(n4119) );
  NAND2_X1 U35120 ( .A1(n4132), .A2(n4119), .ZN(n3789) );
  NAND2_X1 U35130 ( .A1(n4153), .A2(n4137), .ZN(n4108) );
  NAND2_X1 U35140 ( .A1(n3789), .A2(n4108), .ZN(n4088) );
  AOI21_X1 U35150 ( .B1(n3862), .B2(n4088), .A(n3758), .ZN(n3867) );
  NAND2_X1 U35160 ( .A1(n3700), .A2(n3543), .ZN(n3735) );
  NAND2_X1 U35170 ( .A1(n4094), .A2(n4080), .ZN(n3865) );
  INV_X1 U35180 ( .A(n3735), .ZN(n2693) );
  XNOR2_X1 U35190 ( .A(n2694), .B(n4053), .ZN(n2710) );
  NAND2_X1 U35200 ( .A1(n2695), .A2(n2812), .ZN(n3878) );
  NAND2_X1 U35210 ( .A1(n4459), .A2(n3884), .ZN(n2696) );
  INV_X1 U35220 ( .A(n4068), .ZN(n2703) );
  INV_X1 U35230 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U35240 ( .A1(n2697), .A2(REG0_REG_29__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U35250 ( .A1(n3739), .A2(REG1_REG_29__SCAN_IN), .ZN(n2698) );
  OAI211_X1 U35260 ( .C1(n2700), .C2(n3742), .A(n2699), .B(n2698), .ZN(n2701)
         );
  NAND2_X1 U35270 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(
        n2705) );
  NAND2_X1 U35280 ( .A1(n2704), .A2(n2705), .ZN(n2706) );
  XNOR2_X1 U35290 ( .A(n2706), .B(IR_REG_28__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U35300 ( .A1(n2908), .A2(n4467), .ZN(n4311) );
  NOR2_X1 U35310 ( .A1(n3799), .A2(n4311), .ZN(n2709) );
  INV_X1 U35320 ( .A(n4467), .ZN(n2768) );
  NAND2_X1 U35330 ( .A1(n2908), .A2(n2768), .ZN(n4263) );
  INV_X1 U35340 ( .A(n3884), .ZN(n2707) );
  OAI22_X1 U35350 ( .A1(n3700), .A2(n4263), .B1(n3519), .B2(n4262), .ZN(n2708)
         );
  NAND2_X1 U35360 ( .A1(n2712), .A2(n2711), .ZN(n2716) );
  INV_X1 U35370 ( .A(n2716), .ZN(n2714) );
  NAND2_X1 U35380 ( .A1(n2714), .A2(n2713), .ZN(n2720) );
  NAND2_X1 U35390 ( .A1(n2740), .A2(n2739), .ZN(n2717) );
  NAND2_X1 U35400 ( .A1(n2736), .A2(n2735), .ZN(n2722) );
  MUX2_X1 U35410 ( .A(n2736), .B(n2722), .S(B_REG_SCAN_IN), .Z(n2723) );
  INV_X1 U35420 ( .A(D_REG_0__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U35430 ( .A1(n2903), .A2(n2818), .ZN(n2724) );
  INV_X1 U35440 ( .A(n2738), .ZN(n2734) );
  NAND2_X1 U35450 ( .A1(n2734), .A2(n2736), .ZN(n2816) );
  NOR4_X1 U35460 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U35470 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .ZN(n2727)
         );
  NOR4_X1 U35480 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2726) );
  NOR4_X1 U35490 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2725) );
  NAND4_X1 U35500 ( .A1(n4709), .A2(n2727), .A3(n2726), .A4(n2725), .ZN(n2733)
         );
  NOR4_X1 U35510 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2731) );
  NOR4_X1 U35520 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2730) );
  NOR4_X1 U35530 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2729) );
  NOR4_X1 U35540 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2728) );
  NAND4_X1 U35550 ( .A1(n2731), .A2(n2730), .A3(n2729), .A4(n2728), .ZN(n2732)
         );
  NOR2_X1 U35560 ( .A1(n2733), .A2(n2732), .ZN(n2900) );
  NAND2_X1 U35570 ( .A1(n2734), .A2(n2735), .ZN(n2819) );
  OAI21_X1 U35580 ( .B1(n2815), .B2(D_REG_1__SCAN_IN), .A(n2819), .ZN(n2743)
         );
  INV_X1 U35590 ( .A(n2736), .ZN(n2737) );
  XNOR2_X1 U35600 ( .A(n2740), .B(n2739), .ZN(n2973) );
  NAND2_X1 U35610 ( .A1(n4537), .A2(n3800), .ZN(n2920) );
  NAND2_X1 U35620 ( .A1(n4034), .A2(n3874), .ZN(n2741) );
  NAND2_X1 U35630 ( .A1(n2908), .A2(n2741), .ZN(n3024) );
  AND3_X1 U35640 ( .A1(n3026), .A2(n2920), .A3(n3024), .ZN(n2742) );
  OAI211_X1 U35650 ( .C1(n2900), .C2(n2815), .A(n2743), .B(n2742), .ZN(n2753)
         );
  INV_X1 U35660 ( .A(n2744), .ZN(n2752) );
  NAND2_X1 U35670 ( .A1(n3101), .A2(n3100), .ZN(n3099) );
  NOR2_X4 U35680 ( .A1(n3336), .A2(n3384), .ZN(n4298) );
  INV_X1 U35690 ( .A(n2747), .ZN(n4216) );
  NOR2_X4 U35700 ( .A1(n4216), .A2(n3611), .ZN(n4192) );
  NAND2_X1 U35710 ( .A1(n2749), .A2(n4055), .ZN(n2750) );
  NAND2_X1 U35720 ( .A1(n4058), .A2(n2750), .ZN(n3530) );
  NAND2_X1 U35730 ( .A1(n2752), .A2(n2287), .ZN(U3546) );
  INV_X1 U35740 ( .A(n2755), .ZN(n2756) );
  NAND2_X1 U35750 ( .A1(n2756), .A2(n2286), .ZN(U3514) );
  INV_X1 U35760 ( .A(n4517), .ZN(n2757) );
  OR2_X2 U35770 ( .A1(n2759), .A2(n2757), .ZN(n3899) );
  INV_X2 U35780 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  XNOR2_X1 U35790 ( .A(n2704), .B(IR_REG_27__SCAN_IN), .ZN(n4457) );
  AOI21_X1 U35800 ( .B1(n4457), .B2(n2758), .A(n4467), .ZN(n2879) );
  AND2_X1 U35810 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3903) );
  INV_X1 U3582 ( .A(n4457), .ZN(n2780) );
  NAND2_X2 U3583 ( .A1(n2760), .A2(n2759), .ZN(n2932) );
  NAND2_X1 U3584 ( .A1(n3456), .A2(n2923), .ZN(n2761) );
  AND2_X1 U3585 ( .A1(n2762), .A2(n2761), .ZN(n2938) );
  NAND2_X1 U3586 ( .A1(n2938), .A2(n2278), .ZN(n2937) );
  INV_X1 U3587 ( .A(n2937), .ZN(n2767) );
  NAND2_X1 U3588 ( .A1(n2971), .A2(n2671), .ZN(n2766) );
  INV_X1 U3589 ( .A(n2759), .ZN(n2764) );
  AOI22_X1 U3590 ( .A1(n2007), .A2(n2923), .B1(IR_REG_0__SCAN_IN), .B2(n2764), 
        .ZN(n2765) );
  NAND2_X1 U3591 ( .A1(n2766), .A2(n2765), .ZN(n2936) );
  XNOR2_X1 U3592 ( .A(n2767), .B(n2936), .ZN(n2924) );
  NAND2_X1 U3593 ( .A1(n2924), .A2(n2780), .ZN(n2769) );
  OAI211_X1 U3594 ( .C1(n3903), .C2(n2780), .A(n2769), .B(n2768), .ZN(n2770)
         );
  OAI211_X1 U3595 ( .C1(IR_REG_0__SCAN_IN), .C2(n2879), .A(n2770), .B(U4043), 
        .ZN(n3921) );
  INV_X1 U3596 ( .A(n3921), .ZN(n2791) );
  OR2_X1 U3597 ( .A1(n2973), .A2(U3149), .ZN(n3886) );
  INV_X1 U3598 ( .A(n3886), .ZN(n2771) );
  OR2_X1 U3599 ( .A1(n3026), .A2(n2771), .ZN(n2773) );
  AOI21_X1 U3600 ( .B1(n2908), .B2(n2973), .A(n2316), .ZN(n2772) );
  NAND2_X1 U3601 ( .A1(n2878), .A2(n4467), .ZN(n4500) );
  INV_X1 U3602 ( .A(n2772), .ZN(n2774) );
  NAND2_X1 U3603 ( .A1(n4494), .A2(ADDR_REG_4__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3604 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3018) );
  OAI211_X1 U3605 ( .C1(n2828), .C2(n4500), .A(n2775), .B(n3018), .ZN(n2790)
         );
  XNOR2_X1 U3606 ( .A(n2794), .B(REG1_REG_2__SCAN_IN), .ZN(n3911) );
  XNOR2_X1 U3607 ( .A(n2792), .B(REG1_REG_1__SCAN_IN), .ZN(n3904) );
  AND2_X1 U3608 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3905)
         );
  NAND2_X1 U3609 ( .A1(n3904), .A2(n3905), .ZN(n2777) );
  INV_X1 U3610 ( .A(n2792), .ZN(n3900) );
  NAND2_X1 U3611 ( .A1(n3900), .A2(REG1_REG_1__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3612 ( .A1(n2777), .A2(n2776), .ZN(n3912) );
  INV_X1 U3613 ( .A(n2794), .ZN(n3914) );
  AOI22_X1 U3614 ( .A1(n3911), .A2(n3912), .B1(n3914), .B2(REG1_REG_2__SCAN_IN), .ZN(n2778) );
  XNOR2_X1 U3615 ( .A(n2778), .B(n4465), .ZN(n2822) );
  INV_X1 U3616 ( .A(n2778), .ZN(n2779) );
  XNOR2_X1 U3617 ( .A(n2830), .B(REG1_REG_4__SCAN_IN), .ZN(n2788) );
  NOR2_X1 U3618 ( .A1(n4467), .A2(n2780), .ZN(n3881) );
  INV_X1 U3619 ( .A(n4498), .ZN(n4038) );
  NAND2_X1 U3620 ( .A1(n3900), .A2(REG2_REG_1__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U3621 ( .A1(n3901), .A2(n2782), .ZN(n3916) );
  OR2_X1 U3622 ( .A1(n2794), .A2(n2783), .ZN(n2784) );
  INV_X1 U3623 ( .A(n4465), .ZN(n2827) );
  NAND2_X1 U3624 ( .A1(n2785), .A2(n4465), .ZN(n2786) );
  XNOR2_X1 U3625 ( .A(n2831), .B(REG2_REG_4__SCAN_IN), .ZN(n2787) );
  OAI22_X1 U3626 ( .A1(n2788), .A2(n4490), .B1(n4038), .B2(n2787), .ZN(n2789)
         );
  OR3_X1 U3627 ( .A1(n2791), .A2(n2790), .A3(n2789), .ZN(U3244) );
  MUX2_X1 U3628 ( .A(n2792), .B(n2315), .S(U3149), .Z(n2793) );
  INV_X1 U3629 ( .A(n2793), .ZN(U3351) );
  MUX2_X1 U3630 ( .A(n2794), .B(n2340), .S(U3149), .Z(n2795) );
  INV_X1 U3631 ( .A(n2795), .ZN(U3350) );
  INV_X1 U3632 ( .A(DATAI_5_), .ZN(n2796) );
  INV_X1 U3633 ( .A(n2836), .ZN(n2897) );
  MUX2_X1 U3634 ( .A(n2796), .B(n2897), .S(STATE_REG_SCAN_IN), .Z(n2797) );
  INV_X1 U3635 ( .A(n2797), .ZN(U3347) );
  INV_X1 U3636 ( .A(n4009), .ZN(n3998) );
  NAND2_X1 U3637 ( .A1(n3998), .A2(STATE_REG_SCAN_IN), .ZN(n2798) );
  OAI21_X1 U3638 ( .B1(STATE_REG_SCAN_IN), .B2(n2484), .A(n2798), .ZN(U3338)
         );
  MUX2_X1 U3639 ( .A(n2445), .B(n3955), .S(STATE_REG_SCAN_IN), .Z(n2799) );
  INV_X1 U3640 ( .A(n2799), .ZN(U3341) );
  INV_X1 U3641 ( .A(n4006), .ZN(n4028) );
  NAND2_X1 U3642 ( .A1(n4028), .A2(STATE_REG_SCAN_IN), .ZN(n2800) );
  OAI21_X1 U3643 ( .B1(STATE_REG_SCAN_IN), .B2(n2537), .A(n2800), .ZN(U3335)
         );
  MUX2_X1 U3644 ( .A(n2480), .B(n3987), .S(STATE_REG_SCAN_IN), .Z(n2801) );
  INV_X1 U3645 ( .A(n2801), .ZN(U3339) );
  INV_X1 U3646 ( .A(DATAI_10_), .ZN(n2802) );
  MUX2_X1 U3647 ( .A(n3132), .B(n2802), .S(U3149), .Z(n2803) );
  INV_X1 U3648 ( .A(n2803), .ZN(U3342) );
  INV_X1 U3649 ( .A(DATAI_22_), .ZN(n2805) );
  NAND2_X1 U3650 ( .A1(n3884), .A2(STATE_REG_SCAN_IN), .ZN(n2804) );
  OAI21_X1 U3651 ( .B1(STATE_REG_SCAN_IN), .B2(n2805), .A(n2804), .ZN(U3330)
         );
  INV_X1 U3652 ( .A(DATAI_24_), .ZN(n2806) );
  MUX2_X1 U3653 ( .A(n2806), .B(n2736), .S(STATE_REG_SCAN_IN), .Z(n2807) );
  INV_X1 U3654 ( .A(n2807), .ZN(U3328) );
  INV_X1 U3655 ( .A(DATAI_8_), .ZN(n2808) );
  INV_X1 U3656 ( .A(n3124), .ZN(n3130) );
  MUX2_X1 U3657 ( .A(n2808), .B(n3130), .S(STATE_REG_SCAN_IN), .Z(n2809) );
  INV_X1 U3658 ( .A(n2809), .ZN(U3344) );
  INV_X1 U3659 ( .A(DATAI_21_), .ZN(n2811) );
  NAND2_X1 U3660 ( .A1(n2695), .A2(STATE_REG_SCAN_IN), .ZN(n2810) );
  OAI21_X1 U3661 ( .B1(STATE_REG_SCAN_IN), .B2(n2811), .A(n2810), .ZN(U3331)
         );
  INV_X1 U3662 ( .A(DATAI_20_), .ZN(n2814) );
  NAND2_X1 U3663 ( .A1(n2812), .A2(STATE_REG_SCAN_IN), .ZN(n2813) );
  OAI21_X1 U3664 ( .B1(STATE_REG_SCAN_IN), .B2(n2814), .A(n2813), .ZN(U3332)
         );
  INV_X1 U3665 ( .A(n2816), .ZN(n2817) );
  AOI22_X1 U3666 ( .A1(n4562), .A2(n2818), .B1(n2817), .B2(n4517), .ZN(U3458)
         );
  INV_X1 U3667 ( .A(D_REG_1__SCAN_IN), .ZN(n2820) );
  INV_X1 U3668 ( .A(n2819), .ZN(n2901) );
  AOI22_X1 U3669 ( .A1(n4562), .A2(n2820), .B1(n2901), .B2(n4517), .ZN(U3459)
         );
  XNOR2_X1 U3670 ( .A(n2821), .B(n3102), .ZN(n2824) );
  XOR2_X1 U3671 ( .A(REG1_REG_3__SCAN_IN), .B(n2822), .Z(n2823) );
  AOI22_X1 U3672 ( .A1(n4498), .A2(n2824), .B1(n4486), .B2(n2823), .ZN(n2826)
         );
  AOI22_X1 U3673 ( .A1(n4494), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2825) );
  OAI211_X1 U3674 ( .C1(n2827), .C2(n4500), .A(n2826), .B(n2825), .ZN(U3243)
         );
  INV_X1 U3675 ( .A(n2828), .ZN(n4464) );
  MUX2_X1 U3676 ( .A(n2370), .B(REG1_REG_5__SCAN_IN), .S(n2836), .Z(n2890) );
  XNOR2_X1 U3677 ( .A(n2846), .B(REG1_REG_6__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3678 ( .A1(n2832), .A2(n4464), .ZN(n2833) );
  NAND2_X1 U3679 ( .A1(n2834), .A2(n2833), .ZN(n2893) );
  MUX2_X1 U3680 ( .A(REG2_REG_5__SCAN_IN), .B(n2835), .S(n2836), .Z(n2894) );
  NAND2_X1 U3681 ( .A1(n2836), .A2(REG2_REG_5__SCAN_IN), .ZN(n2837) );
  INV_X1 U3682 ( .A(n4463), .ZN(n2839) );
  XOR2_X1 U3683 ( .A(n2849), .B(REG2_REG_6__SCAN_IN), .Z(n2841) );
  AND2_X1 U3684 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3119) );
  AOI21_X1 U3685 ( .B1(n4494), .B2(ADDR_REG_6__SCAN_IN), .A(n3119), .ZN(n2838)
         );
  OAI21_X1 U3686 ( .B1(n2839), .B2(n4500), .A(n2838), .ZN(n2840) );
  AOI21_X1 U3687 ( .B1(n2841), .B2(n4498), .A(n2840), .ZN(n2842) );
  OAI21_X1 U3688 ( .B1(n2843), .B2(n4490), .A(n2842), .ZN(U3246) );
  NOR2_X1 U3689 ( .A1(n4494), .A2(U4043), .ZN(U3148) );
  INV_X1 U3690 ( .A(n2844), .ZN(n2845) );
  XNOR2_X1 U3691 ( .A(n2985), .B(n2399), .ZN(n2847) );
  XNOR2_X1 U3692 ( .A(n2984), .B(n2847), .ZN(n2859) );
  AND2_X1 U3693 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3219) );
  NOR2_X1 U3694 ( .A1(n4500), .A2(n2985), .ZN(n2848) );
  AOI211_X1 U3695 ( .C1(n4494), .C2(ADDR_REG_7__SCAN_IN), .A(n3219), .B(n2848), 
        .ZN(n2858) );
  NAND2_X1 U3696 ( .A1(n2849), .A2(REG2_REG_6__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U3697 ( .A1(n2850), .A2(n4463), .ZN(n2851) );
  NAND2_X1 U3698 ( .A1(n2852), .A2(n2851), .ZN(n2856) );
  MUX2_X1 U3699 ( .A(REG2_REG_7__SCAN_IN), .B(n2398), .S(n2985), .Z(n2853) );
  INV_X1 U3700 ( .A(n2853), .ZN(n2855) );
  MUX2_X1 U3701 ( .A(n2398), .B(REG2_REG_7__SCAN_IN), .S(n2985), .Z(n2854) );
  NAND2_X1 U3702 ( .A1(n2856), .A2(n2854), .ZN(n2983) );
  OAI211_X1 U3703 ( .C1(n2856), .C2(n2855), .A(n2983), .B(n4498), .ZN(n2857)
         );
  OAI211_X1 U3704 ( .C1(n2859), .C2(n4490), .A(n2858), .B(n2857), .ZN(U3247)
         );
  NAND2_X1 U3705 ( .A1(n2671), .A2(n2871), .ZN(n3804) );
  AND2_X1 U3706 ( .A1(n3802), .A2(n3804), .ZN(n3764) );
  INV_X1 U3707 ( .A(n3764), .ZN(n4511) );
  INV_X1 U3708 ( .A(n2751), .ZN(n2860) );
  NOR2_X1 U3709 ( .A1(n2871), .A2(n2860), .ZN(n4509) );
  INV_X1 U3710 ( .A(n4212), .ZN(n3333) );
  NOR2_X1 U3711 ( .A1(n3333), .A2(n4304), .ZN(n2861) );
  OAI22_X1 U3712 ( .A1(n2861), .A2(n3764), .B1(n2319), .B2(n4311), .ZN(n4507)
         );
  AOI211_X1 U3713 ( .C1(n4537), .C2(n4511), .A(n4509), .B(n4507), .ZN(n4525)
         );
  NAND2_X1 U3714 ( .A1(n4559), .A2(REG1_REG_0__SCAN_IN), .ZN(n2862) );
  OAI21_X1 U3715 ( .B1(n4525), .B2(n4559), .A(n2862), .ZN(U3518) );
  NAND2_X1 U3716 ( .A1(n4308), .A2(n2671), .ZN(n2866) );
  NAND2_X1 U3717 ( .A1(n4266), .A2(n3594), .ZN(n2865) );
  OAI211_X1 U3718 ( .C1(n4262), .C2(n2745), .A(n2866), .B(n2865), .ZN(n2867)
         );
  INV_X1 U3719 ( .A(n2867), .ZN(n2870) );
  NAND2_X1 U3720 ( .A1(n2868), .A2(n4304), .ZN(n2869) );
  OAI211_X1 U3721 ( .C1(n3031), .C2(n4212), .A(n2870), .B(n2869), .ZN(n3033)
         );
  INV_X1 U3722 ( .A(n4544), .ZN(n4528) );
  OAI21_X1 U3723 ( .B1(n2871), .B2(n2745), .A(n2962), .ZN(n3037) );
  OAI22_X1 U3724 ( .A1(n3031), .A2(n4529), .B1(n4528), .B2(n3037), .ZN(n2872)
         );
  NOR2_X1 U3725 ( .A1(n3033), .A2(n2872), .ZN(n4526) );
  NAND2_X1 U3726 ( .A1(n4559), .A2(REG1_REG_1__SCAN_IN), .ZN(n2873) );
  OAI21_X1 U3727 ( .B1(n4526), .B2(n4559), .A(n2873), .ZN(U3519) );
  INV_X1 U3728 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U3729 ( .A1(U4043), .A2(n3216), .ZN(n2874) );
  OAI21_X1 U3730 ( .B1(U4043), .B2(n4698), .A(n2874), .ZN(U3558) );
  INV_X1 U3731 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U3732 ( .A1(U4043), .A2(n3205), .ZN(n2875) );
  OAI21_X1 U3733 ( .B1(U4043), .B2(n4616), .A(n2875), .ZN(U3557) );
  INV_X1 U3734 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U3735 ( .A1(U4043), .A2(n4307), .ZN(n2876) );
  OAI21_X1 U3736 ( .B1(U4043), .B2(n4669), .A(n2876), .ZN(U3564) );
  INV_X1 U3737 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U3738 ( .A1(U4043), .A2(n3594), .ZN(n2877) );
  OAI21_X1 U3739 ( .B1(U4043), .B2(n4632), .A(n2877), .ZN(U3552) );
  INV_X1 U3740 ( .A(n2878), .ZN(n2883) );
  OAI21_X1 U3741 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4457), .A(n2879), .ZN(n2880)
         );
  MUX2_X1 U3742 ( .A(n2880), .B(n2879), .S(IR_REG_0__SCAN_IN), .Z(n2882) );
  OAI22_X1 U3743 ( .A1(n2883), .A2(n2882), .B1(STATE_REG_SCAN_IN), .B2(n2881), 
        .ZN(n2885) );
  INV_X1 U3744 ( .A(IR_REG_0__SCAN_IN), .ZN(n4676) );
  NOR3_X1 U3745 ( .A1(n4490), .A2(REG1_REG_0__SCAN_IN), .A3(n4676), .ZN(n2884)
         );
  AOI211_X1 U3746 ( .C1(n4494), .C2(ADDR_REG_0__SCAN_IN), .A(n2885), .B(n2884), 
        .ZN(n2886) );
  INV_X1 U3747 ( .A(n2886), .ZN(U3240) );
  INV_X1 U3748 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U3749 ( .A1(n4265), .A2(U4043), .ZN(n2887) );
  OAI21_X1 U3750 ( .B1(U4043), .B2(n4671), .A(n2887), .ZN(U3568) );
  INV_X1 U3751 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U3752 ( .A1(n3648), .A2(U4043), .ZN(n2888) );
  OAI21_X1 U3753 ( .B1(U4043), .B2(n4579), .A(n2888), .ZN(U3566) );
  AOI211_X1 U3754 ( .C1(n2891), .C2(n2890), .A(n4490), .B(n2889), .ZN(n2899)
         );
  OAI211_X1 U3755 ( .C1(n2894), .C2(n2893), .A(n4498), .B(n2892), .ZN(n2896)
         );
  NOR2_X1 U3756 ( .A1(STATE_REG_SCAN_IN), .A2(n2383), .ZN(n3049) );
  AOI21_X1 U3757 ( .B1(n4494), .B2(ADDR_REG_5__SCAN_IN), .A(n3049), .ZN(n2895)
         );
  OAI211_X1 U3758 ( .C1(n4500), .C2(n2897), .A(n2896), .B(n2895), .ZN(n2898)
         );
  OR2_X1 U3759 ( .A1(n2899), .A2(n2898), .ZN(U3245) );
  NAND2_X1 U3760 ( .A1(n2900), .A2(D_REG_1__SCAN_IN), .ZN(n2902) );
  AOI21_X1 U3761 ( .B1(n2903), .B2(n2902), .A(n2901), .ZN(n3027) );
  NAND2_X1 U3762 ( .A1(n3027), .A2(n2904), .ZN(n2919) );
  NAND2_X1 U3763 ( .A1(n4034), .A2(n3884), .ZN(n2930) );
  INV_X1 U3764 ( .A(n2930), .ZN(n2905) );
  NAND2_X1 U3765 ( .A1(n4517), .A2(n2905), .ZN(n2906) );
  OR2_X1 U3766 ( .A1(n3508), .A2(n2906), .ZN(n2913) );
  OR2_X1 U3767 ( .A1(n2919), .A2(n2913), .ZN(n2947) );
  INV_X1 U3768 ( .A(n2947), .ZN(n2907) );
  INV_X1 U3769 ( .A(n2908), .ZN(n2910) );
  NAND2_X1 U3770 ( .A1(n2751), .A2(n4459), .ZN(n2909) );
  NAND3_X1 U3771 ( .A1(n2910), .A2(n4262), .A3(n2909), .ZN(n2915) );
  NAND2_X1 U3772 ( .A1(n2915), .A2(n4262), .ZN(n2911) );
  NAND2_X1 U3773 ( .A1(n2919), .A2(n2911), .ZN(n2912) );
  NAND2_X1 U3774 ( .A1(n2912), .A2(n3024), .ZN(n2975) );
  INV_X1 U3775 ( .A(n2975), .ZN(n2914) );
  INV_X1 U3776 ( .A(n2913), .ZN(n3882) );
  NAND2_X1 U3777 ( .A1(n2919), .A2(n3882), .ZN(n2976) );
  NAND3_X1 U3778 ( .A1(n2914), .A2(n3026), .A3(n2976), .ZN(n3595) );
  NAND2_X1 U3779 ( .A1(n3595), .A2(REG3_REG_0__SCAN_IN), .ZN(n2926) );
  INV_X1 U3780 ( .A(n2915), .ZN(n2916) );
  NAND2_X1 U3781 ( .A1(n2916), .A2(n3026), .ZN(n2917) );
  NAND2_X1 U3782 ( .A1(n4306), .A2(n3026), .ZN(n2918) );
  OR2_X1 U3783 ( .A1(n2919), .A2(n2918), .ZN(n2922) );
  INV_X1 U3784 ( .A(n2920), .ZN(n2921) );
  AOI22_X1 U3785 ( .A1(n2924), .A2(n3713), .B1(n3719), .B2(n2923), .ZN(n2925)
         );
  OAI211_X1 U3786 ( .C1(n2319), .C2(n3715), .A(n2926), .B(n2925), .ZN(U3229)
         );
  INV_X1 U3787 ( .A(n2929), .ZN(n2931) );
  NAND2_X4 U3788 ( .A1(n2760), .A2(n2930), .ZN(n3506) );
  XNOR2_X1 U3789 ( .A(n2931), .B(n3506), .ZN(n2967) );
  AOI22_X1 U3790 ( .A1(n2011), .A2(n3594), .B1(n2341), .B2(n2007), .ZN(n2968)
         );
  XNOR2_X1 U3791 ( .A(n2967), .B(n2968), .ZN(n2946) );
  NAND2_X1 U3792 ( .A1(n2325), .A2(n3012), .ZN(n2933) );
  NAND2_X1 U3793 ( .A1(n2933), .A2(n2036), .ZN(n2935) );
  AOI22_X1 U3794 ( .A1(n2971), .A2(n2325), .B1(n3596), .B2(n2007), .ZN(n2942)
         );
  NAND2_X1 U3795 ( .A1(n2937), .A2(n2936), .ZN(n2940) );
  NAND2_X1 U3796 ( .A1(n2941), .A2(n3598), .ZN(n3600) );
  OR2_X1 U3797 ( .A1(n2943), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U3798 ( .A1(n3600), .A2(n2944), .ZN(n2945) );
  NOR2_X1 U3799 ( .A1(n2945), .A2(n2946), .ZN(n2970) );
  AOI21_X1 U3800 ( .B1(n2946), .B2(n2945), .A(n2970), .ZN(n2950) );
  NOR2_X2 U3801 ( .A1(n2947), .A2(n4467), .ZN(n3667) );
  AOI22_X1 U3802 ( .A1(n3667), .A2(n2325), .B1(n2341), .B2(n3719), .ZN(n2949)
         );
  AOI22_X1 U3803 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3595), .B1(n3668), .B2(n3898), .ZN(n2948) );
  OAI211_X1 U3804 ( .C1(n2950), .C2(n3706), .A(n2949), .B(n2948), .ZN(U3234)
         );
  INV_X1 U3805 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4670) );
  NAND2_X1 U3806 ( .A1(n4189), .A2(U4043), .ZN(n2951) );
  OAI21_X1 U3807 ( .B1(U4043), .B2(n4670), .A(n2951), .ZN(U3572) );
  OAI21_X1 U3808 ( .B1(n2954), .B2(n2953), .A(n2952), .ZN(n4501) );
  INV_X1 U3809 ( .A(n3898), .ZN(n3019) );
  OAI21_X1 U3810 ( .B1(n3782), .B2(n2956), .A(n2955), .ZN(n2957) );
  NAND2_X1 U3811 ( .A1(n2957), .A2(n4304), .ZN(n2959) );
  AOI22_X1 U3812 ( .A1(n4308), .A2(n2325), .B1(n4306), .B2(n2341), .ZN(n2958)
         );
  OAI211_X1 U3813 ( .C1(n3019), .C2(n4311), .A(n2959), .B(n2958), .ZN(n2960)
         );
  AOI21_X1 U3814 ( .B1(n3333), .B2(n4501), .A(n2960), .ZN(n4506) );
  INV_X1 U3815 ( .A(n4506), .ZN(n2961) );
  AOI21_X1 U3816 ( .B1(n4537), .B2(n4501), .A(n2961), .ZN(n2995) );
  AND2_X1 U3817 ( .A1(n2962), .A2(n2341), .ZN(n2963) );
  NOR2_X1 U3818 ( .A1(n3101), .A2(n2963), .ZN(n4502) );
  INV_X1 U3819 ( .A(n4502), .ZN(n2964) );
  OAI22_X1 U3820 ( .A1(n4453), .A2(n2964), .B1(n4553), .B2(n2327), .ZN(n2965)
         );
  INV_X1 U3821 ( .A(n2965), .ZN(n2966) );
  OAI21_X1 U3822 ( .B1(n2995), .B2(n4552), .A(n2966), .ZN(U3471) );
  OR2_X2 U3823 ( .A1(n2970), .A2(n2969), .ZN(n3011) );
  AOI22_X1 U3824 ( .A1(n2011), .A2(n3898), .B1(n3094), .B2(n2007), .ZN(n3008)
         );
  XNOR2_X1 U3825 ( .A(n2972), .B(n3010), .ZN(n2981) );
  OAI22_X1 U3826 ( .A1(n3717), .A2(n2928), .B1(n3699), .B2(n3100), .ZN(n2979)
         );
  NAND2_X1 U3827 ( .A1(n2759), .A2(n2973), .ZN(n2974) );
  OAI21_X1 U3828 ( .B1(n2975), .B2(n2974), .A(STATE_REG_SCAN_IN), .ZN(n2977)
         );
  MUX2_X1 U3829 ( .A(n3703), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2978) );
  AOI211_X1 U3830 ( .C1(n3668), .C2(n3897), .A(n2979), .B(n2978), .ZN(n2980)
         );
  OAI21_X1 U3831 ( .B1(n2981), .B2(n3706), .A(n2980), .ZN(U3215) );
  OR2_X1 U3832 ( .A1(n2985), .A2(n2398), .ZN(n2982) );
  XNOR2_X1 U3833 ( .A(n3125), .B(n3130), .ZN(n3123) );
  XNOR2_X1 U3834 ( .A(n3123), .B(n3232), .ZN(n2992) );
  INV_X1 U3835 ( .A(n2985), .ZN(n4462) );
  OAI21_X1 U3836 ( .B1(n2399), .B2(n2985), .A(n2984), .ZN(n2986) );
  OAI211_X1 U3837 ( .C1(n2987), .C2(REG1_REG_8__SCAN_IN), .A(n3129), .B(n4486), 
        .ZN(n2990) );
  NAND2_X1 U3838 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3206) );
  INV_X1 U3839 ( .A(n3206), .ZN(n2988) );
  AOI21_X1 U3840 ( .B1(n4494), .B2(ADDR_REG_8__SCAN_IN), .A(n2988), .ZN(n2989)
         );
  OAI211_X1 U3841 ( .C1(n4500), .C2(n3130), .A(n2990), .B(n2989), .ZN(n2991)
         );
  AOI21_X1 U3842 ( .B1(n4498), .B2(n2992), .A(n2991), .ZN(n2993) );
  INV_X1 U3843 ( .A(n2993), .ZN(U3248) );
  INV_X1 U3844 ( .A(n4395), .ZN(n3166) );
  AOI22_X1 U3845 ( .A1(n3166), .A2(n4502), .B1(REG1_REG_2__SCAN_IN), .B2(n4559), .ZN(n2994) );
  OAI21_X1 U3846 ( .B1(n2995), .B2(n4559), .A(n2994), .ZN(U3520) );
  AND2_X1 U3847 ( .A1(n3819), .A2(n3831), .ZN(n3763) );
  XOR2_X1 U3848 ( .A(n2997), .B(n3763), .Z(n3265) );
  XNOR2_X1 U3849 ( .A(n2998), .B(n3763), .ZN(n3001) );
  INV_X1 U3850 ( .A(n3205), .ZN(n3190) );
  AOI22_X1 U3851 ( .A1(n4308), .A2(n3896), .B1(n4306), .B2(n3120), .ZN(n2999)
         );
  OAI21_X1 U3852 ( .B1(n3190), .B2(n4311), .A(n2999), .ZN(n3000) );
  AOI21_X1 U3853 ( .B1(n3001), .B2(n4304), .A(n3000), .ZN(n3273) );
  OAI21_X1 U3854 ( .B1(n3265), .B2(n4539), .A(n3273), .ZN(n3006) );
  NOR2_X1 U3855 ( .A1(n3150), .A2(n3250), .ZN(n3002) );
  OR2_X1 U3856 ( .A1(n3246), .A2(n3002), .ZN(n3269) );
  INV_X1 U3857 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4569) );
  OAI22_X1 U3858 ( .A1(n3269), .A2(n4395), .B1(n4561), .B2(n4569), .ZN(n3003)
         );
  AOI21_X1 U3859 ( .B1(n3006), .B2(n4561), .A(n3003), .ZN(n3004) );
  INV_X1 U3860 ( .A(n3004), .ZN(U3524) );
  OAI22_X1 U3861 ( .A1(n3269), .A2(n4453), .B1(n4553), .B2(n2381), .ZN(n3005)
         );
  AOI21_X1 U3862 ( .B1(n3006), .B2(n4553), .A(n3005), .ZN(n3007) );
  INV_X1 U3863 ( .A(n3007), .ZN(U3479) );
  AOI22_X1 U3864 ( .A1(n2011), .A2(n3897), .B1(n3372), .B2(n3067), .ZN(n3041)
         );
  NAND2_X1 U3865 ( .A1(n3372), .A2(n3897), .ZN(n3014) );
  NAND2_X1 U3866 ( .A1(n3456), .A2(n3067), .ZN(n3013) );
  NAND2_X1 U3867 ( .A1(n3014), .A2(n3013), .ZN(n3015) );
  XNOR2_X1 U3868 ( .A(n3015), .B(n3506), .ZN(n3040) );
  XNOR2_X1 U3869 ( .A(n3041), .B(n3040), .ZN(n3016) );
  OAI211_X1 U3870 ( .C1(n3017), .C2(n3016), .A(n3044), .B(n3713), .ZN(n3023)
         );
  INV_X1 U3871 ( .A(n3018), .ZN(n3021) );
  INV_X1 U3872 ( .A(n3896), .ZN(n3117) );
  OAI22_X1 U3873 ( .A1(n3717), .A2(n3019), .B1(n3117), .B2(n3715), .ZN(n3020)
         );
  AOI211_X1 U3874 ( .C1(n3067), .C2(n3719), .A(n3021), .B(n3020), .ZN(n3022)
         );
  OAI211_X1 U3875 ( .C1(n3722), .C2(n3075), .A(n3023), .B(n3022), .ZN(U3227)
         );
  NAND4_X1 U3876 ( .A1(n3027), .A2(n3026), .A3(n3025), .A4(n3024), .ZN(n3028)
         );
  NAND2_X1 U3877 ( .A1(n3029), .A2(n4459), .ZN(n3140) );
  INV_X1 U3878 ( .A(n3140), .ZN(n3030) );
  INV_X1 U3879 ( .A(n3031), .ZN(n3032) );
  AOI22_X1 U3880 ( .A1(n4512), .A2(n3032), .B1(REG3_REG_1__SCAN_IN), .B2(n4510), .ZN(n3036) );
  MUX2_X1 U3881 ( .A(n3033), .B(REG2_REG_1__SCAN_IN), .S(n4515), .Z(n3034) );
  INV_X1 U3882 ( .A(n3034), .ZN(n3035) );
  OAI211_X1 U3883 ( .C1(n4272), .C2(n3037), .A(n3036), .B(n3035), .ZN(U3289)
         );
  NAND2_X1 U3884 ( .A1(n3899), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3038) );
  OAI21_X1 U3885 ( .B1(n3799), .B2(n3899), .A(n3038), .ZN(U3579) );
  INV_X1 U3886 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U3887 ( .A1(n4094), .A2(U4043), .ZN(n3039) );
  OAI21_X1 U3888 ( .B1(U4043), .B2(n4697), .A(n3039), .ZN(U3577) );
  NAND2_X1 U3889 ( .A1(n3040), .A2(n3042), .ZN(n3043) );
  AOI22_X1 U3890 ( .A1(n2011), .A2(n3896), .B1(n3151), .B2(n2007), .ZN(n3109)
         );
  AOI22_X1 U3891 ( .A1(n3372), .A2(n3896), .B1(n3456), .B2(n3151), .ZN(n3045)
         );
  XNOR2_X1 U3892 ( .A(n3045), .B(n3506), .ZN(n3108) );
  XOR2_X1 U3893 ( .A(n3109), .B(n3108), .Z(n3046) );
  OAI211_X1 U3894 ( .C1(n3047), .C2(n3046), .A(n3113), .B(n3713), .ZN(n3051)
         );
  INV_X1 U3895 ( .A(n3897), .ZN(n3149) );
  INV_X1 U3896 ( .A(n3895), .ZN(n3217) );
  OAI22_X1 U3897 ( .A1(n3717), .A2(n3149), .B1(n3217), .B2(n3715), .ZN(n3048)
         );
  AOI211_X1 U3898 ( .C1(n3151), .C2(n3719), .A(n3049), .B(n3048), .ZN(n3050)
         );
  OAI211_X1 U3899 ( .C1(n3722), .C2(n3152), .A(n3051), .B(n3050), .ZN(U3224)
         );
  NAND2_X1 U3900 ( .A1(n3053), .A2(n3052), .ZN(n3054) );
  AND2_X1 U3901 ( .A1(n3826), .A2(n3824), .ZN(n3771) );
  XNOR2_X1 U3902 ( .A(n3054), .B(n3771), .ZN(n3235) );
  XNOR2_X1 U3903 ( .A(n3055), .B(n3771), .ZN(n3058) );
  AOI22_X1 U3904 ( .A1(n4266), .A2(n3894), .B1(n4306), .B2(n3196), .ZN(n3057)
         );
  NAND2_X1 U3905 ( .A1(n4308), .A2(n3205), .ZN(n3056) );
  OAI211_X1 U3906 ( .C1(n3058), .C2(n4268), .A(n3057), .B(n3056), .ZN(n3230)
         );
  AOI21_X1 U3907 ( .B1(n3235), .B2(n4547), .A(n3230), .ZN(n3062) );
  INV_X1 U3908 ( .A(n3086), .ZN(n3059) );
  AOI21_X1 U3909 ( .B1(n3196), .B2(n3244), .A(n3059), .ZN(n3234) );
  AOI22_X1 U3910 ( .A1(n3234), .A2(n3166), .B1(REG1_REG_8__SCAN_IN), .B2(n4559), .ZN(n3060) );
  OAI21_X1 U3911 ( .B1(n3062), .B2(n4559), .A(n3060), .ZN(U3526) );
  INV_X1 U3912 ( .A(n4453), .ZN(n3164) );
  AOI22_X1 U3913 ( .A1(n3234), .A2(n3164), .B1(REG0_REG_8__SCAN_IN), .B2(n4552), .ZN(n3061) );
  OAI21_X1 U3914 ( .B1(n3062), .B2(n4552), .A(n3061), .ZN(U3483) );
  NAND2_X1 U3915 ( .A1(n3064), .A2(n3778), .ZN(n3065) );
  NAND2_X1 U3916 ( .A1(n3063), .A2(n3065), .ZN(n4533) );
  INV_X1 U3917 ( .A(n4512), .ZN(n3107) );
  XNOR2_X1 U3918 ( .A(n3066), .B(n3778), .ZN(n3071) );
  AOI22_X1 U3919 ( .A1(n4308), .A2(n3898), .B1(n4306), .B2(n3067), .ZN(n3069)
         );
  NAND2_X1 U3920 ( .A1(n4266), .A2(n3896), .ZN(n3068) );
  OAI211_X1 U3921 ( .C1(n4533), .C2(n4212), .A(n3069), .B(n3068), .ZN(n3070)
         );
  AOI21_X1 U3922 ( .B1(n3071), .B2(n4304), .A(n3070), .ZN(n3072) );
  INV_X1 U3923 ( .A(n3072), .ZN(n4535) );
  INV_X1 U3924 ( .A(n3099), .ZN(n3074) );
  OAI211_X1 U3925 ( .C1(n3074), .C2(n3073), .A(n4544), .B(n2025), .ZN(n4534)
         );
  OAI22_X1 U3926 ( .A1(n4534), .A2(n4459), .B1(n4299), .B2(n3075), .ZN(n3076)
         );
  OAI21_X1 U3927 ( .B1(n4535), .B2(n3076), .A(n4313), .ZN(n3078) );
  NAND2_X1 U3928 ( .A1(n4515), .A2(REG2_REG_4__SCAN_IN), .ZN(n3077) );
  OAI211_X1 U3929 ( .C1(n4533), .C2(n3107), .A(n3078), .B(n3077), .ZN(U3286)
         );
  INV_X1 U3930 ( .A(n3079), .ZN(n3841) );
  AND2_X1 U3931 ( .A1(n3841), .A2(n3827), .ZN(n3773) );
  XNOR2_X1 U3932 ( .A(n3080), .B(n3773), .ZN(n3263) );
  XNOR2_X1 U3933 ( .A(n3081), .B(n3773), .ZN(n3085) );
  INV_X1 U3934 ( .A(n3893), .ZN(n3307) );
  OAI22_X1 U3935 ( .A1(n3307), .A2(n4311), .B1(n4262), .B2(n3082), .ZN(n3083)
         );
  AOI21_X1 U3936 ( .B1(n4308), .B2(n3216), .A(n3083), .ZN(n3084) );
  OAI21_X1 U3937 ( .B1(n3085), .B2(n4268), .A(n3084), .ZN(n3260) );
  AOI21_X1 U3938 ( .B1(n3263), .B2(n4547), .A(n3260), .ZN(n3091) );
  AND2_X1 U3939 ( .A1(n3086), .A2(n3310), .ZN(n3087) );
  NOR2_X1 U3940 ( .A1(n3162), .A2(n3087), .ZN(n3258) );
  AOI22_X1 U3941 ( .A1(n3258), .A2(n3164), .B1(REG0_REG_9__SCAN_IN), .B2(n4552), .ZN(n3088) );
  OAI21_X1 U3942 ( .B1(n3091), .B2(n4552), .A(n3088), .ZN(U3485) );
  NAND2_X1 U3943 ( .A1(n4559), .A2(REG1_REG_9__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3944 ( .A1(n3258), .A2(n3166), .ZN(n3089) );
  OAI211_X1 U3945 ( .C1(n3091), .C2(n4559), .A(n3090), .B(n3089), .ZN(U3527)
         );
  XNOR2_X1 U3946 ( .A(n3092), .B(n3781), .ZN(n4530) );
  XNOR2_X1 U3947 ( .A(n3093), .B(n3781), .ZN(n3097) );
  AOI22_X1 U3948 ( .A1(n4308), .A2(n3594), .B1(n4306), .B2(n3094), .ZN(n3095)
         );
  OAI21_X1 U3949 ( .B1(n3149), .B2(n4311), .A(n3095), .ZN(n3096) );
  AOI21_X1 U3950 ( .B1(n3097), .B2(n4304), .A(n3096), .ZN(n3098) );
  OAI21_X1 U3951 ( .B1(n4530), .B2(n4212), .A(n3098), .ZN(n4532) );
  NAND2_X1 U3952 ( .A1(n4532), .A2(n4313), .ZN(n3106) );
  OAI21_X1 U3953 ( .B1(n3101), .B2(n3100), .A(n3099), .ZN(n4527) );
  INV_X1 U3954 ( .A(n4527), .ZN(n3104) );
  OAI22_X1 U3955 ( .A1(n4313), .A2(n3102), .B1(REG3_REG_3__SCAN_IN), .B2(n4299), .ZN(n3103) );
  AOI21_X1 U3956 ( .B1(n4503), .B2(n3104), .A(n3103), .ZN(n3105) );
  OAI211_X1 U3957 ( .C1(n4530), .C2(n3107), .A(n3106), .B(n3105), .ZN(U3287)
         );
  INV_X1 U3958 ( .A(n3108), .ZN(n3111) );
  INV_X1 U3959 ( .A(n3109), .ZN(n3110) );
  AOI22_X1 U3960 ( .A1(n3372), .A2(n3895), .B1(n3456), .B2(n3120), .ZN(n3114)
         );
  XOR2_X1 U3961 ( .A(n3506), .B(n3114), .Z(n3184) );
  INV_X2 U3962 ( .A(n2007), .ZN(n3505) );
  OAI22_X1 U3963 ( .A1(n3509), .A2(n3217), .B1(n3250), .B2(n3505), .ZN(n3185)
         );
  XNOR2_X1 U3964 ( .A(n3184), .B(n3185), .ZN(n3115) );
  XNOR2_X1 U3965 ( .A(n3186), .B(n3115), .ZN(n3116) );
  NAND2_X1 U3966 ( .A1(n3116), .A2(n3713), .ZN(n3122) );
  OAI22_X1 U3967 ( .A1(n3717), .A2(n3117), .B1(n3190), .B2(n3715), .ZN(n3118)
         );
  AOI211_X1 U3968 ( .C1(n3120), .C2(n3719), .A(n3119), .B(n3118), .ZN(n3121)
         );
  OAI211_X1 U3969 ( .C1(n3722), .C2(n3266), .A(n3122), .B(n3121), .ZN(U3236)
         );
  NAND2_X1 U3970 ( .A1(n3125), .A2(n3124), .ZN(n3126) );
  MUX2_X1 U3971 ( .A(REG2_REG_9__SCAN_IN), .B(n3127), .S(n4461), .Z(n3929) );
  NAND2_X1 U3972 ( .A1(n4461), .A2(REG2_REG_9__SCAN_IN), .ZN(n3128) );
  XNOR2_X1 U3973 ( .A(n3941), .B(n3223), .ZN(n3138) );
  XOR2_X1 U3974 ( .A(REG1_REG_9__SCAN_IN), .B(n4461), .Z(n3923) );
  INV_X1 U3975 ( .A(n4461), .ZN(n3925) );
  INV_X1 U3976 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3131) );
  OAI211_X1 U3977 ( .C1(n3133), .C2(REG1_REG_10__SCAN_IN), .A(n3936), .B(n4486), .ZN(n3136) );
  NAND2_X1 U3978 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n3574) );
  INV_X1 U3979 ( .A(n3574), .ZN(n3134) );
  AOI21_X1 U3980 ( .B1(n4494), .B2(ADDR_REG_10__SCAN_IN), .A(n3134), .ZN(n3135) );
  OAI211_X1 U3981 ( .C1(n4500), .C2(n3132), .A(n3136), .B(n3135), .ZN(n3137)
         );
  AOI21_X1 U3982 ( .B1(n4498), .B2(n3138), .A(n3137), .ZN(n3139) );
  INV_X1 U3983 ( .A(n3139), .ZN(U3250) );
  NAND2_X1 U3984 ( .A1(n4212), .A2(n3140), .ZN(n3141) );
  INV_X1 U3985 ( .A(n3816), .ZN(n3142) );
  AND2_X1 U3986 ( .A1(n3142), .A2(n3830), .ZN(n3774) );
  INV_X1 U3987 ( .A(n3774), .ZN(n3144) );
  XNOR2_X1 U3988 ( .A(n3143), .B(n3144), .ZN(n4540) );
  XNOR2_X1 U3989 ( .A(n3145), .B(n3144), .ZN(n3146) );
  NAND2_X1 U3990 ( .A1(n3146), .A2(n4304), .ZN(n3148) );
  AOI22_X1 U3991 ( .A1(n4266), .A2(n3895), .B1(n4306), .B2(n3151), .ZN(n3147)
         );
  OAI211_X1 U3992 ( .C1(n3149), .C2(n4263), .A(n3148), .B(n3147), .ZN(n4542)
         );
  NAND2_X1 U3993 ( .A1(n4542), .A2(n4313), .ZN(n3155) );
  AOI21_X1 U3994 ( .B1(n3151), .B2(n2025), .A(n3150), .ZN(n4543) );
  OAI22_X1 U3995 ( .A1(n4313), .A2(n2835), .B1(n3152), .B2(n4299), .ZN(n3153)
         );
  AOI21_X1 U3996 ( .B1(n4543), .B2(n4503), .A(n3153), .ZN(n3154) );
  OAI211_X1 U3997 ( .C1(n4316), .C2(n4540), .A(n3155), .B(n3154), .ZN(U3285)
         );
  NAND2_X1 U3998 ( .A1(n3838), .A2(n3839), .ZN(n3157) );
  XNOR2_X1 U3999 ( .A(n3156), .B(n3157), .ZN(n3226) );
  INV_X1 U4000 ( .A(n3892), .ZN(n3622) );
  INV_X1 U4001 ( .A(n3157), .ZN(n3761) );
  XNOR2_X1 U4002 ( .A(n3158), .B(n3761), .ZN(n3159) );
  NAND2_X1 U4003 ( .A1(n3159), .A2(n4304), .ZN(n3161) );
  AOI22_X1 U4004 ( .A1(n4308), .A2(n3894), .B1(n4306), .B2(n3348), .ZN(n3160)
         );
  OAI211_X1 U4005 ( .C1(n3622), .C2(n4311), .A(n3161), .B(n3160), .ZN(n3222)
         );
  AOI21_X1 U4006 ( .B1(n4547), .B2(n3226), .A(n3222), .ZN(n3168) );
  INV_X1 U4007 ( .A(n3162), .ZN(n3163) );
  AOI21_X1 U4008 ( .B1(n3348), .B2(n3163), .A(n3177), .ZN(n3225) );
  AOI22_X1 U4009 ( .A1(n3225), .A2(n3164), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4552), .ZN(n3165) );
  OAI21_X1 U4010 ( .B1(n3168), .B2(n4552), .A(n3165), .ZN(U3487) );
  AOI22_X1 U4011 ( .A1(n3225), .A2(n3166), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4559), .ZN(n3167) );
  OAI21_X1 U4012 ( .B1(n3168), .B2(n4559), .A(n3167), .ZN(U3528) );
  XOR2_X1 U4013 ( .A(n3277), .B(n3779), .Z(n3176) );
  NAND2_X1 U4014 ( .A1(n3170), .A2(n3779), .ZN(n3171) );
  NAND2_X1 U4015 ( .A1(n3169), .A2(n3171), .ZN(n3315) );
  INV_X1 U4016 ( .A(n3891), .ZN(n3173) );
  AOI22_X1 U4017 ( .A1(n4308), .A2(n3893), .B1(n4306), .B2(n3353), .ZN(n3172)
         );
  OAI21_X1 U4018 ( .B1(n3173), .B2(n4311), .A(n3172), .ZN(n3174) );
  AOI21_X1 U4019 ( .B1(n3315), .B2(n3333), .A(n3174), .ZN(n3175) );
  OAI21_X1 U4020 ( .B1(n3176), .B2(n4268), .A(n3175), .ZN(n3314) );
  INV_X1 U4021 ( .A(n3314), .ZN(n3183) );
  OR2_X1 U4022 ( .A1(n3177), .A2(n3357), .ZN(n3178) );
  NAND2_X1 U4023 ( .A1(n3283), .A2(n3178), .ZN(n3320) );
  INV_X1 U4024 ( .A(n3179), .ZN(n3359) );
  AOI22_X1 U4025 ( .A1(n4515), .A2(REG2_REG_11__SCAN_IN), .B1(n3359), .B2(
        n4510), .ZN(n3180) );
  OAI21_X1 U4026 ( .B1(n3320), .B2(n4272), .A(n3180), .ZN(n3181) );
  AOI21_X1 U4027 ( .B1(n3315), .B2(n4512), .A(n3181), .ZN(n3182) );
  OAI21_X1 U4028 ( .B1(n3183), .B2(n4515), .A(n3182), .ZN(U3279) );
  NAND2_X1 U4029 ( .A1(n3372), .A2(n3205), .ZN(n3188) );
  NAND2_X1 U4030 ( .A1(n3456), .A2(n3240), .ZN(n3187) );
  NAND2_X1 U4031 ( .A1(n3188), .A2(n3187), .ZN(n3189) );
  XNOR2_X1 U4032 ( .A(n3189), .B(n2934), .ZN(n3195) );
  OR2_X1 U4033 ( .A1(n3509), .A2(n3190), .ZN(n3192) );
  NAND2_X1 U4034 ( .A1(n3372), .A2(n3240), .ZN(n3191) );
  NAND2_X1 U4035 ( .A1(n3192), .A2(n3191), .ZN(n3193) );
  XNOR2_X1 U4036 ( .A(n3195), .B(n3193), .ZN(n3214) );
  INV_X1 U4037 ( .A(n3193), .ZN(n3194) );
  AOI22_X1 U4038 ( .A1(n2011), .A2(n3216), .B1(n2007), .B2(n3196), .ZN(n3201)
         );
  NAND2_X1 U4039 ( .A1(n3372), .A2(n3216), .ZN(n3198) );
  NAND2_X1 U4040 ( .A1(n3456), .A2(n3196), .ZN(n3197) );
  NAND2_X1 U4041 ( .A1(n3198), .A2(n3197), .ZN(n3199) );
  XNOR2_X1 U4042 ( .A(n3199), .B(n2934), .ZN(n3200) );
  INV_X1 U40430 ( .A(n3200), .ZN(n3203) );
  INV_X1 U4044 ( .A(n3201), .ZN(n3202) );
  NAND2_X1 U4045 ( .A1(n3203), .A2(n3202), .ZN(n3302) );
  NAND2_X1 U4046 ( .A1(n2052), .A2(n3302), .ZN(n3204) );
  XNOR2_X1 U4047 ( .A(n3303), .B(n3204), .ZN(n3212) );
  INV_X1 U4048 ( .A(n3231), .ZN(n3210) );
  AOI22_X1 U4049 ( .A1(n3668), .A2(n3894), .B1(n3667), .B2(n3205), .ZN(n3207)
         );
  OAI211_X1 U4050 ( .C1(n3699), .C2(n3208), .A(n3207), .B(n3206), .ZN(n3209)
         );
  AOI21_X1 U4051 ( .B1(n3210), .B2(n3703), .A(n3209), .ZN(n3211) );
  OAI21_X1 U4052 ( .B1(n3212), .B2(n3706), .A(n3211), .ZN(U3218) );
  XOR2_X1 U4053 ( .A(n3214), .B(n3213), .Z(n3215) );
  NAND2_X1 U4054 ( .A1(n3215), .A2(n3713), .ZN(n3221) );
  INV_X1 U4055 ( .A(n3216), .ZN(n3308) );
  OAI22_X1 U4056 ( .A1(n3717), .A2(n3217), .B1(n3308), .B2(n3715), .ZN(n3218)
         );
  AOI211_X1 U4057 ( .C1(n3240), .C2(n3719), .A(n3219), .B(n3218), .ZN(n3220)
         );
  OAI211_X1 U4058 ( .C1(n3722), .C2(n3247), .A(n3221), .B(n3220), .ZN(U3210)
         );
  INV_X1 U4059 ( .A(n3222), .ZN(n3229) );
  OAI22_X1 U4060 ( .A1(n4313), .A2(n3223), .B1(n3573), .B2(n4299), .ZN(n3224)
         );
  AOI21_X1 U4061 ( .B1(n3225), .B2(n4503), .A(n3224), .ZN(n3228) );
  NAND2_X1 U4062 ( .A1(n3226), .A2(n4257), .ZN(n3227) );
  OAI211_X1 U4063 ( .C1(n3229), .C2(n4515), .A(n3228), .B(n3227), .ZN(U3280)
         );
  INV_X1 U4064 ( .A(n3230), .ZN(n3238) );
  OAI22_X1 U4065 ( .A1(n4313), .A2(n3232), .B1(n3231), .B2(n4299), .ZN(n3233)
         );
  AOI21_X1 U4066 ( .B1(n3234), .B2(n4503), .A(n3233), .ZN(n3237) );
  NAND2_X1 U4067 ( .A1(n3235), .A2(n4257), .ZN(n3236) );
  OAI211_X1 U4068 ( .C1(n3238), .C2(n4515), .A(n3237), .B(n3236), .ZN(U3282)
         );
  INV_X1 U4069 ( .A(n3820), .ZN(n3762) );
  XNOR2_X1 U4070 ( .A(n3239), .B(n3762), .ZN(n3243) );
  AOI22_X1 U4071 ( .A1(n4308), .A2(n3895), .B1(n4306), .B2(n3240), .ZN(n3241)
         );
  OAI21_X1 U4072 ( .B1(n3308), .B2(n4311), .A(n3241), .ZN(n3242) );
  AOI21_X1 U4073 ( .B1(n3243), .B2(n4304), .A(n3242), .ZN(n4551) );
  OAI211_X1 U4074 ( .C1(n3246), .C2(n3245), .A(n4544), .B(n3244), .ZN(n4550)
         );
  INV_X1 U4075 ( .A(n4550), .ZN(n3249) );
  OAI22_X1 U4076 ( .A1(n4313), .A2(n2398), .B1(n3247), .B2(n4299), .ZN(n3248)
         );
  AOI21_X1 U4077 ( .B1(n3249), .B2(n4252), .A(n3248), .ZN(n3257) );
  NAND2_X1 U4078 ( .A1(n2997), .A2(n3895), .ZN(n3251) );
  NAND2_X1 U4079 ( .A1(n3251), .A2(n3250), .ZN(n3253) );
  OR2_X1 U4080 ( .A1(n2997), .A2(n3895), .ZN(n3252) );
  AND2_X1 U4081 ( .A1(n3253), .A2(n3252), .ZN(n3254) );
  NAND2_X1 U4082 ( .A1(n3254), .A2(n3820), .ZN(n4548) );
  INV_X1 U4083 ( .A(n3254), .ZN(n3255) );
  NAND2_X1 U4084 ( .A1(n3255), .A2(n3762), .ZN(n4546) );
  NAND3_X1 U4085 ( .A1(n4548), .A2(n4257), .A3(n4546), .ZN(n3256) );
  OAI211_X1 U4086 ( .C1(n4551), .C2(n4515), .A(n3257), .B(n3256), .ZN(U3283)
         );
  INV_X1 U4087 ( .A(n3258), .ZN(n3259) );
  OAI22_X1 U4088 ( .A1(n3259), .A2(n4272), .B1(n3313), .B2(n4299), .ZN(n3262)
         );
  MUX2_X1 U4089 ( .A(REG2_REG_9__SCAN_IN), .B(n3260), .S(n4313), .Z(n3261) );
  AOI211_X1 U4090 ( .C1(n4257), .C2(n3263), .A(n3262), .B(n3261), .ZN(n3264)
         );
  INV_X1 U4091 ( .A(n3264), .ZN(U3281) );
  INV_X1 U4092 ( .A(n3265), .ZN(n3271) );
  INV_X1 U4093 ( .A(n3266), .ZN(n3267) );
  AOI22_X1 U4094 ( .A1(n4515), .A2(REG2_REG_6__SCAN_IN), .B1(n3267), .B2(n4510), .ZN(n3268) );
  OAI21_X1 U4095 ( .B1(n4272), .B2(n3269), .A(n3268), .ZN(n3270) );
  AOI21_X1 U4096 ( .B1(n3271), .B2(n4257), .A(n3270), .ZN(n3272) );
  OAI21_X1 U4097 ( .B1(n4515), .B2(n3273), .A(n3272), .ZN(U3284) );
  NAND2_X1 U4098 ( .A1(n3326), .A2(n3324), .ZN(n3783) );
  INV_X1 U4099 ( .A(n3274), .ZN(n3276) );
  OAI21_X1 U4100 ( .B1(n3277), .B2(n3276), .A(n3275), .ZN(n3327) );
  XOR2_X1 U4101 ( .A(n3783), .B(n3327), .Z(n3281) );
  OAI22_X1 U4102 ( .A1(n3622), .A2(n4263), .B1(n4262), .B2(n3278), .ZN(n3279)
         );
  AOI21_X1 U4103 ( .B1(n4266), .B2(n3890), .A(n3279), .ZN(n3280) );
  OAI21_X1 U4104 ( .B1(n3281), .B2(n4268), .A(n3280), .ZN(n4392) );
  INV_X1 U4105 ( .A(n4392), .ZN(n3289) );
  XNOR2_X1 U4106 ( .A(n3282), .B(n3783), .ZN(n4393) );
  NAND2_X1 U4107 ( .A1(n3283), .A2(n3624), .ZN(n3284) );
  NAND2_X1 U4108 ( .A1(n3334), .A2(n3284), .ZN(n4454) );
  INV_X1 U4109 ( .A(n3627), .ZN(n3285) );
  AOI22_X1 U4110 ( .A1(n4515), .A2(REG2_REG_12__SCAN_IN), .B1(n3285), .B2(
        n4510), .ZN(n3286) );
  OAI21_X1 U4111 ( .B1(n4454), .B2(n4272), .A(n3286), .ZN(n3287) );
  AOI21_X1 U4112 ( .B1(n4393), .B2(n4257), .A(n3287), .ZN(n3288) );
  OAI21_X1 U4113 ( .B1(n3289), .B2(n4515), .A(n3288), .ZN(U3278) );
  XNOR2_X1 U4114 ( .A(n3727), .B(n3294), .ZN(n3292) );
  OAI22_X1 U4115 ( .A1(n3621), .A2(n4263), .B1(n3557), .B2(n4262), .ZN(n3290)
         );
  AOI21_X1 U4116 ( .B1(n4266), .B2(n4291), .A(n3290), .ZN(n3291) );
  OAI21_X1 U4117 ( .B1(n3292), .B2(n4268), .A(n3291), .ZN(n4383) );
  INV_X1 U4118 ( .A(n4383), .ZN(n3301) );
  OAI21_X1 U4119 ( .B1(n3295), .B2(n3294), .A(n3293), .ZN(n4384) );
  INV_X1 U4120 ( .A(n3336), .ZN(n3297) );
  INV_X1 U4121 ( .A(n4298), .ZN(n3296) );
  OAI21_X1 U4122 ( .B1(n3297), .B2(n3557), .A(n3296), .ZN(n4445) );
  AOI22_X1 U4123 ( .A1(n4515), .A2(REG2_REG_14__SCAN_IN), .B1(n3559), .B2(
        n4510), .ZN(n3298) );
  OAI21_X1 U4124 ( .B1(n4445), .B2(n4272), .A(n3298), .ZN(n3299) );
  AOI21_X1 U4125 ( .B1(n4384), .B2(n4257), .A(n3299), .ZN(n3300) );
  OAI21_X1 U4126 ( .B1(n4515), .B2(n3301), .A(n3300), .ZN(U3276) );
  AOI22_X1 U4127 ( .A1(n2007), .A2(n3894), .B1(n3456), .B2(n3310), .ZN(n3304)
         );
  XNOR2_X1 U4128 ( .A(n3304), .B(n3506), .ZN(n3342) );
  AOI22_X1 U4129 ( .A1(n2011), .A2(n3894), .B1(n3310), .B2(n2007), .ZN(n3341)
         );
  XNOR2_X1 U4130 ( .A(n3342), .B(n3341), .ZN(n3343) );
  XNOR2_X1 U4131 ( .A(n3344), .B(n3343), .ZN(n3305) );
  NAND2_X1 U4132 ( .A1(n3305), .A2(n3713), .ZN(n3312) );
  NOR2_X1 U4133 ( .A1(n3306), .A2(STATE_REG_SCAN_IN), .ZN(n3927) );
  OAI22_X1 U4134 ( .A1(n3717), .A2(n3308), .B1(n3307), .B2(n3715), .ZN(n3309)
         );
  AOI211_X1 U4135 ( .C1(n3310), .C2(n3719), .A(n3927), .B(n3309), .ZN(n3311)
         );
  OAI211_X1 U4136 ( .C1(n3722), .C2(n3313), .A(n3312), .B(n3311), .ZN(U3228)
         );
  INV_X1 U4137 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3316) );
  AOI21_X1 U4138 ( .B1(n4537), .B2(n3315), .A(n3314), .ZN(n3318) );
  MUX2_X1 U4139 ( .A(n3316), .B(n3318), .S(n4553), .Z(n3317) );
  OAI21_X1 U4140 ( .B1(n3320), .B2(n4453), .A(n3317), .ZN(U3489) );
  MUX2_X1 U4141 ( .A(n3954), .B(n3318), .S(n4561), .Z(n3319) );
  OAI21_X1 U4142 ( .B1(n4395), .B2(n3320), .A(n3319), .ZN(U3529) );
  AND2_X1 U4143 ( .A1(n3322), .A2(n3321), .ZN(n3772) );
  XNOR2_X1 U4144 ( .A(n3323), .B(n3772), .ZN(n4389) );
  INV_X1 U4145 ( .A(n4307), .ZN(n3716) );
  INV_X1 U4146 ( .A(n3324), .ZN(n3325) );
  AOI21_X1 U4147 ( .B1(n3327), .B2(n3326), .A(n3325), .ZN(n3328) );
  XNOR2_X1 U4148 ( .A(n3328), .B(n3772), .ZN(n3329) );
  NAND2_X1 U4149 ( .A1(n3329), .A2(n4304), .ZN(n3331) );
  AOI22_X1 U4150 ( .A1(n4308), .A2(n3891), .B1(n4306), .B2(n3378), .ZN(n3330)
         );
  OAI211_X1 U4151 ( .C1(n3716), .C2(n4311), .A(n3331), .B(n3330), .ZN(n3332)
         );
  AOI21_X1 U4152 ( .B1(n3333), .B2(n4389), .A(n3332), .ZN(n4387) );
  NAND2_X1 U4153 ( .A1(n3334), .A2(n3378), .ZN(n3335) );
  NAND2_X1 U4154 ( .A1(n3336), .A2(n3335), .ZN(n4449) );
  INV_X1 U4155 ( .A(n3337), .ZN(n3672) );
  AOI22_X1 U4156 ( .A1(n4515), .A2(REG2_REG_13__SCAN_IN), .B1(n3672), .B2(
        n4510), .ZN(n3338) );
  OAI21_X1 U4157 ( .B1(n4449), .B2(n4272), .A(n3338), .ZN(n3339) );
  AOI21_X1 U4158 ( .B1(n4389), .B2(n4512), .A(n3339), .ZN(n3340) );
  OAI21_X1 U4159 ( .B1(n4387), .B2(n4515), .A(n3340), .ZN(U3277) );
  NAND2_X1 U4160 ( .A1(n3372), .A2(n3893), .ZN(n3346) );
  NAND2_X1 U4161 ( .A1(n3456), .A2(n3348), .ZN(n3345) );
  NAND2_X1 U4162 ( .A1(n3346), .A2(n3345), .ZN(n3347) );
  XNOR2_X1 U4163 ( .A(n3347), .B(n3506), .ZN(n3350) );
  AOI22_X1 U4164 ( .A1(n2011), .A2(n3893), .B1(n3348), .B2(n2007), .ZN(n3352)
         );
  XOR2_X1 U4165 ( .A(n3350), .B(n3352), .Z(n3580) );
  INV_X1 U4166 ( .A(n3350), .ZN(n3351) );
  NAND2_X1 U4167 ( .A1(n3577), .A2(n2279), .ZN(n3365) );
  OAI22_X1 U4168 ( .A1(n3509), .A2(n3622), .B1(n3505), .B2(n3357), .ZN(n3364)
         );
  AOI22_X1 U4169 ( .A1(n2007), .A2(n3892), .B1(n3456), .B2(n3353), .ZN(n3354)
         );
  XOR2_X1 U4170 ( .A(n3506), .B(n3354), .Z(n3367) );
  XOR2_X1 U4171 ( .A(n3364), .B(n3367), .Z(n3355) );
  XNOR2_X1 U4172 ( .A(n3365), .B(n3355), .ZN(n3361) );
  AOI22_X1 U4173 ( .A1(n3668), .A2(n3891), .B1(n3667), .B2(n3893), .ZN(n3356)
         );
  NAND2_X1 U4174 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3939) );
  OAI211_X1 U4175 ( .C1(n3699), .C2(n3357), .A(n3356), .B(n3939), .ZN(n3358)
         );
  AOI21_X1 U4176 ( .B1(n3359), .B2(n3703), .A(n3358), .ZN(n3360) );
  OAI21_X1 U4177 ( .B1(n3361), .B2(n3706), .A(n3360), .ZN(U3233) );
  OAI22_X1 U4178 ( .A1(n2548), .A2(n3509), .B1(n3505), .B2(n3362), .ZN(n3417)
         );
  INV_X1 U4179 ( .A(n3417), .ZN(n3685) );
  NOR2_X1 U4180 ( .A1(n3365), .A2(n3364), .ZN(n3363) );
  INV_X1 U4181 ( .A(n3363), .ZN(n3368) );
  NAND2_X1 U4182 ( .A1(n3372), .A2(n3891), .ZN(n3370) );
  NAND2_X1 U4183 ( .A1(n3456), .A2(n3624), .ZN(n3369) );
  NAND2_X1 U4184 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  XNOR2_X1 U4185 ( .A(n3371), .B(n2934), .ZN(n3375) );
  INV_X1 U4186 ( .A(n3375), .ZN(n3374) );
  AOI22_X1 U4187 ( .A1(n2011), .A2(n3891), .B1(n3372), .B2(n3624), .ZN(n3376)
         );
  INV_X1 U4188 ( .A(n3376), .ZN(n3373) );
  AND2_X1 U4189 ( .A1(n3376), .A2(n3375), .ZN(n3617) );
  OAI22_X1 U4190 ( .A1(n3621), .A2(n3505), .B1(n2932), .B2(n3670), .ZN(n3377)
         );
  XNOR2_X1 U4191 ( .A(n3377), .B(n2934), .ZN(n3552) );
  OR2_X1 U4192 ( .A1(n3509), .A2(n3621), .ZN(n3380) );
  NAND2_X1 U4193 ( .A1(n3372), .A2(n3378), .ZN(n3379) );
  NAND2_X1 U4194 ( .A1(n3372), .A2(n4307), .ZN(n3382) );
  NAND2_X1 U4195 ( .A1(n3456), .A2(n3384), .ZN(n3381) );
  NAND2_X1 U4196 ( .A1(n3382), .A2(n3381), .ZN(n3383) );
  XNOR2_X1 U4197 ( .A(n3383), .B(n2934), .ZN(n3397) );
  INV_X1 U4198 ( .A(n3397), .ZN(n3388) );
  OR2_X1 U4199 ( .A1(n3509), .A2(n3716), .ZN(n3386) );
  NAND2_X1 U4200 ( .A1(n3372), .A2(n3384), .ZN(n3385) );
  INV_X1 U4201 ( .A(n3396), .ZN(n3387) );
  NAND2_X1 U4202 ( .A1(n3388), .A2(n3387), .ZN(n3630) );
  OAI21_X1 U4203 ( .B1(n3552), .B2(n3664), .A(n3630), .ZN(n3401) );
  NAND2_X1 U4204 ( .A1(n2011), .A2(n4291), .ZN(n3390) );
  NAND2_X1 U4205 ( .A1(n3372), .A2(n4305), .ZN(n3389) );
  NAND2_X1 U4206 ( .A1(n3390), .A2(n3389), .ZN(n3711) );
  NAND2_X1 U4207 ( .A1(n4291), .A2(n3372), .ZN(n3392) );
  NAND2_X1 U4208 ( .A1(n3456), .A2(n4305), .ZN(n3391) );
  NAND2_X1 U4209 ( .A1(n3392), .A2(n3391), .ZN(n3393) );
  XNOR2_X1 U4210 ( .A(n3393), .B(n3506), .ZN(n3634) );
  OAI22_X1 U4211 ( .A1(n4312), .A2(n3505), .B1(n2932), .B2(n3640), .ZN(n3394)
         );
  XNOR2_X1 U4212 ( .A(n3394), .B(n2934), .ZN(n3402) );
  NOR2_X1 U4213 ( .A1(n3505), .A2(n3640), .ZN(n3395) );
  AOI21_X1 U4214 ( .B1(n3648), .B2(n2011), .A(n3395), .ZN(n3403) );
  NAND2_X1 U4215 ( .A1(n3402), .A2(n3403), .ZN(n3406) );
  NAND2_X1 U4216 ( .A1(n3397), .A2(n3396), .ZN(n3631) );
  OAI211_X1 U4217 ( .C1(n3711), .C2(n3634), .A(n3406), .B(n3631), .ZN(n3398)
         );
  INV_X1 U4218 ( .A(n3398), .ZN(n3400) );
  NAND3_X1 U4219 ( .A1(n3552), .A2(n3630), .A3(n3664), .ZN(n3399) );
  INV_X1 U4220 ( .A(n3402), .ZN(n3405) );
  INV_X1 U4221 ( .A(n3403), .ZN(n3404) );
  AND2_X1 U4222 ( .A1(n3405), .A2(n3404), .ZN(n3628) );
  AOI21_X1 U4223 ( .B1(n3711), .B2(n3634), .A(n3628), .ZN(n3407) );
  INV_X1 U4224 ( .A(n3406), .ZN(n3629) );
  OAI22_X1 U4225 ( .A1(n4294), .A2(n3505), .B1(n2932), .B2(n4271), .ZN(n3409)
         );
  XNOR2_X1 U4226 ( .A(n3409), .B(n2934), .ZN(n3414) );
  OR2_X1 U4227 ( .A1(n4294), .A2(n3509), .ZN(n3412) );
  NAND2_X1 U4228 ( .A1(n3372), .A2(n3410), .ZN(n3411) );
  NOR2_X1 U4229 ( .A1(n3414), .A2(n3413), .ZN(n3645) );
  INV_X1 U4230 ( .A(n3684), .ZN(n3419) );
  AOI22_X1 U4231 ( .A1(n4265), .A2(n3372), .B1(n3456), .B2(n2274), .ZN(n3416)
         );
  XOR2_X1 U4232 ( .A(n3506), .B(n3416), .Z(n3686) );
  INV_X1 U4233 ( .A(n3587), .ZN(n3428) );
  NAND2_X1 U4234 ( .A1(n4244), .A2(n2007), .ZN(n3422) );
  NAND2_X1 U4235 ( .A1(n3456), .A2(n3420), .ZN(n3421) );
  NAND2_X1 U4236 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  XNOR2_X1 U4237 ( .A(n3423), .B(n2934), .ZN(n3426) );
  NOR2_X1 U4238 ( .A1(n3505), .A2(n4235), .ZN(n3424) );
  AOI21_X1 U4239 ( .B1(n4244), .B2(n2011), .A(n3424), .ZN(n3425) );
  NAND2_X1 U4240 ( .A1(n3426), .A2(n3425), .ZN(n3429) );
  OAI21_X1 U4241 ( .B1(n3426), .B2(n3425), .A(n3429), .ZN(n3588) );
  NAND2_X1 U4242 ( .A1(n3428), .A2(n3427), .ZN(n3585) );
  OAI22_X1 U4243 ( .A1(n4187), .A2(n3505), .B1(n2932), .B2(n3659), .ZN(n3430)
         );
  XNOR2_X1 U4244 ( .A(n3430), .B(n3506), .ZN(n3431) );
  OAI22_X1 U4245 ( .A1(n4187), .A2(n3509), .B1(n3505), .B2(n3659), .ZN(n3432)
         );
  NAND2_X1 U4246 ( .A1(n3431), .A2(n3432), .ZN(n3654) );
  INV_X1 U4247 ( .A(n3431), .ZN(n3434) );
  INV_X1 U4248 ( .A(n3432), .ZN(n3433) );
  NAND2_X1 U4249 ( .A1(n3434), .A2(n3433), .ZN(n3656) );
  NAND2_X1 U4250 ( .A1(n4171), .A2(n2007), .ZN(n3436) );
  NAND2_X1 U4251 ( .A1(n3456), .A2(n3611), .ZN(n3435) );
  NAND2_X1 U4252 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  XNOR2_X1 U4253 ( .A(n3437), .B(n2934), .ZN(n3439) );
  NOR2_X1 U4254 ( .A1(n3505), .A2(n4194), .ZN(n3438) );
  AOI21_X1 U4255 ( .B1(n4171), .B2(n2011), .A(n3438), .ZN(n3440) );
  NAND2_X1 U4256 ( .A1(n3439), .A2(n3440), .ZN(n3606) );
  INV_X1 U4257 ( .A(n3439), .ZN(n3442) );
  INV_X1 U4258 ( .A(n3440), .ZN(n3441) );
  NAND2_X1 U4259 ( .A1(n3442), .A2(n3441), .ZN(n3605) );
  OAI22_X1 U4260 ( .A1(n4151), .A2(n3505), .B1(n4179), .B2(n2932), .ZN(n3443)
         );
  XNOR2_X1 U4261 ( .A(n3443), .B(n3506), .ZN(n3446) );
  OAI22_X1 U4262 ( .A1(n4151), .A2(n3509), .B1(n4179), .B2(n3505), .ZN(n3445)
         );
  XNOR2_X1 U4263 ( .A(n3446), .B(n3445), .ZN(n3677) );
  OAI22_X1 U4264 ( .A1(n4173), .A2(n3505), .B1(n2932), .B2(n4156), .ZN(n3444)
         );
  XNOR2_X1 U4265 ( .A(n3444), .B(n3506), .ZN(n3449) );
  OAI22_X1 U4266 ( .A1(n4173), .A2(n3509), .B1(n3505), .B2(n4156), .ZN(n3448)
         );
  XNOR2_X1 U4267 ( .A(n3449), .B(n3448), .ZN(n3563) );
  NOR2_X1 U4268 ( .A1(n3446), .A2(n3445), .ZN(n3564) );
  NOR2_X1 U4269 ( .A1(n3563), .A2(n3564), .ZN(n3447) );
  NAND2_X1 U4270 ( .A1(n3449), .A2(n3448), .ZN(n3452) );
  NOR2_X1 U4271 ( .A1(n3505), .A2(n4137), .ZN(n3450) );
  AOI21_X1 U4272 ( .B1(n4153), .B2(n2011), .A(n3450), .ZN(n3490) );
  NAND2_X1 U4273 ( .A1(n3452), .A2(n3490), .ZN(n3484) );
  INV_X1 U4274 ( .A(n3484), .ZN(n3451) );
  INV_X1 U4275 ( .A(n3472), .ZN(n3454) );
  INV_X1 U4276 ( .A(n3452), .ZN(n3485) );
  INV_X1 U4277 ( .A(n3490), .ZN(n3453) );
  NAND2_X1 U4278 ( .A1(n3454), .A2(n3471), .ZN(n3460) );
  NAND2_X1 U4279 ( .A1(n4153), .A2(n3372), .ZN(n3458) );
  NAND2_X1 U4280 ( .A1(n3456), .A2(n3455), .ZN(n3457) );
  NAND2_X1 U4281 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  XNOR2_X1 U4282 ( .A(n3459), .B(n3506), .ZN(n3493) );
  XNOR2_X1 U4283 ( .A(n3460), .B(n3493), .ZN(n3461) );
  NAND2_X1 U4284 ( .A1(n3461), .A2(n3713), .ZN(n3466) );
  OAI22_X1 U4285 ( .A1(n3699), .A2(n4137), .B1(STATE_REG_SCAN_IN), .B2(n3462), 
        .ZN(n3464) );
  OAI22_X1 U4286 ( .A1(n4092), .A2(n3715), .B1(n4173), .B2(n3717), .ZN(n3463)
         );
  AOI211_X1 U4287 ( .C1(n4139), .C2(n3703), .A(n3464), .B(n3463), .ZN(n3465)
         );
  NAND2_X1 U4288 ( .A1(n3466), .A2(n3465), .ZN(U3226) );
  NAND3_X1 U4289 ( .A1(n3468), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3470) );
  INV_X1 U4290 ( .A(DATAI_31_), .ZN(n3469) );
  OAI22_X1 U4291 ( .A1(n3467), .A2(n3470), .B1(STATE_REG_SCAN_IN), .B2(n3469), 
        .ZN(U3321) );
  INV_X1 U4292 ( .A(n3493), .ZN(n3489) );
  OAI22_X1 U4293 ( .A1(n4092), .A2(n3505), .B1(n2932), .B2(n4119), .ZN(n3473)
         );
  XNOR2_X1 U4294 ( .A(n3473), .B(n3506), .ZN(n3495) );
  NAND2_X1 U4295 ( .A1(n4132), .A2(n2011), .ZN(n3475) );
  OR2_X1 U4296 ( .A1(n3508), .A2(n4119), .ZN(n3474) );
  NAND2_X1 U4297 ( .A1(n3475), .A2(n3474), .ZN(n3488) );
  NAND2_X1 U4298 ( .A1(n3495), .A2(n3488), .ZN(n3487) );
  OAI21_X1 U4299 ( .B1(n3495), .B2(n3488), .A(n3487), .ZN(n3476) );
  XNOR2_X1 U4300 ( .A(n3477), .B(n3476), .ZN(n3478) );
  NAND2_X1 U4301 ( .A1(n3478), .A2(n3713), .ZN(n3483) );
  OAI22_X1 U4302 ( .A1(n3699), .A2(n4119), .B1(STATE_REG_SCAN_IN), .B2(n3479), 
        .ZN(n3481) );
  OAI22_X1 U4303 ( .A1(n4074), .A2(n3715), .B1(n4117), .B2(n3717), .ZN(n3480)
         );
  AOI211_X1 U4304 ( .C1(n4121), .C2(n3703), .A(n3481), .B(n3480), .ZN(n3482)
         );
  NAND2_X1 U4305 ( .A1(n3483), .A2(n3482), .ZN(U3222) );
  OAI21_X1 U4306 ( .B1(n3485), .B2(n3493), .A(n3484), .ZN(n3486) );
  NAND3_X1 U4307 ( .A1(n3565), .A2(n3487), .A3(n3486), .ZN(n3694) );
  INV_X1 U4308 ( .A(n3488), .ZN(n3491) );
  AOI21_X1 U4309 ( .B1(n3489), .B2(n3490), .A(n3491), .ZN(n3494) );
  NAND2_X1 U4310 ( .A1(n3491), .A2(n3490), .ZN(n3492) );
  OAI22_X1 U4311 ( .A1(n3495), .A2(n3494), .B1(n3493), .B2(n3492), .ZN(n3496)
         );
  INV_X1 U4312 ( .A(n3496), .ZN(n3693) );
  OAI22_X1 U4313 ( .A1(n4074), .A2(n3505), .B1(n2932), .B2(n4099), .ZN(n3497)
         );
  XNOR2_X1 U4314 ( .A(n3497), .B(n3506), .ZN(n3502) );
  OAI22_X1 U4315 ( .A1(n4074), .A2(n3509), .B1(n3505), .B2(n4099), .ZN(n3501)
         );
  OR2_X1 U4316 ( .A1(n3502), .A2(n3501), .ZN(n3696) );
  AND2_X1 U4317 ( .A1(n3693), .A2(n3696), .ZN(n3540) );
  OAI22_X1 U4318 ( .A1(n3700), .A2(n3505), .B1(n4080), .B2(n2932), .ZN(n3498)
         );
  XNOR2_X1 U4319 ( .A(n3498), .B(n3506), .ZN(n3513) );
  OAI22_X1 U4320 ( .A1(n3700), .A2(n3509), .B1(n4080), .B2(n3505), .ZN(n3512)
         );
  XNOR2_X1 U4321 ( .A(n3513), .B(n3512), .ZN(n3541) );
  INV_X1 U4322 ( .A(n3541), .ZN(n3499) );
  AND2_X1 U4323 ( .A1(n3540), .A2(n3499), .ZN(n3500) );
  NAND2_X1 U4324 ( .A1(n3694), .A2(n3500), .ZN(n3504) );
  NAND2_X1 U4325 ( .A1(n3502), .A2(n3501), .ZN(n3695) );
  OR2_X1 U4326 ( .A1(n3541), .A2(n3695), .ZN(n3503) );
  NAND2_X1 U4327 ( .A1(n3504), .A2(n3503), .ZN(n3526) );
  INV_X1 U4328 ( .A(n3526), .ZN(n3515) );
  OAI22_X1 U4329 ( .A1(n4066), .A2(n3505), .B1(n2932), .B2(n3519), .ZN(n3507)
         );
  XNOR2_X1 U4330 ( .A(n3507), .B(n3506), .ZN(n3511) );
  OAI22_X1 U4331 ( .A1(n4066), .A2(n3509), .B1(n3508), .B2(n3519), .ZN(n3510)
         );
  XNOR2_X1 U4332 ( .A(n3511), .B(n3510), .ZN(n3525) );
  INV_X1 U4333 ( .A(n3525), .ZN(n3514) );
  NAND2_X1 U4334 ( .A1(n3513), .A2(n3512), .ZN(n3516) );
  NAND4_X1 U4335 ( .A1(n3515), .A2(n3713), .A3(n3514), .A4(n3516), .ZN(n3529)
         );
  INV_X1 U4336 ( .A(n3516), .ZN(n3517) );
  NAND3_X1 U4337 ( .A1(n3525), .A2(n3713), .A3(n3517), .ZN(n3524) );
  INV_X1 U4338 ( .A(n3532), .ZN(n3522) );
  OAI22_X1 U4339 ( .A1(n3699), .A2(n3519), .B1(STATE_REG_SCAN_IN), .B2(n3518), 
        .ZN(n3521) );
  OAI22_X1 U4340 ( .A1(n3799), .A2(n3715), .B1(n3700), .B2(n3717), .ZN(n3520)
         );
  AOI211_X1 U4341 ( .C1(n3522), .C2(n3703), .A(n3521), .B(n3520), .ZN(n3523)
         );
  AND2_X1 U4342 ( .A1(n3524), .A2(n3523), .ZN(n3528) );
  NAND3_X1 U4343 ( .A1(n3526), .A2(n3713), .A3(n3525), .ZN(n3527) );
  NAND3_X1 U4344 ( .A1(n3529), .A2(n3528), .A3(n3527), .ZN(U3217) );
  INV_X1 U4345 ( .A(n3530), .ZN(n3536) );
  INV_X1 U4346 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3531) );
  OAI22_X1 U4347 ( .A1(n3532), .A2(n4299), .B1(n3531), .B2(n4313), .ZN(n3535)
         );
  NOR2_X1 U4348 ( .A1(n3533), .A2(n4515), .ZN(n3534) );
  AOI211_X1 U4349 ( .C1(n4503), .C2(n3536), .A(n3535), .B(n3534), .ZN(n3537)
         );
  OAI21_X1 U4350 ( .B1(n3538), .B2(n4316), .A(n3537), .ZN(U3262) );
  XNOR2_X1 U4351 ( .A(n3542), .B(n3541), .ZN(n3550) );
  NAND2_X1 U4352 ( .A1(n3719), .A2(n3543), .ZN(n3544) );
  OAI21_X1 U4353 ( .B1(STATE_REG_SCAN_IN), .B2(n3545), .A(n3544), .ZN(n3546)
         );
  AOI21_X1 U4354 ( .B1(n4114), .B2(n3667), .A(n3546), .ZN(n3547) );
  OAI21_X1 U4355 ( .B1(n4066), .B2(n3715), .A(n3547), .ZN(n3548) );
  AOI21_X1 U4356 ( .B1(n4081), .B2(n3703), .A(n3548), .ZN(n3549) );
  OAI21_X1 U4357 ( .B1(n3550), .B2(n3706), .A(n3549), .ZN(U3211) );
  NAND2_X1 U4358 ( .A1(n3630), .A2(n3631), .ZN(n3555) );
  INV_X1 U4359 ( .A(n3552), .ZN(n3665) );
  NOR2_X1 U4360 ( .A1(n3551), .A2(n3665), .ZN(n3554) );
  INV_X1 U4361 ( .A(n3551), .ZN(n3553) );
  OAI22_X1 U4362 ( .A1(n3554), .A2(n3664), .B1(n3553), .B2(n3552), .ZN(n3633)
         );
  XOR2_X1 U4363 ( .A(n3555), .B(n3633), .Z(n3561) );
  AOI22_X1 U4364 ( .A1(n3668), .A2(n4291), .B1(n3667), .B2(n3890), .ZN(n3556)
         );
  NAND2_X1 U4365 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n3991) );
  OAI211_X1 U4366 ( .C1(n3699), .C2(n3557), .A(n3556), .B(n3991), .ZN(n3558)
         );
  AOI21_X1 U4367 ( .B1(n3559), .B2(n3703), .A(n3558), .ZN(n3560) );
  OAI21_X1 U4368 ( .B1(n3561), .B2(n3706), .A(n3560), .ZN(U3212) );
  INV_X1 U4369 ( .A(n3562), .ZN(n3676) );
  OAI21_X1 U4370 ( .B1(n3676), .B2(n3564), .A(n3563), .ZN(n3566) );
  NAND3_X1 U4371 ( .A1(n3566), .A2(n3713), .A3(n3565), .ZN(n3572) );
  OAI22_X1 U4372 ( .A1(n3699), .A2(n4156), .B1(STATE_REG_SCAN_IN), .B2(n3567), 
        .ZN(n3569) );
  OAI22_X1 U4373 ( .A1(n4117), .A2(n3715), .B1(n4151), .B2(n3717), .ZN(n3568)
         );
  AOI211_X1 U4374 ( .C1(n3570), .C2(n3703), .A(n3569), .B(n3568), .ZN(n3571)
         );
  NAND2_X1 U4375 ( .A1(n3572), .A2(n3571), .ZN(U3213) );
  INV_X1 U4376 ( .A(n3573), .ZN(n3583) );
  AOI22_X1 U4377 ( .A1(n3668), .A2(n3892), .B1(n3667), .B2(n3894), .ZN(n3575)
         );
  OAI211_X1 U4378 ( .C1(n3699), .C2(n3576), .A(n3575), .B(n3574), .ZN(n3582)
         );
  INV_X1 U4379 ( .A(n3577), .ZN(n3578) );
  AOI211_X1 U4380 ( .C1(n3580), .C2(n3579), .A(n3706), .B(n3578), .ZN(n3581)
         );
  AOI211_X1 U4381 ( .C1(n3583), .C2(n3703), .A(n3582), .B(n3581), .ZN(n3584)
         );
  INV_X1 U4382 ( .A(n3584), .ZN(U3214) );
  INV_X1 U4383 ( .A(n3585), .ZN(n3586) );
  AOI21_X1 U4384 ( .B1(n3588), .B2(n3587), .A(n3586), .ZN(n3593) );
  INV_X1 U4385 ( .A(n4237), .ZN(n3591) );
  AOI22_X1 U4386 ( .A1(n3668), .A2(n4231), .B1(n3667), .B2(n4265), .ZN(n3589)
         );
  NAND2_X1 U4387 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4033) );
  OAI211_X1 U4388 ( .C1(n3699), .C2(n4235), .A(n3589), .B(n4033), .ZN(n3590)
         );
  AOI21_X1 U4389 ( .B1(n3591), .B2(n3703), .A(n3590), .ZN(n3592) );
  OAI21_X1 U4390 ( .B1(n3593), .B2(n3706), .A(n3592), .ZN(U3216) );
  AOI22_X1 U4391 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3595), .B1(n3668), .B2(n3594), .ZN(n3604) );
  AOI22_X1 U4392 ( .A1(n3667), .A2(n2671), .B1(n3596), .B2(n3719), .ZN(n3603)
         );
  INV_X1 U4393 ( .A(n3598), .ZN(n3599) );
  AOI21_X1 U4394 ( .B1(n3597), .B2(n3599), .A(n3706), .ZN(n3601) );
  NAND2_X1 U4395 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  NAND3_X1 U4396 ( .A1(n3604), .A2(n3603), .A3(n3602), .ZN(U3219) );
  NAND2_X1 U4397 ( .A1(n3606), .A2(n3605), .ZN(n3610) );
  INV_X1 U4398 ( .A(n3656), .ZN(n3608) );
  OAI211_X1 U4399 ( .C1(n3607), .C2(n3608), .A(n3654), .B(n3610), .ZN(n3609)
         );
  OAI211_X1 U4400 ( .C1(n2042), .C2(n3610), .A(n3713), .B(n3609), .ZN(n3616)
         );
  AOI22_X1 U4401 ( .A1(n3719), .A2(n3611), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3615) );
  AOI22_X1 U4402 ( .A1(n4189), .A2(n3668), .B1(n3667), .B2(n4231), .ZN(n3614)
         );
  INV_X1 U4403 ( .A(n3612), .ZN(n4195) );
  NAND2_X1 U4404 ( .A1(n3703), .A2(n4195), .ZN(n3613) );
  NAND4_X1 U4405 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(U3220)
         );
  NOR2_X1 U4406 ( .A1(n2069), .A2(n3617), .ZN(n3618) );
  XNOR2_X1 U4407 ( .A(n3619), .B(n3618), .ZN(n3620) );
  NAND2_X1 U4408 ( .A1(n3620), .A2(n3713), .ZN(n3626) );
  AND2_X1 U4409 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3959) );
  OAI22_X1 U4410 ( .A1(n3717), .A2(n3622), .B1(n3621), .B2(n3715), .ZN(n3623)
         );
  AOI211_X1 U4411 ( .C1(n3624), .C2(n3719), .A(n3959), .B(n3623), .ZN(n3625)
         );
  OAI211_X1 U4412 ( .C1(n3722), .C2(n3627), .A(n3626), .B(n3625), .ZN(U3221)
         );
  NOR2_X1 U4413 ( .A1(n3629), .A2(n3628), .ZN(n3638) );
  INV_X1 U4414 ( .A(n3630), .ZN(n3632) );
  OAI21_X1 U4415 ( .B1(n3633), .B2(n3632), .A(n3631), .ZN(n3636) );
  INV_X1 U4416 ( .A(n3634), .ZN(n3635) );
  NOR2_X1 U4417 ( .A1(n3636), .A2(n3635), .ZN(n3708) );
  NAND2_X1 U4418 ( .A1(n3636), .A2(n3635), .ZN(n3709) );
  OAI21_X1 U4419 ( .B1(n3708), .B2(n3711), .A(n3709), .ZN(n3637) );
  XOR2_X1 U4420 ( .A(n3638), .B(n3637), .Z(n3644) );
  INV_X1 U4421 ( .A(n4284), .ZN(n3642) );
  AOI22_X1 U4422 ( .A1(n3668), .A2(n3889), .B1(n3667), .B2(n4291), .ZN(n3639)
         );
  NAND2_X1 U4423 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4479) );
  OAI211_X1 U4424 ( .C1(n3699), .C2(n3640), .A(n3639), .B(n4479), .ZN(n3641)
         );
  AOI21_X1 U4425 ( .B1(n3642), .B2(n3703), .A(n3641), .ZN(n3643) );
  OAI21_X1 U4426 ( .B1(n3644), .B2(n3706), .A(n3643), .ZN(U3223) );
  NOR2_X1 U4427 ( .A1(n3645), .A2(n2288), .ZN(n3646) );
  XNOR2_X1 U4428 ( .A(n3647), .B(n3646), .ZN(n3652) );
  AOI22_X1 U4429 ( .A1(n3668), .A2(n4265), .B1(n3667), .B2(n3648), .ZN(n3649)
         );
  NAND2_X1 U4430 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4021) );
  OAI211_X1 U4431 ( .C1(n3699), .C2(n4271), .A(n3649), .B(n4021), .ZN(n3650)
         );
  AOI21_X1 U4432 ( .B1(n4273), .B2(n3703), .A(n3650), .ZN(n3651) );
  OAI21_X1 U4433 ( .B1(n3652), .B2(n3706), .A(n3651), .ZN(U3225) );
  INV_X1 U4434 ( .A(n3653), .ZN(n3657) );
  AOI21_X1 U4435 ( .B1(n3654), .B2(n3656), .A(n3607), .ZN(n3655) );
  AOI21_X1 U4436 ( .B1(n3657), .B2(n3656), .A(n3655), .ZN(n3663) );
  OAI22_X1 U4437 ( .A1(n3699), .A2(n3659), .B1(STATE_REG_SCAN_IN), .B2(n3658), 
        .ZN(n3661) );
  OAI22_X1 U4438 ( .A1(n3717), .A2(n3688), .B1(n4208), .B2(n3715), .ZN(n3660)
         );
  AOI211_X1 U4439 ( .C1(n4217), .C2(n3703), .A(n3661), .B(n3660), .ZN(n3662)
         );
  OAI21_X1 U4440 ( .B1(n3663), .B2(n3706), .A(n3662), .ZN(U3230) );
  XNOR2_X1 U4441 ( .A(n3665), .B(n3664), .ZN(n3666) );
  XNOR2_X1 U4442 ( .A(n3551), .B(n3666), .ZN(n3674) );
  AOI22_X1 U4443 ( .A1(n3668), .A2(n4307), .B1(n3667), .B2(n3891), .ZN(n3669)
         );
  NAND2_X1 U4444 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3976) );
  OAI211_X1 U4445 ( .C1(n3699), .C2(n3670), .A(n3669), .B(n3976), .ZN(n3671)
         );
  AOI21_X1 U4446 ( .B1(n3672), .B2(n3703), .A(n3671), .ZN(n3673) );
  OAI21_X1 U4447 ( .B1(n3674), .B2(n3706), .A(n3673), .ZN(U3231) );
  AOI21_X1 U4448 ( .B1(n3677), .B2(n3675), .A(n3676), .ZN(n3683) );
  INV_X1 U4449 ( .A(n4177), .ZN(n3681) );
  OAI22_X1 U4450 ( .A1(n3699), .A2(n4179), .B1(STATE_REG_SCAN_IN), .B2(n3678), 
        .ZN(n3680) );
  OAI22_X1 U4451 ( .A1(n4173), .A2(n3715), .B1(n4208), .B2(n3717), .ZN(n3679)
         );
  AOI211_X1 U4452 ( .C1(n3681), .C2(n3703), .A(n3680), .B(n3679), .ZN(n3682)
         );
  OAI21_X1 U4453 ( .B1(n3683), .B2(n3706), .A(n3682), .ZN(U3232) );
  XNOR2_X1 U4454 ( .A(n3686), .B(n3685), .ZN(n3687) );
  XNOR2_X1 U4455 ( .A(n3684), .B(n3687), .ZN(n3692) );
  AND2_X1 U4456 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4493) );
  OAI22_X1 U4457 ( .A1(n3717), .A2(n4294), .B1(n3688), .B2(n3715), .ZN(n3689)
         );
  AOI211_X1 U4458 ( .C1(n2274), .C2(n3719), .A(n4493), .B(n3689), .ZN(n3691)
         );
  NAND2_X1 U4459 ( .A1(n3703), .A2(n4253), .ZN(n3690) );
  OAI211_X1 U4460 ( .C1(n3692), .C2(n3706), .A(n3691), .B(n3690), .ZN(U3235)
         );
  NAND2_X1 U4461 ( .A1(n3694), .A2(n3693), .ZN(n3698) );
  NAND2_X1 U4462 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  XNOR2_X1 U4463 ( .A(n3698), .B(n3697), .ZN(n3707) );
  INV_X1 U4464 ( .A(n4102), .ZN(n3704) );
  OAI22_X1 U4465 ( .A1(n3699), .A2(n4099), .B1(STATE_REG_SCAN_IN), .B2(n4705), 
        .ZN(n3702) );
  OAI22_X1 U4466 ( .A1(n3700), .A2(n3715), .B1(n4092), .B2(n3717), .ZN(n3701)
         );
  AOI211_X1 U4467 ( .C1(n3704), .C2(n3703), .A(n3702), .B(n3701), .ZN(n3705)
         );
  OAI21_X1 U4468 ( .B1(n3707), .B2(n3706), .A(n3705), .ZN(U3237) );
  INV_X1 U4469 ( .A(n3708), .ZN(n3710) );
  NAND2_X1 U4470 ( .A1(n3710), .A2(n3709), .ZN(n3712) );
  XNOR2_X1 U4471 ( .A(n3712), .B(n3711), .ZN(n3714) );
  NAND2_X1 U4472 ( .A1(n3714), .A2(n3713), .ZN(n3721) );
  AND2_X1 U4473 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4472) );
  OAI22_X1 U4474 ( .A1(n3717), .A2(n3716), .B1(n4312), .B2(n3715), .ZN(n3718)
         );
  AOI211_X1 U4475 ( .C1(n4305), .C2(n3719), .A(n4472), .B(n3718), .ZN(n3720)
         );
  OAI211_X1 U4476 ( .C1(n3722), .C2(n4300), .A(n3721), .B(n3720), .ZN(U3238)
         );
  NAND2_X1 U4477 ( .A1(n3726), .A2(n3723), .ZN(n3845) );
  NAND2_X1 U4478 ( .A1(n3725), .A2(n3724), .ZN(n3829) );
  NAND2_X1 U4479 ( .A1(n3829), .A2(n3726), .ZN(n3844) );
  OAI21_X1 U4480 ( .B1(n3727), .B2(n3845), .A(n3844), .ZN(n3729) );
  INV_X1 U4481 ( .A(n3851), .ZN(n3728) );
  AOI211_X1 U4482 ( .C1(n3729), .C2(n3849), .A(n3728), .B(n3854), .ZN(n3730)
         );
  INV_X1 U4483 ( .A(n3730), .ZN(n3731) );
  AOI21_X1 U4484 ( .B1(n3731), .B2(n3853), .A(n3856), .ZN(n3733) );
  OAI21_X1 U4485 ( .B1(n3733), .B2(n3858), .A(n3732), .ZN(n3734) );
  AOI21_X1 U4486 ( .B1(n3734), .B2(n3861), .A(n4088), .ZN(n3752) );
  NAND2_X1 U4487 ( .A1(n3736), .A2(n3735), .ZN(n4060) );
  INV_X1 U4488 ( .A(n4060), .ZN(n3745) );
  NAND2_X1 U4489 ( .A1(n2009), .A2(DATAI_29_), .ZN(n3798) );
  INV_X1 U4490 ( .A(n3798), .ZN(n4062) );
  INV_X1 U4491 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4666) );
  INV_X1 U4492 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4678) );
  OR2_X1 U4493 ( .A1(n2357), .A2(n4678), .ZN(n3738) );
  NAND2_X1 U4494 ( .A1(n3739), .A2(REG1_REG_31__SCAN_IN), .ZN(n3737) );
  OAI211_X1 U4495 ( .C1(n3742), .C2(n4666), .A(n3738), .B(n3737), .ZN(n4041)
         );
  NAND2_X1 U4496 ( .A1(n2010), .A2(DATAI_31_), .ZN(n4042) );
  NAND2_X1 U4497 ( .A1(n4041), .A2(n4042), .ZN(n3871) );
  INV_X1 U4498 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U4499 ( .A1(n3739), .A2(REG1_REG_30__SCAN_IN), .ZN(n3741) );
  INV_X1 U4500 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4400) );
  OR2_X1 U4501 ( .A1(n2357), .A2(n4400), .ZN(n3740) );
  OAI211_X1 U4502 ( .C1(n3742), .C2(n4646), .A(n3741), .B(n3740), .ZN(n4063)
         );
  NAND2_X1 U4503 ( .A1(n2009), .A2(DATAI_30_), .ZN(n4048) );
  OR2_X1 U4504 ( .A1(n4063), .A2(n4048), .ZN(n3744) );
  NAND2_X1 U4505 ( .A1(n3871), .A2(n3744), .ZN(n3776) );
  AOI21_X1 U4506 ( .B1(n3799), .B2(n4062), .A(n3776), .ZN(n3748) );
  NAND3_X1 U4507 ( .A1(n3745), .A2(n3862), .A3(n3748), .ZN(n3751) );
  OR2_X1 U4508 ( .A1(n3799), .A2(n4062), .ZN(n3746) );
  AND2_X1 U4509 ( .A1(n4059), .A2(n3746), .ZN(n3866) );
  INV_X1 U4510 ( .A(n3866), .ZN(n3747) );
  NOR3_X1 U4511 ( .A1(n3747), .A2(n4076), .A3(n3758), .ZN(n3750) );
  NAND2_X1 U4512 ( .A1(n3866), .A2(n4060), .ZN(n3749) );
  NAND2_X1 U4513 ( .A1(n3749), .A2(n3748), .ZN(n3869) );
  OAI22_X1 U4514 ( .A1(n3752), .A2(n3751), .B1(n3750), .B2(n3869), .ZN(n3757)
         );
  INV_X1 U4515 ( .A(n4041), .ZN(n3754) );
  INV_X1 U4516 ( .A(n4048), .ZN(n3753) );
  NAND2_X1 U4517 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  NAND2_X1 U4518 ( .A1(n4063), .A2(n4048), .ZN(n3775) );
  AOI21_X1 U4519 ( .B1(n3775), .B2(n4041), .A(n4042), .ZN(n3755) );
  AOI21_X1 U4520 ( .B1(n3757), .B2(n3756), .A(n3755), .ZN(n3879) );
  INV_X1 U4521 ( .A(n3758), .ZN(n3760) );
  NAND2_X1 U4522 ( .A1(n3760), .A2(n3759), .ZN(n4090) );
  INV_X1 U4523 ( .A(n3857), .ZN(n4145) );
  NAND2_X1 U4524 ( .A1(n4145), .A2(n4146), .ZN(n4185) );
  NAND4_X1 U4525 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3768)
         );
  INV_X1 U4526 ( .A(n4249), .ZN(n3766) );
  INV_X1 U4527 ( .A(n4224), .ZN(n3765) );
  AND2_X1 U4528 ( .A1(n3765), .A2(n4223), .ZN(n4260) );
  NAND3_X1 U4529 ( .A1(n3766), .A2(n4260), .A3(n4288), .ZN(n3767) );
  NOR4_X1 U4530 ( .A1(n4164), .A2(n4185), .A3(n3768), .A4(n3767), .ZN(n3788)
         );
  XNOR2_X1 U4531 ( .A(n4187), .B(n4214), .ZN(n4200) );
  INV_X1 U4532 ( .A(n4200), .ZN(n4205) );
  NAND2_X1 U4533 ( .A1(n3770), .A2(n3769), .ZN(n4229) );
  NAND4_X1 U4534 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3777)
         );
  OAI21_X1 U4535 ( .B1(n4041), .B2(n4042), .A(n3775), .ZN(n3870) );
  NOR4_X1 U4536 ( .A1(n4229), .A2(n3777), .A3(n3776), .A4(n3870), .ZN(n3787)
         );
  NAND4_X1 U4537 ( .A1(n2049), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3785)
         );
  NAND2_X1 U4538 ( .A1(n3782), .A2(n3781), .ZN(n3784) );
  NAND4_X1 U4539 ( .A1(n3788), .A2(n4205), .A3(n3787), .A4(n3786), .ZN(n3792)
         );
  NAND2_X1 U4540 ( .A1(n4087), .A2(n3789), .ZN(n4110) );
  INV_X1 U4541 ( .A(n3790), .ZN(n4127) );
  NAND2_X1 U4542 ( .A1(n4127), .A2(n3791), .ZN(n4149) );
  NOR4_X1 U4543 ( .A1(n4090), .A2(n3792), .A3(n4110), .A4(n4149), .ZN(n3797)
         );
  INV_X1 U4544 ( .A(n4053), .ZN(n3796) );
  INV_X1 U4545 ( .A(n4076), .ZN(n3795) );
  INV_X1 U4546 ( .A(n4108), .ZN(n3793) );
  NOR2_X1 U4547 ( .A1(n3794), .A2(n3793), .ZN(n4130) );
  NAND4_X1 U4548 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n4130), .ZN(n3801)
         );
  XNOR2_X1 U4549 ( .A(n3799), .B(n3798), .ZN(n4323) );
  INV_X1 U4550 ( .A(n4323), .ZN(n4326) );
  OAI21_X1 U4551 ( .B1(n3801), .B2(n4326), .A(n3800), .ZN(n3876) );
  INV_X1 U4552 ( .A(n3802), .ZN(n3805) );
  OAI211_X1 U4553 ( .C1(n3805), .C2(n2695), .A(n3804), .B(n3803), .ZN(n3808)
         );
  NAND3_X1 U4554 ( .A1(n3808), .A2(n3807), .A3(n3806), .ZN(n3811) );
  NAND3_X1 U4555 ( .A1(n3811), .A2(n3810), .A3(n3809), .ZN(n3814) );
  NAND3_X1 U4556 ( .A1(n3814), .A2(n3813), .A3(n3812), .ZN(n3823) );
  INV_X1 U4557 ( .A(n3831), .ZN(n3818) );
  INV_X1 U4558 ( .A(n3815), .ZN(n3817) );
  NOR3_X1 U4559 ( .A1(n3818), .A2(n3817), .A3(n3816), .ZN(n3822) );
  INV_X1 U4560 ( .A(n3819), .ZN(n3821) );
  AOI211_X1 U4561 ( .C1(n3823), .C2(n3822), .A(n3821), .B(n3820), .ZN(n3828)
         );
  NAND2_X1 U4562 ( .A1(n3825), .A2(n3824), .ZN(n3833) );
  OAI211_X1 U4563 ( .C1(n3828), .C2(n3833), .A(n3827), .B(n3826), .ZN(n3837)
         );
  INV_X1 U4564 ( .A(n3829), .ZN(n3836) );
  INV_X1 U4565 ( .A(n3830), .ZN(n3832) );
  NAND2_X1 U4566 ( .A1(n3832), .A2(n3831), .ZN(n3834) );
  OAI21_X1 U4567 ( .B1(n3834), .B2(n3833), .A(n3838), .ZN(n3835) );
  AOI22_X1 U4568 ( .A1(n3837), .A2(n3836), .B1(n3844), .B2(n3835), .ZN(n3848)
         );
  INV_X1 U4569 ( .A(n3838), .ZN(n3842) );
  OAI211_X1 U4570 ( .C1(n3842), .C2(n3841), .A(n3840), .B(n3839), .ZN(n3847)
         );
  OAI21_X1 U4571 ( .B1(n2157), .B2(n3845), .A(n3844), .ZN(n3846) );
  OAI21_X1 U4572 ( .B1(n3848), .B2(n3847), .A(n3846), .ZN(n3852) );
  INV_X1 U4573 ( .A(n3849), .ZN(n3850) );
  AOI21_X1 U4574 ( .B1(n3852), .B2(n3851), .A(n3850), .ZN(n3855) );
  OAI21_X1 U4575 ( .B1(n3855), .B2(n3854), .A(n3853), .ZN(n3860) );
  NOR2_X1 U4576 ( .A1(n3857), .A2(n3856), .ZN(n3859) );
  AOI21_X1 U4577 ( .B1(n3860), .B2(n3859), .A(n3858), .ZN(n3864) );
  OAI211_X1 U4578 ( .C1(n3864), .C2(n3863), .A(n3862), .B(n3861), .ZN(n3868)
         );
  NAND4_X1 U4579 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3873)
         );
  INV_X1 U4580 ( .A(n3869), .ZN(n3872) );
  AOI22_X1 U4581 ( .A1(n3873), .A2(n3872), .B1(n3871), .B2(n3870), .ZN(n3875)
         );
  MUX2_X1 U4582 ( .A(n3876), .B(n3875), .S(n3874), .Z(n3877) );
  OAI21_X1 U4583 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n3880) );
  XNOR2_X1 U4584 ( .A(n3880), .B(n4034), .ZN(n3887) );
  NAND2_X1 U4585 ( .A1(n3882), .A2(n3881), .ZN(n3883) );
  OAI211_X1 U4586 ( .C1(n3884), .C2(n3886), .A(n3883), .B(B_REG_SCAN_IN), .ZN(
        n3885) );
  OAI21_X1 U4587 ( .B1(n3887), .B2(n3886), .A(n3885), .ZN(U3239) );
  MUX2_X1 U4588 ( .A(n4041), .B(DATAO_REG_31__SCAN_IN), .S(n3899), .Z(U3581)
         );
  MUX2_X1 U4589 ( .A(n4063), .B(DATAO_REG_30__SCAN_IN), .S(n3899), .Z(U3580)
         );
  MUX2_X1 U4590 ( .A(n4079), .B(DATAO_REG_28__SCAN_IN), .S(n3899), .Z(U3578)
         );
  MUX2_X1 U4591 ( .A(n4114), .B(DATAO_REG_26__SCAN_IN), .S(n3899), .Z(U3576)
         );
  MUX2_X1 U4592 ( .A(n4132), .B(DATAO_REG_25__SCAN_IN), .S(n3899), .Z(U3575)
         );
  MUX2_X1 U4593 ( .A(n4153), .B(DATAO_REG_24__SCAN_IN), .S(n3899), .Z(U3574)
         );
  MUX2_X1 U4594 ( .A(n3888), .B(DATAO_REG_23__SCAN_IN), .S(n3899), .Z(U3573)
         );
  MUX2_X1 U4595 ( .A(n4171), .B(DATAO_REG_21__SCAN_IN), .S(n3899), .Z(U3571)
         );
  MUX2_X1 U4596 ( .A(n4231), .B(DATAO_REG_20__SCAN_IN), .S(n3899), .Z(U3570)
         );
  MUX2_X1 U4597 ( .A(n4244), .B(DATAO_REG_19__SCAN_IN), .S(n3899), .Z(U3569)
         );
  MUX2_X1 U4598 ( .A(DATAO_REG_17__SCAN_IN), .B(n3889), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4599 ( .A(n4291), .B(DATAO_REG_15__SCAN_IN), .S(n3899), .Z(U3565)
         );
  MUX2_X1 U4600 ( .A(DATAO_REG_13__SCAN_IN), .B(n3890), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4601 ( .A(n3891), .B(DATAO_REG_12__SCAN_IN), .S(n3899), .Z(U3562)
         );
  MUX2_X1 U4602 ( .A(n3892), .B(DATAO_REG_11__SCAN_IN), .S(n3899), .Z(U3561)
         );
  MUX2_X1 U4603 ( .A(n3893), .B(DATAO_REG_10__SCAN_IN), .S(n3899), .Z(U3560)
         );
  MUX2_X1 U4604 ( .A(n3894), .B(DATAO_REG_9__SCAN_IN), .S(n3899), .Z(U3559) );
  MUX2_X1 U4605 ( .A(n3895), .B(DATAO_REG_6__SCAN_IN), .S(n3899), .Z(U3556) );
  MUX2_X1 U4606 ( .A(n3896), .B(DATAO_REG_5__SCAN_IN), .S(n3899), .Z(U3555) );
  MUX2_X1 U4607 ( .A(n3897), .B(DATAO_REG_4__SCAN_IN), .S(n3899), .Z(U3554) );
  MUX2_X1 U4608 ( .A(n3898), .B(DATAO_REG_3__SCAN_IN), .S(n3899), .Z(U3553) );
  MUX2_X1 U4609 ( .A(n2325), .B(DATAO_REG_1__SCAN_IN), .S(n3899), .Z(U3551) );
  MUX2_X1 U4610 ( .A(n2671), .B(DATAO_REG_0__SCAN_IN), .S(n3899), .Z(U3550) );
  INV_X1 U4611 ( .A(n4500), .ZN(n4005) );
  NAND2_X1 U4612 ( .A1(n4005), .A2(n3900), .ZN(n3910) );
  OAI211_X1 U4613 ( .C1(n3903), .C2(n3902), .A(n4498), .B(n3901), .ZN(n3909)
         );
  AOI22_X1 U4614 ( .A1(n4494), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3908) );
  XOR2_X1 U4615 ( .A(n3905), .B(n3904), .Z(n3906) );
  NAND2_X1 U4616 ( .A1(n4486), .A2(n3906), .ZN(n3907) );
  NAND4_X1 U4617 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(U3241)
         );
  AOI22_X1 U4618 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4494), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3920) );
  XOR2_X1 U4619 ( .A(n3912), .B(n3911), .Z(n3913) );
  AOI22_X1 U4620 ( .A1(n4005), .A2(n3914), .B1(n4486), .B2(n3913), .ZN(n3919)
         );
  OAI211_X1 U4621 ( .C1(n3917), .C2(n3916), .A(n4498), .B(n3915), .ZN(n3918)
         );
  NAND4_X1 U4622 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(U3242)
         );
  OAI211_X1 U4623 ( .C1(n3924), .C2(n3923), .A(n3922), .B(n4486), .ZN(n3933)
         );
  NOR2_X1 U4624 ( .A1(n4500), .A2(n3925), .ZN(n3926) );
  AOI211_X1 U4625 ( .C1(n4494), .C2(ADDR_REG_9__SCAN_IN), .A(n3927), .B(n3926), 
        .ZN(n3932) );
  OAI211_X1 U4626 ( .C1(n3930), .C2(n3929), .A(n3928), .B(n4498), .ZN(n3931)
         );
  NAND3_X1 U4627 ( .A1(n3933), .A2(n3932), .A3(n3931), .ZN(U3249) );
  INV_X1 U4628 ( .A(n3934), .ZN(n3935) );
  XNOR2_X1 U4629 ( .A(n3955), .B(REG1_REG_11__SCAN_IN), .ZN(n3937) );
  OAI211_X1 U4630 ( .C1(n3938), .C2(n3937), .A(n3957), .B(n4486), .ZN(n3950)
         );
  INV_X1 U4631 ( .A(n3939), .ZN(n3940) );
  AOI21_X1 U4632 ( .B1(n4494), .B2(ADDR_REG_11__SCAN_IN), .A(n3940), .ZN(n3949) );
  MUX2_X1 U4633 ( .A(n3951), .B(REG2_REG_11__SCAN_IN), .S(n3955), .Z(n3945) );
  OAI211_X1 U4634 ( .C1(n3946), .C2(n3945), .A(n3953), .B(n4498), .ZN(n3948)
         );
  OR2_X1 U4635 ( .A1(n4500), .A2(n3955), .ZN(n3947) );
  NAND4_X1 U4636 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(U3251)
         );
  OR2_X1 U4637 ( .A1(n3955), .A2(n3951), .ZN(n3952) );
  INV_X1 U4638 ( .A(n4460), .ZN(n3972) );
  XOR2_X1 U4639 ( .A(REG2_REG_12__SCAN_IN), .B(n3965), .Z(n3963) );
  OAI211_X1 U4640 ( .C1(n3958), .C2(REG1_REG_12__SCAN_IN), .A(n3971), .B(n4486), .ZN(n3961) );
  AOI21_X1 U4641 ( .B1(n4494), .B2(ADDR_REG_12__SCAN_IN), .A(n3959), .ZN(n3960) );
  OAI211_X1 U4642 ( .C1(n4500), .C2(n3972), .A(n3961), .B(n3960), .ZN(n3962)
         );
  AOI21_X1 U4643 ( .B1(n4498), .B2(n3963), .A(n3962), .ZN(n3964) );
  INV_X1 U4644 ( .A(n3964), .ZN(U3252) );
  NAND2_X1 U4645 ( .A1(n3965), .A2(REG2_REG_12__SCAN_IN), .ZN(n3968) );
  NAND2_X1 U4646 ( .A1(n3966), .A2(n4460), .ZN(n3967) );
  NOR2_X1 U4647 ( .A1(n3987), .A2(n3986), .ZN(n3984) );
  AOI21_X1 U4648 ( .B1(n3986), .B2(n3987), .A(n3984), .ZN(n3969) );
  XNOR2_X1 U4649 ( .A(n3985), .B(n3969), .ZN(n3980) );
  XNOR2_X1 U4650 ( .A(n3987), .B(REG1_REG_13__SCAN_IN), .ZN(n3973) );
  OAI211_X1 U4651 ( .C1(n3974), .C2(n3973), .A(n3982), .B(n4486), .ZN(n3979)
         );
  NAND2_X1 U4652 ( .A1(n4494), .A2(ADDR_REG_13__SCAN_IN), .ZN(n3975) );
  OAI211_X1 U4653 ( .C1(n4500), .C2(n3987), .A(n3976), .B(n3975), .ZN(n3977)
         );
  INV_X1 U4654 ( .A(n3977), .ZN(n3978) );
  OAI211_X1 U4655 ( .C1(n3980), .C2(n4038), .A(n3979), .B(n3978), .ZN(U3253)
         );
  INV_X1 U4656 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4390) );
  OAI211_X1 U4657 ( .C1(n3983), .C2(REG1_REG_14__SCAN_IN), .A(n4008), .B(n4486), .ZN(n3995) );
  NAND2_X1 U4658 ( .A1(n3987), .A2(n3986), .ZN(n3988) );
  AOI211_X1 U4659 ( .C1(n2485), .C2(n3989), .A(n4038), .B(n3997), .ZN(n3993)
         );
  NAND2_X1 U4660 ( .A1(n4494), .A2(ADDR_REG_14__SCAN_IN), .ZN(n3990) );
  OAI211_X1 U4661 ( .C1(n4500), .C2(n4009), .A(n3991), .B(n3990), .ZN(n3992)
         );
  NOR2_X1 U4662 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  NAND2_X1 U4663 ( .A1(n3995), .A2(n3994), .ZN(U3254) );
  XNOR2_X1 U4664 ( .A(n4006), .B(REG2_REG_17__SCAN_IN), .ZN(n4003) );
  INV_X1 U4665 ( .A(n3996), .ZN(n3999) );
  INV_X1 U4666 ( .A(n4013), .ZN(n4523) );
  AOI22_X1 U4667 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4523), .B1(n4013), .B2(
        n4301), .ZN(n4475) );
  NAND2_X1 U4668 ( .A1(n4000), .A2(n4521), .ZN(n4001) );
  OAI21_X1 U4669 ( .B1(n4003), .B2(n4002), .A(n4024), .ZN(n4004) );
  AOI22_X1 U4670 ( .A1(n4005), .A2(n4028), .B1(n4498), .B2(n4004), .ZN(n4022)
         );
  XNOR2_X1 U4671 ( .A(n4006), .B(REG1_REG_17__SCAN_IN), .ZN(n4017) );
  INV_X1 U4672 ( .A(n4007), .ZN(n4010) );
  OAI21_X1 U4673 ( .B1(n4010), .B2(n4009), .A(n4008), .ZN(n4011) );
  INV_X1 U4674 ( .A(n4011), .ZN(n4470) );
  AOI22_X1 U4675 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4523), .B1(n4013), .B2(
        n4012), .ZN(n4469) );
  NAND2_X1 U4676 ( .A1(n2038), .A2(n4521), .ZN(n4015) );
  OAI21_X1 U4677 ( .B1(n4017), .B2(n4016), .A(n4027), .ZN(n4018) );
  NAND2_X1 U4678 ( .A1(n4486), .A2(n4018), .ZN(n4020) );
  NAND2_X1 U4679 ( .A1(n4494), .A2(ADDR_REG_17__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U4680 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(U3257)
         );
  MUX2_X1 U4681 ( .A(n4238), .B(REG2_REG_19__SCAN_IN), .S(n4034), .Z(n4025) );
  NAND2_X1 U4682 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4029), .ZN(n4023) );
  OAI21_X1 U4683 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4029), .A(n4023), .ZN(n4497) );
  INV_X1 U4684 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4685 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4519), .B1(n4029), .B2(
        n4026), .ZN(n4492) );
  XNOR2_X1 U4686 ( .A(n4034), .B(REG1_REG_19__SCAN_IN), .ZN(n4030) );
  XNOR2_X1 U4687 ( .A(n4031), .B(n4030), .ZN(n4036) );
  NAND2_X1 U4688 ( .A1(n4494), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4032) );
  OAI211_X1 U4689 ( .C1(n4500), .C2(n4034), .A(n4033), .B(n4032), .ZN(n4035)
         );
  AOI21_X1 U4690 ( .B1(n4036), .B2(n4486), .A(n4035), .ZN(n4037) );
  OAI21_X1 U4691 ( .B1(n4039), .B2(n4038), .A(n4037), .ZN(U3259) );
  NAND2_X1 U4692 ( .A1(n4057), .A2(n4048), .ZN(n4046) );
  XOR2_X1 U4693 ( .A(n4042), .B(n4046), .Z(n4399) );
  AND2_X1 U4694 ( .A1(n4457), .A2(B_REG_SCAN_IN), .ZN(n4040) );
  NOR2_X1 U4695 ( .A1(n4311), .A2(n4040), .ZN(n4064) );
  NAND2_X1 U4696 ( .A1(n4064), .A2(n4041), .ZN(n4050) );
  OR2_X1 U4697 ( .A1(n4262), .A2(n4042), .ZN(n4043) );
  NAND2_X1 U4698 ( .A1(n4050), .A2(n4043), .ZN(n4396) );
  NAND2_X1 U4699 ( .A1(n4313), .A2(n4396), .ZN(n4045) );
  NAND2_X1 U4700 ( .A1(n4515), .A2(REG2_REG_31__SCAN_IN), .ZN(n4044) );
  OAI211_X1 U4701 ( .C1(n4399), .C2(n4272), .A(n4045), .B(n4044), .ZN(U3260)
         );
  OAI21_X1 U4702 ( .B1(n4057), .B2(n4048), .A(n4046), .ZN(n4404) );
  INV_X1 U4703 ( .A(n4404), .ZN(n4047) );
  NAND2_X1 U4704 ( .A1(n4047), .A2(n4503), .ZN(n4052) );
  OR2_X1 U4705 ( .A1(n4262), .A2(n4048), .ZN(n4049) );
  NAND2_X1 U4706 ( .A1(n4050), .A2(n4049), .ZN(n4402) );
  NAND2_X1 U4707 ( .A1(n4313), .A2(n4402), .ZN(n4051) );
  OAI211_X1 U4708 ( .C1(n4313), .C2(n4646), .A(n4052), .B(n4051), .ZN(U3261)
         );
  NAND2_X1 U4709 ( .A1(n4079), .A2(n4055), .ZN(n4325) );
  NAND2_X1 U4710 ( .A1(n4327), .A2(n4325), .ZN(n4056) );
  XOR2_X1 U4711 ( .A(n4323), .B(n4056), .Z(n4072) );
  AOI22_X1 U4712 ( .A1(n4322), .A2(n4503), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4515), .ZN(n4071) );
  OAI21_X1 U4713 ( .B1(n4075), .B2(n4060), .A(n4059), .ZN(n4061) );
  AOI22_X1 U4714 ( .A1(n4064), .A2(n4063), .B1(n4306), .B2(n4062), .ZN(n4065)
         );
  OAI21_X1 U4715 ( .B1(n4066), .B2(n4263), .A(n4065), .ZN(n4067) );
  OAI21_X1 U4716 ( .B1(n4068), .B2(n4299), .A(n4330), .ZN(n4069) );
  NAND2_X1 U4717 ( .A1(n4069), .A2(n4313), .ZN(n4070) );
  OAI211_X1 U4718 ( .C1(n4072), .C2(n4316), .A(n4071), .B(n4070), .ZN(U3354)
         );
  XNOR2_X1 U4719 ( .A(n4073), .B(n4076), .ZN(n4332) );
  INV_X1 U4720 ( .A(n4332), .ZN(n4086) );
  OAI22_X1 U4721 ( .A1(n4074), .A2(n4263), .B1(n4080), .B2(n4262), .ZN(n4078)
         );
  INV_X1 U4722 ( .A(n4333), .ZN(n4084) );
  OAI21_X1 U4723 ( .B1(n4097), .B2(n4080), .A(n2749), .ZN(n4334) );
  AOI22_X1 U4724 ( .A1(n4081), .A2(n4510), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4515), .ZN(n4082) );
  OAI21_X1 U4725 ( .B1(n4334), .B2(n4272), .A(n4082), .ZN(n4083) );
  AOI21_X1 U4726 ( .B1(n4084), .B2(n4313), .A(n4083), .ZN(n4085) );
  OAI21_X1 U4727 ( .B1(n4086), .B2(n4316), .A(n4085), .ZN(U3263) );
  INV_X1 U4728 ( .A(n4336), .ZN(n4106) );
  INV_X1 U4729 ( .A(n4109), .ZN(n4089) );
  OAI21_X1 U4730 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4091) );
  XNOR2_X1 U4731 ( .A(n4091), .B(n4090), .ZN(n4096) );
  OAI22_X1 U4732 ( .A1(n4092), .A2(n4263), .B1(n4099), .B2(n4262), .ZN(n4093)
         );
  AOI21_X1 U4733 ( .B1(n4266), .B2(n4094), .A(n4093), .ZN(n4095) );
  OAI21_X1 U4734 ( .B1(n4096), .B2(n4268), .A(n4095), .ZN(n4335) );
  INV_X1 U4735 ( .A(n4118), .ZN(n4100) );
  INV_X1 U4736 ( .A(n4097), .ZN(n4098) );
  NOR2_X1 U4737 ( .A1(n4409), .A2(n4272), .ZN(n4104) );
  INV_X1 U4738 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4101) );
  OAI22_X1 U4739 ( .A1(n4102), .A2(n4299), .B1(n4101), .B2(n4313), .ZN(n4103)
         );
  AOI211_X1 U4740 ( .C1(n4335), .C2(n4313), .A(n4104), .B(n4103), .ZN(n4105)
         );
  OAI21_X1 U4741 ( .B1(n4106), .B2(n4316), .A(n4105), .ZN(U3264) );
  XNOR2_X1 U4742 ( .A(n4107), .B(n4110), .ZN(n4340) );
  INV_X1 U4743 ( .A(n4340), .ZN(n4125) );
  NAND2_X1 U4744 ( .A1(n4109), .A2(n4108), .ZN(n4111) );
  XNOR2_X1 U4745 ( .A(n4111), .B(n4110), .ZN(n4112) );
  NAND2_X1 U4746 ( .A1(n4112), .A2(n4304), .ZN(n4116) );
  AOI22_X1 U4747 ( .A1(n4114), .A2(n4266), .B1(n4306), .B2(n4113), .ZN(n4115)
         );
  OAI211_X1 U4748 ( .C1(n4117), .C2(n4263), .A(n4116), .B(n4115), .ZN(n4339)
         );
  INV_X1 U4749 ( .A(n4136), .ZN(n4120) );
  OAI21_X1 U4750 ( .B1(n4120), .B2(n4119), .A(n4118), .ZN(n4413) );
  AOI22_X1 U4751 ( .A1(n4121), .A2(n4510), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4515), .ZN(n4122) );
  OAI21_X1 U4752 ( .B1(n4413), .B2(n4272), .A(n4122), .ZN(n4123) );
  AOI21_X1 U4753 ( .B1(n4339), .B2(n4313), .A(n4123), .ZN(n4124) );
  OAI21_X1 U4754 ( .B1(n4125), .B2(n4316), .A(n4124), .ZN(U3265) );
  XOR2_X1 U4755 ( .A(n4130), .B(n4126), .Z(n4344) );
  INV_X1 U4756 ( .A(n4344), .ZN(n4143) );
  NAND2_X1 U4757 ( .A1(n4128), .A2(n4127), .ZN(n4129) );
  XOR2_X1 U4758 ( .A(n4130), .B(n4129), .Z(n4134) );
  OAI22_X1 U4759 ( .A1(n4173), .A2(n4263), .B1(n4137), .B2(n4262), .ZN(n4131)
         );
  AOI21_X1 U4760 ( .B1(n4266), .B2(n4132), .A(n4131), .ZN(n4133) );
  OAI21_X1 U4761 ( .B1(n4134), .B2(n4268), .A(n4133), .ZN(n4343) );
  INV_X1 U4762 ( .A(n4135), .ZN(n4138) );
  OAI21_X1 U4763 ( .B1(n4138), .B2(n4137), .A(n4136), .ZN(n4417) );
  AOI22_X1 U4764 ( .A1(n4139), .A2(n4510), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4515), .ZN(n4140) );
  OAI21_X1 U4765 ( .B1(n4417), .B2(n4272), .A(n4140), .ZN(n4141) );
  AOI21_X1 U4766 ( .B1(n4343), .B2(n4313), .A(n4141), .ZN(n4142) );
  OAI21_X1 U4767 ( .B1(n4143), .B2(n4316), .A(n4142), .ZN(U3266) );
  XOR2_X1 U4768 ( .A(n4149), .B(n4144), .Z(n4348) );
  INV_X1 U4769 ( .A(n4348), .ZN(n4162) );
  NAND2_X1 U4770 ( .A1(n4186), .A2(n4145), .ZN(n4147) );
  NAND2_X1 U4771 ( .A1(n4147), .A2(n4146), .ZN(n4167) );
  INV_X1 U4772 ( .A(n4164), .ZN(n4166) );
  NAND2_X1 U4773 ( .A1(n4167), .A2(n4166), .ZN(n4169) );
  NAND2_X1 U4774 ( .A1(n4169), .A2(n4148), .ZN(n4150) );
  XNOR2_X1 U4775 ( .A(n4150), .B(n4149), .ZN(n4155) );
  OAI22_X1 U4776 ( .A1(n4151), .A2(n4263), .B1(n4262), .B2(n4156), .ZN(n4152)
         );
  AOI21_X1 U4777 ( .B1(n4266), .B2(n4153), .A(n4152), .ZN(n4154) );
  OAI21_X1 U4778 ( .B1(n4155), .B2(n4268), .A(n4154), .ZN(n4347) );
  OAI21_X1 U4779 ( .B1(n4352), .B2(n4156), .A(n4135), .ZN(n4421) );
  NOR2_X1 U4780 ( .A1(n4421), .A2(n4272), .ZN(n4160) );
  OAI22_X1 U4781 ( .A1(n4158), .A2(n4299), .B1(n4157), .B2(n4313), .ZN(n4159)
         );
  AOI211_X1 U4782 ( .C1(n4347), .C2(n4313), .A(n4160), .B(n4159), .ZN(n4161)
         );
  OAI21_X1 U4783 ( .B1(n4162), .B2(n4316), .A(n4161), .ZN(U3267) );
  OAI21_X1 U4784 ( .B1(n4165), .B2(n4164), .A(n4163), .ZN(n4355) );
  OR2_X1 U4785 ( .A1(n4167), .A2(n4166), .ZN(n4168) );
  NAND2_X1 U4786 ( .A1(n4169), .A2(n4168), .ZN(n4175) );
  NOR2_X1 U4787 ( .A1(n4262), .A2(n4179), .ZN(n4170) );
  AOI21_X1 U4788 ( .B1(n4171), .B2(n4308), .A(n4170), .ZN(n4172) );
  OAI21_X1 U4789 ( .B1(n4173), .B2(n4311), .A(n4172), .ZN(n4174) );
  AOI21_X1 U4790 ( .B1(n4175), .B2(n4304), .A(n4174), .ZN(n4354) );
  OAI22_X1 U4791 ( .A1(n4177), .A2(n4299), .B1(n4313), .B2(n4176), .ZN(n4178)
         );
  INV_X1 U4792 ( .A(n4178), .ZN(n4181) );
  NOR2_X1 U4793 ( .A1(n4192), .A2(n4179), .ZN(n4351) );
  OR3_X1 U4794 ( .A1(n4352), .A2(n4351), .A3(n4272), .ZN(n4180) );
  OAI211_X1 U4795 ( .C1(n4354), .C2(n4515), .A(n4181), .B(n4180), .ZN(n4182)
         );
  INV_X1 U4796 ( .A(n4182), .ZN(n4183) );
  OAI21_X1 U4797 ( .B1(n4355), .B2(n4316), .A(n4183), .ZN(U3268) );
  XNOR2_X1 U4798 ( .A(n4184), .B(n4185), .ZN(n4357) );
  INV_X1 U4799 ( .A(n4357), .ZN(n4199) );
  XNOR2_X1 U4800 ( .A(n4186), .B(n4185), .ZN(n4191) );
  OAI22_X1 U4801 ( .A1(n4187), .A2(n4263), .B1(n4194), .B2(n4262), .ZN(n4188)
         );
  AOI21_X1 U4802 ( .B1(n4189), .B2(n4266), .A(n4188), .ZN(n4190) );
  OAI21_X1 U4803 ( .B1(n4191), .B2(n4268), .A(n4190), .ZN(n4356) );
  INV_X1 U4804 ( .A(n4192), .ZN(n4193) );
  OAI21_X1 U4805 ( .B1(n2747), .B2(n4194), .A(n4193), .ZN(n4426) );
  AOI22_X1 U4806 ( .A1(n4515), .A2(REG2_REG_21__SCAN_IN), .B1(n4195), .B2(
        n4510), .ZN(n4196) );
  OAI21_X1 U4807 ( .B1(n4426), .B2(n4272), .A(n4196), .ZN(n4197) );
  AOI21_X1 U4808 ( .B1(n4356), .B2(n4313), .A(n4197), .ZN(n4198) );
  OAI21_X1 U4809 ( .B1(n4199), .B2(n4316), .A(n4198), .ZN(U3269) );
  XNOR2_X1 U4810 ( .A(n4201), .B(n4200), .ZN(n4213) );
  INV_X1 U4811 ( .A(n4202), .ZN(n4203) );
  NAND2_X1 U4812 ( .A1(n4204), .A2(n4203), .ZN(n4206) );
  XNOR2_X1 U4813 ( .A(n4206), .B(n4205), .ZN(n4210) );
  AOI22_X1 U4814 ( .A1(n4244), .A2(n4308), .B1(n4214), .B2(n4306), .ZN(n4207)
         );
  OAI21_X1 U4815 ( .B1(n4208), .B2(n4311), .A(n4207), .ZN(n4209) );
  AOI21_X1 U4816 ( .B1(n4210), .B2(n4304), .A(n4209), .ZN(n4211) );
  OAI21_X1 U4817 ( .B1(n4213), .B2(n4212), .A(n4211), .ZN(n4359) );
  INV_X1 U4818 ( .A(n4359), .ZN(n4221) );
  INV_X1 U4819 ( .A(n4213), .ZN(n4360) );
  NAND2_X1 U4820 ( .A1(n4234), .A2(n4214), .ZN(n4215) );
  NAND2_X1 U4821 ( .A1(n4216), .A2(n4215), .ZN(n4430) );
  AOI22_X1 U4822 ( .A1(n4515), .A2(REG2_REG_20__SCAN_IN), .B1(n4217), .B2(
        n4510), .ZN(n4218) );
  OAI21_X1 U4823 ( .B1(n4430), .B2(n4272), .A(n4218), .ZN(n4219) );
  AOI21_X1 U4824 ( .B1(n4360), .B2(n4512), .A(n4219), .ZN(n4220) );
  OAI21_X1 U4825 ( .B1(n4221), .B2(n4515), .A(n4220), .ZN(U3270) );
  XNOR2_X1 U4826 ( .A(n4222), .B(n4229), .ZN(n4364) );
  INV_X1 U4827 ( .A(n4364), .ZN(n4242) );
  OAI21_X1 U4828 ( .B1(n4261), .B2(n4224), .A(n4223), .ZN(n4243) );
  INV_X1 U4829 ( .A(n4225), .ZN(n4227) );
  OAI21_X1 U4830 ( .B1(n4243), .B2(n4227), .A(n4226), .ZN(n4228) );
  XOR2_X1 U4831 ( .A(n4229), .B(n4228), .Z(n4233) );
  OAI22_X1 U4832 ( .A1(n2548), .A2(n4263), .B1(n4262), .B2(n4235), .ZN(n4230)
         );
  AOI21_X1 U4833 ( .B1(n4231), .B2(n4266), .A(n4230), .ZN(n4232) );
  OAI21_X1 U4834 ( .B1(n4233), .B2(n4268), .A(n4232), .ZN(n4363) );
  OAI21_X1 U4835 ( .B1(n4236), .B2(n4235), .A(n4234), .ZN(n4434) );
  NOR2_X1 U4836 ( .A1(n4434), .A2(n4272), .ZN(n4240) );
  OAI22_X1 U4837 ( .A1(n4313), .A2(n4238), .B1(n4237), .B2(n4299), .ZN(n4239)
         );
  AOI211_X1 U4838 ( .C1(n4363), .C2(n4313), .A(n4240), .B(n4239), .ZN(n4241)
         );
  OAI21_X1 U4839 ( .B1(n4242), .B2(n4316), .A(n4241), .ZN(U3271) );
  XOR2_X1 U4840 ( .A(n4249), .B(n4243), .Z(n4247) );
  AOI22_X1 U4841 ( .A1(n4244), .A2(n4266), .B1(n2274), .B2(n4306), .ZN(n4245)
         );
  OAI21_X1 U4842 ( .B1(n4294), .B2(n4263), .A(n4245), .ZN(n4246) );
  AOI21_X1 U4843 ( .B1(n4247), .B2(n4304), .A(n4246), .ZN(n4369) );
  OAI21_X1 U4844 ( .B1(n4250), .B2(n4249), .A(n4248), .ZN(n4367) );
  XNOR2_X1 U4845 ( .A(n4270), .B(n2274), .ZN(n4251) );
  NAND2_X1 U4846 ( .A1(n4251), .A2(n4544), .ZN(n4368) );
  INV_X1 U4847 ( .A(n4252), .ZN(n4255) );
  AOI22_X1 U4848 ( .A1(n4515), .A2(REG2_REG_18__SCAN_IN), .B1(n4253), .B2(
        n4510), .ZN(n4254) );
  OAI21_X1 U4849 ( .B1(n4368), .B2(n4255), .A(n4254), .ZN(n4256) );
  AOI21_X1 U4850 ( .B1(n4367), .B2(n4257), .A(n4256), .ZN(n4258) );
  OAI21_X1 U4851 ( .B1(n4515), .B2(n4369), .A(n4258), .ZN(U3272) );
  XNOR2_X1 U4852 ( .A(n2064), .B(n4260), .ZN(n4372) );
  INV_X1 U4853 ( .A(n4372), .ZN(n4279) );
  XNOR2_X1 U4854 ( .A(n4261), .B(n4260), .ZN(n4269) );
  OAI22_X1 U4855 ( .A1(n4312), .A2(n4263), .B1(n4262), .B2(n4271), .ZN(n4264)
         );
  AOI21_X1 U4856 ( .B1(n4266), .B2(n4265), .A(n4264), .ZN(n4267) );
  OAI21_X1 U4857 ( .B1(n4269), .B2(n4268), .A(n4267), .ZN(n4371) );
  OAI21_X1 U4858 ( .B1(n2023), .B2(n4271), .A(n2275), .ZN(n4439) );
  NOR2_X1 U4859 ( .A1(n4439), .A2(n4272), .ZN(n4277) );
  INV_X1 U4860 ( .A(n4273), .ZN(n4274) );
  OAI22_X1 U4861 ( .A1(n4313), .A2(n4275), .B1(n4274), .B2(n4299), .ZN(n4276)
         );
  AOI211_X1 U4862 ( .C1(n4371), .C2(n4313), .A(n4277), .B(n4276), .ZN(n4278)
         );
  OAI21_X1 U4863 ( .B1(n4279), .B2(n4316), .A(n4278), .ZN(U3273) );
  OAI21_X1 U4864 ( .B1(n4282), .B2(n4281), .A(n4280), .ZN(n4378) );
  AOI21_X1 U4865 ( .B1(n4290), .B2(n4283), .A(n2023), .ZN(n4376) );
  OAI22_X1 U4866 ( .A1(n4313), .A2(n4285), .B1(n4284), .B2(n4299), .ZN(n4286)
         );
  AOI21_X1 U4867 ( .B1(n4376), .B2(n4503), .A(n4286), .ZN(n4296) );
  OAI211_X1 U4868 ( .C1(n4289), .C2(n4288), .A(n4287), .B(n4304), .ZN(n4293)
         );
  AOI22_X1 U4869 ( .A1(n4291), .A2(n4308), .B1(n4306), .B2(n4290), .ZN(n4292)
         );
  OAI211_X1 U4870 ( .C1(n4294), .C2(n4311), .A(n4293), .B(n4292), .ZN(n4375)
         );
  NAND2_X1 U4871 ( .A1(n4375), .A2(n4313), .ZN(n4295) );
  OAI211_X1 U4872 ( .C1(n4378), .C2(n4316), .A(n4296), .B(n4295), .ZN(U3274)
         );
  XNOR2_X1 U4873 ( .A(n4297), .B(n2049), .ZN(n4382) );
  XNOR2_X1 U4874 ( .A(n4298), .B(n4305), .ZN(n4380) );
  OAI22_X1 U4875 ( .A1(n4313), .A2(n4301), .B1(n4300), .B2(n4299), .ZN(n4302)
         );
  AOI21_X1 U4876 ( .B1(n4380), .B2(n4503), .A(n4302), .ZN(n4315) );
  OAI211_X1 U4877 ( .C1(n2039), .C2(n2049), .A(n4304), .B(n4303), .ZN(n4310)
         );
  AOI22_X1 U4878 ( .A1(n4308), .A2(n4307), .B1(n4306), .B2(n4305), .ZN(n4309)
         );
  OAI211_X1 U4879 ( .C1(n4312), .C2(n4311), .A(n4310), .B(n4309), .ZN(n4379)
         );
  NAND2_X1 U4880 ( .A1(n4379), .A2(n4313), .ZN(n4314) );
  OAI211_X1 U4881 ( .C1(n4382), .C2(n4316), .A(n4315), .B(n4314), .ZN(U3275)
         );
  NAND2_X1 U4882 ( .A1(n4561), .A2(n4396), .ZN(n4318) );
  NAND2_X1 U4883 ( .A1(n4559), .A2(REG1_REG_31__SCAN_IN), .ZN(n4317) );
  OAI211_X1 U4884 ( .C1(n4399), .C2(n4395), .A(n4318), .B(n4317), .ZN(U3549)
         );
  NAND2_X1 U4885 ( .A1(n4561), .A2(n4402), .ZN(n4320) );
  NAND2_X1 U4886 ( .A1(n4559), .A2(REG1_REG_30__SCAN_IN), .ZN(n4319) );
  OAI211_X1 U4887 ( .C1(n4404), .C2(n4395), .A(n4320), .B(n4319), .ZN(U3548)
         );
  NOR2_X1 U4888 ( .A1(n4325), .A2(n4539), .ZN(n4321) );
  AOI22_X1 U4889 ( .A1(n4322), .A2(n4544), .B1(n4323), .B2(n4321), .ZN(n4331)
         );
  INV_X1 U4890 ( .A(n4327), .ZN(n4324) );
  NAND3_X1 U4891 ( .A1(n4324), .A2(n4323), .A3(n4547), .ZN(n4329) );
  NAND4_X1 U4892 ( .A1(n4327), .A2(n4547), .A3(n4326), .A4(n4325), .ZN(n4328)
         );
  MUX2_X1 U4893 ( .A(REG1_REG_29__SCAN_IN), .B(n4405), .S(n4561), .Z(U3547) );
  MUX2_X1 U4894 ( .A(REG1_REG_27__SCAN_IN), .B(n4406), .S(n4561), .Z(U3545) );
  INV_X1 U4895 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4337) );
  AOI21_X1 U4896 ( .B1(n4336), .B2(n4547), .A(n4335), .ZN(n4407) );
  MUX2_X1 U4897 ( .A(n4337), .B(n4407), .S(n4561), .Z(n4338) );
  INV_X1 U4898 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4341) );
  AOI21_X1 U4899 ( .B1(n4340), .B2(n4547), .A(n4339), .ZN(n4410) );
  MUX2_X1 U4900 ( .A(n4341), .B(n4410), .S(n4561), .Z(n4342) );
  OAI21_X1 U4901 ( .B1(n4395), .B2(n4413), .A(n4342), .ZN(U3543) );
  INV_X1 U4902 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4345) );
  AOI21_X1 U4903 ( .B1(n4344), .B2(n4547), .A(n4343), .ZN(n4414) );
  MUX2_X1 U4904 ( .A(n4345), .B(n4414), .S(n4561), .Z(n4346) );
  OAI21_X1 U4905 ( .B1(n4395), .B2(n4417), .A(n4346), .ZN(U3542) );
  INV_X1 U4906 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4349) );
  AOI21_X1 U4907 ( .B1(n4348), .B2(n4547), .A(n4347), .ZN(n4418) );
  MUX2_X1 U4908 ( .A(n4349), .B(n4418), .S(n4561), .Z(n4350) );
  OAI21_X1 U4909 ( .B1(n4395), .B2(n4421), .A(n4350), .ZN(U3541) );
  OR3_X1 U4910 ( .A1(n4352), .A2(n4351), .A3(n4528), .ZN(n4353) );
  OAI211_X1 U4911 ( .C1(n4355), .C2(n4539), .A(n4354), .B(n4353), .ZN(n4422)
         );
  MUX2_X1 U4912 ( .A(REG1_REG_22__SCAN_IN), .B(n4422), .S(n4561), .Z(U3540) );
  AOI21_X1 U4913 ( .B1(n4357), .B2(n4547), .A(n4356), .ZN(n4423) );
  MUX2_X1 U4914 ( .A(n4680), .B(n4423), .S(n4561), .Z(n4358) );
  OAI21_X1 U4915 ( .B1(n4395), .B2(n4426), .A(n4358), .ZN(U3539) );
  INV_X1 U4916 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4361) );
  AOI21_X1 U4917 ( .B1(n4537), .B2(n4360), .A(n4359), .ZN(n4427) );
  MUX2_X1 U4918 ( .A(n4361), .B(n4427), .S(n4561), .Z(n4362) );
  OAI21_X1 U4919 ( .B1(n4395), .B2(n4430), .A(n4362), .ZN(U3538) );
  INV_X1 U4920 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4365) );
  AOI21_X1 U4921 ( .B1(n4364), .B2(n4547), .A(n4363), .ZN(n4431) );
  MUX2_X1 U4922 ( .A(n4365), .B(n4431), .S(n4561), .Z(n4366) );
  OAI21_X1 U4923 ( .B1(n4395), .B2(n4434), .A(n4366), .ZN(U3537) );
  INV_X1 U4924 ( .A(n4367), .ZN(n4370) );
  OAI211_X1 U4925 ( .C1(n4370), .C2(n4539), .A(n4369), .B(n4368), .ZN(n4435)
         );
  MUX2_X1 U4926 ( .A(REG1_REG_18__SCAN_IN), .B(n4435), .S(n4561), .Z(U3536) );
  AOI21_X1 U4927 ( .B1(n4372), .B2(n4547), .A(n4371), .ZN(n4436) );
  MUX2_X1 U4928 ( .A(n4373), .B(n4436), .S(n4561), .Z(n4374) );
  OAI21_X1 U4929 ( .B1(n4395), .B2(n4439), .A(n4374), .ZN(U3535) );
  AOI21_X1 U4930 ( .B1(n4544), .B2(n4376), .A(n4375), .ZN(n4377) );
  OAI21_X1 U4931 ( .B1(n4378), .B2(n4539), .A(n4377), .ZN(n4440) );
  MUX2_X1 U4932 ( .A(REG1_REG_16__SCAN_IN), .B(n4440), .S(n4561), .Z(U3534) );
  AOI21_X1 U4933 ( .B1(n4544), .B2(n4380), .A(n4379), .ZN(n4381) );
  OAI21_X1 U4934 ( .B1(n4382), .B2(n4539), .A(n4381), .ZN(n4441) );
  MUX2_X1 U4935 ( .A(REG1_REG_15__SCAN_IN), .B(n4441), .S(n4561), .Z(U3533) );
  AOI21_X1 U4936 ( .B1(n4384), .B2(n4547), .A(n4383), .ZN(n4442) );
  MUX2_X1 U4937 ( .A(n4385), .B(n4442), .S(n4561), .Z(n4386) );
  OAI21_X1 U4938 ( .B1(n4395), .B2(n4445), .A(n4386), .ZN(U3532) );
  INV_X1 U4939 ( .A(n4387), .ZN(n4388) );
  AOI21_X1 U4940 ( .B1(n4537), .B2(n4389), .A(n4388), .ZN(n4446) );
  MUX2_X1 U4941 ( .A(n4390), .B(n4446), .S(n4561), .Z(n4391) );
  OAI21_X1 U4942 ( .B1(n4395), .B2(n4449), .A(n4391), .ZN(U3531) );
  AOI21_X1 U4943 ( .B1(n4547), .B2(n4393), .A(n4392), .ZN(n4450) );
  MUX2_X1 U4944 ( .A(n2121), .B(n4450), .S(n4561), .Z(n4394) );
  OAI21_X1 U4945 ( .B1(n4395), .B2(n4454), .A(n4394), .ZN(U3530) );
  NAND2_X1 U4946 ( .A1(n4553), .A2(n4396), .ZN(n4398) );
  NAND2_X1 U4947 ( .A1(n4552), .A2(REG0_REG_31__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U4948 ( .C1(n4399), .C2(n4453), .A(n4398), .B(n4397), .ZN(U3517)
         );
  NOR2_X1 U4949 ( .A1(n4553), .A2(n4400), .ZN(n4401) );
  AOI21_X1 U4950 ( .B1(n4553), .B2(n4402), .A(n4401), .ZN(n4403) );
  OAI21_X1 U4951 ( .B1(n4404), .B2(n4453), .A(n4403), .ZN(U3516) );
  MUX2_X1 U4952 ( .A(REG0_REG_29__SCAN_IN), .B(n4405), .S(n4553), .Z(U3515) );
  MUX2_X1 U4953 ( .A(REG0_REG_27__SCAN_IN), .B(n4406), .S(n4553), .Z(U3513) );
  MUX2_X1 U4954 ( .A(n4679), .B(n4407), .S(n4553), .Z(n4408) );
  INV_X1 U4955 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U4956 ( .A(n4411), .B(n4410), .S(n4553), .Z(n4412) );
  OAI21_X1 U4957 ( .B1(n4413), .B2(n4453), .A(n4412), .ZN(U3511) );
  INV_X1 U4958 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4415) );
  MUX2_X1 U4959 ( .A(n4415), .B(n4414), .S(n4553), .Z(n4416) );
  OAI21_X1 U4960 ( .B1(n4417), .B2(n4453), .A(n4416), .ZN(U3510) );
  INV_X1 U4961 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4419) );
  MUX2_X1 U4962 ( .A(n4419), .B(n4418), .S(n4553), .Z(n4420) );
  OAI21_X1 U4963 ( .B1(n4421), .B2(n4453), .A(n4420), .ZN(U3509) );
  MUX2_X1 U4964 ( .A(REG0_REG_22__SCAN_IN), .B(n4422), .S(n4553), .Z(U3508) );
  INV_X1 U4965 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4424) );
  MUX2_X1 U4966 ( .A(n4424), .B(n4423), .S(n4553), .Z(n4425) );
  OAI21_X1 U4967 ( .B1(n4426), .B2(n4453), .A(n4425), .ZN(U3507) );
  INV_X1 U4968 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4428) );
  MUX2_X1 U4969 ( .A(n4428), .B(n4427), .S(n4553), .Z(n4429) );
  OAI21_X1 U4970 ( .B1(n4430), .B2(n4453), .A(n4429), .ZN(U3506) );
  INV_X1 U4971 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4432) );
  MUX2_X1 U4972 ( .A(n4432), .B(n4431), .S(n4553), .Z(n4433) );
  OAI21_X1 U4973 ( .B1(n4434), .B2(n4453), .A(n4433), .ZN(U3505) );
  MUX2_X1 U4974 ( .A(REG0_REG_18__SCAN_IN), .B(n4435), .S(n4553), .Z(U3503) );
  INV_X1 U4975 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4437) );
  MUX2_X1 U4976 ( .A(n4437), .B(n4436), .S(n4553), .Z(n4438) );
  OAI21_X1 U4977 ( .B1(n4439), .B2(n4453), .A(n4438), .ZN(U3501) );
  MUX2_X1 U4978 ( .A(REG0_REG_16__SCAN_IN), .B(n4440), .S(n4553), .Z(U3499) );
  MUX2_X1 U4979 ( .A(REG0_REG_15__SCAN_IN), .B(n4441), .S(n4553), .Z(U3497) );
  MUX2_X1 U4980 ( .A(n4443), .B(n4442), .S(n4553), .Z(n4444) );
  OAI21_X1 U4981 ( .B1(n4445), .B2(n4453), .A(n4444), .ZN(U3495) );
  MUX2_X1 U4982 ( .A(n4447), .B(n4446), .S(n4553), .Z(n4448) );
  OAI21_X1 U4983 ( .B1(n4449), .B2(n4453), .A(n4448), .ZN(U3493) );
  MUX2_X1 U4984 ( .A(n4451), .B(n4450), .S(n4553), .Z(n4452) );
  OAI21_X1 U4985 ( .B1(n4454), .B2(n4453), .A(n4452), .ZN(U3491) );
  MUX2_X1 U4986 ( .A(DATAI_30_), .B(n4455), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4987 ( .A(n4456), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4988 ( .A(n4457), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4989 ( .A(n2738), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4990 ( .A(DATAI_25_), .B(n4458), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4991 ( .A(n4459), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4992 ( .A(DATAI_12_), .B(n4460), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U4993 ( .A(n4461), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4994 ( .A(DATAI_7_), .B(n4462), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4995 ( .A(n4463), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4996 ( .A(n4464), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U4997 ( .A(n4465), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  INV_X1 U4998 ( .A(DATAI_28_), .ZN(n4466) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n4467), .B1(n4466), .B2(U3149), 
        .ZN(U3324) );
  AOI211_X1 U5000 ( .C1(n4470), .C2(n4469), .A(n4468), .B(n4490), .ZN(n4471)
         );
  AOI211_X1 U5001 ( .C1(n4494), .C2(ADDR_REG_15__SCAN_IN), .A(n4472), .B(n4471), .ZN(n4478) );
  AOI21_X1 U5002 ( .B1(n4475), .B2(n4474), .A(n4473), .ZN(n4476) );
  NAND2_X1 U5003 ( .A1(n4498), .A2(n4476), .ZN(n4477) );
  OAI211_X1 U5004 ( .C1(n4500), .C2(n4523), .A(n4478), .B(n4477), .ZN(U3255)
         );
  INV_X1 U5005 ( .A(n4479), .ZN(n4480) );
  AOI21_X1 U5006 ( .B1(n4494), .B2(ADDR_REG_16__SCAN_IN), .A(n4480), .ZN(n4489) );
  OAI21_X1 U5007 ( .B1(n4482), .B2(n4285), .A(n4481), .ZN(n4487) );
  AOI22_X1 U5008 ( .A1(n4498), .A2(n4487), .B1(n4486), .B2(n4485), .ZN(n4488)
         );
  OAI211_X1 U5009 ( .C1(n4521), .C2(n4500), .A(n4489), .B(n4488), .ZN(U3256)
         );
  OAI211_X1 U5010 ( .C1(n4500), .C2(n4519), .A(n2046), .B(n4499), .ZN(U3258)
         );
  AOI22_X1 U5011 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4515), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4510), .ZN(n4505) );
  AOI22_X1 U5012 ( .A1(n4503), .A2(n4502), .B1(n4512), .B2(n4501), .ZN(n4504)
         );
  OAI211_X1 U5013 ( .C1(n4515), .C2(n4506), .A(n4505), .B(n4504), .ZN(U3288)
         );
  AOI21_X1 U5014 ( .B1(n4509), .B2(n4508), .A(n4507), .ZN(n4514) );
  AOI22_X1 U5015 ( .A1(n4512), .A2(n4511), .B1(REG3_REG_0__SCAN_IN), .B2(n4510), .ZN(n4513) );
  OAI221_X1 U5016 ( .B1(n4515), .B2(n4514), .C1(n4313), .C2(n2758), .A(n4513), 
        .ZN(U3290) );
  AND2_X1 U5017 ( .A1(D_REG_31__SCAN_IN), .A2(n4562), .ZN(U3291) );
  AND2_X1 U5018 ( .A1(D_REG_30__SCAN_IN), .A2(n4562), .ZN(U3292) );
  AND2_X1 U5019 ( .A1(D_REG_29__SCAN_IN), .A2(n4562), .ZN(U3293) );
  INV_X1 U5020 ( .A(D_REG_28__SCAN_IN), .ZN(n4620) );
  NOR2_X1 U5021 ( .A1(n4516), .A2(n4620), .ZN(U3294) );
  AND2_X1 U5022 ( .A1(D_REG_27__SCAN_IN), .A2(n4562), .ZN(U3295) );
  AND2_X1 U5023 ( .A1(D_REG_26__SCAN_IN), .A2(n4562), .ZN(U3296) );
  AND2_X1 U5024 ( .A1(D_REG_25__SCAN_IN), .A2(n4562), .ZN(U3297) );
  INV_X1 U5025 ( .A(D_REG_24__SCAN_IN), .ZN(n4656) );
  NOR2_X1 U5026 ( .A1(n4516), .A2(n4656), .ZN(U3298) );
  AND2_X1 U5027 ( .A1(D_REG_23__SCAN_IN), .A2(n4562), .ZN(U3299) );
  AND2_X1 U5028 ( .A1(D_REG_22__SCAN_IN), .A2(n4562), .ZN(U3300) );
  INV_X1 U5029 ( .A(D_REG_21__SCAN_IN), .ZN(n4653) );
  NOR2_X1 U5030 ( .A1(n4516), .A2(n4653), .ZN(U3301) );
  INV_X1 U5031 ( .A(D_REG_20__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U5032 ( .A1(n4516), .A2(n4606), .ZN(U3302) );
  AND2_X1 U5033 ( .A1(D_REG_19__SCAN_IN), .A2(n4562), .ZN(U3303) );
  AND2_X1 U5034 ( .A1(D_REG_18__SCAN_IN), .A2(n4562), .ZN(U3304) );
  AND2_X1 U5035 ( .A1(D_REG_17__SCAN_IN), .A2(n4562), .ZN(U3305) );
  AND2_X1 U5036 ( .A1(D_REG_16__SCAN_IN), .A2(n4562), .ZN(U3306) );
  AND2_X1 U5037 ( .A1(D_REG_15__SCAN_IN), .A2(n4562), .ZN(U3307) );
  INV_X1 U5038 ( .A(D_REG_14__SCAN_IN), .ZN(n4602) );
  NOR2_X1 U5039 ( .A1(n4516), .A2(n4602), .ZN(U3308) );
  INV_X1 U5040 ( .A(D_REG_13__SCAN_IN), .ZN(n4622) );
  NOR2_X1 U5041 ( .A1(n4516), .A2(n4622), .ZN(U3309) );
  AND2_X1 U5042 ( .A1(D_REG_12__SCAN_IN), .A2(n4562), .ZN(U3310) );
  AND2_X1 U5043 ( .A1(D_REG_11__SCAN_IN), .A2(n4562), .ZN(U3311) );
  INV_X1 U5044 ( .A(D_REG_9__SCAN_IN), .ZN(n4652) );
  NOR2_X1 U5045 ( .A1(n4516), .A2(n4652), .ZN(U3313) );
  INV_X1 U5046 ( .A(D_REG_8__SCAN_IN), .ZN(n4655) );
  NOR2_X1 U5047 ( .A1(n4516), .A2(n4655), .ZN(U3314) );
  INV_X1 U5048 ( .A(D_REG_7__SCAN_IN), .ZN(n4601) );
  NOR2_X1 U5049 ( .A1(n4516), .A2(n4601), .ZN(U3315) );
  AND2_X1 U5050 ( .A1(D_REG_6__SCAN_IN), .A2(n4562), .ZN(U3316) );
  AND2_X1 U5051 ( .A1(D_REG_5__SCAN_IN), .A2(n4562), .ZN(U3317) );
  AND2_X1 U5052 ( .A1(D_REG_4__SCAN_IN), .A2(n4562), .ZN(U3318) );
  AND2_X1 U5053 ( .A1(D_REG_3__SCAN_IN), .A2(n4562), .ZN(U3319) );
  AND2_X1 U5054 ( .A1(D_REG_2__SCAN_IN), .A2(n4562), .ZN(U3320) );
  INV_X1 U5055 ( .A(DATAI_23_), .ZN(n4518) );
  AOI21_X1 U5056 ( .B1(U3149), .B2(n4518), .A(n4517), .ZN(U3329) );
  AOI22_X1 U5057 ( .A1(STATE_REG_SCAN_IN), .A2(n4519), .B1(n2547), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5058 ( .A(DATAI_16_), .ZN(n4520) );
  AOI22_X1 U5059 ( .A1(STATE_REG_SCAN_IN), .A2(n4521), .B1(n4520), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5060 ( .A(DATAI_15_), .ZN(n4522) );
  AOI22_X1 U5061 ( .A1(STATE_REG_SCAN_IN), .A2(n4523), .B1(n4522), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5062 ( .A(DATAI_0_), .ZN(n4524) );
  AOI22_X1 U5063 ( .A1(STATE_REG_SCAN_IN), .A2(n4676), .B1(n4524), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5064 ( .A1(n4553), .A2(n4525), .B1(n2322), .B2(n4552), .ZN(U3467)
         );
  AOI22_X1 U5065 ( .A1(n4553), .A2(n4526), .B1(n2307), .B2(n4552), .ZN(U3469)
         );
  OAI22_X1 U5066 ( .A1(n4530), .A2(n4529), .B1(n4528), .B2(n4527), .ZN(n4531)
         );
  NOR2_X1 U5067 ( .A1(n4532), .A2(n4531), .ZN(n4555) );
  AOI22_X1 U5068 ( .A1(n4553), .A2(n4555), .B1(n2343), .B2(n4552), .ZN(U3473)
         );
  INV_X1 U5069 ( .A(n4533), .ZN(n4538) );
  INV_X1 U5070 ( .A(n4534), .ZN(n4536) );
  AOI211_X1 U5071 ( .C1(n4538), .C2(n4537), .A(n4536), .B(n4535), .ZN(n4557)
         );
  AOI22_X1 U5072 ( .A1(n4553), .A2(n4557), .B1(n2358), .B2(n4552), .ZN(U3475)
         );
  NOR2_X1 U5073 ( .A1(n4540), .A2(n4539), .ZN(n4541) );
  AOI211_X1 U5074 ( .C1(n4544), .C2(n4543), .A(n4542), .B(n4541), .ZN(n4558)
         );
  INV_X1 U5075 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5076 ( .A1(n4553), .A2(n4558), .B1(n4545), .B2(n4552), .ZN(U3477)
         );
  NAND3_X1 U5077 ( .A1(n4548), .A2(n4547), .A3(n4546), .ZN(n4549) );
  AND3_X1 U5078 ( .A1(n4551), .A2(n4550), .A3(n4549), .ZN(n4560) );
  AOI22_X1 U5079 ( .A1(n4553), .A2(n4560), .B1(n2400), .B2(n4552), .ZN(U3481)
         );
  INV_X1 U5080 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5081 ( .A1(n4561), .A2(n4555), .B1(n4554), .B2(n4559), .ZN(U3521)
         );
  INV_X1 U5082 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5083 ( .A1(n4561), .A2(n4557), .B1(n4556), .B2(n4559), .ZN(U3522)
         );
  AOI22_X1 U5084 ( .A1(n4561), .A2(n4558), .B1(n2370), .B2(n4559), .ZN(U3523)
         );
  AOI22_X1 U5085 ( .A1(n4561), .A2(n4560), .B1(n2399), .B2(n4559), .ZN(U3525)
         );
  NAND2_X1 U5086 ( .A1(n4562), .A2(D_REG_10__SCAN_IN), .ZN(n4715) );
  XOR2_X1 U5087 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput13), .Z(n4568) );
  XNOR2_X1 U5088 ( .A(n4563), .B(keyinput12), .ZN(n4567) );
  XNOR2_X1 U5089 ( .A(n2652), .B(keyinput38), .ZN(n4566) );
  XNOR2_X1 U5090 ( .A(n4564), .B(keyinput46), .ZN(n4565) );
  NOR4_X1 U5091 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), .ZN(n4573)
         );
  XOR2_X1 U5092 ( .A(n4569), .B(keyinput14), .Z(n4572) );
  XNOR2_X1 U5093 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput59), .ZN(n4571) );
  XNOR2_X1 U5094 ( .A(DATAI_30_), .B(keyinput47), .ZN(n4570) );
  NAND4_X1 U5095 ( .A1(n4573), .A2(n4572), .A3(n4571), .A4(n4570), .ZN(n4600)
         );
  AOI22_X1 U5096 ( .A1(n4575), .A2(keyinput20), .B1(keyinput23), .B2(n4678), 
        .ZN(n4574) );
  OAI221_X1 U5097 ( .B1(n4575), .B2(keyinput20), .C1(n4678), .C2(keyinput23), 
        .A(n4574), .ZN(n4599) );
  AOI22_X1 U5098 ( .A1(n4674), .A2(keyinput43), .B1(n4676), .B2(keyinput34), 
        .ZN(n4576) );
  OAI221_X1 U5099 ( .B1(n4674), .B2(keyinput43), .C1(n4676), .C2(keyinput34), 
        .A(n4576), .ZN(n4598) );
  AOI22_X1 U5100 ( .A1(n4698), .A2(keyinput15), .B1(n4578), .B2(keyinput27), 
        .ZN(n4577) );
  OAI221_X1 U5101 ( .B1(n4698), .B2(keyinput15), .C1(n4578), .C2(keyinput27), 
        .A(n4577), .ZN(n4596) );
  INV_X1 U5102 ( .A(IR_REG_5__SCAN_IN), .ZN(n4677) );
  XOR2_X1 U5103 ( .A(n4677), .B(keyinput5), .Z(n4584) );
  XOR2_X1 U5104 ( .A(n4579), .B(keyinput53), .Z(n4583) );
  INV_X1 U5105 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4580) );
  XOR2_X1 U5106 ( .A(n4580), .B(keyinput2), .Z(n4582) );
  XOR2_X1 U5107 ( .A(n2383), .B(keyinput6), .Z(n4581) );
  NAND4_X1 U5108 ( .A1(n4584), .A2(n4583), .A3(n4582), .A4(n4581), .ZN(n4595)
         );
  XNOR2_X1 U5109 ( .A(IR_REG_25__SCAN_IN), .B(keyinput31), .ZN(n4588) );
  XNOR2_X1 U5110 ( .A(IR_REG_9__SCAN_IN), .B(keyinput44), .ZN(n4587) );
  XNOR2_X1 U5111 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput32), .ZN(n4586) );
  XNOR2_X1 U5112 ( .A(DATAI_7_), .B(keyinput30), .ZN(n4585) );
  NAND4_X1 U5113 ( .A1(n4588), .A2(n4587), .A3(n4586), .A4(n4585), .ZN(n4594)
         );
  XNOR2_X1 U5114 ( .A(IR_REG_11__SCAN_IN), .B(keyinput9), .ZN(n4592) );
  XNOR2_X1 U5115 ( .A(IR_REG_3__SCAN_IN), .B(keyinput63), .ZN(n4591) );
  XNOR2_X1 U5116 ( .A(IR_REG_28__SCAN_IN), .B(keyinput48), .ZN(n4590) );
  XNOR2_X1 U5117 ( .A(IR_REG_26__SCAN_IN), .B(keyinput24), .ZN(n4589) );
  NAND4_X1 U5118 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(n4593)
         );
  OR4_X1 U5119 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(n4597) );
  NOR4_X1 U5120 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4613)
         );
  XOR2_X1 U5121 ( .A(keyinput40), .B(n4601), .Z(n4612) );
  XOR2_X1 U5122 ( .A(keyinput41), .B(n4602), .Z(n4611) );
  INV_X1 U5123 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5124 ( .A1(n4604), .A2(keyinput57), .B1(n3232), .B2(keyinput10), 
        .ZN(n4603) );
  OAI221_X1 U5125 ( .B1(n4604), .B2(keyinput57), .C1(n3232), .C2(keyinput10), 
        .A(n4603), .ZN(n4609) );
  AOI22_X1 U5126 ( .A1(n2445), .A2(keyinput60), .B1(n2335), .B2(keyinput52), 
        .ZN(n4605) );
  OAI221_X1 U5127 ( .B1(n2445), .B2(keyinput60), .C1(n2335), .C2(keyinput52), 
        .A(n4605), .ZN(n4608) );
  XNOR2_X1 U5128 ( .A(n4606), .B(keyinput29), .ZN(n4607) );
  NOR3_X1 U5129 ( .A1(n4609), .A2(n4608), .A3(n4607), .ZN(n4610) );
  NAND4_X1 U5130 ( .A1(n4613), .A2(n4612), .A3(n4611), .A4(n4610), .ZN(n4640)
         );
  AOI22_X1 U5131 ( .A1(n2783), .A2(keyinput11), .B1(n2398), .B2(keyinput45), 
        .ZN(n4614) );
  OAI221_X1 U5132 ( .B1(n2783), .B2(keyinput11), .C1(n2398), .C2(keyinput45), 
        .A(n4614), .ZN(n4618) );
  AOI22_X1 U5133 ( .A1(n4616), .A2(keyinput39), .B1(keyinput55), .B2(n4671), 
        .ZN(n4615) );
  OAI221_X1 U5134 ( .B1(n4616), .B2(keyinput39), .C1(n4671), .C2(keyinput55), 
        .A(n4615), .ZN(n4617) );
  NOR2_X1 U5135 ( .A1(n4618), .A2(n4617), .ZN(n4638) );
  AOI22_X1 U5136 ( .A1(n4697), .A2(keyinput17), .B1(n4620), .B2(keyinput8), 
        .ZN(n4619) );
  OAI221_X1 U5137 ( .B1(n4697), .B2(keyinput17), .C1(n4620), .C2(keyinput8), 
        .A(n4619), .ZN(n4624) );
  AOI22_X1 U5138 ( .A1(n4670), .A2(keyinput49), .B1(n4622), .B2(keyinput50), 
        .ZN(n4621) );
  OAI221_X1 U5139 ( .B1(n4670), .B2(keyinput49), .C1(n4622), .C2(keyinput50), 
        .A(n4621), .ZN(n4623) );
  NOR2_X1 U5140 ( .A1(n4624), .A2(n4623), .ZN(n4637) );
  AOI22_X1 U5141 ( .A1(n2603), .A2(keyinput22), .B1(n4285), .B2(keyinput62), 
        .ZN(n4625) );
  OAI221_X1 U5142 ( .B1(n2603), .B2(keyinput22), .C1(n4285), .C2(keyinput62), 
        .A(n4625), .ZN(n4629) );
  INV_X1 U5143 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5144 ( .A1(n3223), .A2(keyinput35), .B1(keyinput37), .B2(n4627), 
        .ZN(n4626) );
  OAI221_X1 U5145 ( .B1(n3223), .B2(keyinput35), .C1(n4627), .C2(keyinput37), 
        .A(n4626), .ZN(n4628) );
  NOR2_X1 U5146 ( .A1(n4629), .A2(n4628), .ZN(n4636) );
  AOI22_X1 U5147 ( .A1(n2381), .A2(keyinput1), .B1(n2400), .B2(keyinput0), 
        .ZN(n4630) );
  OAI221_X1 U5148 ( .B1(n2381), .B2(keyinput1), .C1(n2400), .C2(keyinput0), 
        .A(n4630), .ZN(n4634) );
  AOI22_X1 U5149 ( .A1(n4669), .A2(keyinput58), .B1(n4632), .B2(keyinput61), 
        .ZN(n4631) );
  OAI221_X1 U5150 ( .B1(n4669), .B2(keyinput58), .C1(n4632), .C2(keyinput61), 
        .A(n4631), .ZN(n4633) );
  NOR2_X1 U5151 ( .A1(n4634), .A2(n4633), .ZN(n4635) );
  NAND4_X1 U5152 ( .A1(n4638), .A2(n4637), .A3(n4636), .A4(n4635), .ZN(n4639)
         );
  NOR2_X1 U5153 ( .A1(n4640), .A2(n4639), .ZN(n4665) );
  INV_X1 U5154 ( .A(keyinput36), .ZN(n4642) );
  XNOR2_X1 U5155 ( .A(REG2_REG_17__SCAN_IN), .B(keyinput42), .ZN(n4641) );
  OAI21_X1 U5156 ( .B1(IR_REG_4__SCAN_IN), .B2(n4642), .A(n4641), .ZN(n4650)
         );
  AOI22_X1 U5157 ( .A1(n2881), .A2(keyinput21), .B1(n2700), .B2(keyinput25), 
        .ZN(n4643) );
  OAI221_X1 U5158 ( .B1(n2881), .B2(keyinput21), .C1(n2700), .C2(keyinput25), 
        .A(n4643), .ZN(n4649) );
  INV_X1 U5159 ( .A(B_REG_SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5160 ( .A1(n4705), .A2(keyinput54), .B1(n4683), .B2(keyinput19), 
        .ZN(n4644) );
  OAI221_X1 U5161 ( .B1(n4705), .B2(keyinput54), .C1(n4683), .C2(keyinput19), 
        .A(n4644), .ZN(n4648) );
  AOI22_X1 U5162 ( .A1(n4666), .A2(keyinput51), .B1(n4646), .B2(keyinput7), 
        .ZN(n4645) );
  OAI221_X1 U5163 ( .B1(n4666), .B2(keyinput51), .C1(n4646), .C2(keyinput7), 
        .A(n4645), .ZN(n4647) );
  NOR4_X1 U5164 ( .A1(n4650), .A2(n4649), .A3(n4648), .A4(n4647), .ZN(n4664)
         );
  AOI22_X1 U5165 ( .A1(n4653), .A2(keyinput18), .B1(keyinput28), .B2(n4652), 
        .ZN(n4651) );
  OAI221_X1 U5166 ( .B1(n4653), .B2(keyinput18), .C1(n4652), .C2(keyinput28), 
        .A(n4651), .ZN(n4662) );
  AOI22_X1 U5167 ( .A1(n4656), .A2(keyinput16), .B1(keyinput4), .B2(n4655), 
        .ZN(n4654) );
  OAI221_X1 U5168 ( .B1(n4656), .B2(keyinput16), .C1(n4655), .C2(keyinput4), 
        .A(n4654), .ZN(n4661) );
  AOI22_X1 U5169 ( .A1(n4680), .A2(keyinput26), .B1(n4679), .B2(keyinput56), 
        .ZN(n4657) );
  OAI221_X1 U5170 ( .B1(n4680), .B2(keyinput26), .C1(n4679), .C2(keyinput56), 
        .A(n4657), .ZN(n4660) );
  AOI22_X1 U5171 ( .A1(n4667), .A2(keyinput3), .B1(n4668), .B2(keyinput33), 
        .ZN(n4658) );
  OAI221_X1 U5172 ( .B1(n4667), .B2(keyinput3), .C1(n4668), .C2(keyinput33), 
        .A(n4658), .ZN(n4659) );
  NOR4_X1 U5173 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4663)
         );
  NAND3_X1 U5174 ( .A1(n4665), .A2(n4664), .A3(n4663), .ZN(n4713) );
  NOR4_X1 U5175 ( .A1(REG2_REG_16__SCAN_IN), .A2(REG2_REG_30__SCAN_IN), .A3(
        n2603), .A4(n4666), .ZN(n4704) );
  AND4_X1 U5176 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(n4668), 
        .A4(n4667), .ZN(n4672) );
  AND4_X1 U5177 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4703)
         );
  INV_X1 U5178 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4673) );
  NAND4_X1 U5179 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(REG1_REG_0__SCAN_IN), .ZN(n4691) );
  NAND4_X1 U5180 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .A3(n4677), 
        .A4(n4676), .ZN(n4682) );
  NAND4_X1 U5181 ( .A1(REG1_REG_27__SCAN_IN), .A2(n4680), .A3(n4679), .A4(
        n4678), .ZN(n4681) );
  NOR2_X1 U5182 ( .A1(n4682), .A2(n4681), .ZN(n4686) );
  NOR4_X1 U5183 ( .A1(REG0_REG_7__SCAN_IN), .A2(REG2_REG_7__SCAN_IN), .A3(
        REG0_REG_6__SCAN_IN), .A4(n2383), .ZN(n4685) );
  AND4_X1 U5184 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .A3(
        IR_REG_26__SCAN_IN), .A4(n4683), .ZN(n4684) );
  AND4_X1 U5185 ( .A1(n4686), .A2(n2783), .A3(n4685), .A4(n4684), .ZN(n4687)
         );
  NAND4_X1 U5186 ( .A1(n4689), .A2(n4688), .A3(REG3_REG_11__SCAN_IN), .A4(
        n4687), .ZN(n4690) );
  NOR2_X1 U5187 ( .A1(n4691), .A2(n4690), .ZN(n4696) );
  NAND4_X1 U5188 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(REG3_REG_7__SCAN_IN), .ZN(n4694) );
  INV_X1 U5189 ( .A(DATAI_30_), .ZN(n4692) );
  NAND4_X1 U5190 ( .A1(n4627), .A2(n4692), .A3(DATAO_REG_16__SCAN_IN), .A4(
        ADDR_REG_16__SCAN_IN), .ZN(n4693) );
  NOR2_X1 U5191 ( .A1(n4694), .A2(n4693), .ZN(n4695) );
  AND2_X1 U5192 ( .A1(n4696), .A2(n4695), .ZN(n4702) );
  NAND4_X1 U5193 ( .A1(REG3_REG_4__SCAN_IN), .A2(DATAI_7_), .A3(
        DATAO_REG_2__SCAN_IN), .A4(n2445), .ZN(n4700) );
  NAND4_X1 U5194 ( .A1(REG3_REG_16__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        n4698), .A4(n4697), .ZN(n4699) );
  NOR2_X1 U5195 ( .A1(n4700), .A2(n4699), .ZN(n4701) );
  AND4_X1 U5196 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), .ZN(n4708)
         );
  NOR4_X1 U5197 ( .A1(REG1_REG_6__SCAN_IN), .A2(REG2_REG_8__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(n3223), .ZN(n4707) );
  NOR4_X1 U5198 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG2_REG_17__SCAN_IN), .A3(
        n4705), .A4(n2881), .ZN(n4706) );
  NAND4_X1 U5199 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n4711)
         );
  AOI21_X1 U5200 ( .B1(n4711), .B2(n4710), .A(keyinput36), .ZN(n4712) );
  NOR2_X1 U5201 ( .A1(n4713), .A2(n4712), .ZN(n4714) );
  XNOR2_X1 U5202 ( .A(n4715), .B(n4714), .ZN(U3312) );
  OR2_X1 U2260 ( .A1(n2871), .A2(n2671), .ZN(n3802) );
  CLKBUF_X1 U2473 ( .A(n2369), .Z(n2646) );
  CLKBUF_X1 U2887 ( .A(n4259), .Z(n2064) );
  AND4_X1 U3029 ( .A1(n2366), .A2(n2297), .A3(n2296), .A4(n4689), .ZN(n4718)
         );
endmodule

