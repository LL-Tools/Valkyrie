

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9597, n9598, n9600, n9603, n9605, n9606, n9607, n9608, n9609, n9610,
         n9612, n9613, n9615, n9616, n9617, n9618, n9619, n9620, n9622, n9623,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472;

  OR2_X1 U11041 ( .A1(n16281), .A2(n19668), .ZN(n9810) );
  INV_X1 U11042 ( .A(n18264), .ZN(n18558) );
  INV_X1 U11043 ( .A(n18100), .ZN(n18118) );
  MUX2_X1 U11044 ( .A(n12603), .B(n12602), .S(n12601), .Z(n12604) );
  INV_X1 U11045 ( .A(n17599), .ZN(n17581) );
  CLKBUF_X2 U11046 ( .A(n15046), .Z(n9623) );
  AND2_X1 U11047 ( .A1(n12378), .A2(n15818), .ZN(n15482) );
  AND4_X1 U11049 ( .A1(n10075), .A2(n10078), .A3(n10084), .A4(n10076), .ZN(
        n10072) );
  NOR2_X1 U11050 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  AOI22_X1 U11051 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19843), .B1(
        n19685), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12420) );
  INV_X1 U11052 ( .A(n10570), .ZN(n9821) );
  NOR2_X1 U11053 ( .A1(n19517), .A2(n19518), .ZN(n13470) );
  BUF_X2 U11054 ( .A(n10453), .Z(n10561) );
  INV_X2 U11055 ( .A(n17931), .ZN(n17799) );
  NOR2_X1 U11056 ( .A1(n12777), .A2(n16142), .ZN(n12780) );
  INV_X1 U11057 ( .A(n16942), .ZN(n17932) );
  NOR2_X1 U11058 ( .A1(n19562), .A2(n16219), .ZN(n19534) );
  INV_X4 U11059 ( .A(n12281), .ZN(n12282) );
  INV_X2 U11060 ( .A(n17950), .ZN(n17858) );
  CLKBUF_X2 U11061 ( .A(n10447), .Z(n13411) );
  AND2_X1 U11062 ( .A1(n10414), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10479) );
  CLKBUF_X2 U11063 ( .A(n12365), .Z(n16554) );
  MUX2_X1 U11064 ( .A(n17084), .B(n11241), .S(n21084), .Z(n10430) );
  AND2_X2 U11065 ( .A1(n13077), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12058) );
  AND2_X2 U11066 ( .A1(n13076), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12126) );
  CLKBUF_X2 U11067 ( .A(n13266), .Z(n14305) );
  NAND2_X1 U11068 ( .A1(n13946), .A2(n10432), .ZN(n13824) );
  MUX2_X1 U11069 ( .A(n11789), .B(n12066), .S(n16546), .Z(n11790) );
  INV_X4 U11070 ( .A(n9754), .ZN(n17036) );
  NOR2_X1 U11071 ( .A1(n12759), .A2(n16236), .ZN(n12761) );
  AND2_X1 U11072 ( .A1(n10597), .A2(n14116), .ZN(n10312) );
  INV_X2 U11073 ( .A(n11252), .ZN(n17941) );
  INV_X4 U11074 ( .A(n9668), .ZN(n17020) );
  NAND3_X1 U11075 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12759) );
  CLKBUF_X2 U11076 ( .A(n10525), .Z(n13404) );
  CLKBUF_X2 U11077 ( .A(n10466), .Z(n11220) );
  CLKBUF_X2 U11078 ( .A(n10402), .Z(n13405) );
  CLKBUF_X2 U11079 ( .A(n10446), .Z(n11123) );
  CLKBUF_X2 U11080 ( .A(n10532), .Z(n9615) );
  CLKBUF_X2 U11081 ( .A(n11759), .Z(n16542) );
  CLKBUF_X2 U11083 ( .A(n9600), .Z(n10467) );
  CLKBUF_X2 U11084 ( .A(n9626), .Z(n10454) );
  NAND2_X1 U11086 ( .A1(n11743), .A2(n11744), .ZN(n12309) );
  AND2_X1 U11087 ( .A1(n11747), .A2(n16566), .ZN(n12045) );
  INV_X1 U11088 ( .A(n16558), .ZN(n13646) );
  AND4_X1 U11089 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10349) );
  AND4_X1 U11090 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10350) );
  NAND2_X1 U11091 ( .A1(n10042), .A2(n10041), .ZN(n11753) );
  AND2_X2 U11092 ( .A1(n10323), .A2(n15370), .ZN(n10533) );
  AND2_X1 U11093 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15365) );
  AND2_X1 U11094 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15370) );
  AND2_X2 U11095 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14273) );
  NAND2_X1 U11097 ( .A1(n9873), .A2(n12425), .ZN(n12426) );
  AND2_X1 U11098 ( .A1(n9873), .A2(n9748), .ZN(n10012) );
  NAND4_X1 U11099 ( .A1(n10069), .A2(n10068), .A3(n10072), .A4(n9669), .ZN(
        n9873) );
  NOR2_X2 U11100 ( .A1(n15578), .A2(n15579), .ZN(n15567) );
  XNOR2_X2 U11101 ( .A(n12755), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12946) );
  NAND2_X2 U11102 ( .A1(n16249), .A2(n16250), .ZN(n16252) );
  CLKBUF_X3 U11103 ( .A(n12403), .Z(n16572) );
  NAND4_X1 U11104 ( .A1(n9958), .A2(n9957), .A3(n9837), .A4(n9956), .ZN(n9597)
         );
  NAND2_X1 U11105 ( .A1(n9636), .A2(n9630), .ZN(n9598) );
  AND2_X2 U11107 ( .A1(n9598), .A2(n21471), .ZN(n12610) );
  AND2_X2 U11108 ( .A1(n10322), .A2(n9989), .ZN(n9600) );
  NAND3_X1 U11110 ( .A1(n10427), .A2(n21472), .A3(n10426), .ZN(n9817) );
  NAND2_X2 U11112 ( .A1(n15045), .A2(n10704), .ZN(n9603) );
  AND2_X1 U11113 ( .A1(n10322), .A2(n9989), .ZN(n10556) );
  NAND2_X1 U11114 ( .A1(n15045), .A2(n10704), .ZN(n10062) );
  MUX2_X2 U11115 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12946), .S(
        n17153), .Z(n19559) );
  NOR2_X1 U11117 ( .A1(n12065), .A2(n16566), .ZN(n11743) );
  INV_X1 U11118 ( .A(n11904), .ZN(n11899) );
  NAND2_X1 U11119 ( .A1(n16663), .A2(n13923), .ZN(n11593) );
  AND4_X1 U11120 ( .A1(n15051), .A2(n15057), .A3(n10703), .A4(n15053), .ZN(
        n10704) );
  AND2_X1 U11121 ( .A1(n9688), .A2(n10311), .ZN(n14116) );
  AND2_X1 U11122 ( .A1(n12482), .A2(n12483), .ZN(n12485) );
  AND3_X1 U11123 ( .A1(n11809), .A2(n11805), .A3(n11808), .ZN(n11810) );
  INV_X1 U11124 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16519) );
  AND2_X1 U11125 ( .A1(n11620), .A2(n10144), .ZN(n11623) );
  INV_X1 U11126 ( .A(n11447), .ZN(n11436) );
  NAND2_X1 U11127 ( .A1(n11042), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11157) );
  AND2_X1 U11128 ( .A1(n15103), .A2(n10700), .ZN(n15051) );
  INV_X1 U11129 ( .A(n15049), .ZN(n15046) );
  INV_X1 U11131 ( .A(n12309), .ZN(n12311) );
  AND4_X1 U11132 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12354) );
  AND2_X1 U11133 ( .A1(n12570), .A2(n10196), .ZN(n10195) );
  INV_X2 U11134 ( .A(n12354), .ZN(n12644) );
  INV_X2 U11136 ( .A(n17941), .ZN(n17898) );
  INV_X1 U11137 ( .A(n17891), .ZN(n17878) );
  NOR2_X2 U11138 ( .A1(n18301), .A2(n18339), .ZN(n11620) );
  AND2_X1 U11139 ( .A1(n16930), .A2(n11253), .ZN(n11465) );
  CLKBUF_X3 U11140 ( .A(n14305), .Z(n13361) );
  INV_X2 U11141 ( .A(n10431), .ZN(n13946) );
  AND2_X1 U11142 ( .A1(n14955), .A2(n9645), .ZN(n14398) );
  NAND2_X1 U11143 ( .A1(n11669), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11676) );
  OR2_X1 U11144 ( .A1(n13747), .A2(n13820), .ZN(n13891) );
  OR2_X1 U11145 ( .A1(n12400), .A2(n12399), .ZN(n12402) );
  OAI21_X1 U11146 ( .B1(n10052), .B2(n10051), .A(n10049), .ZN(n16100) );
  XNOR2_X1 U11147 ( .A(n9597), .B(n16469), .ZN(n16214) );
  NOR2_X1 U11149 ( .A1(n18899), .A2(n18896), .ZN(n11520) );
  INV_X1 U11150 ( .A(n18417), .ZN(n18402) );
  NOR2_X1 U11151 ( .A1(n11460), .A2(n11459), .ZN(n11531) );
  INV_X1 U11152 ( .A(n14772), .ZN(n13435) );
  AND2_X1 U11153 ( .A1(n14644), .A2(n13316), .ZN(n14631) );
  NAND2_X1 U11154 ( .A1(n14202), .A2(n14217), .ZN(n14216) );
  INV_X1 U11155 ( .A(n10432), .ZN(n10476) );
  INV_X1 U11157 ( .A(n15772), .ZN(n15773) );
  NOR2_X2 U11158 ( .A1(n13891), .A2(n13890), .ZN(n13893) );
  NAND2_X1 U11159 ( .A1(n12742), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16174) );
  INV_X1 U11160 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20318) );
  INV_X1 U11161 ( .A(n17595), .ZN(n17525) );
  INV_X1 U11162 ( .A(n18873), .ZN(n18133) );
  AND2_X1 U11163 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18562), .ZN(n18417) );
  NAND2_X1 U11164 ( .A1(n15683), .A2(n19563), .ZN(n15772) );
  INV_X2 U11165 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13875) );
  NAND2_X1 U11166 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17573), .ZN(n17595) );
  AND4_X1 U11168 ( .A1(n11803), .A2(n11802), .A3(n15432), .A4(n11801), .ZN(
        n9605) );
  AND2_X1 U11169 ( .A1(n9769), .A2(n12413), .ZN(n9606) );
  AND2_X2 U11170 ( .A1(n10324), .A2(n15370), .ZN(n9626) );
  AND4_X1 U11171 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n9607) );
  AND2_X2 U11172 ( .A1(n10323), .A2(n15370), .ZN(n9627) );
  NOR2_X2 U11174 ( .A1(n14553), .A2(n14555), .ZN(n14542) );
  BUF_X4 U11175 ( .A(n11737), .Z(n13207) );
  NAND2_X2 U11176 ( .A1(n14208), .A2(n10696), .ZN(n10698) );
  AND4_X2 U11177 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10339) );
  NOR2_X2 U11178 ( .A1(n9663), .A2(n12714), .ZN(n12715) );
  NOR2_X2 U11179 ( .A1(n11539), .A2(n11538), .ZN(n11543) );
  AND2_X4 U11180 ( .A1(n11701), .A2(n11700), .ZN(n12065) );
  NOR2_X2 U11181 ( .A1(n16636), .A2(n18495), .ZN(n12900) );
  NAND2_X2 U11182 ( .A1(n14167), .A2(n10548), .ZN(n13729) );
  NAND2_X1 U11183 ( .A1(n16127), .A2(n16101), .ZN(n16126) );
  AOI21_X1 U11184 ( .B1(n15799), .B2(n10200), .A(n15794), .ZN(n15787) );
  AOI21_X1 U11185 ( .B1(n15804), .B2(n13150), .A(n13149), .ZN(n13167) );
  AND2_X1 U11186 ( .A1(n10259), .A2(n16186), .ZN(n10255) );
  AND2_X1 U11187 ( .A1(n16724), .A2(n9746), .ZN(n16707) );
  XNOR2_X1 U11188 ( .A(n12693), .B(n12290), .ZN(n14462) );
  AND2_X1 U11189 ( .A1(n11405), .A2(n9920), .ZN(n16706) );
  NAND2_X1 U11190 ( .A1(n9800), .A2(n12610), .ZN(n12642) );
  XNOR2_X1 U11191 ( .A(n14309), .B(n14308), .ZN(n14404) );
  NAND2_X1 U11192 ( .A1(n12257), .A2(n12256), .ZN(n15635) );
  NAND2_X1 U11193 ( .A1(n11635), .A2(n11634), .ZN(n18462) );
  NAND2_X1 U11194 ( .A1(n11159), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11198) );
  OR2_X1 U11195 ( .A1(n10813), .A2(n10973), .ZN(n10820) );
  INV_X4 U11196 ( .A(n18484), .ZN(n18557) );
  AND2_X2 U11197 ( .A1(n9769), .A2(n12414), .ZN(n9641) );
  AND2_X2 U11198 ( .A1(n12415), .A2(n9769), .ZN(n20037) );
  NAND2_X1 U11199 ( .A1(n11063), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11066) );
  NAND2_X1 U11200 ( .A1(n9821), .A2(n10604), .ZN(n14162) );
  OR2_X1 U11201 ( .A1(n13921), .A2(n10030), .ZN(n18070) );
  NOR2_X2 U11202 ( .A1(n19300), .A2(n18851), .ZN(n18736) );
  NAND2_X1 U11203 ( .A1(n10770), .A2(n10769), .ZN(n14173) );
  NOR2_X2 U11204 ( .A1(n12480), .A2(n12353), .ZN(n12482) );
  BUF_X1 U11205 ( .A(n11804), .Z(n11814) );
  NOR2_X2 U11206 ( .A1(n18910), .A2(n11531), .ZN(n11544) );
  NAND2_X4 U11207 ( .A1(n13274), .A2(n14305), .ZN(n14307) );
  INV_X2 U11208 ( .A(n19471), .ZN(n13916) );
  INV_X1 U11209 ( .A(n12090), .ZN(n12280) );
  NOR2_X1 U11210 ( .A1(n11501), .A2(n11500), .ZN(n11517) );
  CLKBUF_X2 U11211 ( .A(n11951), .Z(n12004) );
  BUF_X1 U11212 ( .A(n11753), .Z(n16549) );
  INV_X4 U11213 ( .A(n11436), .ZN(n17877) );
  INV_X4 U11214 ( .A(n9666), .ZN(n17921) );
  INV_X4 U11215 ( .A(n17943), .ZN(n9608) );
  INV_X2 U11216 ( .A(n11411), .ZN(n17939) );
  INV_X1 U11217 ( .A(n16574), .ZN(n9609) );
  INV_X4 U11218 ( .A(n17747), .ZN(n11322) );
  NAND4_X2 U11219 ( .A1(n9896), .A2(n11253), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17747) );
  INV_X2 U11220 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16900) );
  NAND2_X1 U11221 ( .A1(n10007), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14415) );
  OAI21_X1 U11222 ( .B1(n16345), .B2(n14265), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9793) );
  INV_X1 U11223 ( .A(n14260), .ZN(n9970) );
  OR2_X1 U11224 ( .A1(n16174), .A2(n16141), .ZN(n16147) );
  AOI211_X1 U11225 ( .C1(n16342), .C2(n19672), .A(n16341), .B(n16340), .ZN(
        n16343) );
  XNOR2_X1 U11226 ( .A(n10057), .B(n10056), .ZN(n16085) );
  AND2_X1 U11227 ( .A1(n9804), .A2(n9801), .ZN(n16020) );
  NAND2_X1 U11228 ( .A1(n16049), .A2(n12581), .ZN(n16314) );
  NOR2_X1 U11229 ( .A1(n11247), .A2(n11246), .ZN(n11248) );
  XNOR2_X1 U11230 ( .A(n14313), .B(n14312), .ZN(n14432) );
  NOR2_X1 U11231 ( .A1(n12339), .A2(n12338), .ZN(n12654) );
  NAND2_X1 U11232 ( .A1(n17291), .A2(n17290), .ZN(n17289) );
  AND2_X1 U11233 ( .A1(n9798), .A2(n9720), .ZN(n9876) );
  XNOR2_X1 U11234 ( .A(n14467), .B(n13432), .ZN(n14443) );
  AND2_X1 U11235 ( .A1(n9785), .A2(n12646), .ZN(n10089) );
  OR2_X1 U11236 ( .A1(n15080), .A2(n15077), .ZN(n15076) );
  NOR2_X1 U11237 ( .A1(n13167), .A2(n13166), .ZN(n15793) );
  CLKBUF_X1 U11238 ( .A(n14466), .Z(n14480) );
  NAND2_X1 U11239 ( .A1(n17298), .A2(n17300), .ZN(n17299) );
  AOI21_X1 U11240 ( .B1(n14579), .B2(n14570), .A(n14569), .ZN(n15018) );
  AND2_X1 U11241 ( .A1(n14569), .A2(n14509), .ZN(n14526) );
  NOR2_X1 U11242 ( .A1(n10260), .A2(n10088), .ZN(n9799) );
  NAND2_X1 U11243 ( .A1(n16707), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16673) );
  INV_X1 U11244 ( .A(n14551), .ZN(n14569) );
  NOR2_X1 U11245 ( .A1(n14614), .A2(n14596), .ZN(n14595) );
  NAND2_X1 U11246 ( .A1(n16197), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10260) );
  OR2_X1 U11247 ( .A1(n14551), .A2(n14552), .ZN(n14549) );
  XNOR2_X1 U11248 ( .A(n12643), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16186) );
  AND2_X1 U11249 ( .A1(n15805), .A2(n15809), .ZN(n13149) );
  AND2_X1 U11250 ( .A1(n12490), .A2(n10278), .ZN(n10048) );
  AND3_X1 U11251 ( .A1(n16159), .A2(n16202), .A3(n16189), .ZN(n12490) );
  NAND2_X1 U11252 ( .A1(n14629), .A2(n14508), .ZN(n14551) );
  NOR2_X1 U11253 ( .A1(n14671), .A2(n14656), .ZN(n14655) );
  AND2_X1 U11254 ( .A1(n13145), .A2(n13144), .ZN(n15805) );
  NAND2_X1 U11255 ( .A1(n10256), .A2(n16451), .ZN(n10259) );
  INV_X1 U11256 ( .A(n10256), .ZN(n16197) );
  NAND2_X1 U11257 ( .A1(n14629), .A2(n14615), .ZN(n14614) );
  NAND2_X1 U11258 ( .A1(n10006), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10066) );
  XNOR2_X1 U11259 ( .A(n12642), .B(n12354), .ZN(n10256) );
  INV_X1 U11260 ( .A(n12642), .ZN(n12645) );
  NOR2_X1 U11261 ( .A1(n12581), .A2(n9869), .ZN(n9868) );
  NAND2_X1 U11262 ( .A1(n17320), .A2(n17321), .ZN(n17319) );
  NAND4_X1 U11263 ( .A1(n9958), .A2(n9957), .A3(n9837), .A4(n9956), .ZN(n9771)
         );
  AND2_X1 U11264 ( .A1(n14729), .A2(n9719), .ZN(n14507) );
  NAND2_X1 U11265 ( .A1(n12635), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12637) );
  AND2_X1 U11266 ( .A1(n14729), .A2(n10115), .ZN(n14690) );
  OAI21_X1 U11267 ( .B1(n15472), .B2(n16025), .A(n19563), .ZN(n15462) );
  NAND2_X1 U11268 ( .A1(n12630), .A2(n12629), .ZN(n16239) );
  NOR2_X1 U11269 ( .A1(n10061), .A2(n9755), .ZN(n10060) );
  NOR2_X1 U11270 ( .A1(n14197), .A2(n14240), .ZN(n14238) );
  AND2_X1 U11271 ( .A1(n12864), .A2(n16071), .ZN(n14283) );
  AND2_X1 U11272 ( .A1(n15089), .A2(n10699), .ZN(n15103) );
  OR2_X1 U11273 ( .A1(n15054), .A2(n9653), .ZN(n10061) );
  NAND2_X1 U11274 ( .A1(n9877), .A2(n12467), .ZN(n12481) );
  NOR2_X2 U11275 ( .A1(n20094), .A2(n19942), .ZN(n19965) );
  NAND2_X1 U11276 ( .A1(n9812), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10697) );
  NOR2_X2 U11277 ( .A1(n19881), .A2(n20156), .ZN(n10291) );
  NOR2_X2 U11278 ( .A1(n20073), .A2(n20156), .ZN(n20204) );
  NOR2_X2 U11279 ( .A1(n19840), .A2(n20304), .ZN(n19770) );
  NAND2_X1 U11280 ( .A1(n10135), .A2(n18263), .ZN(n17351) );
  AND2_X1 U11281 ( .A1(n15098), .A2(n10694), .ZN(n14209) );
  AND2_X1 U11282 ( .A1(n10674), .A2(n10673), .ZN(n17101) );
  AND2_X1 U11283 ( .A1(n11399), .A2(n16748), .ZN(n10160) );
  AND4_X1 U11284 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(n9880)
         );
  NAND2_X1 U11285 ( .A1(n10820), .A2(n10819), .ZN(n14003) );
  AND2_X1 U11286 ( .A1(n10812), .A2(n10811), .ZN(n14054) );
  NOR2_X1 U11287 ( .A1(n16463), .A2(n12331), .ZN(n10023) );
  AND2_X1 U11288 ( .A1(n17581), .A2(n12932), .ZN(n17328) );
  AOI22_X1 U11289 ( .A1(n20037), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n19718), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12419) );
  NOR2_X2 U11290 ( .A1(n18552), .A2(n16771), .ZN(n18436) );
  NAND2_X1 U11291 ( .A1(n13773), .A2(n12967), .ZN(n13784) );
  NAND2_X2 U11292 ( .A1(n17257), .A2(n11614), .ZN(n18547) );
  NAND2_X1 U11293 ( .A1(n9992), .A2(n10634), .ZN(n14058) );
  OR2_X1 U11294 ( .A1(n10805), .A2(n10973), .ZN(n10812) );
  NAND2_X1 U11295 ( .A1(n9808), .A2(n9807), .ZN(n12526) );
  AND2_X1 U11296 ( .A1(n12416), .A2(n12413), .ZN(n12461) );
  NAND2_X1 U11297 ( .A1(n9993), .A2(n10640), .ZN(n15413) );
  NAND2_X1 U11298 ( .A1(n18472), .A2(n11387), .ZN(n11394) );
  NAND2_X1 U11299 ( .A1(n15407), .A2(n9821), .ZN(n9993) );
  INV_X1 U11300 ( .A(n12524), .ZN(n9808) );
  XNOR2_X1 U11301 ( .A(n12966), .B(n12964), .ZN(n13769) );
  NAND2_X1 U11302 ( .A1(n17380), .A2(n18305), .ZN(n17379) );
  NAND3_X1 U11303 ( .A1(n10570), .A2(n10248), .A3(n10631), .ZN(n10642) );
  OR2_X1 U11304 ( .A1(n19295), .A2(n11580), .ZN(n9894) );
  NOR2_X1 U11305 ( .A1(n11608), .A2(n11607), .ZN(n18469) );
  AOI21_X1 U11306 ( .B1(n9775), .B2(n13674), .A(n12963), .ZN(n13770) );
  INV_X2 U11307 ( .A(n19575), .ZN(n19570) );
  INV_X2 U11308 ( .A(n13981), .ZN(n20512) );
  NAND2_X1 U11309 ( .A1(n17391), .A2(n18320), .ZN(n17392) );
  XNOR2_X1 U11310 ( .A(n13644), .B(n12961), .ZN(n13674) );
  NAND2_X1 U11311 ( .A1(n9919), .A2(n10148), .ZN(n11386) );
  NAND2_X1 U11312 ( .A1(n20452), .A2(n14444), .ZN(n14835) );
  CLKBUF_X1 U11313 ( .A(n20691), .Z(n9622) );
  NOR2_X1 U11314 ( .A1(n16486), .A2(n19643), .ZN(n12413) );
  OAI21_X1 U11315 ( .B1(n16486), .B2(n15428), .A(n12957), .ZN(n13675) );
  AND2_X2 U11316 ( .A1(n18736), .A2(n18746), .ZN(n18773) );
  AND2_X1 U11317 ( .A1(n16486), .A2(n15779), .ZN(n12415) );
  AND2_X1 U11318 ( .A1(n17051), .A2(n12927), .ZN(n19293) );
  NAND2_X1 U11319 ( .A1(n12926), .A2(n16914), .ZN(n17051) );
  NAND2_X1 U11320 ( .A1(n12542), .A2(n12492), .ZN(n12538) );
  OAI21_X1 U11321 ( .B1(n11378), .B2(n10150), .A(n11382), .ZN(n10149) );
  OR2_X1 U11322 ( .A1(n12497), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12533) );
  XNOR2_X1 U11323 ( .A(n10615), .B(n10780), .ZN(n21093) );
  NAND2_X1 U11324 ( .A1(n12482), .A2(n9699), .ZN(n12492) );
  NAND2_X1 U11325 ( .A1(n11782), .A2(n11781), .ZN(n11783) );
  OR2_X1 U11326 ( .A1(n10970), .A2(n14662), .ZN(n10943) );
  NAND4_X1 U11327 ( .A1(n10254), .A2(n11769), .A3(n10253), .A4(n9635), .ZN(
        n11813) );
  NAND2_X1 U11328 ( .A1(n10172), .A2(n10173), .ZN(n12480) );
  AND2_X1 U11329 ( .A1(n10544), .A2(n10543), .ZN(n14168) );
  INV_X1 U11330 ( .A(n12444), .ZN(n10173) );
  NAND2_X1 U11331 ( .A1(n9605), .A2(n11810), .ZN(n12399) );
  NAND2_X1 U11332 ( .A1(n10018), .A2(n18189), .ZN(n11542) );
  NAND2_X1 U11333 ( .A1(n12429), .A2(n12430), .ZN(n12444) );
  NAND2_X1 U11334 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10253) );
  AOI22_X1 U11335 ( .A1(n12038), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12392), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11777) );
  NAND2_X1 U11336 ( .A1(n18539), .A2(n11364), .ZN(n11367) );
  NOR2_X1 U11337 ( .A1(n10439), .A2(n9819), .ZN(n9818) );
  NAND2_X1 U11338 ( .A1(n11793), .A2(n11792), .ZN(n16506) );
  AND2_X1 U11339 ( .A1(n10417), .A2(n10416), .ZN(n10427) );
  AND2_X1 U11340 ( .A1(n10440), .A2(n9718), .ZN(n9819) );
  NAND2_X1 U11341 ( .A1(n9871), .A2(n9805), .ZN(n12430) );
  AND2_X1 U11342 ( .A1(n10247), .A2(n10780), .ZN(n10246) );
  OR2_X1 U11343 ( .A1(n9618), .A2(n11800), .ZN(n11803) );
  NAND2_X1 U11344 ( .A1(n9806), .A2(n12341), .ZN(n12433) );
  AND2_X1 U11345 ( .A1(n12442), .A2(n12447), .ZN(n10172) );
  AND2_X1 U11346 ( .A1(n10889), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10890) );
  MUX2_X1 U11347 ( .A(n20034), .B(n12068), .S(n20318), .Z(n13850) );
  NAND2_X1 U11348 ( .A1(n11771), .A2(n12311), .ZN(n11904) );
  AOI21_X1 U11349 ( .B1(n10440), .B2(n10411), .A(n10410), .ZN(n10417) );
  CLKBUF_X1 U11350 ( .A(n12304), .Z(n15430) );
  INV_X1 U11351 ( .A(n11790), .ZN(n11793) );
  INV_X4 U11352 ( .A(n18031), .ZN(n18910) );
  AND2_X1 U11353 ( .A1(n11770), .A2(n12024), .ZN(n11771) );
  AND2_X1 U11354 ( .A1(n10498), .A2(n14266), .ZN(n14130) );
  OAI21_X1 U11355 ( .B1(n12280), .B2(n20232), .A(n12053), .ZN(n12069) );
  NAND2_X1 U11356 ( .A1(n11763), .A2(n12045), .ZN(n9784) );
  AND2_X1 U11357 ( .A1(n11944), .A2(n12024), .ZN(n12312) );
  AND2_X1 U11358 ( .A1(n12045), .A2(n11763), .ZN(n11775) );
  AND2_X1 U11359 ( .A1(n12345), .A2(n12344), .ZN(n12438) );
  AND2_X1 U11360 ( .A1(n13824), .A2(n14305), .ZN(n13652) );
  INV_X1 U11361 ( .A(n13824), .ZN(n14770) );
  OR2_X1 U11362 ( .A1(n11360), .A2(n11359), .ZN(n16667) );
  NAND2_X2 U11363 ( .A1(n9665), .A2(n9914), .ZN(n13923) );
  NOR2_X1 U11364 ( .A1(n10554), .A2(n10692), .ZN(n10482) );
  AND2_X2 U11365 ( .A1(n11786), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11770) );
  INV_X1 U11366 ( .A(n12523), .ZN(n9807) );
  AND2_X1 U11367 ( .A1(n9926), .A2(n14116), .ZN(n15378) );
  INV_X2 U11368 ( .A(n11951), .ZN(n15806) );
  AND2_X1 U11369 ( .A1(n11716), .A2(n11759), .ZN(n12024) );
  AND4_X1 U11370 ( .A1(n11746), .A2(n11753), .A3(n11759), .A4(n16546), .ZN(
        n11763) );
  AND2_X1 U11371 ( .A1(n11951), .A2(n16535), .ZN(n11944) );
  AND3_X1 U11372 ( .A1(n12365), .A2(n16535), .A3(n13646), .ZN(n11788) );
  INV_X1 U11373 ( .A(n11677), .ZN(n11744) );
  CLKBUF_X1 U11374 ( .A(n10436), .Z(n14101) );
  AND2_X2 U11375 ( .A1(n10476), .A2(n10479), .ZN(n10757) );
  AND2_X1 U11376 ( .A1(n11752), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15425) );
  NOR2_X2 U11377 ( .A1(n11418), .A2(n11417), .ZN(n18873) );
  OR2_X1 U11378 ( .A1(n11981), .A2(n11980), .ZN(n13732) );
  INV_X1 U11379 ( .A(n11753), .ZN(n11962) );
  NAND2_X2 U11380 ( .A1(n11713), .A2(n11712), .ZN(n16546) );
  OR2_X1 U11381 ( .A1(n10460), .A2(n10459), .ZN(n10684) );
  INV_X1 U11382 ( .A(n12065), .ZN(n12365) );
  NAND2_X2 U11383 ( .A1(n9676), .A2(n9607), .ZN(n20611) );
  OR2_X1 U11385 ( .A1(n10473), .A2(n10472), .ZN(n10609) );
  NAND2_X1 U11386 ( .A1(n11688), .A2(n11687), .ZN(n11759) );
  AND4_X2 U11387 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10432) );
  NAND2_X1 U11388 ( .A1(n11674), .A2(n13875), .ZN(n11675) );
  NOR2_X1 U11389 ( .A1(n18394), .A2(n10137), .ZN(n10136) );
  NAND2_X1 U11390 ( .A1(n11616), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18394) );
  INV_X2 U11391 ( .A(n17891), .ZN(n9625) );
  AND4_X1 U11392 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10386) );
  AND4_X1 U11393 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10385) );
  AND4_X1 U11394 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10384) );
  AND2_X2 U11395 ( .A1(n12005), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13067) );
  NAND2_X2 U11396 ( .A1(n13559), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21268) );
  INV_X2 U11397 ( .A(n19379), .ZN(n9610) );
  CLKBUF_X2 U11398 ( .A(n10483), .Z(n10531) );
  NAND2_X2 U11399 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20347), .ZN(n20281) );
  NAND2_X2 U11400 ( .A1(n20347), .A2(n20231), .ZN(n20284) );
  BUF_X2 U11401 ( .A(n10461), .Z(n13410) );
  NAND2_X2 U11402 ( .A1(n19434), .A2(n19375), .ZN(n19421) );
  AND3_X1 U11403 ( .A1(n11690), .A2(n11689), .A3(n13875), .ZN(n11694) );
  AND3_X1 U11405 ( .A1(n11696), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11695), .ZN(n11699) );
  AND2_X1 U11406 ( .A1(n16902), .A2(n11261), .ZN(n11252) );
  NAND2_X1 U11407 ( .A1(n16902), .A2(n11260), .ZN(n16942) );
  NAND2_X2 U11409 ( .A1(n11259), .A2(n16902), .ZN(n17891) );
  AND2_X2 U11410 ( .A1(n13082), .A2(n13875), .ZN(n13866) );
  NAND2_X1 U11411 ( .A1(n16904), .A2(n11260), .ZN(n17818) );
  CLKBUF_X1 U11412 ( .A(n13082), .Z(n16574) );
  BUF_X2 U11413 ( .A(n10530), .Z(n9613) );
  INV_X2 U11414 ( .A(n11691), .ZN(n11723) );
  INV_X2 U11415 ( .A(n17244), .ZN(n17246) );
  AND2_X2 U11416 ( .A1(n9989), .A2(n15365), .ZN(n10483) );
  AND2_X2 U11417 ( .A1(n11909), .A2(n13875), .ZN(n9673) );
  AND2_X2 U11418 ( .A1(n17046), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16930) );
  AND2_X2 U11419 ( .A1(n16900), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16911) );
  AND2_X1 U11420 ( .A1(n9896), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16904) );
  AND2_X1 U11421 ( .A1(n11253), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11258) );
  INV_X2 U11422 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10317) );
  NOR2_X1 U11423 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10324) );
  AND2_X1 U11424 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11643) );
  AND2_X1 U11425 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11260) );
  AND2_X1 U11426 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17046) );
  INV_X1 U11427 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16909) );
  NOR2_X1 U11428 ( .A1(n9839), .A2(n9961), .ZN(n9838) );
  OR2_X2 U11429 ( .A1(n9961), .A2(n12426), .ZN(n12630) );
  INV_X1 U11430 ( .A(n10668), .ZN(n9887) );
  INV_X1 U11431 ( .A(n12631), .ZN(n16241) );
  AND2_X1 U11433 ( .A1(n11951), .A2(n11754), .ZN(n12308) );
  NOR2_X2 U11434 ( .A1(n10814), .A2(n20393), .ZN(n10821) );
  AND2_X1 U11435 ( .A1(n9989), .A2(n15365), .ZN(n9616) );
  INV_X2 U11436 ( .A(n10414), .ZN(n10445) );
  AND2_X2 U11438 ( .A1(n15361), .A2(n14273), .ZN(n10447) );
  OR2_X1 U11439 ( .A1(n10408), .A2(n10407), .ZN(n9617) );
  AND2_X2 U11440 ( .A1(n12428), .A2(n12628), .ZN(n16249) );
  INV_X2 U11441 ( .A(n12042), .ZN(n11951) );
  NAND2_X1 U11442 ( .A1(n17299), .A2(n17508), .ZN(n17291) );
  NAND2_X2 U11443 ( .A1(n10012), .A2(n9965), .ZN(n12628) );
  NAND2_X1 U11444 ( .A1(n9965), .A2(n9659), .ZN(n9961) );
  NOR2_X1 U11445 ( .A1(n10317), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10323) );
  OAI21_X2 U11446 ( .B1(n14162), .B2(n14068), .A(n10607), .ZN(n14079) );
  NAND2_X1 U11447 ( .A1(n11771), .A2(n12311), .ZN(n9618) );
  NAND2_X1 U11448 ( .A1(n11771), .A2(n12311), .ZN(n9619) );
  AND2_X1 U11449 ( .A1(n13861), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9620) );
  NAND2_X1 U11450 ( .A1(n10570), .A2(n10631), .ZN(n10640) );
  OAI21_X1 U11451 ( .B1(n9886), .B2(n10775), .A(n10510), .ZN(n10603) );
  AND2_X2 U11452 ( .A1(n10302), .A2(n13361), .ZN(n13347) );
  OR2_X1 U11453 ( .A1(n13376), .A2(n13361), .ZN(n13338) );
  NAND2_X2 U11454 ( .A1(n11776), .A2(n12291), .ZN(n12038) );
  AND2_X2 U11455 ( .A1(n12831), .A2(n12028), .ZN(n12291) );
  NOR2_X2 U11456 ( .A1(n14494), .A2(n14495), .ZN(n14479) );
  NAND2_X2 U11457 ( .A1(n15001), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10712) );
  OAI21_X2 U11458 ( .B1(n10062), .B2(n9990), .A(n9927), .ZN(n15001) );
  NOR2_X2 U11460 ( .A1(n14398), .A2(n9717), .ZN(n14329) );
  OR2_X2 U11461 ( .A1(n11432), .A2(n11431), .ZN(n19471) );
  NAND2_X2 U11462 ( .A1(n10622), .A2(n10689), .ZN(n10509) );
  AND2_X2 U11463 ( .A1(n9817), .A2(n9816), .ZN(n10503) );
  AOI21_X2 U11464 ( .B1(n10517), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10501), .ZN(n10502) );
  XNOR2_X1 U11465 ( .A(n10512), .B(n10502), .ZN(n20722) );
  OR2_X1 U11466 ( .A1(n17257), .A2(n19471), .ZN(n18484) );
  XNOR2_X1 U11467 ( .A(n10775), .B(n9886), .ZN(n20691) );
  AOI21_X2 U11468 ( .B1(n11521), .B2(n13919), .A(n11542), .ZN(n16914) );
  NAND2_X1 U11469 ( .A1(n12705), .A2(n12704), .ZN(n9804) );
  NOR2_X1 U11470 ( .A1(n10597), .A2(n10414), .ZN(n10367) );
  NAND3_X1 U11471 ( .A1(n11694), .A2(n11693), .A3(n11692), .ZN(n11701) );
  INV_X1 U11472 ( .A(n9868), .ZN(n9867) );
  AND2_X1 U11473 ( .A1(n9940), .A2(n13828), .ZN(n14134) );
  OR2_X1 U11474 ( .A1(n14106), .A2(n14116), .ZN(n9943) );
  OR2_X1 U11475 ( .A1(n15621), .A2(n15622), .ZN(n9628) );
  AOI21_X1 U11476 ( .B1(n12037), .B2(n12036), .A(n17160), .ZN(n12651) );
  NOR2_X1 U11477 ( .A1(n12673), .A2(n12035), .ZN(n12036) );
  OR2_X1 U11478 ( .A1(n10725), .A2(n9929), .ZN(n10718) );
  INV_X1 U11479 ( .A(n10721), .ZN(n9929) );
  AND2_X1 U11480 ( .A1(n10724), .A2(n10723), .ZN(n10728) );
  NAND4_X1 U11481 ( .A1(n9792), .A2(n9791), .A3(n9790), .A4(n9789), .ZN(n11804) );
  NAND2_X1 U11482 ( .A1(n11762), .A2(n9648), .ZN(n9792) );
  NAND2_X1 U11483 ( .A1(n9889), .A2(n9888), .ZN(n10668) );
  INV_X1 U11484 ( .A(n10595), .ZN(n9888) );
  NOR2_X1 U11485 ( .A1(n10554), .A2(n10684), .ZN(n10477) );
  AND2_X2 U11486 ( .A1(n10314), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10100) );
  INV_X1 U11487 ( .A(n12573), .ZN(n10169) );
  NAND2_X1 U11488 ( .A1(n11757), .A2(n11756), .ZN(n11807) );
  AND2_X1 U11489 ( .A1(n12296), .A2(n11755), .ZN(n11756) );
  NAND2_X1 U11490 ( .A1(n11784), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10254) );
  NAND2_X1 U11491 ( .A1(n12401), .A2(n11783), .ZN(n9952) );
  INV_X1 U11492 ( .A(n13431), .ZN(n13425) );
  INV_X1 U11493 ( .A(n10783), .ZN(n11233) );
  INV_X1 U11494 ( .A(n14305), .ZN(n13360) );
  INV_X1 U11495 ( .A(n14006), .ZN(n13286) );
  AND2_X1 U11496 ( .A1(n10476), .A2(n10431), .ZN(n10302) );
  INV_X1 U11497 ( .A(n10428), .ZN(n10244) );
  OAI21_X1 U11498 ( .B1(n10431), .B2(n13385), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10428) );
  OR2_X1 U11499 ( .A1(n11995), .A2(n11994), .ZN(n10161) );
  NAND2_X1 U11500 ( .A1(n12383), .A2(n10169), .ZN(n10166) );
  NAND2_X1 U11501 ( .A1(n10169), .A2(n10168), .ZN(n10167) );
  INV_X1 U11502 ( .A(n12364), .ZN(n10168) );
  AND2_X2 U11503 ( .A1(n12042), .A2(n11752), .ZN(n11786) );
  NAND2_X1 U11504 ( .A1(n16297), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14372) );
  NAND2_X1 U11505 ( .A1(n10195), .A2(n10197), .ZN(n10193) );
  NOR2_X2 U11506 ( .A1(n15635), .A2(n10234), .ZN(n13252) );
  NAND2_X1 U11507 ( .A1(n12262), .A2(n10235), .ZN(n10234) );
  NOR2_X1 U11508 ( .A1(n10236), .A2(n13253), .ZN(n10235) );
  NOR2_X1 U11509 ( .A1(n10284), .A2(n12731), .ZN(n9844) );
  INV_X1 U11510 ( .A(n16090), .ZN(n10286) );
  AND4_X1 U11511 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12144) );
  AND4_X1 U11512 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12142) );
  AND4_X1 U11513 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12141) );
  OAI21_X1 U11514 ( .B1(n20342), .B2(n12650), .A(n12020), .ZN(n12673) );
  NOR2_X2 U11515 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11261) );
  OR2_X1 U11516 ( .A1(n11373), .A2(n18114), .ZN(n11380) );
  NOR2_X1 U11517 ( .A1(n13917), .A2(n19299), .ZN(n16883) );
  INV_X2 U11518 ( .A(n11233), .ZN(n14311) );
  NAND2_X1 U11519 ( .A1(n13379), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13384) );
  INV_X1 U11520 ( .A(n13378), .ZN(n13379) );
  AND2_X1 U11521 ( .A1(n14479), .A2(n10106), .ZN(n14313) );
  NOR2_X1 U11522 ( .A1(n10109), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U11523 ( .A1(n10114), .A2(n10110), .ZN(n10109) );
  INV_X1 U11524 ( .A(n10111), .ZN(n10110) );
  NOR2_X1 U11525 ( .A1(n14194), .A2(n14054), .ZN(n10101) );
  INV_X1 U11526 ( .A(n14055), .ZN(n10102) );
  INV_X1 U11527 ( .A(n14955), .ZN(n10714) );
  NAND2_X1 U11528 ( .A1(n10065), .A2(n14962), .ZN(n14955) );
  AND2_X1 U11529 ( .A1(n20547), .A2(n14349), .ZN(n15257) );
  OR2_X1 U11530 ( .A1(n20546), .A2(n20573), .ZN(n15293) );
  NAND2_X1 U11531 ( .A1(n20582), .A2(n20572), .ZN(n20546) );
  INV_X1 U11532 ( .A(n20611), .ZN(n9926) );
  OR2_X1 U11533 ( .A1(n10767), .A2(n10766), .ZN(n10770) );
  AND2_X1 U11534 ( .A1(n13372), .A2(n10765), .ZN(n10766) );
  AND2_X1 U11535 ( .A1(n16591), .A2(n16626), .ZN(n12832) );
  NAND2_X1 U11536 ( .A1(n12382), .A2(n15828), .ZN(n12386) );
  NAND2_X1 U11537 ( .A1(n15453), .A2(n12660), .ZN(n12694) );
  AND2_X2 U11538 ( .A1(n15506), .A2(n10231), .ZN(n15453) );
  AND2_X1 U11539 ( .A1(n9658), .A2(n14416), .ZN(n10231) );
  AND2_X1 U11540 ( .A1(n15453), .A2(n15452), .ZN(n15455) );
  AND2_X1 U11541 ( .A1(n19586), .A2(n13231), .ZN(n13741) );
  AND2_X1 U11542 ( .A1(n19586), .A2(n12045), .ZN(n15985) );
  INV_X1 U11543 ( .A(n10219), .ZN(n10217) );
  NOR3_X1 U11544 ( .A1(n12699), .A2(n12336), .A3(n12649), .ZN(n10026) );
  NAND2_X1 U11545 ( .A1(n9711), .A2(n9770), .ZN(n12711) );
  INV_X1 U11546 ( .A(n16020), .ZN(n9770) );
  NAND2_X1 U11547 ( .A1(n11889), .A2(n10212), .ZN(n10211) );
  AND2_X1 U11548 ( .A1(n14366), .A2(n14365), .ZN(n11889) );
  NAND2_X1 U11549 ( .A1(n9878), .A2(n10255), .ZN(n10087) );
  NAND2_X1 U11550 ( .A1(n10255), .A2(n10257), .ZN(n9785) );
  INV_X1 U11551 ( .A(n10260), .ZN(n10257) );
  NAND2_X1 U11552 ( .A1(n9970), .A2(n9972), .ZN(n14289) );
  INV_X1 U11553 ( .A(n16365), .ZN(n9875) );
  NAND2_X1 U11554 ( .A1(n13769), .A2(n13770), .ZN(n13773) );
  NAND2_X1 U11555 ( .A1(n11966), .A2(n11965), .ZN(n16592) );
  NAND2_X1 U11556 ( .A1(n20323), .A2(n19782), .ZN(n20072) );
  NAND2_X1 U11557 ( .A1(n20323), .A2(n20308), .ZN(n20156) );
  OR2_X1 U11558 ( .A1(n11332), .A2(n11331), .ZN(n11605) );
  INV_X1 U11559 ( .A(n18104), .ZN(n16771) );
  INV_X1 U11560 ( .A(n14932), .ZN(n14935) );
  INV_X1 U11561 ( .A(n19547), .ZN(n19529) );
  INV_X1 U11562 ( .A(n16085), .ZN(n10055) );
  INV_X1 U11563 ( .A(n19642), .ZN(n16222) );
  INV_X1 U11564 ( .A(n9975), .ZN(n9974) );
  OAI211_X1 U11565 ( .C1(n14382), .C2(n17133), .A(n12698), .B(n9976), .ZN(
        n9975) );
  NAND2_X1 U11566 ( .A1(n13248), .A2(n19665), .ZN(n9976) );
  AND2_X1 U11567 ( .A1(n16087), .A2(n19669), .ZN(n10086) );
  AND2_X1 U11568 ( .A1(n13824), .A2(n10721), .ZN(n10737) );
  INV_X1 U11569 ( .A(n10757), .ZN(n10754) );
  NAND2_X1 U11570 ( .A1(n9619), .A2(n11785), .ZN(n11787) );
  NAND2_X1 U11571 ( .A1(n16517), .A2(n13862), .ZN(n11691) );
  INV_X1 U11572 ( .A(n14717), .ZN(n10117) );
  NOR2_X1 U11573 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  INV_X1 U11574 ( .A(n10303), .ZN(n10120) );
  AND2_X1 U11575 ( .A1(n10665), .A2(n10664), .ZN(n10667) );
  INV_X1 U11576 ( .A(n10639), .ZN(n10248) );
  AND2_X1 U11577 ( .A1(n10435), .A2(n10445), .ZN(n10292) );
  OR2_X1 U11578 ( .A1(n10493), .A2(n10492), .ZN(n10610) );
  NAND2_X1 U11579 ( .A1(n10418), .A2(n10414), .ZN(n10420) );
  NAND2_X1 U11580 ( .A1(n10500), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U11581 ( .A1(n10432), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10553) );
  OR2_X1 U11582 ( .A1(n10731), .A2(n10730), .ZN(n9939) );
  NAND2_X1 U11583 ( .A1(n9934), .A2(n10761), .ZN(n9933) );
  INV_X1 U11584 ( .A(n9936), .ZN(n9934) );
  AOI21_X1 U11585 ( .B1(n9685), .B2(n10739), .A(n9937), .ZN(n9936) );
  NOR2_X1 U11586 ( .A1(n10764), .A2(n10752), .ZN(n9937) );
  INV_X1 U11587 ( .A(n10760), .ZN(n9935) );
  NAND2_X1 U11588 ( .A1(n11753), .A2(n16558), .ZN(n11677) );
  INV_X1 U11589 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11785) );
  AOI21_X1 U11590 ( .B1(n13188), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(n9764), .ZN(n13190) );
  INV_X1 U11591 ( .A(n12641), .ZN(n9800) );
  AND2_X1 U11592 ( .A1(n12610), .A2(n12354), .ZN(n9959) );
  XNOR2_X1 U11593 ( .A(n12641), .B(n12610), .ZN(n12632) );
  INV_X1 U11594 ( .A(n9784), .ZN(n12023) );
  NOR2_X1 U11595 ( .A1(n11920), .A2(n11919), .ZN(n12421) );
  INV_X1 U11596 ( .A(n18488), .ZN(n10150) );
  AND2_X1 U11597 ( .A1(n11592), .A2(n18126), .ZN(n11590) );
  INV_X1 U11598 ( .A(n10792), .ZN(n10105) );
  AND2_X1 U11599 ( .A1(n14115), .A2(n10774), .ZN(n13718) );
  NAND2_X1 U11600 ( .A1(n9824), .A2(n9822), .ZN(n14953) );
  NAND2_X1 U11601 ( .A1(n9823), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9822) );
  INV_X1 U11602 ( .A(n15183), .ZN(n9823) );
  AND2_X1 U11603 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  INV_X1 U11604 ( .A(n14597), .ZN(n10128) );
  AND2_X1 U11605 ( .A1(n10130), .A2(n14632), .ZN(n10129) );
  AND2_X1 U11606 ( .A1(n14234), .A2(n10133), .ZN(n10132) );
  INV_X1 U11607 ( .A(n14735), .ZN(n10133) );
  AND2_X1 U11608 ( .A1(n10697), .A2(n9672), .ZN(n9811) );
  OR2_X1 U11609 ( .A1(n10567), .A2(n10566), .ZN(n10643) );
  NAND2_X1 U11610 ( .A1(n10445), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U11611 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10364) );
  OR2_X2 U11612 ( .A1(n10330), .A2(n10329), .ZN(n10597) );
  XNOR2_X1 U11613 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11983) );
  OAI21_X1 U11614 ( .B1(n12609), .B2(n12421), .A(n9872), .ZN(n12346) );
  NAND2_X1 U11615 ( .A1(n12609), .A2(n12011), .ZN(n9872) );
  AOI21_X1 U11616 ( .B1(n19559), .B2(n10182), .A(n10181), .ZN(n10180) );
  INV_X1 U11617 ( .A(n15479), .ZN(n10182) );
  INV_X1 U11618 ( .A(n15471), .ZN(n10181) );
  NAND2_X1 U11619 ( .A1(n12708), .A2(n12492), .ZN(n12377) );
  INV_X1 U11620 ( .A(n12520), .ZN(n12546) );
  CLKBUF_X1 U11621 ( .A(n11908), .Z(n13188) );
  CLKBUF_X1 U11622 ( .A(n13083), .Z(n13206) );
  INV_X1 U11623 ( .A(n14371), .ZN(n10232) );
  NAND2_X1 U11624 ( .A1(n10204), .A2(n10202), .ZN(n14154) );
  NOR2_X1 U11625 ( .A1(n9724), .A2(n10203), .ZN(n10202) );
  INV_X1 U11626 ( .A(n14155), .ZN(n10203) );
  NOR2_X1 U11627 ( .A1(n12115), .A2(n12114), .ZN(n12478) );
  INV_X1 U11628 ( .A(n12065), .ZN(n11747) );
  INV_X1 U11629 ( .A(n14044), .ZN(n10223) );
  NAND2_X1 U11630 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U11631 ( .A1(n11807), .A2(n11770), .ZN(n10010) );
  INV_X1 U11632 ( .A(n15432), .ZN(n12392) );
  NOR2_X1 U11633 ( .A1(n10213), .A2(n10215), .ZN(n10212) );
  AND2_X1 U11634 ( .A1(n15519), .A2(n12644), .ZN(n12582) );
  OR2_X1 U11635 ( .A1(n15546), .A2(n12354), .ZN(n12578) );
  NAND2_X1 U11636 ( .A1(n10237), .A2(n14295), .ZN(n10236) );
  INV_X1 U11637 ( .A(n14156), .ZN(n10237) );
  NAND2_X1 U11638 ( .A1(n9855), .A2(n12553), .ZN(n9856) );
  NOR2_X1 U11639 ( .A1(n9857), .A2(n12354), .ZN(n9855) );
  NAND2_X1 U11640 ( .A1(n10255), .A2(n9799), .ZN(n9798) );
  NAND2_X1 U11641 ( .A1(n16241), .A2(n10066), .ZN(n10014) );
  BUF_X1 U11642 ( .A(n12632), .Z(n12638) );
  OAI211_X1 U11643 ( .C1(n9619), .C2(n12347), .A(n11816), .B(n11815), .ZN(
        n12393) );
  AND2_X1 U11644 ( .A1(n12304), .A2(n11791), .ZN(n11792) );
  AND2_X1 U11645 ( .A1(n12045), .A2(n12979), .ZN(n11760) );
  AND2_X2 U11646 ( .A1(n12416), .A2(n12414), .ZN(n19934) );
  AND2_X1 U11647 ( .A1(n9702), .A2(n12402), .ZN(n12406) );
  INV_X1 U11648 ( .A(n9952), .ZN(n9951) );
  OR2_X1 U11649 ( .A1(n11957), .A2(n11958), .ZN(n12009) );
  AND4_X1 U11650 ( .A1(n11293), .A2(n11292), .A3(n11291), .A4(n11290), .ZN(
        n11297) );
  NOR2_X1 U11651 ( .A1(n18880), .A2(n11533), .ZN(n11523) );
  INV_X1 U11652 ( .A(n10142), .ZN(n10138) );
  NAND2_X1 U11653 ( .A1(n10305), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10142) );
  NAND2_X1 U11654 ( .A1(n11289), .A2(n18126), .ZN(n11369) );
  OAI21_X1 U11655 ( .B1(n13923), .B2(n16663), .A(n11593), .ZN(n11362) );
  NAND2_X1 U11656 ( .A1(n16706), .A2(n16813), .ZN(n16671) );
  OAI21_X1 U11657 ( .B1(n11536), .B2(n18910), .A(n18889), .ZN(n11537) );
  NOR2_X1 U11658 ( .A1(n11541), .A2(n13799), .ZN(n13919) );
  AND2_X1 U11659 ( .A1(n9667), .A2(n13375), .ZN(n20399) );
  AND2_X1 U11660 ( .A1(n21294), .A2(n13374), .ZN(n13375) );
  AND2_X1 U11661 ( .A1(n14675), .A2(n14687), .ZN(n13310) );
  AND2_X1 U11662 ( .A1(n13285), .A2(n13284), .ZN(n14006) );
  NAND2_X1 U11663 ( .A1(n13838), .A2(n10795), .ZN(n13885) );
  INV_X1 U11664 ( .A(n10858), .ZN(n14310) );
  NAND2_X1 U11665 ( .A1(n13432), .A2(n10112), .ZN(n10111) );
  INV_X1 U11666 ( .A(n14468), .ZN(n10112) );
  INV_X1 U11667 ( .A(n13433), .ZN(n10114) );
  OR2_X1 U11668 ( .A1(n14969), .A2(n13431), .ZN(n11180) );
  NAND2_X1 U11669 ( .A1(n10986), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10970) );
  INV_X1 U11670 ( .A(n10888), .ZN(n10889) );
  INV_X1 U11671 ( .A(n10826), .ZN(n10827) );
  INV_X1 U11672 ( .A(n14199), .ZN(n10832) );
  OR2_X1 U11673 ( .A1(n14173), .A2(n20348), .ZN(n13792) );
  NAND2_X1 U11674 ( .A1(n14993), .A2(n14940), .ZN(n14943) );
  OR2_X1 U11675 ( .A1(n14352), .A2(n14399), .ZN(n9949) );
  OAI21_X1 U11676 ( .B1(n14974), .B2(n10711), .A(n15049), .ZN(n14962) );
  NAND2_X1 U11677 ( .A1(n10712), .A2(n10249), .ZN(n14974) );
  AOI21_X1 U11678 ( .B1(n15010), .B2(n15049), .A(n10250), .ZN(n10249) );
  INV_X1 U11679 ( .A(n10251), .ZN(n10250) );
  AOI21_X1 U11680 ( .B1(n15049), .B2(n10710), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10251) );
  NAND2_X1 U11681 ( .A1(n10712), .A2(n15002), .ZN(n14993) );
  NAND2_X1 U11682 ( .A1(n15076), .A2(n15057), .ZN(n15068) );
  AND2_X1 U11683 ( .A1(n13303), .A2(n13302), .ZN(n14703) );
  NAND2_X1 U11684 ( .A1(n10123), .A2(n14203), .ZN(n10122) );
  NAND2_X1 U11685 ( .A1(n10125), .A2(n13286), .ZN(n17116) );
  INV_X1 U11686 ( .A(n20558), .ZN(n20547) );
  NAND2_X1 U11687 ( .A1(n10430), .A2(n10429), .ZN(n9816) );
  OAI211_X1 U11688 ( .C1(n10616), .C2(n10476), .A(n10481), .B(n10480), .ZN(
        n10780) );
  NAND2_X1 U11689 ( .A1(n10516), .A2(n20658), .ZN(n14171) );
  INV_X1 U11690 ( .A(n20653), .ZN(n20763) );
  OR3_X1 U11691 ( .A1(n13724), .A2(n13827), .A3(n13723), .ZN(n17063) );
  INV_X1 U11692 ( .A(n20694), .ZN(n20967) );
  NOR2_X1 U11693 ( .A1(n15413), .A2(n15408), .ZN(n20994) );
  INV_X1 U11694 ( .A(n21089), .ZN(n21094) );
  NOR2_X1 U11695 ( .A1(n20763), .A2(n20964), .ZN(n21138) );
  INV_X1 U11697 ( .A(n21184), .ZN(n21186) );
  NAND2_X1 U11698 ( .A1(n11959), .A2(n11958), .ZN(n12015) );
  OAI21_X1 U11699 ( .B1(n10161), .B2(n12609), .A(n11997), .ZN(n12340) );
  NAND2_X1 U11700 ( .A1(n12348), .A2(n12346), .ZN(n9982) );
  INV_X1 U11701 ( .A(n15439), .ZN(n15461) );
  NAND2_X1 U11702 ( .A1(n15482), .A2(n15485), .ZN(n12708) );
  OR2_X1 U11703 ( .A1(n10167), .A2(n10165), .ZN(n10164) );
  NAND2_X1 U11704 ( .A1(n10163), .A2(n12579), .ZN(n10162) );
  INV_X1 U11705 ( .A(n12579), .ZN(n10165) );
  AND3_X1 U11706 ( .A1(n12103), .A2(n12102), .A3(n12101), .ZN(n13457) );
  NOR2_X1 U11707 ( .A1(n12956), .A2(n12979), .ZN(n13846) );
  INV_X1 U11708 ( .A(n15637), .ZN(n12256) );
  INV_X1 U11709 ( .A(n14145), .ZN(n12257) );
  AND3_X1 U11710 ( .A1(n12187), .A2(n12186), .A3(n12185), .ZN(n13890) );
  AND2_X1 U11711 ( .A1(n12744), .A2(n12745), .ZN(n15541) );
  AND2_X1 U11712 ( .A1(n12788), .A2(n9750), .ZN(n12796) );
  INV_X1 U11713 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16152) );
  AOI21_X1 U11714 ( .B1(n10270), .B2(n10272), .A(n9740), .ZN(n10267) );
  OAI211_X1 U11715 ( .C1(n12628), .C2(n10046), .A(n10045), .B(n10270), .ZN(
        n10268) );
  AND2_X1 U11716 ( .A1(n12673), .A2(n12672), .ZN(n12689) );
  OAI21_X1 U11717 ( .B1(n14462), .B2(n19648), .A(n10028), .ZN(n10027) );
  INV_X1 U11718 ( .A(n12945), .ZN(n10028) );
  NOR2_X1 U11719 ( .A1(n16044), .A2(n10263), .ZN(n12674) );
  NOR2_X1 U11720 ( .A1(n14372), .A2(n10004), .ZN(n16272) );
  AND2_X1 U11721 ( .A1(n9660), .A2(n12334), .ZN(n10002) );
  AND2_X1 U11722 ( .A1(n9660), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10003) );
  NAND2_X1 U11723 ( .A1(n12501), .A2(n12507), .ZN(n10196) );
  NAND2_X1 U11724 ( .A1(n10096), .A2(n10099), .ZN(n10095) );
  OR2_X1 U11725 ( .A1(n14293), .A2(n14294), .ZN(n14291) );
  NAND2_X1 U11726 ( .A1(n16158), .A2(n12490), .ZN(n12503) );
  NOR2_X1 U11727 ( .A1(n17135), .A2(n12322), .ZN(n16411) );
  AND2_X1 U11728 ( .A1(n12506), .A2(n12505), .ZN(n16175) );
  NAND2_X1 U11729 ( .A1(n10275), .A2(n16476), .ZN(n10274) );
  INV_X1 U11730 ( .A(n16245), .ZN(n10275) );
  NAND2_X1 U11731 ( .A1(n16245), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10273) );
  AOI21_X1 U11732 ( .B1(n19683), .B2(n19682), .A(n12320), .ZN(n9985) );
  OR2_X1 U11733 ( .A1(n10047), .A2(n10044), .ZN(n10043) );
  INV_X1 U11734 ( .A(n12628), .ZN(n10044) );
  INV_X1 U11735 ( .A(n15740), .ZN(n12085) );
  NAND2_X1 U11736 ( .A1(n12960), .A2(n12959), .ZN(n13644) );
  AND2_X1 U11737 ( .A1(n12317), .A2(n12316), .ZN(n16571) );
  NAND2_X1 U11738 ( .A1(n16526), .A2(n20095), .ZN(n16531) );
  OR3_X1 U11739 ( .A1(n20204), .A2(n19711), .A3(n20313), .ZN(n16526) );
  NAND2_X1 U11740 ( .A1(n19692), .A2(n20330), .ZN(n19840) );
  NAND2_X1 U11741 ( .A1(n19692), .A2(n19691), .ZN(n19881) );
  NAND2_X1 U11742 ( .A1(n20309), .A2(n20330), .ZN(n20094) );
  OR2_X1 U11743 ( .A1(n19692), .A2(n20330), .ZN(n20073) );
  INV_X1 U11744 ( .A(n20101), .ZN(n20152) );
  AND2_X1 U11745 ( .A1(n11576), .A2(n11575), .ZN(n19294) );
  OR2_X1 U11746 ( .A1(n11568), .A2(n11567), .ZN(n19299) );
  INV_X1 U11747 ( .A(n11520), .ZN(n16886) );
  AND2_X1 U11748 ( .A1(n9646), .A2(n10145), .ZN(n10144) );
  INV_X1 U11749 ( .A(n18248), .ZN(n10145) );
  INV_X1 U11750 ( .A(n18429), .ZN(n11616) );
  NAND2_X1 U11751 ( .A1(n10174), .A2(n18776), .ZN(n18368) );
  INV_X1 U11752 ( .A(n11394), .ZN(n10174) );
  XNOR2_X1 U11753 ( .A(n13923), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18550) );
  NAND2_X1 U11754 ( .A1(n10308), .A2(n18550), .ZN(n18549) );
  NAND2_X1 U11755 ( .A1(n16671), .A2(n16673), .ZN(n16694) );
  NAND2_X1 U11756 ( .A1(n9686), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16796) );
  INV_X1 U11757 ( .A(n11380), .ZN(n11333) );
  NAND2_X1 U11758 ( .A1(n10160), .A2(n18299), .ZN(n16747) );
  NAND2_X1 U11759 ( .A1(n10156), .A2(n11396), .ZN(n10155) );
  INV_X1 U11760 ( .A(n18286), .ZN(n10156) );
  INV_X1 U11761 ( .A(n18343), .ZN(n10151) );
  INV_X1 U11762 ( .A(n11396), .ZN(n10157) );
  NAND2_X1 U11763 ( .A1(n18343), .A2(n18369), .ZN(n18299) );
  NAND2_X1 U11764 ( .A1(n9922), .A2(n9921), .ZN(n18343) );
  INV_X1 U11765 ( .A(n18342), .ZN(n9922) );
  AOI21_X1 U11766 ( .B1(n18660), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U11767 ( .A1(n16766), .A2(n11612), .ZN(n18373) );
  OR2_X1 U11768 ( .A1(n18497), .A2(n11604), .ZN(n9907) );
  NOR2_X1 U11769 ( .A1(n18114), .A2(n11589), .ZN(n18481) );
  NAND2_X1 U11770 ( .A1(n18501), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18500) );
  NOR2_X1 U11771 ( .A1(n18499), .A2(n18498), .ZN(n18497) );
  INV_X1 U11772 ( .A(n18528), .ZN(n9903) );
  NOR2_X1 U11773 ( .A1(n18538), .A2(n18537), .ZN(n18536) );
  INV_X1 U11774 ( .A(n20392), .ZN(n20433) );
  AOI22_X1 U11775 ( .A1(n13364), .A2(n13363), .B1(n13362), .B2(n13361), .ZN(
        n13366) );
  NOR2_X2 U11776 ( .A1(n14433), .A2(n14869), .ZN(n14912) );
  OR2_X1 U11777 ( .A1(n14433), .A2(n14430), .ZN(n14915) );
  AND2_X1 U11778 ( .A1(n13829), .A2(n13828), .ZN(n14932) );
  OR2_X1 U11779 ( .A1(n13827), .A2(n13826), .ZN(n13829) );
  NAND2_X1 U11780 ( .A1(n9945), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14400) );
  NAND2_X1 U11781 ( .A1(n9947), .A2(n9946), .ZN(n9945) );
  OR2_X1 U11782 ( .A1(n14401), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9944) );
  NAND2_X1 U11783 ( .A1(n9712), .A2(n9931), .ZN(n15213) );
  INV_X1 U11784 ( .A(n15237), .ZN(n9931) );
  AND2_X1 U11785 ( .A1(n14134), .A2(n14132), .ZN(n20544) );
  INV_X1 U11786 ( .A(n20416), .ZN(n20580) );
  NAND2_X1 U11787 ( .A1(n21246), .A2(n21041), .ZN(n21184) );
  CLKBUF_X1 U11788 ( .A(n14171), .Z(n14172) );
  NAND2_X1 U11789 ( .A1(n15408), .A2(n15407), .ZN(n20866) );
  INV_X1 U11790 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21041) );
  OR2_X1 U11791 ( .A1(n14462), .A2(n19551), .ZN(n12861) );
  OR2_X1 U11792 ( .A1(n12826), .A2(n19537), .ZN(n10184) );
  OR2_X1 U11793 ( .A1(n14382), .A2(n19555), .ZN(n12850) );
  NAND2_X1 U11794 ( .A1(n15441), .A2(n15772), .ZN(n15449) );
  OAI21_X1 U11795 ( .B1(n15461), .B2(n15440), .A(n19563), .ZN(n15441) );
  NAND2_X1 U11796 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  INV_X1 U11797 ( .A(n12552), .ZN(n9857) );
  INV_X1 U11798 ( .A(n12553), .ZN(n9854) );
  AND2_X1 U11799 ( .A1(n15434), .A2(n12839), .ZN(n19554) );
  AND2_X1 U11800 ( .A1(n12844), .A2(n16622), .ZN(n19547) );
  INV_X1 U11801 ( .A(n19513), .ZN(n19548) );
  NAND2_X1 U11802 ( .A1(n19559), .A2(n19563), .ZN(n15784) );
  NAND2_X1 U11803 ( .A1(n9681), .A2(n10216), .ZN(n14463) );
  OAI21_X1 U11804 ( .B1(n9662), .B2(n10218), .A(n11907), .ZN(n10216) );
  NAND2_X1 U11805 ( .A1(n12678), .A2(n12677), .ZN(n14382) );
  OR2_X1 U11806 ( .A1(n9662), .A2(n10218), .ZN(n12678) );
  OR2_X1 U11807 ( .A1(n12676), .A2(n12675), .ZN(n12677) );
  OR2_X1 U11808 ( .A1(n15455), .A2(n12659), .ZN(n12661) );
  OR2_X1 U11809 ( .A1(n15455), .A2(n15454), .ZN(n16275) );
  AND2_X1 U11810 ( .A1(n13741), .A2(n16533), .ZN(n15984) );
  AND2_X1 U11811 ( .A1(n13741), .A2(n13618), .ZN(n15983) );
  AND2_X1 U11812 ( .A1(n13228), .A2(n16626), .ZN(n19586) );
  INV_X1 U11813 ( .A(n20330), .ZN(n19691) );
  NAND2_X1 U11814 ( .A1(n19625), .A2(n15435), .ZN(n19592) );
  OR2_X1 U11815 ( .A1(n12676), .A2(n12666), .ZN(n15791) );
  AND2_X1 U11816 ( .A1(n9632), .A2(n14367), .ZN(n15812) );
  AOI21_X1 U11817 ( .B1(n12746), .B2(n14291), .A(n15541), .ZN(n15845) );
  OAI21_X1 U11818 ( .B1(n14260), .B2(n12741), .A(n16306), .ZN(n9971) );
  INV_X1 U11819 ( .A(n16264), .ZN(n16234) );
  NAND2_X1 U11820 ( .A1(n16237), .A2(n19633), .ZN(n16264) );
  AND2_X1 U11821 ( .A1(n16237), .A2(n12680), .ZN(n19642) );
  NOR2_X1 U11822 ( .A1(n12687), .A2(n10092), .ZN(n10091) );
  NAND2_X1 U11823 ( .A1(n10093), .A2(n12685), .ZN(n10092) );
  NAND2_X1 U11824 ( .A1(n10262), .A2(n10261), .ZN(n10264) );
  NOR2_X1 U11825 ( .A1(n10263), .A2(n12335), .ZN(n10261) );
  OAI211_X1 U11826 ( .C1(n12658), .C2(n9863), .A(n9859), .B(n9858), .ZN(n12702) );
  NAND2_X1 U11827 ( .A1(n12688), .A2(n12686), .ZN(n9863) );
  NAND2_X1 U11828 ( .A1(n12658), .A2(n9700), .ZN(n9858) );
  OAI21_X1 U11829 ( .B1(n10198), .B2(n9861), .A(n9860), .ZN(n9859) );
  NOR3_X1 U11830 ( .A1(n16270), .A2(n12335), .A3(n9737), .ZN(n12699) );
  XNOR2_X1 U11831 ( .A(n12674), .B(n12335), .ZN(n12701) );
  XNOR2_X1 U11832 ( .A(n9955), .B(n16022), .ZN(n16278) );
  INV_X1 U11833 ( .A(n12711), .ZN(n10007) );
  NAND2_X1 U11834 ( .A1(n12711), .A2(n16019), .ZN(n14414) );
  NAND2_X1 U11835 ( .A1(n10005), .A2(n14369), .ZN(n14379) );
  OAI21_X1 U11836 ( .B1(n10087), .B2(n10001), .A(n9999), .ZN(n10005) );
  INV_X1 U11837 ( .A(n10000), .ZN(n9999) );
  OAI21_X1 U11838 ( .B1(n10089), .B2(n10001), .A(n14374), .ZN(n10000) );
  NAND2_X1 U11839 ( .A1(n9852), .A2(n16044), .ZN(n16301) );
  NAND2_X1 U11840 ( .A1(n9846), .A2(n14286), .ZN(n12735) );
  OAI21_X1 U11841 ( .B1(n16089), .B2(n9843), .A(n9840), .ZN(n9846) );
  AOI22_X1 U11842 ( .A1(n14260), .A2(n9679), .B1(n12886), .B2(n9968), .ZN(
        n9966) );
  NAND2_X1 U11843 ( .A1(n19657), .A2(n9969), .ZN(n9968) );
  NAND2_X1 U11844 ( .A1(n12741), .A2(n16306), .ZN(n9969) );
  AOI21_X1 U11845 ( .B1(n9842), .B2(n10281), .A(n10280), .ZN(n10279) );
  INV_X1 U11846 ( .A(n14251), .ZN(n10056) );
  INV_X1 U11847 ( .A(n14252), .ZN(n10057) );
  NOR2_X1 U11848 ( .A1(n14258), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10085) );
  NAND2_X1 U11849 ( .A1(n9795), .A2(n9794), .ZN(n16345) );
  AND2_X1 U11850 ( .A1(n16361), .A2(n9749), .ZN(n9794) );
  NAND2_X1 U11851 ( .A1(n14260), .A2(n9796), .ZN(n9795) );
  AND2_X1 U11852 ( .A1(n12651), .A2(n12040), .ZN(n19669) );
  INV_X1 U11853 ( .A(n19669), .ZN(n17133) );
  NAND2_X1 U11854 ( .A1(n19683), .A2(n14264), .ZN(n9986) );
  INV_X1 U11855 ( .A(n9986), .ZN(n16408) );
  INV_X1 U11856 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20335) );
  AND2_X1 U11857 ( .A1(n13774), .A2(n13773), .ZN(n20323) );
  INV_X1 U11858 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20317) );
  XNOR2_X1 U11859 ( .A(n13676), .B(n13675), .ZN(n20308) );
  INV_X1 U11860 ( .A(n13674), .ZN(n13676) );
  INV_X1 U11861 ( .A(n19692), .ZN(n20309) );
  NOR2_X1 U11862 ( .A1(n17294), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n12930) );
  XNOR2_X1 U11863 ( .A(n17280), .B(n12923), .ZN(n12924) );
  OR2_X1 U11864 ( .A1(n11346), .A2(n11345), .ZN(n18104) );
  OR2_X1 U11865 ( .A1(n13921), .A2(n10033), .ZN(n18105) );
  INV_X1 U11866 ( .A(n18123), .ZN(n18128) );
  NOR2_X1 U11867 ( .A1(n16886), .A2(n13921), .ZN(n18127) );
  NOR2_X1 U11868 ( .A1(n19472), .A2(n19349), .ZN(n19469) );
  NAND2_X1 U11869 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9884) );
  NOR2_X1 U11870 ( .A1(n10768), .A2(n10716), .ZN(n10725) );
  AOI22_X1 U11871 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12458), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U11872 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12458), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12473) );
  AND2_X2 U11873 ( .A1(n10315), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9989) );
  AOI21_X1 U11874 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n9729), .ZN(n13101) );
  AOI21_X1 U11875 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(n9741), .ZN(n13096) );
  NAND3_X1 U11876 ( .A1(n9965), .A2(n9960), .A3(n9877), .ZN(n12641) );
  NOR2_X1 U11877 ( .A1(n12426), .A2(n9962), .ZN(n9960) );
  NAND2_X1 U11878 ( .A1(n9659), .A2(n12467), .ZN(n9962) );
  NAND2_X1 U11879 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10083) );
  NAND2_X1 U11880 ( .A1(n10077), .A2(n10266), .ZN(n10070) );
  NAND2_X1 U11881 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10077) );
  NAND2_X1 U11882 ( .A1(n19843), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10084) );
  NAND2_X1 U11883 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10075) );
  NAND2_X1 U11884 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10076) );
  NAND2_X1 U11885 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10078) );
  NAND2_X1 U11886 ( .A1(n12454), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10079) );
  NAND2_X1 U11887 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10073) );
  INV_X1 U11888 ( .A(n16558), .ZN(n11746) );
  AND2_X1 U11889 ( .A1(n10746), .A2(n10747), .ZN(n10753) );
  NAND2_X1 U11890 ( .A1(n10475), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10247) );
  INV_X1 U11891 ( .A(n10482), .ZN(n10689) );
  INV_X1 U11892 ( .A(n10597), .ZN(n10497) );
  AOI21_X1 U11893 ( .B1(n10517), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10518), .ZN(n10544) );
  AOI22_X1 U11894 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U11895 ( .A1(n10532), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U11896 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10402), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U11897 ( .A1(n10453), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10532), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U11898 ( .A1(n10757), .A2(n13715), .ZN(n10764) );
  NOR2_X2 U11899 ( .A1(n12433), .A2(n12438), .ZN(n12429) );
  AOI21_X1 U11900 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n9761), .ZN(n13158) );
  AOI21_X1 U11901 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A(n9760), .ZN(n13153) );
  AOI21_X1 U11902 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n9745), .ZN(n13138) );
  AOI21_X1 U11903 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(n9744), .ZN(n13133) );
  AOI21_X1 U11904 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n9743), .ZN(n13123) );
  AOI21_X1 U11905 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(n9742), .ZN(n13118) );
  AOI21_X1 U11906 ( .B1(n13188), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(n9657), .ZN(n13085) );
  AOI21_X1 U11907 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n9728), .ZN(n13089) );
  NOR2_X1 U11908 ( .A1(n12042), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U11909 ( .A1(n11746), .A2(n12065), .ZN(n11754) );
  NAND2_X1 U11910 ( .A1(n10193), .A2(n12585), .ZN(n9864) );
  AOI22_X1 U11911 ( .A1(n12052), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U11912 ( .A1(n12066), .A2(n11962), .ZN(n12296) );
  XNOR2_X1 U11913 ( .A(n13646), .B(n12065), .ZN(n12022) );
  NAND2_X1 U11914 ( .A1(n11955), .A2(n9981), .ZN(n9980) );
  NAND2_X1 U11915 ( .A1(n9982), .A2(n12609), .ZN(n9981) );
  AND3_X1 U11916 ( .A1(n11950), .A2(n11949), .A3(n11948), .ZN(n11954) );
  INV_X1 U11917 ( .A(n16546), .ZN(n11716) );
  AND3_X1 U11918 ( .A1(n11683), .A2(n11682), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U11919 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U11920 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11710) );
  AND3_X1 U11921 ( .A1(n11646), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11645), .ZN(n11648) );
  AND2_X1 U11922 ( .A1(n13083), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11642) );
  XNOR2_X1 U11923 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11937) );
  NAND2_X1 U11924 ( .A1(n11924), .A2(n11923), .ZN(n11938) );
  AND2_X1 U11925 ( .A1(n11545), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11554) );
  INV_X1 U11926 ( .A(n11534), .ZN(n11536) );
  NAND2_X1 U11927 ( .A1(n18899), .A2(n9893), .ZN(n11534) );
  INV_X1 U11928 ( .A(n18896), .ZN(n9893) );
  NAND2_X1 U11929 ( .A1(n18873), .A2(n18031), .ZN(n11516) );
  NAND2_X1 U11930 ( .A1(n10437), .A2(n10597), .ZN(n10442) );
  AND2_X1 U11931 ( .A1(n11154), .A2(n14568), .ZN(n14508) );
  INV_X1 U11932 ( .A(n13428), .ZN(n11235) );
  AND2_X1 U11933 ( .A1(n11118), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U11934 ( .A1(n14425), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13428) );
  AND2_X1 U11935 ( .A1(n10116), .A2(n9747), .ZN(n10115) );
  OR2_X1 U11936 ( .A1(n10118), .A2(n9735), .ZN(n10116) );
  NAND2_X1 U11937 ( .A1(n14729), .A2(n10118), .ZN(n14688) );
  NOR2_X1 U11938 ( .A1(n10539), .A2(n10538), .ZN(n10605) );
  OR2_X1 U11939 ( .A1(n9886), .A2(n13946), .ZN(n10614) );
  INV_X1 U11940 ( .A(n14523), .ZN(n10121) );
  INV_X1 U11941 ( .A(n14543), .ZN(n13334) );
  NAND2_X1 U11942 ( .A1(n9603), .A2(n10060), .ZN(n15010) );
  INV_X1 U11943 ( .A(n10684), .ZN(n10692) );
  AND2_X1 U11944 ( .A1(n13286), .A2(n10124), .ZN(n10123) );
  INV_X1 U11945 ( .A(n17117), .ZN(n10124) );
  OR2_X1 U11946 ( .A1(n10663), .A2(n10662), .ZN(n10682) );
  OR2_X1 U11947 ( .A1(n20515), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U11948 ( .A1(n20515), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9828) );
  OR2_X1 U11949 ( .A1(n10592), .A2(n10591), .ZN(n10670) );
  INV_X1 U11950 ( .A(n13347), .ZN(n13337) );
  NAND2_X1 U11951 ( .A1(n14058), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10635) );
  OR2_X1 U11952 ( .A1(n10580), .A2(n10579), .ZN(n10645) );
  AOI21_X1 U11953 ( .B1(n13347), .B2(n13268), .A(n9678), .ZN(n13269) );
  NAND2_X1 U11954 ( .A1(n9942), .A2(n14116), .ZN(n9941) );
  INV_X1 U11955 ( .A(n14105), .ZN(n9942) );
  OAI211_X1 U11956 ( .C1(n10507), .C2(n10553), .A(n10495), .B(n10494), .ZN(
        n10508) );
  NAND2_X1 U11957 ( .A1(n10569), .A2(n10568), .ZN(n10631) );
  AND2_X1 U11958 ( .A1(n10497), .A2(n15378), .ZN(n14266) );
  NAND2_X1 U11959 ( .A1(n10503), .A2(n10505), .ZN(n10506) );
  AOI22_X1 U11960 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10556), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U11961 ( .A1(n10554), .A2(n10553), .ZN(n10768) );
  AOI21_X1 U11962 ( .B1(n9938), .B2(n9689), .A(n9932), .ZN(n10767) );
  NAND2_X1 U11963 ( .A1(n9935), .A2(n9933), .ZN(n9932) );
  INV_X1 U11964 ( .A(n10166), .ZN(n10163) );
  NAND2_X1 U11965 ( .A1(n9809), .A2(n12362), .ZN(n12524) );
  INV_X1 U11966 ( .A(n12517), .ZN(n9809) );
  NOR2_X1 U11967 ( .A1(n10171), .A2(n12544), .ZN(n10170) );
  NAND2_X1 U11968 ( .A1(n12485), .A2(n12359), .ZN(n12542) );
  AND2_X1 U11969 ( .A1(n12486), .A2(n12358), .ZN(n12359) );
  NAND2_X1 U11970 ( .A1(n16554), .A2(n12347), .ZN(n9871) );
  NAND2_X1 U11971 ( .A1(n9782), .A2(n9781), .ZN(n11811) );
  INV_X1 U11972 ( .A(n11781), .ZN(n9781) );
  INV_X1 U11973 ( .A(n11782), .ZN(n9782) );
  CLKBUF_X1 U11974 ( .A(n13076), .Z(n13210) );
  CLKBUF_X1 U11975 ( .A(n13077), .Z(n13212) );
  CLKBUF_X1 U11976 ( .A(n13078), .Z(n13211) );
  AOI21_X1 U11977 ( .B1(n13207), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A(n9759), .ZN(n13184) );
  AOI21_X1 U11978 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n9763), .ZN(n13176) );
  AOI21_X1 U11979 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(n9762), .ZN(n13171) );
  INV_X1 U11980 ( .A(n15854), .ZN(n10206) );
  INV_X1 U11981 ( .A(n14011), .ZN(n10205) );
  OR2_X1 U11982 ( .A1(n13479), .A2(n14089), .ZN(n14086) );
  NOR2_X1 U11983 ( .A1(n10220), .A2(n15457), .ZN(n10219) );
  NOR2_X1 U11984 ( .A1(n12802), .A2(n12801), .ZN(n12800) );
  NOR2_X1 U11985 ( .A1(n12779), .A2(n12783), .ZN(n12782) );
  AND2_X1 U11986 ( .A1(n10208), .A2(n13902), .ZN(n10207) );
  INV_X1 U11987 ( .A(n16239), .ZN(n10006) );
  INV_X1 U11988 ( .A(n15738), .ZN(n10046) );
  INV_X1 U11989 ( .A(n10273), .ZN(n10272) );
  INV_X1 U11990 ( .A(n10271), .ZN(n10270) );
  OAI21_X1 U11991 ( .B1(n10274), .B2(n10272), .A(n16229), .ZN(n10271) );
  NAND2_X1 U11992 ( .A1(n10254), .A2(n11758), .ZN(n11773) );
  NAND2_X1 U11993 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  XNOR2_X1 U11994 ( .A(n12601), .B(n12649), .ZN(n12599) );
  INV_X1 U11995 ( .A(n15491), .ZN(n10233) );
  AND2_X1 U11996 ( .A1(n11887), .A2(n15509), .ZN(n15494) );
  INV_X1 U11997 ( .A(n10212), .ZN(n10210) );
  AND2_X1 U11998 ( .A1(n15582), .A2(n12644), .ZN(n12558) );
  NAND2_X1 U11999 ( .A1(n10214), .A2(n15604), .ZN(n10213) );
  INV_X1 U12000 ( .A(n14254), .ZN(n10214) );
  INV_X1 U12001 ( .A(n10050), .ZN(n10049) );
  OAI21_X1 U12002 ( .B1(n10276), .B2(n10051), .A(n12725), .ZN(n10050) );
  INV_X1 U12003 ( .A(n16139), .ZN(n10051) );
  INV_X1 U12004 ( .A(n13907), .ZN(n10225) );
  INV_X1 U12005 ( .A(n19531), .ZN(n9956) );
  NAND2_X1 U12006 ( .A1(n9959), .A2(n12630), .ZN(n9957) );
  AND2_X1 U12007 ( .A1(n11822), .A2(n10209), .ZN(n10208) );
  INV_X1 U12008 ( .A(n13454), .ZN(n10209) );
  INV_X1 U12009 ( .A(n11902), .ZN(n11884) );
  INV_X1 U12010 ( .A(n16231), .ZN(n11823) );
  NAND2_X1 U12011 ( .A1(n16252), .A2(n12626), .ZN(n12631) );
  NAND2_X1 U12012 ( .A1(n9965), .A2(n12422), .ZN(n12427) );
  NAND2_X1 U12013 ( .A1(n12428), .A2(n12354), .ZN(n10047) );
  NAND2_X1 U12015 ( .A1(n12004), .A2(n16542), .ZN(n9783) );
  INV_X1 U12016 ( .A(n12421), .ZN(n12081) );
  NAND2_X1 U12017 ( .A1(n12953), .A2(n20318), .ZN(n12972) );
  NOR2_X2 U12018 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16579) );
  INV_X1 U12019 ( .A(n12015), .ZN(n11964) );
  NAND2_X1 U12020 ( .A1(n9978), .A2(n9977), .ZN(n11966) );
  NAND2_X1 U12021 ( .A1(n17153), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9977) );
  NAND2_X1 U12022 ( .A1(n9979), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U12023 ( .A1(n9980), .A2(n11961), .ZN(n9979) );
  AOI22_X1 U12024 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11705) );
  NOR2_X1 U12025 ( .A1(n20101), .A2(n20303), .ZN(n16534) );
  AOI22_X1 U12026 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11721) );
  OR2_X1 U12027 ( .A1(n11561), .A2(n11577), .ZN(n11570) );
  OAI211_X1 U12028 ( .C1(n10153), .C2(n18343), .A(n10154), .B(n10152), .ZN(
        n11401) );
  AOI21_X1 U12029 ( .B1(n10160), .B2(n18367), .A(n18267), .ZN(n10154) );
  NAND2_X1 U12030 ( .A1(n10155), .A2(n9725), .ZN(n10152) );
  NOR2_X1 U12031 ( .A1(n10160), .A2(n10155), .ZN(n10153) );
  NAND2_X1 U12032 ( .A1(n9906), .A2(n9905), .ZN(n11608) );
  NAND2_X1 U12033 ( .A1(n9907), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9905) );
  OAI21_X1 U12034 ( .B1(n9907), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n9644), .ZN(n9906) );
  INV_X1 U12035 ( .A(n10149), .ZN(n10148) );
  NOR2_X1 U12036 ( .A1(n10150), .A2(n9918), .ZN(n9917) );
  NOR4_X1 U12037 ( .A1(n18885), .A2(n18889), .A3(n11516), .A4(n11534), .ZN(
        n11540) );
  NOR2_X1 U12038 ( .A1(n19471), .A2(n11516), .ZN(n11521) );
  INV_X1 U12039 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U12040 ( .A1(n11487), .A2(n11486), .ZN(n13809) );
  INV_X1 U12041 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20393) );
  XNOR2_X1 U12042 ( .A(n13729), .B(n21030), .ZN(n14166) );
  INV_X1 U12043 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14773) );
  AND2_X1 U12044 ( .A1(n13273), .A2(n13272), .ZN(n13841) );
  NOR2_X1 U12045 ( .A1(n14055), .A2(n14054), .ZN(n14004) );
  NAND2_X1 U12046 ( .A1(n10796), .A2(n10983), .ZN(n10804) );
  INV_X1 U12047 ( .A(n11066), .ZN(n10996) );
  AND2_X1 U12048 ( .A1(n11102), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11083) );
  AND2_X1 U12049 ( .A1(n10942), .A2(n10941), .ZN(n10986) );
  NAND2_X1 U12050 ( .A1(n10890), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10940) );
  INV_X1 U12051 ( .A(n10873), .ZN(n10874) );
  NAND2_X1 U12052 ( .A1(n10857), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10873) );
  INV_X1 U12053 ( .A(n10856), .ZN(n10857) );
  AND3_X1 U12054 ( .A1(n10845), .A2(n10844), .A3(n10843), .ZN(n14240) );
  CLKBUF_X1 U12055 ( .A(n14238), .Z(n14239) );
  AOI21_X1 U12056 ( .B1(n10831), .B2(n10983), .A(n10830), .ZN(n14199) );
  AOI21_X1 U12057 ( .B1(n10825), .B2(n10983), .A(n10824), .ZN(n14194) );
  NAND2_X1 U12058 ( .A1(n14004), .A2(n14003), .ZN(n14193) );
  NAND2_X1 U12059 ( .A1(n10806), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10814) );
  NAND2_X1 U12060 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10797) );
  AND2_X1 U12061 ( .A1(n10793), .A2(n10795), .ZN(n10289) );
  NOR2_X1 U12062 ( .A1(n10105), .A2(n9738), .ZN(n10104) );
  NAND2_X1 U12063 ( .A1(n9821), .A2(n9643), .ZN(n10103) );
  NAND2_X1 U12064 ( .A1(n10794), .A2(n10289), .ZN(n13838) );
  AND2_X1 U12065 ( .A1(n10240), .A2(n14328), .ZN(n10239) );
  AND2_X1 U12066 ( .A1(n9645), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9825) );
  NOR2_X1 U12067 ( .A1(n10064), .A2(n10241), .ZN(n10063) );
  INV_X1 U12068 ( .A(n14962), .ZN(n10064) );
  NOR2_X2 U12069 ( .A1(n14469), .A2(n13355), .ZN(n14472) );
  NAND2_X1 U12070 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  AOI21_X1 U12071 ( .B1(n15293), .B2(n15163), .A(n14353), .ZN(n9948) );
  NAND2_X1 U12072 ( .A1(n15201), .A2(n9703), .ZN(n15179) );
  NOR2_X1 U12073 ( .A1(n15213), .A2(n9930), .ZN(n15201) );
  AND2_X1 U12074 ( .A1(n20573), .A2(n15203), .ZN(n9930) );
  NAND2_X1 U12075 ( .A1(n14542), .A2(n13334), .ZN(n14545) );
  NAND2_X1 U12076 ( .A1(n9890), .A2(n15049), .ZN(n15002) );
  AOI21_X1 U12077 ( .B1(n10061), .B2(n9928), .A(n15049), .ZN(n9927) );
  INV_X1 U12078 ( .A(n9990), .ZN(n9928) );
  NAND2_X1 U12079 ( .A1(n15038), .A2(n9991), .ZN(n9990) );
  AND2_X1 U12080 ( .A1(n10127), .A2(n14583), .ZN(n10126) );
  AND2_X1 U12081 ( .A1(n13324), .A2(n13323), .ZN(n14597) );
  NAND2_X1 U12082 ( .A1(n14631), .A2(n10129), .ZN(n14618) );
  INV_X1 U12083 ( .A(n10061), .ZN(n10707) );
  INV_X1 U12084 ( .A(n15058), .ZN(n9833) );
  NAND2_X1 U12085 ( .A1(n15052), .A2(n9705), .ZN(n15056) );
  NOR2_X2 U12086 ( .A1(n14216), .A2(n10131), .ZN(n14704) );
  NAND2_X1 U12087 ( .A1(n10132), .A2(n9693), .ZN(n10131) );
  NAND2_X1 U12088 ( .A1(n10134), .A2(n10132), .ZN(n14719) );
  INV_X1 U12089 ( .A(n14209), .ZN(n9812) );
  AND2_X1 U12090 ( .A1(n10638), .A2(n10637), .ZN(n20517) );
  INV_X1 U12091 ( .A(n10436), .ZN(n21298) );
  OR2_X1 U12092 ( .A1(n14134), .A2(n20580), .ZN(n14135) );
  NAND2_X1 U12093 ( .A1(n10782), .A2(n20351), .ZN(n10245) );
  INV_X1 U12094 ( .A(n10631), .ZN(n15407) );
  INV_X1 U12095 ( .A(n14162), .ZN(n15408) );
  INV_X1 U12096 ( .A(n10441), .ZN(n14425) );
  INV_X1 U12097 ( .A(n20994), .ZN(n21004) );
  NAND2_X1 U12098 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20653), .ZN(n20589) );
  AND2_X1 U12099 ( .A1(n21180), .A2(n15409), .ZN(n21089) );
  INV_X1 U12100 ( .A(n14116), .ZN(n14187) );
  AND2_X1 U12101 ( .A1(n9622), .A2(n21093), .ZN(n21126) );
  INV_X1 U12102 ( .A(n20589), .ZN(n20648) );
  AND2_X1 U12103 ( .A1(n9622), .A2(n14163), .ZN(n20993) );
  NAND2_X1 U12104 ( .A1(n20519), .A2(n14430), .ZN(n20646) );
  NOR2_X1 U12105 ( .A1(n15409), .A2(n20900), .ZN(n21179) );
  NOR2_X1 U12106 ( .A1(n14162), .A2(n15407), .ZN(n21180) );
  AOI21_X1 U12107 ( .B1(n21084), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20763), 
        .ZN(n21182) );
  AOI221_X2 U12108 ( .B1(n21296), .B2(n17056), .C1(n17131), .C2(n17056), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n20653) );
  AND2_X1 U12109 ( .A1(n15388), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17084) );
  NAND2_X1 U12110 ( .A1(n11765), .A2(n12609), .ZN(n12304) );
  AND4_X1 U12111 ( .A1(n16566), .A2(n12065), .A3(n16546), .A4(n11759), .ZN(
        n11745) );
  NAND2_X1 U12112 ( .A1(n12821), .A2(n16025), .ZN(n15439) );
  NAND2_X1 U12113 ( .A1(n10179), .A2(n10178), .ZN(n12821) );
  AOI21_X1 U12114 ( .B1(n10180), .B2(n15683), .A(n15683), .ZN(n10178) );
  INV_X1 U12115 ( .A(n12386), .ZN(n12378) );
  OAI21_X1 U12116 ( .B1(n12551), .B2(n10167), .A(n10166), .ZN(n12571) );
  NAND2_X1 U12117 ( .A1(n19559), .A2(n9675), .ZN(n10188) );
  INV_X1 U12118 ( .A(n15559), .ZN(n10187) );
  NOR2_X1 U12119 ( .A1(n15628), .A2(n12790), .ZN(n15609) );
  AND2_X1 U12120 ( .A1(n12522), .A2(n12530), .ZN(n15660) );
  AND2_X1 U12121 ( .A1(n13470), .A2(n16134), .ZN(n15657) );
  OR2_X1 U12122 ( .A1(n13487), .A2(n16154), .ZN(n19517) );
  INV_X1 U12123 ( .A(n12763), .ZN(n10191) );
  INV_X1 U12124 ( .A(n15784), .ZN(n15733) );
  NAND2_X1 U12125 ( .A1(n13935), .A2(n13934), .ZN(n13937) );
  NOR2_X1 U12126 ( .A1(n16504), .A2(n15765), .ZN(n15767) );
  CLKBUF_X1 U12127 ( .A(n11786), .Z(n12836) );
  NAND2_X1 U12128 ( .A1(n10219), .A2(n12675), .ZN(n10218) );
  NAND2_X1 U12129 ( .A1(n10224), .A2(n9639), .ZN(n14046) );
  AND2_X2 U12130 ( .A1(n15453), .A2(n12287), .ZN(n12693) );
  AOI21_X1 U12131 ( .B1(n13207), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A(n9767), .ZN(n13202) );
  AOI21_X1 U12132 ( .B1(n16574), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n9766), .ZN(n13208) );
  INV_X1 U12133 ( .A(n13166), .ZN(n10199) );
  CLKBUF_X1 U12134 ( .A(n15837), .Z(n15838) );
  NAND2_X1 U12135 ( .A1(n13019), .A2(n13018), .ZN(n15859) );
  AND2_X1 U12136 ( .A1(n12259), .A2(n12258), .ZN(n14156) );
  CLKBUF_X1 U12137 ( .A(n14154), .Z(n15861) );
  NOR2_X1 U12138 ( .A1(n14010), .A2(n9724), .ZN(n15870) );
  AND3_X1 U12139 ( .A1(n12174), .A2(n12173), .A3(n12172), .ZN(n13820) );
  AND3_X1 U12140 ( .A1(n12159), .A2(n12158), .A3(n12157), .ZN(n13749) );
  NAND2_X1 U12141 ( .A1(n10230), .A2(n12145), .ZN(n13757) );
  AOI21_X1 U12142 ( .B1(n9642), .B2(n9629), .A(n10229), .ZN(n10228) );
  OR2_X1 U12143 ( .A1(n15739), .A2(n15995), .ZN(n15997) );
  INV_X1 U12144 ( .A(n13593), .ZN(n19628) );
  NOR2_X1 U12145 ( .A1(n12831), .A2(n12833), .ZN(n13563) );
  INV_X1 U12146 ( .A(n12832), .ZN(n12833) );
  NAND2_X1 U12147 ( .A1(n12798), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12802) );
  AND2_X1 U12148 ( .A1(n12796), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U12149 ( .A1(n12788), .A2(n9656), .ZN(n12794) );
  AND2_X1 U12150 ( .A1(n12782), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12788) );
  NOR2_X1 U12151 ( .A1(n13994), .A2(n10221), .ZN(n15655) );
  NAND2_X1 U12152 ( .A1(n9639), .A2(n10222), .ZN(n10221) );
  INV_X1 U12153 ( .A(n13477), .ZN(n10222) );
  NAND2_X1 U12154 ( .A1(n10185), .A2(n9649), .ZN(n12777) );
  INV_X1 U12155 ( .A(n12772), .ZN(n10185) );
  OR2_X1 U12156 ( .A1(n15700), .A2(n13995), .ZN(n13994) );
  NAND2_X1 U12157 ( .A1(n10190), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10189) );
  INV_X1 U12158 ( .A(n10192), .ZN(n10190) );
  NAND2_X1 U12159 ( .A1(n11837), .A2(n11836), .ZN(n15700) );
  INV_X1 U12160 ( .A(n15698), .ZN(n11836) );
  INV_X1 U12161 ( .A(n13879), .ZN(n11837) );
  XNOR2_X1 U12162 ( .A(n12394), .B(n12393), .ZN(n12395) );
  AND2_X1 U12163 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12760) );
  INV_X1 U12164 ( .A(n12599), .ZN(n10093) );
  NAND2_X1 U12165 ( .A1(n12648), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U12166 ( .A1(n10198), .A2(n12686), .ZN(n9860) );
  NOR2_X1 U12167 ( .A1(n12656), .A2(n9862), .ZN(n9861) );
  INV_X1 U12168 ( .A(n12686), .ZN(n9862) );
  NAND2_X1 U12169 ( .A1(n9682), .A2(n12644), .ZN(n16021) );
  NAND2_X1 U12170 ( .A1(n9804), .A2(n9803), .ZN(n9802) );
  INV_X1 U12171 ( .A(n16016), .ZN(n9801) );
  INV_X1 U12172 ( .A(n10003), .ZN(n10001) );
  NAND2_X1 U12173 ( .A1(n12333), .A2(n16296), .ZN(n16283) );
  NAND2_X1 U12174 ( .A1(n15506), .A2(n9726), .ZN(n15493) );
  AND2_X1 U12175 ( .A1(n16411), .A2(n9984), .ZN(n16297) );
  NOR2_X1 U12176 ( .A1(n12325), .A2(n16308), .ZN(n9984) );
  NAND2_X1 U12177 ( .A1(n9631), .A2(n10021), .ZN(n16296) );
  INV_X1 U12178 ( .A(n10022), .ZN(n10021) );
  OAI21_X1 U12179 ( .B1(n16408), .B2(n12647), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U12180 ( .A1(n9709), .A2(n9870), .ZN(n16049) );
  NAND2_X1 U12181 ( .A1(n12503), .A2(n10195), .ZN(n9870) );
  AND2_X1 U12182 ( .A1(n12270), .A2(n12269), .ZN(n15522) );
  NAND2_X1 U12183 ( .A1(n13252), .A2(n12268), .ZN(n15545) );
  INV_X1 U12184 ( .A(n13252), .ZN(n15543) );
  NAND2_X1 U12185 ( .A1(n12742), .A2(n13255), .ZN(n16061) );
  NOR2_X1 U12186 ( .A1(n9683), .A2(n9841), .ZN(n9840) );
  AND2_X1 U12187 ( .A1(n9842), .A2(n9844), .ZN(n9841) );
  INV_X1 U12188 ( .A(n9844), .ZN(n9843) );
  INV_X1 U12189 ( .A(n12741), .ZN(n10097) );
  NOR2_X1 U12190 ( .A1(n14290), .A2(n16306), .ZN(n10098) );
  NAND2_X1 U12191 ( .A1(n9856), .A2(n14290), .ZN(n14285) );
  INV_X1 U12192 ( .A(n9856), .ZN(n12566) );
  NOR2_X1 U12193 ( .A1(n12741), .A2(n16306), .ZN(n9972) );
  INV_X1 U12194 ( .A(n16071), .ZN(n10280) );
  NAND2_X1 U12195 ( .A1(n16089), .A2(n10285), .ZN(n9845) );
  NOR2_X1 U12196 ( .A1(n15635), .A2(n14156), .ZN(n15591) );
  OR2_X1 U12197 ( .A1(n14261), .A2(n19657), .ZN(n9796) );
  AND3_X1 U12198 ( .A1(n12225), .A2(n12224), .A3(n12223), .ZN(n13986) );
  AOI21_X1 U12199 ( .B1(n10278), .B2(n12501), .A(n10277), .ZN(n10276) );
  INV_X1 U12200 ( .A(n16149), .ZN(n10277) );
  NOR2_X1 U12201 ( .A1(n13994), .A2(n13907), .ZN(n13908) );
  NAND2_X1 U12202 ( .A1(n12645), .A2(n12644), .ZN(n12643) );
  NAND2_X1 U12203 ( .A1(n12639), .A2(n12638), .ZN(n9847) );
  AOI21_X1 U12204 ( .B1(n15725), .B2(n12644), .A(n13456), .ZN(n10009) );
  NAND2_X1 U12205 ( .A1(n11823), .A2(n11822), .ZN(n16233) );
  NOR2_X1 U12206 ( .A1(n16506), .A2(n12294), .ZN(n16594) );
  INV_X1 U12207 ( .A(n13675), .ZN(n9775) );
  CLKBUF_X1 U12208 ( .A(n13861), .Z(n16518) );
  NAND2_X1 U12209 ( .A1(n12312), .A2(n11760), .ZN(n11776) );
  CLKBUF_X1 U12210 ( .A(n11914), .Z(n13864) );
  OAI21_X1 U12211 ( .B1(n16531), .B2(n16529), .A(n9780), .ZN(n9779) );
  NAND2_X1 U12212 ( .A1(n20144), .A2(n20145), .ZN(n9780) );
  INV_X1 U12213 ( .A(n12458), .ZN(n19751) );
  OR2_X1 U12214 ( .A1(n12459), .A2(n19873), .ZN(n19877) );
  INV_X1 U12215 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20034) );
  NAND2_X1 U12216 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20152), .ZN(n16553) );
  NAND2_X1 U12217 ( .A1(n16534), .A2(n16533), .ZN(n16563) );
  NAND2_X1 U12218 ( .A1(n13618), .A2(n16534), .ZN(n16564) );
  AND2_X1 U12219 ( .A1(n12015), .A2(n12014), .ZN(n16591) );
  NAND2_X1 U12220 ( .A1(n18873), .A2(n19471), .ZN(n11526) );
  NAND2_X1 U12221 ( .A1(n11540), .A2(n18880), .ZN(n17249) );
  INV_X1 U12222 ( .A(n11542), .ZN(n12927) );
  INV_X1 U12223 ( .A(n12913), .ZN(n12916) );
  NAND2_X1 U12224 ( .A1(n17425), .A2(n17508), .ZN(n17410) );
  NAND2_X1 U12225 ( .A1(n12920), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12922) );
  AOI21_X1 U12226 ( .B1(n17858), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n10037), .ZN(n10036) );
  INV_X1 U12227 ( .A(n11435), .ZN(n10038) );
  NOR2_X1 U12228 ( .A1(n18137), .A2(n18205), .ZN(n10024) );
  INV_X1 U12229 ( .A(n18899), .ZN(n17990) );
  NAND2_X1 U12230 ( .A1(n10032), .A2(n18071), .ZN(n10030) );
  NAND2_X1 U12231 ( .A1(n10034), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n10033) );
  INV_X1 U12232 ( .A(n18109), .ZN(n10034) );
  OR2_X1 U12233 ( .A1(n11303), .A2(n11302), .ZN(n11587) );
  AOI21_X1 U12234 ( .B1(n13919), .B2(n13918), .A(n16883), .ZN(n16937) );
  NOR2_X1 U12235 ( .A1(n18243), .A2(n12911), .ZN(n12914) );
  INV_X1 U12236 ( .A(n18278), .ZN(n10146) );
  OR2_X1 U12237 ( .A1(n11618), .A2(n12903), .ZN(n12907) );
  NAND2_X1 U12238 ( .A1(n10138), .A2(n11617), .ZN(n10137) );
  INV_X1 U12239 ( .A(n18351), .ZN(n11617) );
  NOR2_X1 U12240 ( .A1(n18394), .A2(n10142), .ZN(n10141) );
  NAND2_X1 U12241 ( .A1(n10139), .A2(n10140), .ZN(n18380) );
  NOR2_X1 U12242 ( .A1(n18394), .A2(n10143), .ZN(n10139) );
  OR2_X1 U12243 ( .A1(n18277), .A2(n18561), .ZN(n11622) );
  INV_X1 U12244 ( .A(n18440), .ZN(n11615) );
  NAND2_X1 U12245 ( .A1(n12900), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16762) );
  NAND2_X1 U12246 ( .A1(n18547), .A2(n18519), .ZN(n18478) );
  NOR2_X1 U12247 ( .A1(n16670), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9920) );
  NAND2_X1 U12248 ( .A1(n11405), .A2(n16854), .ZN(n16829) );
  AND2_X1 U12249 ( .A1(n16835), .A2(n9909), .ZN(n9908) );
  INV_X1 U12250 ( .A(n18241), .ZN(n9909) );
  OR2_X1 U12251 ( .A1(n18286), .A2(n18333), .ZN(n18312) );
  AND2_X1 U12252 ( .A1(n18369), .A2(n18635), .ZN(n18329) );
  NAND2_X1 U12253 ( .A1(n18299), .A2(n18286), .ZN(n18334) );
  OAI21_X1 U12254 ( .B1(n18368), .B2(n9758), .A(n18369), .ZN(n18348) );
  NOR2_X2 U12255 ( .A1(n19485), .A2(n13917), .ZN(n19300) );
  OAI21_X1 U12256 ( .B1(n9892), .B2(n9891), .A(n11543), .ZN(n16906) );
  NAND2_X1 U12257 ( .A1(n18189), .A2(n9651), .ZN(n9891) );
  AOI21_X1 U12258 ( .B1(n18724), .B2(n18661), .A(n16834), .ZN(n16851) );
  XNOR2_X1 U12259 ( .A(n11386), .B(n11384), .ZN(n18473) );
  OAI21_X1 U12260 ( .B1(n18536), .B2(n9901), .A(n9900), .ZN(n18518) );
  NAND2_X1 U12261 ( .A1(n9677), .A2(n9902), .ZN(n9901) );
  NAND2_X1 U12262 ( .A1(n18528), .A2(n9677), .ZN(n9900) );
  INV_X1 U12263 ( .A(n11599), .ZN(n9902) );
  OR2_X1 U12264 ( .A1(n19295), .A2(n18834), .ZN(n16772) );
  NOR3_X1 U12265 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n17254), .ZN(n19159) );
  INV_X1 U12266 ( .A(n13809), .ZN(n18880) );
  INV_X1 U12267 ( .A(n11517), .ZN(n18889) );
  NAND2_X1 U12268 ( .A1(n19475), .A2(n18872), .ZN(n18914) );
  NAND2_X1 U12269 ( .A1(n9895), .A2(n9894), .ZN(n19301) );
  NAND2_X1 U12270 ( .A1(n19298), .A2(n11569), .ZN(n9895) );
  INV_X1 U12271 ( .A(n13658), .ZN(n9988) );
  NAND2_X1 U12272 ( .A1(n14779), .A2(n13387), .ZN(n20392) );
  INV_X1 U12273 ( .A(n20425), .ZN(n20408) );
  AND2_X1 U12275 ( .A1(n14779), .A2(n13377), .ZN(n20425) );
  INV_X1 U12276 ( .A(n20430), .ZN(n20394) );
  INV_X1 U12277 ( .A(n14835), .ZN(n20448) );
  AND2_X2 U12278 ( .A1(n13767), .A2(n13828), .ZN(n20452) );
  AND2_X1 U12279 ( .A1(n14932), .A2(n14445), .ZN(n14911) );
  INV_X1 U12280 ( .A(n14931), .ZN(n14936) );
  INV_X1 U12281 ( .A(n14917), .ZN(n14938) );
  INV_X1 U12282 ( .A(n20484), .ZN(n20453) );
  NAND2_X1 U12283 ( .A1(n13380), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13381) );
  NOR2_X1 U12284 ( .A1(n10111), .A2(n10107), .ZN(n10108) );
  NAND2_X1 U12285 ( .A1(n15052), .A2(n15051), .ZN(n9835) );
  INV_X2 U12286 ( .A(n15122), .ZN(n20519) );
  XNOR2_X1 U12287 ( .A(n9826), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14412) );
  NAND2_X1 U12288 ( .A1(n10242), .A2(n9827), .ZN(n9826) );
  NAND2_X1 U12289 ( .A1(n14955), .A2(n9825), .ZN(n9827) );
  NAND2_X1 U12290 ( .A1(n10714), .A2(n10239), .ZN(n10242) );
  INV_X1 U12291 ( .A(n9947), .ZN(n15157) );
  NAND2_X1 U12292 ( .A1(n14955), .A2(n9634), .ZN(n14326) );
  NAND2_X1 U12293 ( .A1(n10714), .A2(n10713), .ZN(n14327) );
  XNOR2_X1 U12294 ( .A(n9994), .B(n14945), .ZN(n15170) );
  NAND2_X1 U12295 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  OAI21_X1 U12296 ( .B1(n14943), .B2(n14941), .A(n9623), .ZN(n9995) );
  NAND2_X1 U12297 ( .A1(n14944), .A2(n15049), .ZN(n9996) );
  INV_X1 U12298 ( .A(n9949), .ZN(n15174) );
  XNOR2_X1 U12299 ( .A(n9923), .B(n14956), .ZN(n15178) );
  NAND2_X1 U12300 ( .A1(n9925), .A2(n9924), .ZN(n9923) );
  NAND2_X1 U12301 ( .A1(n14954), .A2(n9623), .ZN(n9924) );
  NAND2_X1 U12302 ( .A1(n14955), .A2(n15049), .ZN(n9925) );
  NAND2_X1 U12303 ( .A1(n15257), .A2(n14350), .ZN(n15237) );
  XNOR2_X1 U12304 ( .A(n9831), .B(n15283), .ZN(n15288) );
  NAND2_X1 U12305 ( .A1(n9834), .A2(n9832), .ZN(n9831) );
  NAND2_X1 U12306 ( .A1(n15076), .A2(n9833), .ZN(n9832) );
  NAND2_X1 U12307 ( .A1(n15068), .A2(n15058), .ZN(n9834) );
  NAND2_X1 U12308 ( .A1(n17099), .A2(n10675), .ZN(n10059) );
  INV_X1 U12309 ( .A(n20576), .ZN(n20550) );
  AND2_X1 U12310 ( .A1(n14212), .A2(n14128), .ZN(n20540) );
  AND2_X1 U12311 ( .A1(n14134), .A2(n15367), .ZN(n20573) );
  INV_X1 U12312 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15388) );
  AND2_X1 U12314 ( .A1(n13727), .A2(n13726), .ZN(n21281) );
  AND2_X1 U12315 ( .A1(n14177), .A2(n14176), .ZN(n20613) );
  OR2_X1 U12316 ( .A1(n14180), .A2(n14179), .ZN(n14184) );
  INV_X1 U12317 ( .A(n20613), .ZN(n20655) );
  AND2_X1 U12318 ( .A1(n20727), .A2(n20667), .ZN(n20714) );
  AND2_X1 U12319 ( .A1(n20727), .A2(n21126), .ZN(n20748) );
  OAI21_X1 U12320 ( .B1(n20782), .B2(n20764), .A(n21138), .ZN(n20785) );
  OAI211_X1 U12321 ( .C1(n20922), .C2(n21041), .A(n20967), .B(n20903), .ZN(
        n20925) );
  OR2_X1 U12322 ( .A1(n20902), .A2(n20901), .ZN(n20903) );
  OAI21_X1 U12323 ( .B1(n20971), .B2(n20970), .A(n20969), .ZN(n20989) );
  OAI211_X1 U12324 ( .C1(n21042), .C2(n21041), .A(n21138), .B(n21040), .ZN(
        n21079) );
  AOI22_X1 U12325 ( .A1(n21039), .A2(n21032), .B1(n21129), .B2(n21036), .ZN(
        n21083) );
  OAI211_X1 U12326 ( .C1(n21165), .C2(n21139), .A(n21138), .B(n21137), .ZN(
        n21168) );
  AND2_X1 U12327 ( .A1(n20653), .A2(n20591), .ZN(n21177) );
  AND2_X1 U12328 ( .A1(n10431), .A2(n20648), .ZN(n21191) );
  AND2_X1 U12329 ( .A1(n20653), .A2(n20600), .ZN(n21192) );
  AND2_X1 U12330 ( .A1(n20611), .A2(n20648), .ZN(n21206) );
  AND2_X1 U12331 ( .A1(n10414), .A2(n20648), .ZN(n21212) );
  AND2_X1 U12332 ( .A1(n20653), .A2(n20622), .ZN(n21213) );
  AND2_X1 U12333 ( .A1(n20629), .A2(n20648), .ZN(n21218) );
  AND2_X1 U12334 ( .A1(n20653), .A2(n20631), .ZN(n21219) );
  AND2_X1 U12335 ( .A1(n20653), .A2(n20639), .ZN(n21227) );
  AND2_X1 U12336 ( .A1(n20649), .A2(n20648), .ZN(n21232) );
  NAND2_X1 U12337 ( .A1(n21180), .A2(n20993), .ZN(n21241) );
  INV_X1 U12338 ( .A(n21224), .ZN(n21237) );
  AND2_X1 U12339 ( .A1(n20653), .A2(n20652), .ZN(n21235) );
  OR2_X1 U12340 ( .A1(n14173), .A2(n21041), .ZN(n17056) );
  INV_X1 U12341 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n13525) );
  INV_X1 U12342 ( .A(n21265), .ZN(n13559) );
  INV_X1 U12343 ( .A(n9982), .ZN(n12000) );
  AND2_X1 U12344 ( .A1(n12387), .A2(n12386), .ZN(n15519) );
  OR2_X1 U12345 ( .A1(n19554), .A2(n20318), .ZN(n19513) );
  NAND2_X1 U12346 ( .A1(n10204), .A2(n14011), .ZN(n14048) );
  OR2_X1 U12347 ( .A1(n12184), .A2(n12183), .ZN(n13912) );
  INV_X1 U12348 ( .A(n20308), .ZN(n19782) );
  AND2_X1 U12349 ( .A1(n13649), .A2(n16626), .ZN(n19575) );
  NAND2_X1 U12350 ( .A1(n10227), .A2(n9629), .ZN(n13753) );
  OR2_X1 U12351 ( .A1(n15739), .A2(n9642), .ZN(n10227) );
  OR2_X1 U12352 ( .A1(n15985), .A2(n13741), .ZN(n19577) );
  INV_X1 U12353 ( .A(n15981), .ZN(n19578) );
  INV_X1 U12354 ( .A(n19577), .ZN(n14151) );
  OAI21_X1 U12355 ( .B1(n13681), .B2(n13680), .A(n13679), .ZN(n13682) );
  INV_X2 U12356 ( .A(n19592), .ZN(n19622) );
  NOR2_X1 U12357 ( .A1(n12894), .A2(n19640), .ZN(n12895) );
  AOI21_X1 U12358 ( .B1(n16303), .B2(n19642), .A(n16045), .ZN(n9788) );
  INV_X1 U12359 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16236) );
  CLKBUF_X1 U12360 ( .A(n13865), .Z(n16257) );
  NAND2_X1 U12361 ( .A1(n10029), .A2(n10025), .ZN(n12338) );
  NAND2_X1 U12362 ( .A1(n16272), .A2(n12337), .ZN(n10029) );
  AND2_X1 U12363 ( .A1(n12742), .A2(n10003), .ZN(n16031) );
  OAI21_X1 U12364 ( .B1(n12503), .B2(n10197), .A(n10195), .ZN(n16057) );
  NAND2_X1 U12365 ( .A1(n12503), .A2(n12502), .ZN(n10194) );
  INV_X1 U12366 ( .A(n16411), .ZN(n16438) );
  OAI21_X1 U12367 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n12742), .A(
        n16174), .ZN(n16449) );
  NOR2_X1 U12368 ( .A1(n19661), .A2(n12321), .ZN(n16464) );
  NAND2_X1 U12369 ( .A1(n16244), .A2(n10274), .ZN(n10269) );
  NAND2_X1 U12370 ( .A1(n9687), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19661) );
  NAND2_X1 U12371 ( .A1(n16509), .A2(n13647), .ZN(n20330) );
  OR2_X1 U12372 ( .A1(n20313), .A2(n16495), .ZN(n20303) );
  INV_X1 U12373 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20325) );
  INV_X1 U12374 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16621) );
  INV_X1 U12375 ( .A(n13644), .ZN(n16509) );
  AND2_X1 U12376 ( .A1(n16592), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17152) );
  INV_X1 U12377 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16605) );
  AND2_X1 U12378 ( .A1(n13640), .A2(n13639), .ZN(n20301) );
  OAI21_X1 U12379 ( .B1(n16567), .B2(n16532), .A(n20152), .ZN(n16562) );
  NAND2_X1 U12380 ( .A1(n9777), .A2(n9776), .ZN(n16570) );
  OR2_X1 U12381 ( .A1(n16531), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12382 ( .A1(n9779), .A2(n9778), .ZN(n9777) );
  INV_X1 U12383 ( .A(n16567), .ZN(n9778) );
  NOR2_X1 U12384 ( .A1(n19942), .A2(n19881), .ZN(n19708) );
  OR2_X1 U12385 ( .A1(n19840), .A2(n20072), .ZN(n19783) );
  OAI21_X1 U12386 ( .B1(n19816), .B2(n19815), .A(n19814), .ZN(n19834) );
  OAI211_X1 U12387 ( .C1(n19848), .C2(n19847), .A(n19846), .B(n20152), .ZN(
        n19867) );
  INV_X1 U12388 ( .A(n19863), .ZN(n19866) );
  NOR2_X1 U12389 ( .A1(n20156), .A2(n19840), .ZN(n19882) );
  INV_X1 U12390 ( .A(n19886), .ZN(n19901) );
  OAI21_X1 U12391 ( .B1(n19928), .B2(n19913), .A(n20152), .ZN(n19929) );
  OAI211_X1 U12392 ( .C1(n19941), .C2(n19940), .A(n20152), .B(n19939), .ZN(
        n19966) );
  NOR2_X1 U12393 ( .A1(n20073), .A2(n19942), .ZN(n19974) );
  NOR2_X1 U12394 ( .A1(n20073), .A2(n20304), .ZN(n20039) );
  NOR2_X1 U12395 ( .A1(n20094), .A2(n20072), .ZN(n20064) );
  OAI22_X1 U12396 ( .A1(n20588), .A2(n16564), .B1(n17232), .B2(n16563), .ZN(
        n20102) );
  OAI22_X1 U12397 ( .A1(n20628), .A2(n16564), .B1(n17237), .B2(n16563), .ZN(
        n20127) );
  OAI21_X1 U12398 ( .B1(n20107), .B2(n20106), .A(n20105), .ZN(n20138) );
  NOR2_X2 U12399 ( .A1(n20073), .A2(n20072), .ZN(n20137) );
  NOR2_X1 U12400 ( .A1(n20094), .A2(n20156), .ZN(n20143) );
  OAI22_X1 U12401 ( .A1(n20645), .A2(n16564), .B1(n17240), .B2(n16563), .ZN(
        n20136) );
  AND2_X1 U12402 ( .A1(n20152), .A2(n16525), .ZN(n20150) );
  INV_X1 U12403 ( .A(n20102), .ZN(n20162) );
  AND2_X1 U12404 ( .A1(n15806), .A2(n16565), .ZN(n20163) );
  INV_X1 U12405 ( .A(n19948), .ZN(n20164) );
  INV_X1 U12406 ( .A(n20111), .ZN(n20168) );
  AND2_X1 U12407 ( .A1(n20152), .A2(n16541), .ZN(n20170) );
  INV_X1 U12408 ( .A(n20115), .ZN(n20174) );
  AND2_X1 U12409 ( .A1(n16546), .A2(n16565), .ZN(n20175) );
  INV_X1 U12410 ( .A(n19954), .ZN(n20176) );
  INV_X1 U12411 ( .A(n20119), .ZN(n20180) );
  AND2_X1 U12412 ( .A1(n20152), .A2(n19576), .ZN(n20182) );
  INV_X1 U12413 ( .A(n19960), .ZN(n20188) );
  INV_X1 U12414 ( .A(n20127), .ZN(n20192) );
  AND2_X1 U12415 ( .A1(n20152), .A2(n16557), .ZN(n20194) );
  INV_X1 U12416 ( .A(n20131), .ZN(n20198) );
  INV_X1 U12417 ( .A(n20158), .ZN(n20205) );
  NOR2_X1 U12418 ( .A1(n20151), .A2(n20148), .ZN(n20202) );
  AND2_X1 U12419 ( .A1(n20152), .A2(n16561), .ZN(n20201) );
  INV_X1 U12420 ( .A(n20143), .ZN(n20208) );
  INV_X1 U12421 ( .A(n20136), .ZN(n20209) );
  INV_X1 U12422 ( .A(n19487), .ZN(n19486) );
  NAND2_X1 U12423 ( .A1(n17310), .A2(n17312), .ZN(n17311) );
  NAND2_X1 U12424 ( .A1(n17331), .A2(n17508), .ZN(n17320) );
  NAND2_X1 U12425 ( .A1(n17340), .A2(n17342), .ZN(n17341) );
  NAND2_X1 U12426 ( .A1(n17359), .A2(n17508), .ZN(n10135) );
  NAND2_X1 U12427 ( .A1(n17392), .A2(n17508), .ZN(n17380) );
  NAND2_X1 U12428 ( .A1(n17402), .A2(n18325), .ZN(n17403) );
  INV_X1 U12429 ( .A(n17493), .ZN(n17450) );
  AND2_X1 U12430 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17672), .ZN(n17666) );
  NOR2_X1 U12431 ( .A1(n17608), .A2(n17667), .ZN(n17672) );
  NOR2_X1 U12432 ( .A1(n17606), .A2(n17695), .ZN(n17673) );
  NOR3_X1 U12433 ( .A1(n17928), .A2(n17953), .A3(n17954), .ZN(n17927) );
  INV_X1 U12434 ( .A(n17959), .ZN(n17954) );
  NOR2_X1 U12435 ( .A1(n17962), .A2(n17957), .ZN(n17959) );
  NOR3_X1 U12436 ( .A1(n17564), .A2(n17984), .A3(n17968), .ZN(n17967) );
  INV_X1 U12437 ( .A(n17998), .ZN(n17994) );
  NAND2_X1 U12438 ( .A1(n18011), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n18006) );
  NOR2_X1 U12439 ( .A1(n18140), .A2(n18016), .ZN(n18011) );
  INV_X1 U12440 ( .A(n18022), .ZN(n18017) );
  NAND2_X1 U12441 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18017), .ZN(n18016) );
  NOR2_X1 U12442 ( .A1(n18026), .A2(n18031), .ZN(n18023) );
  NAND2_X1 U12443 ( .A1(n18023), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18022) );
  NOR2_X1 U12444 ( .A1(n18154), .A2(n18058), .ZN(n18049) );
  INV_X1 U12445 ( .A(n18038), .ZN(n18064) );
  NOR2_X1 U12446 ( .A1(n13921), .A2(n10031), .ZN(n18099) );
  INV_X1 U12447 ( .A(n18127), .ZN(n18120) );
  OR2_X1 U12448 ( .A1(n11288), .A2(n11287), .ZN(n18126) );
  NOR2_X1 U12449 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  NOR2_X1 U12450 ( .A1(n18188), .A2(n18132), .ZN(n18171) );
  CLKBUF_X1 U12451 ( .A(n18175), .Z(n18183) );
  NAND2_X1 U12452 ( .A1(n18220), .A2(n19471), .ZN(n18230) );
  INV_X1 U12453 ( .A(n18230), .ZN(n18237) );
  AND2_X1 U12454 ( .A1(n11620), .A2(n9684), .ZN(n18261) );
  INV_X1 U12455 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18548) );
  INV_X1 U12456 ( .A(n18478), .ZN(n18562) );
  INV_X1 U12457 ( .A(n16865), .ZN(n9912) );
  NOR2_X1 U12458 ( .A1(n10159), .A2(n10158), .ZN(n16749) );
  INV_X1 U12459 ( .A(n11399), .ZN(n10158) );
  OAI21_X1 U12460 ( .B1(n10151), .B2(n9725), .A(n10155), .ZN(n18258) );
  INV_X1 U12461 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19472) );
  NAND2_X1 U12462 ( .A1(n18373), .A2(n16835), .ZN(n18671) );
  INV_X1 U12463 ( .A(n9907), .ZN(n18480) );
  NAND2_X1 U12464 ( .A1(n18489), .A2(n18488), .ZN(n18487) );
  NAND2_X1 U12465 ( .A1(n18500), .A2(n11378), .ZN(n18489) );
  INV_X1 U12466 ( .A(n9904), .ZN(n18529) );
  OR2_X1 U12467 ( .A1(n18536), .A2(n11599), .ZN(n9904) );
  AND2_X1 U12468 ( .A1(n19298), .A2(n18813), .ZN(n18845) );
  INV_X1 U12469 ( .A(n18839), .ZN(n18848) );
  INV_X1 U12470 ( .A(n17052), .ZN(n16931) );
  INV_X1 U12471 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17054) );
  OR4_X1 U12472 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), 
        .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n16879), .ZN(n19355) );
  INV_X1 U12473 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19373) );
  NAND2_X1 U12474 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19373), .ZN(n19482) );
  CLKBUF_X1 U12475 ( .A(n17227), .Z(n17241) );
  NOR2_X1 U12476 ( .A1(n17204), .A2(n17164), .ZN(n17201) );
  AND4_X1 U12477 ( .A1(n20379), .A2(n20378), .A3(n20416), .A4(n20377), .ZN(
        n20380) );
  NAND2_X1 U12478 ( .A1(n14432), .A2(n14431), .ZN(n14435) );
  NAND2_X1 U12479 ( .A1(n14400), .A2(n9944), .ZN(n14355) );
  NAND2_X1 U12480 ( .A1(n12855), .A2(n12854), .ZN(n12863) );
  AND2_X1 U12481 ( .A1(n12861), .A2(n12860), .ZN(n12862) );
  INV_X1 U12482 ( .A(n14463), .ZN(n12855) );
  AND2_X1 U12483 ( .A1(n12850), .A2(n12849), .ZN(n12851) );
  OAI21_X1 U12484 ( .B1(n12827), .B2(n19537), .A(n9650), .ZN(n10183) );
  AOI21_X1 U12485 ( .B1(n15449), .B2(n12827), .A(n15448), .ZN(n15450) );
  AOI211_X1 U12486 ( .C1(n19532), .C2(n9682), .A(n15464), .B(n15463), .ZN(
        n15465) );
  NOR2_X1 U12487 ( .A1(n9857), .A2(n9854), .ZN(n15574) );
  AOI211_X1 U12488 ( .C1(n15984), .C2(BUF2_REG_28__SCAN_IN), .A(n15908), .B(
        n15907), .ZN(n15909) );
  INV_X1 U12489 ( .A(n12949), .ZN(n12951) );
  INV_X1 U12490 ( .A(n16026), .ZN(n9953) );
  NAND2_X1 U12491 ( .A1(n16278), .A2(n16263), .ZN(n9954) );
  INV_X1 U12492 ( .A(n12721), .ZN(n12722) );
  OAI211_X1 U12493 ( .C1(n19640), .C2(n14381), .A(n10177), .B(n10176), .ZN(
        P2_U2988) );
  AOI21_X1 U12494 ( .B1(n15812), .B2(n19642), .A(n14370), .ZN(n10176) );
  OR2_X1 U12495 ( .A1(n14379), .A2(n16253), .ZN(n10177) );
  NAND2_X1 U12496 ( .A1(n10011), .A2(n9786), .ZN(P2_U2990) );
  NAND2_X1 U12497 ( .A1(n9637), .A2(n16263), .ZN(n10011) );
  INV_X1 U12498 ( .A(n9787), .ZN(n9786) );
  OAI21_X1 U12499 ( .B1(n16301), .B2(n16253), .A(n9788), .ZN(n9787) );
  NAND2_X1 U12500 ( .A1(n12743), .A2(n19636), .ZN(n12752) );
  AND2_X1 U12501 ( .A1(n9964), .A2(n12872), .ZN(n12873) );
  OAI211_X1 U12502 ( .C1(n16088), .C2(n16253), .A(n10054), .B(n10053), .ZN(
        P2_U2997) );
  AOI21_X1 U12503 ( .B1(n16087), .B2(n19642), .A(n16086), .ZN(n10053) );
  NAND2_X1 U12504 ( .A1(n10055), .A2(n16263), .ZN(n10054) );
  AOI21_X1 U12505 ( .B1(n12701), .B2(n19657), .A(n9973), .ZN(n12703) );
  OAI21_X1 U12506 ( .B1(n12700), .B2(n12699), .A(n9974), .ZN(n9973) );
  NOR2_X1 U12507 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  OAI21_X1 U12508 ( .B1(n14381), .B2(n19653), .A(n9773), .ZN(P2_U3020) );
  INV_X1 U12509 ( .A(n9774), .ZN(n9773) );
  OAI21_X1 U12510 ( .B1(n14379), .B2(n19668), .A(n9652), .ZN(n9774) );
  NOR2_X1 U12511 ( .A1(n16302), .A2(n9851), .ZN(n9850) );
  NAND2_X1 U12512 ( .A1(n9637), .A2(n19672), .ZN(n9849) );
  AND2_X1 U12513 ( .A1(n16303), .A2(n19669), .ZN(n9851) );
  NAND2_X1 U12514 ( .A1(n9967), .A2(n9966), .ZN(n12887) );
  NAND2_X1 U12515 ( .A1(n9970), .A2(n9680), .ZN(n9967) );
  OAI211_X1 U12516 ( .C1(n19653), .C2(n16085), .A(n9797), .B(n9793), .ZN(
        P2_U3029) );
  NOR2_X1 U12517 ( .A1(n9647), .A2(n9708), .ZN(n9797) );
  OR2_X1 U12518 ( .A1(n16437), .A2(n19653), .ZN(n9879) );
  NAND2_X1 U12519 ( .A1(n12924), .A2(n17558), .ZN(n12943) );
  OR2_X1 U12520 ( .A1(n17279), .A2(n12930), .ZN(n12941) );
  NOR2_X1 U12521 ( .A1(n13921), .A2(n18109), .ZN(n18106) );
  OAI21_X1 U12522 ( .B1(n9913), .B2(n18834), .A(n9910), .ZN(P3_U2836) );
  INV_X1 U12523 ( .A(n9911), .ZN(n9910) );
  AOI22_X1 U12524 ( .A1(n16863), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n16862), .B2(n18590), .ZN(n9913) );
  OAI21_X1 U12525 ( .B1(n16866), .B2(n18753), .A(n9912), .ZN(n9911) );
  NAND2_X2 U12526 ( .A1(n11258), .A2(n16911), .ZN(n9754) );
  OR2_X1 U12527 ( .A1(n12478), .A2(n12116), .ZN(n9629) );
  AND4_X1 U12528 ( .A1(n12472), .A2(n12473), .A3(n12476), .A4(n12471), .ZN(
        n9630) );
  XNOR2_X1 U12529 ( .A(n12922), .B(n10147), .ZN(n12902) );
  AND2_X1 U12530 ( .A1(n10023), .A2(n9694), .ZN(n9631) );
  AND2_X1 U12531 ( .A1(n12046), .A2(n12045), .ZN(n12090) );
  OR2_X1 U12532 ( .A1(n9628), .A2(n10211), .ZN(n9632) );
  OR2_X1 U12533 ( .A1(n9619), .A2(n13775), .ZN(n9633) );
  NAND2_X1 U12534 ( .A1(n10134), .A2(n14234), .ZN(n14233) );
  NAND2_X1 U12535 ( .A1(n15558), .A2(n15559), .ZN(n15547) );
  AND2_X1 U12536 ( .A1(n9623), .A2(n15154), .ZN(n9634) );
  AND2_X1 U12537 ( .A1(n9633), .A2(n11758), .ZN(n9635) );
  AND4_X1 U12538 ( .A1(n12477), .A2(n12474), .A3(n12475), .A4(n12470), .ZN(
        n9636) );
  XNOR2_X1 U12539 ( .A(n16041), .B(n16040), .ZN(n9637) );
  AND2_X1 U12540 ( .A1(n10225), .A2(n13494), .ZN(n9638) );
  AND2_X1 U12541 ( .A1(n9638), .A2(n10223), .ZN(n9639) );
  NOR2_X1 U12542 ( .A1(n9628), .A2(n10213), .ZN(n9640) );
  AND2_X1 U12543 ( .A1(n14542), .A2(n9733), .ZN(n14511) );
  NAND2_X1 U12544 ( .A1(n10191), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12765) );
  OR2_X1 U12545 ( .A1(n15995), .A2(n13457), .ZN(n9642) );
  AND2_X1 U12546 ( .A1(n10604), .A2(n10983), .ZN(n9643) );
  NAND2_X1 U12547 ( .A1(n10052), .A2(n10276), .ZN(n16137) );
  XNOR2_X1 U12548 ( .A(n18110), .B(n18481), .ZN(n9644) );
  NAND2_X1 U12549 ( .A1(n17330), .A2(n18244), .ZN(n17331) );
  AND2_X1 U12550 ( .A1(n9634), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9645) );
  AND2_X1 U12551 ( .A1(n9684), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9646) );
  AND2_X1 U12552 ( .A1(n9874), .A2(n10085), .ZN(n9647) );
  AND2_X1 U12553 ( .A1(n16535), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9648) );
  NOR2_X1 U12554 ( .A1(n16152), .A2(n15675), .ZN(n9649) );
  AND2_X1 U12555 ( .A1(n15772), .A2(n10184), .ZN(n9650) );
  NOR2_X1 U12556 ( .A1(n11544), .A2(n13916), .ZN(n9651) );
  NOR2_X1 U12557 ( .A1(n14380), .A2(n9714), .ZN(n9652) );
  AND2_X1 U12558 ( .A1(n15049), .A2(n9756), .ZN(n9653) );
  AND2_X1 U12559 ( .A1(n10060), .A2(n10252), .ZN(n9654) );
  INV_X2 U12560 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U12561 ( .A1(n10224), .A2(n9638), .ZN(n13493) );
  AND2_X1 U12562 ( .A1(n13019), .A2(n9732), .ZN(n15843) );
  AND2_X1 U12563 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9655) );
  AND2_X1 U12564 ( .A1(n9655), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9656) );
  AND2_X1 U12565 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n9657)
         );
  NAND2_X1 U12566 ( .A1(n17358), .A2(n18281), .ZN(n17359) );
  AND2_X1 U12567 ( .A1(n9726), .A2(n10232), .ZN(n9658) );
  AND2_X1 U12568 ( .A1(n12451), .A2(n12422), .ZN(n9659) );
  AND2_X1 U12569 ( .A1(n12647), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9660) );
  AND2_X1 U12570 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9661) );
  OR2_X1 U12571 ( .A1(n9632), .A2(n12713), .ZN(n9662) );
  AND2_X2 U12572 ( .A1(n13076), .A2(n13875), .ZN(n11974) );
  INV_X1 U12573 ( .A(n11467), .ZN(n11434) );
  NAND2_X1 U12574 ( .A1(n15037), .A2(n15038), .ZN(n15009) );
  OR2_X1 U12575 ( .A1(n12812), .A2(n12816), .ZN(n9663) );
  NAND2_X1 U12576 ( .A1(n10245), .A2(n10475), .ZN(n10615) );
  NAND2_X1 U12577 ( .A1(n11811), .A2(n11783), .ZN(n9664) );
  AND2_X1 U12578 ( .A1(n11273), .A2(n9898), .ZN(n9665) );
  NAND2_X1 U12579 ( .A1(n11259), .A2(n16911), .ZN(n9666) );
  INV_X1 U12580 ( .A(n14481), .ZN(n10107) );
  NAND2_X1 U12581 ( .A1(n12983), .A2(n12982), .ZN(n13845) );
  OR2_X1 U12582 ( .A1(n13792), .A2(n9988), .ZN(n9667) );
  NAND2_X2 U12583 ( .A1(n16911), .A2(n11260), .ZN(n9668) );
  NOR2_X1 U12584 ( .A1(n12763), .A2(n10192), .ZN(n12768) );
  AND2_X1 U12585 ( .A1(n14238), .A2(n14743), .ZN(n14729) );
  AND3_X1 U12586 ( .A1(n10265), .A2(n10079), .A3(n10073), .ZN(n9669) );
  AND2_X1 U12587 ( .A1(n14729), .A2(n14728), .ZN(n9670) );
  AND2_X1 U12588 ( .A1(n12818), .A2(n15479), .ZN(n9671) );
  OR2_X1 U12589 ( .A1(n15098), .A2(n15352), .ZN(n9672) );
  INV_X1 U12590 ( .A(n10023), .ZN(n17142) );
  NAND2_X1 U12591 ( .A1(n12823), .A2(n15440), .ZN(n12827) );
  AND2_X1 U12592 ( .A1(n18011), .A2(n10024), .ZN(n9674) );
  OR2_X1 U12593 ( .A1(n12799), .A2(n10187), .ZN(n9675) );
  INV_X1 U12594 ( .A(n10284), .ZN(n10283) );
  OAI21_X1 U12595 ( .B1(n14251), .B2(n12564), .A(n12730), .ZN(n10284) );
  AND4_X1 U12596 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n9676) );
  OR2_X1 U12597 ( .A1(n18805), .A2(n11600), .ZN(n9677) );
  NOR2_X1 U12598 ( .A1(n15545), .A2(n15522), .ZN(n15506) );
  NOR3_X1 U12599 ( .A1(n15635), .A2(n10238), .A3(n14156), .ZN(n12877) );
  AND2_X1 U12600 ( .A1(n13360), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n9678) );
  INV_X1 U12601 ( .A(n14399), .ZN(n9946) );
  AND2_X1 U12602 ( .A1(n12886), .A2(n16306), .ZN(n9679) );
  AND2_X1 U12603 ( .A1(n12886), .A2(n9972), .ZN(n9680) );
  OR3_X1 U12604 ( .A1(n9662), .A2(n11907), .A3(n10218), .ZN(n9681) );
  NOR2_X1 U12605 ( .A1(n16163), .A2(n16175), .ZN(n12507) );
  INV_X1 U12606 ( .A(n12507), .ZN(n10197) );
  AND2_X1 U12607 ( .A1(n12594), .A2(n12375), .ZN(n9682) );
  NAND2_X1 U12608 ( .A1(n10268), .A2(n10267), .ZN(n13463) );
  NAND2_X1 U12609 ( .A1(n10269), .A2(n10273), .ZN(n16228) );
  NAND2_X1 U12610 ( .A1(n10698), .A2(n10697), .ZN(n14224) );
  NAND2_X1 U12611 ( .A1(n10059), .A2(n10677), .ZN(n17093) );
  NAND2_X1 U12612 ( .A1(n12468), .A2(n12469), .ZN(n16213) );
  NAND2_X1 U12613 ( .A1(n14285), .A2(n14283), .ZN(n9683) );
  NOR2_X1 U12614 ( .A1(n12763), .A2(n10189), .ZN(n12770) );
  AND2_X1 U12615 ( .A1(n11619), .A2(n10146), .ZN(n9684) );
  NAND2_X1 U12616 ( .A1(n10754), .A2(n13369), .ZN(n9685) );
  AND2_X1 U12617 ( .A1(n18373), .A2(n9908), .ZN(n9686) );
  AND2_X1 U12618 ( .A1(n9986), .A2(n9985), .ZN(n9687) );
  AND2_X1 U12619 ( .A1(n12981), .A2(n12978), .ZN(n13783) );
  INV_X2 U12620 ( .A(n12116), .ZN(n12041) );
  AND4_X1 U12621 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n9688) );
  NOR2_X1 U12622 ( .A1(n10432), .A2(n9617), .ZN(n10436) );
  NAND2_X1 U12623 ( .A1(n9603), .A2(n10707), .ZN(n15037) );
  AND2_X1 U12624 ( .A1(n12538), .A2(n10170), .ZN(n12520) );
  XNOR2_X1 U12625 ( .A(n13167), .B(n10199), .ZN(n15798) );
  AND3_X1 U12626 ( .A1(n10740), .A2(n9685), .A3(n10761), .ZN(n9689) );
  NOR2_X1 U12627 ( .A1(n14251), .A2(n10286), .ZN(n10285) );
  INV_X1 U12628 ( .A(n10285), .ZN(n9842) );
  NAND2_X1 U12629 ( .A1(n12538), .A2(n12541), .ZN(n12540) );
  NAND2_X1 U12630 ( .A1(n16137), .A2(n16139), .ZN(n16138) );
  OR3_X1 U12631 ( .A1(n15635), .A2(n10238), .A3(n10236), .ZN(n9690) );
  AND2_X1 U12632 ( .A1(n12684), .A2(n12686), .ZN(n9691) );
  AND2_X1 U12633 ( .A1(n9845), .A2(n9844), .ZN(n9692) );
  INV_X1 U12634 ( .A(n16017), .ZN(n9803) );
  AND2_X1 U12635 ( .A1(n14703), .A2(n14718), .ZN(n9693) );
  OR2_X1 U12636 ( .A1(n16408), .A2(n16450), .ZN(n9694) );
  XOR2_X1 U12637 ( .A(n10264), .B(n12649), .Z(n9695) );
  NAND2_X1 U12638 ( .A1(n16213), .A2(n16214), .ZN(n16158) );
  AND3_X1 U12639 ( .A1(n12455), .A2(n9880), .A3(n12456), .ZN(n9696) );
  OR2_X1 U12640 ( .A1(n9619), .A2(n12343), .ZN(n9697) );
  OR2_X1 U12641 ( .A1(n14260), .A2(n12741), .ZN(n9698) );
  AND2_X1 U12642 ( .A1(n12483), .A2(n12342), .ZN(n9699) );
  AND2_X1 U12643 ( .A1(n10198), .A2(n12656), .ZN(n9700) );
  AND2_X1 U12644 ( .A1(n10170), .A2(n12361), .ZN(n9701) );
  AND2_X1 U12645 ( .A1(n9951), .A2(n11811), .ZN(n9702) );
  NAND2_X1 U12646 ( .A1(n9617), .A2(n20611), .ZN(n13266) );
  OR2_X1 U12647 ( .A1(n20566), .A2(n15180), .ZN(n9703) );
  NOR2_X1 U12648 ( .A1(n12572), .A2(n12383), .ZN(n9704) );
  AND2_X1 U12649 ( .A1(n15051), .A2(n15053), .ZN(n9705) );
  NOR2_X1 U12650 ( .A1(n14313), .A2(n10113), .ZN(n14839) );
  INV_X1 U12651 ( .A(n19643), .ZN(n15779) );
  AND2_X1 U12652 ( .A1(n12401), .A2(n12402), .ZN(n19643) );
  AND3_X1 U12653 ( .A1(n10102), .A2(n10101), .A3(n14003), .ZN(n14198) );
  AND2_X1 U12654 ( .A1(n9784), .A2(n15425), .ZN(n9706) );
  INV_X1 U12655 ( .A(n10241), .ZN(n10240) );
  NAND2_X1 U12656 ( .A1(n10713), .A2(n14353), .ZN(n10241) );
  OR2_X1 U12657 ( .A1(n10507), .A2(n10554), .ZN(n9707) );
  OR2_X1 U12658 ( .A1(n10086), .A2(n14259), .ZN(n9708) );
  NOR2_X1 U12659 ( .A1(n9628), .A2(n14254), .ZN(n14253) );
  NAND2_X1 U12660 ( .A1(n12538), .A2(n9701), .ZN(n12517) );
  AND2_X1 U12661 ( .A1(n12577), .A2(n10193), .ZN(n9709) );
  AND2_X1 U12662 ( .A1(n15506), .A2(n9658), .ZN(n9710) );
  AND2_X1 U12663 ( .A1(n12710), .A2(n9803), .ZN(n9711) );
  INV_X1 U12664 ( .A(n12688), .ZN(n10198) );
  NAND2_X1 U12665 ( .A1(n15293), .A2(n14351), .ZN(n9712) );
  INV_X1 U12666 ( .A(n9874), .ZN(n16350) );
  OAI21_X1 U12667 ( .B1(n16114), .B2(n19668), .A(n9875), .ZN(n9874) );
  NAND2_X1 U12668 ( .A1(n12377), .A2(n12706), .ZN(n12373) );
  NAND2_X1 U12669 ( .A1(n15506), .A2(n15507), .ZN(n15490) );
  INV_X1 U12670 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16201) );
  NAND2_X1 U12671 ( .A1(n10194), .A2(n12507), .ZN(n16148) );
  AND2_X1 U12672 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n9713)
         );
  AND2_X1 U12673 ( .A1(n15812), .A2(n19669), .ZN(n9714) );
  AND2_X1 U12674 ( .A1(n12704), .A2(n16016), .ZN(n9715) );
  OR2_X1 U12675 ( .A1(n17249), .A2(n11526), .ZN(n10018) );
  INV_X1 U12676 ( .A(n10018), .ZN(n9892) );
  AND2_X1 U12677 ( .A1(n10255), .A2(n12737), .ZN(n9716) );
  NOR2_X1 U12678 ( .A1(n12724), .A2(n10197), .ZN(n10278) );
  AND2_X1 U12679 ( .A1(n10065), .A2(n10063), .ZN(n9717) );
  AND2_X1 U12680 ( .A1(n10441), .A2(n10431), .ZN(n9718) );
  AND2_X1 U12681 ( .A1(n10115), .A2(n10993), .ZN(n9719) );
  INV_X1 U12682 ( .A(n12646), .ZN(n10090) );
  NAND2_X1 U12683 ( .A1(n10090), .A2(n12737), .ZN(n9720) );
  OR2_X1 U12684 ( .A1(n14173), .A2(n9941), .ZN(n9721) );
  AND2_X1 U12685 ( .A1(n19643), .A2(n9664), .ZN(n12414) );
  INV_X1 U12686 ( .A(n16762), .ZN(n10140) );
  NAND2_X1 U12687 ( .A1(n11775), .A2(n11752), .ZN(n12831) );
  NAND2_X1 U12688 ( .A1(n10173), .A2(n12442), .ZN(n12441) );
  NAND2_X1 U12689 ( .A1(n12715), .A2(n9661), .ZN(n12754) );
  AND2_X1 U12690 ( .A1(n10125), .A2(n10123), .ZN(n9722) );
  NAND2_X1 U12691 ( .A1(n19559), .A2(n12799), .ZN(n15558) );
  AND2_X1 U12692 ( .A1(n14631), .A2(n10127), .ZN(n9723) );
  NAND2_X1 U12693 ( .A1(n12780), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12779) );
  NAND2_X1 U12694 ( .A1(n12788), .A2(n9655), .ZN(n12791) );
  BUF_X1 U12695 ( .A(n10423), .Z(n13661) );
  OR2_X1 U12696 ( .A1(n12997), .A2(n10205), .ZN(n9724) );
  OR2_X1 U12697 ( .A1(n18367), .A2(n10157), .ZN(n9725) );
  AND2_X1 U12698 ( .A1(n10233), .A2(n15507), .ZN(n9726) );
  NOR2_X1 U12699 ( .A1(n14005), .A2(n10122), .ZN(n14202) );
  NAND2_X1 U12700 ( .A1(n10832), .A2(n14198), .ZN(n14197) );
  AND2_X1 U12701 ( .A1(n14631), .A2(n10126), .ZN(n14564) );
  NAND2_X1 U12702 ( .A1(n13893), .A2(n12253), .ZN(n14145) );
  AND2_X1 U12703 ( .A1(n12651), .A2(n20341), .ZN(n19657) );
  INV_X1 U12704 ( .A(n19672), .ZN(n19653) );
  AND2_X1 U12705 ( .A1(n12651), .A2(n20339), .ZN(n19672) );
  NOR2_X1 U12706 ( .A1(n9622), .A2(n14163), .ZN(n9727) );
  AND2_X1 U12707 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n9728) );
  AND2_X1 U12708 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n9729) );
  NAND3_X1 U12709 ( .A1(n9814), .A2(n17094), .A3(n9813), .ZN(n14208) );
  NAND2_X1 U12710 ( .A1(n10653), .A2(n10652), .ZN(n17099) );
  NAND2_X1 U12711 ( .A1(n10043), .A2(n15738), .ZN(n16244) );
  AND2_X1 U12712 ( .A1(n13018), .A2(n10206), .ZN(n9730) );
  AND2_X1 U12713 ( .A1(n13840), .A2(n13841), .ZN(n13839) );
  AND2_X1 U12714 ( .A1(n12715), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12819) );
  AND2_X1 U12715 ( .A1(n12788), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12787) );
  AND2_X1 U12716 ( .A1(n11823), .A2(n10207), .ZN(n9731) );
  AND2_X1 U12717 ( .A1(n9730), .A2(n15849), .ZN(n9732) );
  AND2_X1 U12718 ( .A1(n13334), .A2(n10121), .ZN(n9733) );
  INV_X2 U12719 ( .A(n11824), .ZN(n11906) );
  INV_X1 U12720 ( .A(n12541), .ZN(n10171) );
  AND2_X1 U12721 ( .A1(n20629), .A2(n10431), .ZN(n13715) );
  AND2_X1 U12722 ( .A1(n10141), .A2(n10140), .ZN(n9734) );
  AND2_X1 U12723 ( .A1(n13019), .A2(n9730), .ZN(n15848) );
  NAND2_X1 U12724 ( .A1(n14631), .A2(n14632), .ZN(n14616) );
  NAND2_X1 U12725 ( .A1(n10437), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10973) );
  AND2_X1 U12726 ( .A1(n14728), .A2(n10117), .ZN(n9735) );
  INV_X1 U12727 ( .A(n13994), .ZN(n10224) );
  NAND2_X1 U12728 ( .A1(n13845), .A2(n12985), .ZN(n14010) );
  INV_X1 U12730 ( .A(n14216), .ZN(n10134) );
  AND2_X1 U12731 ( .A1(n9986), .A2(n12696), .ZN(n9737) );
  INV_X1 U12732 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20351) );
  AND2_X1 U12733 ( .A1(n10791), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9738) );
  AND2_X1 U12734 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  NAND2_X1 U12735 ( .A1(n9784), .A2(n11748), .ZN(n9739) );
  AND2_X1 U12736 ( .A1(n13327), .A2(n13326), .ZN(n14583) );
  INV_X1 U12737 ( .A(n13760), .ZN(n10794) );
  AND2_X1 U12738 ( .A1(n12446), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9740) );
  AND2_X1 U12739 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n9741)
         );
  AND2_X1 U12740 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n9742)
         );
  AND2_X1 U12741 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n9743) );
  AND2_X1 U12742 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n9744)
         );
  AND2_X1 U12743 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n9745) );
  INV_X1 U12744 ( .A(n12262), .ZN(n10238) );
  OR2_X1 U12745 ( .A1(n11936), .A2(n11935), .ZN(n12451) );
  INV_X1 U12746 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17153) );
  AND2_X1 U12747 ( .A1(n18367), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9746) );
  AND2_X1 U12748 ( .A1(n15655), .A2(n15654), .ZN(n15640) );
  AND2_X1 U12749 ( .A1(n14701), .A2(n14689), .ZN(n9747) );
  AND2_X1 U12750 ( .A1(n12425), .A2(n12422), .ZN(n9748) );
  OR2_X1 U12751 ( .A1(n14264), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9749) );
  AND2_X1 U12752 ( .A1(n9656), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9750) );
  AND2_X1 U12753 ( .A1(n9733), .A2(n14512), .ZN(n9751) );
  AND2_X1 U12754 ( .A1(n9732), .A2(n15844), .ZN(n9752) );
  INV_X1 U12755 ( .A(n10282), .ZN(n10281) );
  NAND2_X1 U12756 ( .A1(n10283), .A2(n16070), .ZN(n10282) );
  AND2_X1 U12757 ( .A1(n11823), .A2(n10208), .ZN(n9753) );
  NAND2_X1 U12758 ( .A1(n10709), .A2(n10708), .ZN(n9755) );
  NAND2_X1 U12759 ( .A1(n11620), .A2(n11619), .ZN(n18274) );
  NOR2_X1 U12760 ( .A1(n12899), .A2(n17285), .ZN(n16681) );
  INV_X1 U12761 ( .A(n16263), .ZN(n19640) );
  AND2_X1 U12762 ( .A1(n12689), .A2(n15806), .ZN(n16263) );
  INV_X1 U12763 ( .A(n13752), .ZN(n10229) );
  INV_X1 U12764 ( .A(n14617), .ZN(n10130) );
  AND2_X1 U12765 ( .A1(n13814), .A2(n19469), .ZN(n18813) );
  INV_X1 U12766 ( .A(n18813), .ZN(n18834) );
  NAND2_X1 U12767 ( .A1(n11620), .A2(n9646), .ZN(n16752) );
  AOI21_X1 U12768 ( .B1(n13768), .B2(n10302), .A(n13270), .ZN(n13840) );
  NAND2_X1 U12769 ( .A1(n11623), .A2(n10298), .ZN(n12899) );
  AND2_X1 U12770 ( .A1(n16681), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12920) );
  NOR2_X1 U12771 ( .A1(n13711), .A2(n10432), .ZN(n13664) );
  OR2_X1 U12772 ( .A1(n15048), .A2(n10706), .ZN(n9756) );
  INV_X1 U12773 ( .A(n14005), .ZN(n10125) );
  AND2_X1 U12774 ( .A1(n9904), .A2(n9903), .ZN(n9757) );
  OR2_X1 U12775 ( .A1(n11391), .A2(n11392), .ZN(n9758) );
  AND2_X1 U12776 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n9759)
         );
  AND2_X1 U12777 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n9760)
         );
  AND2_X1 U12778 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n9761) );
  AND2_X1 U12779 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n9762)
         );
  AND2_X1 U12780 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n9763) );
  AND2_X1 U12781 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n9764) );
  INV_X1 U12782 ( .A(n10032), .ZN(n10031) );
  NOR2_X1 U12783 ( .A1(n10033), .A2(n18170), .ZN(n10032) );
  AND2_X1 U12784 ( .A1(n9661), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9765) );
  INV_X1 U12785 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9918) );
  INV_X1 U12786 ( .A(n19537), .ZN(n19563) );
  NAND2_X1 U12787 ( .A1(n16634), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16636) );
  NOR2_X1 U12788 ( .A1(n16762), .A2(n18394), .ZN(n17471) );
  AND2_X1 U12789 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16634) );
  INV_X1 U12790 ( .A(n15227), .ZN(n9991) );
  INV_X1 U12791 ( .A(n10710), .ZN(n10252) );
  INV_X1 U12792 ( .A(n12737), .ZN(n10088) );
  AND2_X1 U12793 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n9766) );
  AND2_X1 U12794 ( .A1(n9983), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n9767)
         );
  INV_X1 U12795 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10147) );
  INV_X1 U12796 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16652) );
  INV_X1 U12797 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U12798 ( .A1(n10098), .A2(n10097), .ZN(n10096) );
  AND2_X1 U12799 ( .A1(n10024), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9768) );
  INV_X1 U12800 ( .A(n12334), .ZN(n10004) );
  NOR2_X2 U12801 ( .A1(n17990), .A2(n18118), .ZN(n18063) );
  NOR3_X2 U12802 ( .A1(n19163), .A2(n19311), .A3(n18999), .ZN(n18972) );
  OAI22_X2 U12803 ( .A1(n20620), .A2(n20644), .B1(n20619), .B2(n20646), .ZN(
        n21155) );
  OAI22_X2 U12804 ( .A1(n20598), .A2(n20644), .B1(n20597), .B2(n20646), .ZN(
        n21142) );
  NAND2_X1 U12805 ( .A1(n20519), .A2(n14869), .ZN(n20644) );
  NOR3_X2 U12806 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19163), .A3(
        n19244), .ZN(n19062) );
  NAND2_X2 U12807 ( .A1(n21265), .A2(n13519), .ZN(n21271) );
  INV_X1 U12808 ( .A(n14465), .ZN(n21265) );
  AND2_X2 U12809 ( .A1(n9769), .A2(n12406), .ZN(n12453) );
  AND2_X2 U12810 ( .A1(n13865), .A2(n12404), .ZN(n9769) );
  NAND2_X1 U12811 ( .A1(n9771), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16159) );
  NAND3_X1 U12812 ( .A1(n9838), .A2(n9772), .A3(n12640), .ZN(n9837) );
  INV_X1 U12813 ( .A(n12481), .ZN(n9772) );
  XNOR2_X2 U12814 ( .A(n12396), .B(n12395), .ZN(n13865) );
  XNOR2_X2 U12815 ( .A(n9664), .B(n12401), .ZN(n16486) );
  XNOR2_X2 U12816 ( .A(n13783), .B(n13784), .ZN(n19692) );
  OAI21_X1 U12817 ( .B1(n12023), .B2(n12004), .A(n9783), .ZN(n12034) );
  NAND2_X1 U12818 ( .A1(n12742), .A2(n12647), .ZN(n9853) );
  NAND2_X4 U12819 ( .A1(n10087), .A2(n10089), .ZN(n12742) );
  NAND2_X1 U12820 ( .A1(n11762), .A2(n16535), .ZN(n12028) );
  NAND3_X1 U12821 ( .A1(n12312), .A2(n11760), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9791) );
  NAND3_X1 U12822 ( .A1(n11768), .A2(n11788), .A3(n12304), .ZN(n9789) );
  INV_X2 U12823 ( .A(n11786), .ZN(n12609) );
  NAND3_X1 U12824 ( .A1(n11764), .A2(n11752), .A3(n11775), .ZN(n9790) );
  NAND2_X1 U12825 ( .A1(n12705), .A2(n9715), .ZN(n12710) );
  NAND2_X1 U12826 ( .A1(n9802), .A2(n16016), .ZN(n16018) );
  NAND2_X1 U12827 ( .A1(n12340), .A2(n12342), .ZN(n9806) );
  NAND2_X1 U12828 ( .A1(n12346), .A2(n12342), .ZN(n9805) );
  NAND2_X1 U12829 ( .A1(n12616), .A2(n12342), .ZN(n12345) );
  NOR2_X2 U12830 ( .A1(n12526), .A2(n12514), .ZN(n12510) );
  NAND3_X1 U12831 ( .A1(n16279), .A2(n16280), .A3(n9810), .ZN(P2_U3018) );
  NAND3_X1 U12832 ( .A1(n9867), .A2(n10195), .A3(n12503), .ZN(n9866) );
  NAND2_X2 U12833 ( .A1(n10698), .A2(n9811), .ZN(n15045) );
  NAND2_X1 U12834 ( .A1(n10058), .A2(n17095), .ZN(n9813) );
  NAND3_X1 U12835 ( .A1(n17099), .A2(n17095), .A3(n10675), .ZN(n9814) );
  NAND2_X1 U12837 ( .A1(n13652), .A2(n10443), .ZN(n9815) );
  NAND3_X1 U12838 ( .A1(n10427), .A2(n10426), .A3(n10243), .ZN(n10517) );
  XNOR2_X2 U12839 ( .A(n10503), .B(n10504), .ZN(n10782) );
  AND2_X2 U12840 ( .A1(n9820), .A2(n9818), .ZN(n10504) );
  AND2_X2 U12841 ( .A1(n9836), .A2(n10601), .ZN(n10570) );
  NAND3_X1 U12842 ( .A1(n10712), .A2(n15002), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9824) );
  INV_X1 U12843 ( .A(n14993), .ZN(n14963) );
  OAI21_X2 U12844 ( .B1(n10805), .B2(n14068), .A(n10648), .ZN(n20515) );
  NAND2_X1 U12845 ( .A1(n9828), .A2(n14129), .ZN(n10651) );
  NAND2_X1 U12846 ( .A1(n16211), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9848) );
  NAND2_X1 U12847 ( .A1(n10013), .A2(n10066), .ZN(n13459) );
  NAND2_X1 U12848 ( .A1(n11736), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10020) );
  INV_X1 U12849 ( .A(n18268), .ZN(n16758) );
  INV_X1 U12850 ( .A(n11438), .ZN(n10037) );
  AOI211_X1 U12851 ( .C1(n18889), .C2(n16886), .A(n11519), .B(n11518), .ZN(
        n13800) );
  NAND2_X1 U12852 ( .A1(n10188), .A2(n16064), .ZN(n15530) );
  OR2_X2 U12853 ( .A1(n10408), .A2(n10407), .ZN(n10431) );
  NAND2_X1 U12854 ( .A1(n12811), .A2(n16043), .ZN(n15498) );
  NAND2_X1 U12855 ( .A1(n12807), .A2(n16047), .ZN(n15514) );
  NAND2_X1 U12856 ( .A1(n12815), .A2(n16035), .ZN(n15478) );
  NAND2_X1 U12857 ( .A1(n12818), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U12858 ( .A1(n9853), .A2(n12388), .ZN(n9852) );
  NAND2_X1 U12859 ( .A1(n9696), .A2(n10306), .ZN(n9877) );
  NAND2_X1 U12860 ( .A1(n11742), .A2(n13875), .ZN(n10019) );
  NAND2_X1 U12861 ( .A1(n14953), .A2(n14973), .ZN(n10065) );
  INV_X1 U12862 ( .A(n10642), .ZN(n9889) );
  INV_X1 U12863 ( .A(n10603), .ZN(n9836) );
  INV_X1 U12864 ( .A(n9829), .ZN(n9830) );
  OAI21_X1 U12865 ( .B1(n14094), .B2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10637), .ZN(n9829) );
  NAND3_X1 U12866 ( .A1(n9830), .A2(n10649), .A3(n10638), .ZN(n10653) );
  NAND2_X1 U12867 ( .A1(n9835), .A2(n15089), .ZN(n15091) );
  NAND2_X1 U12868 ( .A1(n15045), .A2(n15047), .ZN(n15131) );
  OR2_X1 U12869 ( .A1(n12426), .A2(n12644), .ZN(n9839) );
  NAND2_X1 U12870 ( .A1(n9845), .A2(n10283), .ZN(n16073) );
  NAND2_X2 U12871 ( .A1(n9848), .A2(n9847), .ZN(n9878) );
  OAI211_X1 U12872 ( .C1(n16301), .C2(n19668), .A(n9850), .B(n9849), .ZN(
        P2_U3022) );
  NAND2_X1 U12873 ( .A1(n12658), .A2(n12656), .ZN(n12687) );
  OR2_X1 U12874 ( .A1(n12702), .A2(n19653), .ZN(n10297) );
  NAND2_X1 U12875 ( .A1(n9864), .A2(n9867), .ZN(n9865) );
  INV_X1 U12876 ( .A(n12585), .ZN(n9869) );
  OAI211_X2 U12877 ( .C1(n12577), .C2(n9868), .A(n9866), .B(n9865), .ZN(n12705) );
  NAND2_X2 U12878 ( .A1(n12510), .A2(n12511), .ZN(n12551) );
  NAND2_X2 U12879 ( .A1(n16113), .A2(n14256), .ZN(n16114) );
  NAND2_X2 U12880 ( .A1(n9963), .A2(n9876), .ZN(n16113) );
  NAND2_X1 U12881 ( .A1(n9878), .A2(n10259), .ZN(n10258) );
  NAND2_X1 U12882 ( .A1(n9716), .A2(n9878), .ZN(n9963) );
  XNOR2_X1 U12883 ( .A(n9878), .B(n16198), .ZN(n17145) );
  NAND2_X1 U12884 ( .A1(n16436), .A2(n9879), .ZN(P2_U3036) );
  NAND2_X1 U12885 ( .A1(n20037), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n9883) );
  NAND2_X1 U12886 ( .A1(n16529), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n9881) );
  AND2_X2 U12887 ( .A1(n12411), .A2(n12415), .ZN(n16529) );
  NAND2_X1 U12888 ( .A1(n19685), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n9882) );
  AND2_X2 U12889 ( .A1(n12411), .A2(n12414), .ZN(n19685) );
  NAND2_X1 U12890 ( .A1(n9885), .A2(n10424), .ZN(n10433) );
  AND2_X2 U12891 ( .A1(n9885), .A2(n10496), .ZN(n13719) );
  AND2_X2 U12892 ( .A1(n10421), .A2(n10422), .ZN(n9885) );
  OAI21_X2 U12893 ( .B1(n14171), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9707), 
        .ZN(n9886) );
  NAND2_X2 U12895 ( .A1(n9887), .A2(n10666), .ZN(n10691) );
  NAND2_X1 U12896 ( .A1(n9654), .A2(n9603), .ZN(n9890) );
  NOR2_X2 U12897 ( .A1(n18360), .A2(n16873), .ZN(n18268) );
  NAND2_X2 U12898 ( .A1(n18462), .A2(n16835), .ZN(n18360) );
  OR2_X2 U12899 ( .A1(n11515), .A2(n11514), .ZN(n18899) );
  NAND2_X2 U12900 ( .A1(n19301), .A2(n19469), .ZN(n17257) );
  NAND2_X2 U12901 ( .A1(n18773), .A2(n13807), .ZN(n19295) );
  AND2_X2 U12902 ( .A1(n18773), .A2(n13916), .ZN(n19298) );
  INV_X2 U12903 ( .A(n16942), .ZN(n17867) );
  AND2_X2 U12904 ( .A1(n9897), .A2(n9896), .ZN(n16902) );
  INV_X2 U12905 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9896) );
  NAND2_X2 U12906 ( .A1(n16902), .A2(n11258), .ZN(n17943) );
  NOR2_X1 U12907 ( .A1(n9899), .A2(n9713), .ZN(n9898) );
  OAI21_X1 U12908 ( .B1(n17950), .B2(n17909), .A(n11268), .ZN(n9899) );
  NAND3_X1 U12909 ( .A1(n11271), .A2(n11269), .A3(n11270), .ZN(n9915) );
  NAND3_X1 U12910 ( .A1(n11274), .A2(n11272), .A3(n11275), .ZN(n9916) );
  NAND2_X1 U12911 ( .A1(n18501), .A2(n9917), .ZN(n9919) );
  XNOR2_X2 U12912 ( .A(n11377), .B(n11375), .ZN(n18501) );
  OAI21_X2 U12913 ( .B1(n16734), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11404), .ZN(n11405) );
  INV_X2 U12914 ( .A(n15098), .ZN(n15049) );
  NAND2_X2 U12915 ( .A1(n10691), .A2(n10690), .ZN(n15098) );
  NAND2_X1 U12916 ( .A1(n15049), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9987) );
  NAND2_X1 U12917 ( .A1(n10729), .A2(n9939), .ZN(n9938) );
  NAND3_X1 U12918 ( .A1(n14109), .A2(n9943), .A3(n9721), .ZN(n9940) );
  NAND3_X1 U12919 ( .A1(n10017), .A2(n12636), .A3(n10016), .ZN(n16211) );
  NAND2_X1 U12920 ( .A1(n9952), .A2(n11811), .ZN(n12398) );
  NAND2_X2 U12921 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  NAND2_X2 U12922 ( .A1(n9950), .A2(n11798), .ZN(n12400) );
  AND2_X2 U12923 ( .A1(n11799), .A2(n10307), .ZN(n9950) );
  INV_X1 U12924 ( .A(n16486), .ZN(n16516) );
  AND2_X2 U12925 ( .A1(n12411), .A2(n12413), .ZN(n19718) );
  AND2_X2 U12926 ( .A1(n13785), .A2(n16572), .ZN(n12411) );
  INV_X1 U12927 ( .A(n13865), .ZN(n13785) );
  NAND2_X2 U12928 ( .A1(n12742), .A2(n9660), .ZN(n16044) );
  NAND2_X1 U12929 ( .A1(n12398), .A2(n11812), .ZN(n10201) );
  OAI211_X1 U12930 ( .C1(n16253), .C2(n16281), .A(n9954), .B(n9953), .ZN(
        P2_U2986) );
  OAI21_X2 U12931 ( .B1(n16020), .B2(n16019), .A(n16018), .ZN(n9955) );
  INV_X1 U12932 ( .A(n12610), .ZN(n12640) );
  NAND2_X1 U12933 ( .A1(n9959), .A2(n12481), .ZN(n9958) );
  NAND2_X1 U12934 ( .A1(n19718), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10081) );
  NAND2_X2 U12935 ( .A1(n16113), .A2(n12740), .ZN(n14260) );
  NAND3_X1 U12936 ( .A1(n14289), .A2(n9971), .A3(n19636), .ZN(n9964) );
  NAND2_X2 U12937 ( .A1(n9998), .A2(n9997), .ZN(n9965) );
  CLKBUF_X1 U12938 ( .A(n11909), .Z(n9983) );
  AND2_X2 U12939 ( .A1(n11909), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U12940 ( .A1(n14166), .A2(n20351), .ZN(n10569) );
  NAND2_X2 U12941 ( .A1(n10516), .A2(n10515), .ZN(n14167) );
  NAND2_X1 U12942 ( .A1(n15089), .A2(n9987), .ZN(n15054) );
  NAND2_X1 U12943 ( .A1(n14964), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15089) );
  AND2_X2 U12944 ( .A1(n13664), .A2(n20649), .ZN(n13658) );
  AND2_X2 U12945 ( .A1(n9989), .A2(n15361), .ZN(n10446) );
  AND2_X2 U12946 ( .A1(n10100), .A2(n9989), .ZN(n10555) );
  NAND3_X1 U12947 ( .A1(n9993), .A2(n10640), .A3(n13715), .ZN(n9992) );
  AND4_X2 U12948 ( .A1(n12420), .A2(n12410), .A3(n12417), .A4(n12418), .ZN(
        n9997) );
  AND4_X2 U12949 ( .A1(n12419), .A2(n12409), .A3(n12408), .A4(n12407), .ZN(
        n9998) );
  NAND2_X2 U12950 ( .A1(n12742), .A2(n10002), .ZN(n14369) );
  NAND2_X1 U12951 ( .A1(n12634), .A2(n15725), .ZN(n10008) );
  XNOR2_X2 U12952 ( .A(n12481), .B(n12630), .ZN(n12634) );
  NAND2_X1 U12953 ( .A1(n10008), .A2(n10009), .ZN(n12468) );
  NAND2_X1 U12954 ( .A1(n11784), .A2(n11787), .ZN(n11799) );
  NAND2_X2 U12955 ( .A1(n11805), .A2(n10010), .ZN(n11784) );
  AND3_X2 U12956 ( .A1(n11750), .A2(n11749), .A3(n11751), .ZN(n11805) );
  NAND3_X1 U12957 ( .A1(n12633), .A2(n13460), .A3(n13459), .ZN(n10016) );
  NAND2_X1 U12958 ( .A1(n12631), .A2(n10067), .ZN(n10013) );
  NAND2_X1 U12959 ( .A1(n10014), .A2(n10067), .ZN(n10015) );
  NAND3_X1 U12960 ( .A1(n10015), .A2(n12637), .A3(n12638), .ZN(n10017) );
  NAND2_X2 U12961 ( .A1(n10020), .A2(n10019), .ZN(n12042) );
  NAND2_X1 U12962 ( .A1(n18011), .A2(n9768), .ZN(n17998) );
  NOR2_X1 U12963 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  INV_X1 U12964 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11253) );
  OR2_X2 U12965 ( .A1(n10035), .A2(n11444), .ZN(n18031) );
  NAND3_X1 U12966 ( .A1(n10038), .A2(n11437), .A3(n10036), .ZN(n10035) );
  NAND2_X1 U12967 ( .A1(n11658), .A2(n13875), .ZN(n10040) );
  NAND2_X1 U12968 ( .A1(n11664), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10039) );
  NAND2_X2 U12969 ( .A1(n10040), .A2(n10039), .ZN(n16558) );
  NAND3_X1 U12970 ( .A1(n10294), .A2(n11653), .A3(n11652), .ZN(n10041) );
  NAND3_X1 U12971 ( .A1(n11647), .A2(n11649), .A3(n11648), .ZN(n10042) );
  NAND2_X1 U12972 ( .A1(n10047), .A2(n15738), .ZN(n10045) );
  NAND2_X1 U12973 ( .A1(n16158), .A2(n10048), .ZN(n10052) );
  INV_X1 U12974 ( .A(n10677), .ZN(n10058) );
  NAND2_X1 U12975 ( .A1(n9706), .A2(n11748), .ZN(n11749) );
  NAND2_X1 U12976 ( .A1(n16239), .A2(n19660), .ZN(n10067) );
  NAND2_X1 U12977 ( .A1(n19934), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10074) );
  NAND2_X1 U12978 ( .A1(n12458), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10082) );
  NAND2_X1 U12979 ( .A1(n16529), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10080) );
  AND4_X2 U12980 ( .A1(n10081), .A2(n12424), .A3(n10082), .A4(n10080), .ZN(
        n10068) );
  NAND3_X1 U12981 ( .A1(n10074), .A2(n12423), .A3(n10083), .ZN(n10071) );
  NOR2_X2 U12982 ( .A1(n12608), .A2(n10091), .ZN(n12944) );
  NAND2_X2 U12983 ( .A1(n10175), .A2(n12592), .ZN(n12658) );
  NAND3_X1 U12984 ( .A1(n10094), .A2(n16061), .A3(n10095), .ZN(n13251) );
  NAND2_X1 U12985 ( .A1(n14260), .A2(n10099), .ZN(n10094) );
  NOR2_X1 U12986 ( .A1(n14260), .A2(n10096), .ZN(n14288) );
  INV_X1 U12987 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10099) );
  AND2_X2 U12988 ( .A1(n10100), .A2(n14273), .ZN(n10525) );
  AND2_X4 U12989 ( .A1(n10100), .A2(n14272), .ZN(n13414) );
  AND2_X2 U12990 ( .A1(n10316), .A2(n10100), .ZN(n10530) );
  NAND2_X1 U12991 ( .A1(n10103), .A2(n10104), .ZN(n10793) );
  NAND2_X1 U12992 ( .A1(n14479), .A2(n14481), .ZN(n14466) );
  AOI21_X1 U12993 ( .B1(n14479), .B2(n10108), .A(n10114), .ZN(n10113) );
  NOR2_X2 U12994 ( .A1(n14466), .A2(n14468), .ZN(n14467) );
  INV_X1 U12995 ( .A(n14728), .ZN(n10119) );
  NAND2_X1 U12996 ( .A1(n14542), .A2(n9751), .ZN(n14496) );
  INV_X1 U12997 ( .A(n14496), .ZN(n13346) );
  OAI211_X1 U12998 ( .C1(n10135), .C2(n18263), .A(n17351), .B(n17558), .ZN(
        n17352) );
  NAND2_X1 U12999 ( .A1(n10140), .A2(n10136), .ZN(n18301) );
  INV_X1 U13000 ( .A(n10305), .ZN(n10143) );
  INV_X2 U13001 ( .A(n12902), .ZN(n17508) );
  INV_X1 U13002 ( .A(n18299), .ZN(n10159) );
  INV_X1 U13003 ( .A(n10161), .ZN(n12619) );
  NOR2_X2 U13004 ( .A1(n11405), .A2(n16854), .ZN(n16724) );
  NOR2_X1 U13005 ( .A1(n12551), .A2(n12364), .ZN(n12572) );
  OAI21_X2 U13006 ( .B1(n12551), .B2(n10164), .A(n10162), .ZN(n12382) );
  NAND3_X1 U13007 ( .A1(n12705), .A2(n12704), .A3(n12391), .ZN(n10175) );
  AND2_X2 U13008 ( .A1(n16909), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11259) );
  OAI21_X1 U13009 ( .B1(n12818), .B2(n15683), .A(n10180), .ZN(n15460) );
  NAND2_X1 U13010 ( .A1(n12828), .A2(n10183), .ZN(n12852) );
  NAND2_X1 U13011 ( .A1(n12715), .A2(n9765), .ZN(n12755) );
  NAND2_X1 U13012 ( .A1(n12813), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12812) );
  NOR2_X2 U13013 ( .A1(n12809), .A2(n12808), .ZN(n12813) );
  INV_X1 U13014 ( .A(n15793), .ZN(n10200) );
  NAND2_X1 U13015 ( .A1(n15798), .A2(n15800), .ZN(n15799) );
  NAND2_X2 U13016 ( .A1(n10201), .A2(n11813), .ZN(n12396) );
  INV_X1 U13017 ( .A(n14010), .ZN(n10204) );
  NAND2_X1 U13018 ( .A1(n13019), .A2(n9752), .ZN(n15837) );
  NAND3_X1 U13019 ( .A1(n11823), .A2(n10207), .A3(n13880), .ZN(n13879) );
  NOR2_X2 U13020 ( .A1(n9628), .A2(n10210), .ZN(n12744) );
  INV_X1 U13021 ( .A(n12869), .ZN(n10215) );
  NOR2_X1 U13022 ( .A1(n9662), .A2(n10217), .ZN(n12676) );
  NOR2_X1 U13023 ( .A1(n9662), .A2(n15457), .ZN(n15456) );
  INV_X1 U13024 ( .A(n12665), .ZN(n10220) );
  NAND2_X1 U13025 ( .A1(n15739), .A2(n9629), .ZN(n10226) );
  NAND2_X1 U13026 ( .A1(n10226), .A2(n10228), .ZN(n10230) );
  NOR2_X4 U13027 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14272) );
  AND2_X2 U13028 ( .A1(n14272), .A2(n15365), .ZN(n10532) );
  NAND3_X1 U13029 ( .A1(n10244), .A2(n20649), .A3(n13664), .ZN(n10243) );
  OAI21_X2 U13030 ( .B1(n10782), .B2(n10474), .A(n10246), .ZN(n10622) );
  NAND2_X1 U13031 ( .A1(n10641), .A2(n10642), .ZN(n10805) );
  NAND2_X1 U13032 ( .A1(n11774), .A2(n11813), .ZN(n12397) );
  NAND3_X1 U13033 ( .A1(n10253), .A2(n11769), .A3(n9633), .ZN(n11772) );
  NAND2_X1 U13034 ( .A1(n10258), .A2(n10260), .ZN(n16185) );
  INV_X1 U13035 ( .A(n16044), .ZN(n10262) );
  AOI21_X1 U13036 ( .B1(n20037), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n11951), .ZN(n10265) );
  NAND2_X1 U13037 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10266) );
  AND2_X2 U13038 ( .A1(n12416), .A2(n12406), .ZN(n12452) );
  AND2_X2 U13039 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13861) );
  AND2_X4 U13040 ( .A1(n13861), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13082) );
  AOI21_X1 U13041 ( .B1(n16089), .B2(n16090), .A(n12728), .ZN(n14252) );
  OAI21_X1 U13042 ( .B1(n16089), .B2(n10282), .A(n10279), .ZN(n12867) );
  NOR2_X1 U13043 ( .A1(n13251), .A2(n19668), .ZN(n13263) );
  NAND2_X1 U13044 ( .A1(n12761), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12763) );
  AOI21_X1 U13045 ( .B1(n14357), .B2(n20544), .A(n14356), .ZN(n14358) );
  NAND2_X1 U13046 ( .A1(n20722), .A2(n10506), .ZN(n20658) );
  NAND2_X1 U13047 ( .A1(n14507), .A2(n11156), .ZN(n14494) );
  OAI21_X1 U13048 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n10514), .A(
        n10513), .ZN(n10515) );
  OAI21_X1 U13049 ( .B1(n12720), .B2(n16015), .A(n12719), .ZN(n12721) );
  INV_X1 U13050 ( .A(n17508), .ZN(n17519) );
  INV_X1 U13051 ( .A(n12800), .ZN(n12805) );
  NAND2_X1 U13052 ( .A1(n12800), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12809) );
  AND2_X2 U13053 ( .A1(n10322), .A2(n14273), .ZN(n10466) );
  AOI22_X1 U13054 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U13055 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10379) );
  AOI22_X1 U13056 ( .A1(n10312), .A2(n10419), .B1(n10420), .B2(n14429), .ZN(
        n10421) );
  AOI21_X1 U13057 ( .B1(n13248), .B2(n19542), .A(n12848), .ZN(n12849) );
  XNOR2_X1 U13058 ( .A(n14329), .B(n14328), .ZN(n14359) );
  OR2_X1 U13059 ( .A1(n10509), .A2(n10508), .ZN(n10510) );
  AOI22_X1 U13060 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U13061 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U13062 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U13063 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11651) );
  INV_X1 U13064 ( .A(n19559), .ZN(n15683) );
  AND2_X2 U13065 ( .A1(n16517), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11659) );
  INV_X1 U13066 ( .A(n12052), .ZN(n12279) );
  AND2_X1 U13067 ( .A1(n16500), .A2(n16499), .ZN(n20101) );
  OR2_X1 U13068 ( .A1(n15720), .A2(n15719), .ZN(P2_U2848) );
  OR2_X1 U13069 ( .A1(n15710), .A2(n15709), .ZN(P2_U2847) );
  INV_X1 U13070 ( .A(n17281), .ZN(n12923) );
  NAND2_X1 U13071 ( .A1(n17369), .A2(n18289), .ZN(n17370) );
  NOR2_X1 U13072 ( .A1(n20963), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10290) );
  AND2_X1 U13073 ( .A1(n14286), .A2(n14285), .ZN(n10293) );
  INV_X1 U13074 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12766) );
  AOI21_X1 U13075 ( .B1(n12368), .B2(n12365), .A(n12383), .ZN(n12369) );
  AND3_X1 U13076 ( .A1(n11651), .A2(n13875), .A3(n11650), .ZN(n10294) );
  AND3_X1 U13077 ( .A1(n11679), .A2(n13875), .A3(n11678), .ZN(n10295) );
  AND2_X1 U13078 ( .A1(n16104), .A2(n16101), .ZN(n10296) );
  AND3_X1 U13079 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10298) );
  AND3_X1 U13080 ( .A1(n14403), .A2(n14408), .A3(n14402), .ZN(n10299) );
  OR2_X1 U13081 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10300) );
  INV_X1 U13082 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12649) );
  XNOR2_X1 U13083 ( .A(n12398), .B(n12397), .ZN(n12403) );
  OR2_X1 U13084 ( .A1(n17430), .A2(n18363), .ZN(n10301) );
  OR2_X1 U13085 ( .A1(n13539), .A2(n15806), .ZN(n16253) );
  INV_X1 U13086 ( .A(n16253), .ZN(n19636) );
  NAND2_X1 U13087 ( .A1(n10895), .A2(n10894), .ZN(n10303) );
  INV_X1 U13088 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16107) );
  INV_X1 U13089 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14328) );
  INV_X1 U13090 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18865) );
  INV_X2 U13091 ( .A(n17985), .ZN(n17980) );
  INV_X1 U13092 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10709) );
  OR2_X1 U13093 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10304) );
  AND2_X1 U13094 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10305) );
  INV_X1 U13095 ( .A(n19555), .ZN(n12854) );
  INV_X1 U13096 ( .A(n10973), .ZN(n10983) );
  AND2_X2 U13097 ( .A1(n15151), .A2(n11238), .ZN(n17105) );
  AND4_X1 U13098 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n10306) );
  INV_X1 U13099 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n21437) );
  INV_X1 U13100 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16142) );
  NAND2_X1 U13101 ( .A1(n12392), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10307) );
  INV_X1 U13102 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17478) );
  OR2_X1 U13103 ( .A1(n12249), .A2(n12248), .ZN(n14011) );
  INV_X1 U13104 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19311) );
  NOR2_X1 U13105 ( .A1(n13792), .A2(n17079), .ZN(n20518) );
  INV_X2 U13106 ( .A(n11488), .ZN(n17872) );
  AND2_X1 U13107 ( .A1(n16667), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10308) );
  INV_X1 U13108 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10708) );
  INV_X2 U13109 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21246) );
  INV_X1 U13110 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15379) );
  INV_X1 U13111 ( .A(n11945), .ZN(n11947) );
  INV_X1 U13112 ( .A(n12853), .ZN(n12828) );
  INV_X1 U13113 ( .A(n11814), .ZN(n11824) );
  INV_X1 U13114 ( .A(n20509), .ZN(n13985) );
  OR2_X1 U13115 ( .A1(n18189), .A2(n13916), .ZN(n10309) );
  INV_X1 U13117 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19452) );
  AND4_X1 U13118 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n10310) );
  AND4_X1 U13119 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10311) );
  OR2_X1 U13120 ( .A1(n15681), .A2(n15680), .ZN(P2_U2845) );
  AND2_X1 U13121 ( .A1(n10441), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10411) );
  AND2_X1 U13122 ( .A1(n10582), .A2(n10581), .ZN(n10639) );
  INV_X1 U13123 ( .A(n10423), .ZN(n10412) );
  INV_X1 U13124 ( .A(n11593), .ZN(n11289) );
  AND2_X1 U13125 ( .A1(n21084), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10733) );
  INV_X1 U13126 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13268) );
  INV_X1 U13127 ( .A(n11157), .ZN(n11158) );
  INV_X1 U13128 ( .A(n10940), .ZN(n10942) );
  NOR2_X1 U13129 ( .A1(n20649), .A2(n21246), .ZN(n10783) );
  NAND2_X1 U13130 ( .A1(n10445), .A2(n10597), .ZN(n10423) );
  AOI22_X1 U13131 ( .A1(n10532), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10402), .ZN(n10404) );
  AOI22_X1 U13132 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10338) );
  INV_X1 U13133 ( .A(n10610), .ZN(n10507) );
  INV_X1 U13134 ( .A(n12479), .ZN(n12353) );
  AOI21_X1 U13135 ( .B1(n11723), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n11642), .ZN(n11649) );
  INV_X1 U13136 ( .A(n12024), .ZN(n12303) );
  AOI21_X1 U13137 ( .B1(n17071), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10753), .ZN(n10763) );
  NAND2_X1 U13138 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10375) );
  INV_X1 U13139 ( .A(n11140), .ZN(n10995) );
  INV_X1 U13140 ( .A(n20410), .ZN(n13281) );
  INV_X1 U13141 ( .A(n14168), .ZN(n10548) );
  INV_X1 U13142 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17071) );
  INV_X1 U13143 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15675) );
  NOR2_X1 U13144 ( .A1(n13163), .A2(n12975), .ZN(n12976) );
  NAND2_X1 U13145 ( .A1(n15806), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12956) );
  AND3_X1 U13146 ( .A1(n12084), .A2(n12083), .A3(n12082), .ZN(n15740) );
  INV_X1 U13147 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16980) );
  INV_X1 U13148 ( .A(n11618), .ZN(n11619) );
  AND2_X1 U13149 ( .A1(n18252), .A2(n11403), .ZN(n11404) );
  INV_X1 U13150 ( .A(n11537), .ZN(n11538) );
  AOI221_X1 U13151 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10763), 
        .C1(n15392), .C2(n10763), .A(n10762), .ZN(n13372) );
  AND4_X1 U13152 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10387) );
  INV_X1 U13153 ( .A(n13384), .ZN(n13380) );
  AND2_X1 U13154 ( .A1(n11155), .A2(n14508), .ZN(n11156) );
  AND4_X1 U13155 ( .A1(n14643), .A2(n14628), .A3(n14627), .A4(n14670), .ZN(
        n10993) );
  INV_X1 U13156 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14662) );
  NAND2_X1 U13157 ( .A1(n10874), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10888) );
  NOR2_X1 U13158 ( .A1(n9623), .A2(n15162), .ZN(n10713) );
  NAND2_X1 U13159 ( .A1(n10552), .A2(n10551), .ZN(n21030) );
  INV_X1 U13160 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10743) );
  INV_X1 U13161 ( .A(n10609), .ZN(n10616) );
  OR2_X1 U13162 ( .A1(n11957), .A2(n11956), .ZN(n11959) );
  AND2_X1 U13163 ( .A1(n11888), .A2(n15494), .ZN(n14365) );
  OR2_X1 U13164 ( .A1(n12156), .A2(n12155), .ZN(n13991) );
  OR2_X1 U13165 ( .A1(n13481), .A2(n13986), .ZN(n13479) );
  INV_X1 U13166 ( .A(n13749), .ZN(n12160) );
  AND3_X1 U13167 ( .A1(n12089), .A2(n12088), .A3(n12087), .ZN(n15995) );
  NAND2_X1 U13168 ( .A1(n12599), .A2(n9691), .ZN(n12606) );
  AND2_X1 U13169 ( .A1(n11886), .A2(n15524), .ZN(n15509) );
  OR2_X1 U13170 ( .A1(n19514), .A2(n12354), .ZN(n12555) );
  NOR2_X1 U13171 ( .A1(n16204), .A2(n16160), .ZN(n16206) );
  NAND2_X1 U13172 ( .A1(n19643), .A2(n12968), .ZN(n12960) );
  NAND2_X1 U13173 ( .A1(n15425), .A2(n11964), .ZN(n11965) );
  INV_X1 U13174 ( .A(n11509), .ZN(n17918) );
  INV_X1 U13175 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17711) );
  NAND2_X1 U13176 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18351) );
  AND2_X1 U13177 ( .A1(n18242), .A2(n16844), .ZN(n16846) );
  OR2_X1 U13178 ( .A1(n18660), .A2(n18627), .ZN(n18286) );
  INV_X1 U13179 ( .A(n18723), .ZN(n18661) );
  OR3_X1 U13180 ( .A1(n11452), .A2(n11451), .A3(n11450), .ZN(n11460) );
  OR2_X1 U13181 ( .A1(n19342), .A2(n19356), .ZN(n18872) );
  NAND2_X1 U13182 ( .A1(n11083), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U13183 ( .A1(n21246), .A2(n20900), .ZN(n13431) );
  NOR2_X1 U13184 ( .A1(n20399), .A2(n21246), .ZN(n14779) );
  AND2_X1 U13185 ( .A1(n20392), .A2(n20428), .ZN(n14798) );
  OR2_X1 U13186 ( .A1(n13354), .A2(n14483), .ZN(n13355) );
  INV_X1 U13187 ( .A(n14542), .ZN(n14554) );
  OR2_X1 U13188 ( .A1(n14537), .A2(n14552), .ZN(n14525) );
  OR3_X1 U13189 ( .A1(n15210), .A2(n15183), .A3(n15182), .ZN(n15171) );
  AND2_X1 U13190 ( .A1(n15065), .A2(n15081), .ZN(n15057) );
  AND2_X1 U13191 ( .A1(n14120), .A2(n14108), .ZN(n15367) );
  AND2_X1 U13192 ( .A1(n14170), .A2(n13729), .ZN(n21031) );
  INV_X1 U13193 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21033) );
  OR2_X1 U13194 ( .A1(n20866), .A2(n20936), .ZN(n20844) );
  OR2_X1 U13195 ( .A1(n20866), .A2(n20960), .ZN(n20852) );
  OR2_X1 U13196 ( .A1(n9622), .A2(n21093), .ZN(n20936) );
  INV_X1 U13197 ( .A(n21126), .ZN(n20960) );
  INV_X1 U13198 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21084) );
  NAND2_X1 U13199 ( .A1(n15640), .A2(n15641), .ZN(n15621) );
  AND2_X1 U13200 ( .A1(n12255), .A2(n12254), .ZN(n15637) );
  NAND2_X1 U13201 ( .A1(n13539), .A2(n12679), .ZN(n16237) );
  INV_X1 U13202 ( .A(n19648), .ZN(n19665) );
  AND2_X1 U13203 ( .A1(n19692), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19872) );
  OR2_X1 U13204 ( .A1(n20323), .A2(n20308), .ZN(n19942) );
  OR2_X1 U13205 ( .A1(n20323), .A2(n19782), .ZN(n20304) );
  NAND2_X1 U13206 ( .A1(n17152), .A2(n17153), .ZN(n16500) );
  INV_X1 U13207 ( .A(n16553), .ZN(n16565) );
  NOR2_X1 U13208 ( .A1(n18278), .A2(n12907), .ZN(n12910) );
  NOR2_X1 U13209 ( .A1(n19486), .A2(n18873), .ZN(n12928) );
  NOR2_X1 U13210 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16656), .ZN(n17562) );
  INV_X1 U13211 ( .A(n11488), .ZN(n17894) );
  INV_X1 U13212 ( .A(n18369), .ZN(n18367) );
  NAND2_X1 U13213 ( .A1(n18547), .A2(n18396), .ZN(n18277) );
  INV_X1 U13214 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18339) );
  NAND2_X1 U13215 ( .A1(n11333), .A2(n11605), .ZN(n16830) );
  INV_X1 U13216 ( .A(n16835), .ZN(n16850) );
  AND2_X1 U13217 ( .A1(n18386), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18663) );
  OR2_X1 U13218 ( .A1(n19295), .A2(n18104), .ZN(n18723) );
  INV_X1 U13219 ( .A(n19158), .ZN(n19135) );
  AND2_X1 U13220 ( .A1(n13449), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14866)
         );
  XNOR2_X1 U13221 ( .A(n13381), .B(n14314), .ZN(n14409) );
  INV_X1 U13222 ( .A(n14798), .ZN(n20397) );
  AND2_X1 U13223 ( .A1(n14409), .A2(n13382), .ZN(n20426) );
  AND2_X1 U13224 ( .A1(n10946), .A2(n10945), .ZN(n14643) );
  AND2_X1 U13225 ( .A1(n14932), .A2(n14444), .ZN(n14431) );
  INV_X1 U13226 ( .A(n14915), .ZN(n14905) );
  AND2_X1 U13227 ( .A1(n13790), .A2(n17058), .ZN(n13791) );
  NAND2_X1 U13228 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  AND2_X1 U13229 ( .A1(n11053), .A2(n11052), .ZN(n14528) );
  NAND2_X1 U13230 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n10827), .ZN(
        n10856) );
  NAND2_X1 U13231 ( .A1(n10821), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10826) );
  INV_X1 U13232 ( .A(n17105), .ZN(n15112) );
  AND2_X1 U13233 ( .A1(n20546), .A2(n14127), .ZN(n20553) );
  AND2_X1 U13234 ( .A1(n13719), .A2(n10431), .ZN(n17060) );
  NOR2_X1 U13235 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21278) );
  NAND2_X1 U13236 ( .A1(n14184), .A2(n14183), .ZN(n20654) );
  AND2_X1 U13237 ( .A1(n15413), .A2(n14162), .ZN(n20727) );
  OAI21_X1 U13238 ( .B1(n20698), .B2(n20697), .A(n20696), .ZN(n20715) );
  INV_X1 U13239 ( .A(n20732), .ZN(n20749) );
  AND2_X1 U13240 ( .A1(n20727), .A2(n20993), .ZN(n20784) );
  INV_X1 U13241 ( .A(n20866), .ZN(n20753) );
  INV_X1 U13242 ( .A(n20844), .ZN(n20854) );
  INV_X1 U13243 ( .A(n20852), .ZN(n20889) );
  INV_X1 U13244 ( .A(n20904), .ZN(n20924) );
  OAI21_X1 U13245 ( .B1(n20935), .B2(n20934), .A(n21182), .ZN(n20956) );
  NOR2_X2 U13246 ( .A1(n21004), .A2(n20936), .ZN(n20988) );
  NOR2_X2 U13247 ( .A1(n21004), .A2(n20960), .ZN(n21025) );
  INV_X1 U13248 ( .A(n21043), .ZN(n21078) );
  NOR2_X2 U13249 ( .A1(n21094), .A2(n21093), .ZN(n21167) );
  INV_X1 U13250 ( .A(n21034), .ZN(n21176) );
  AND2_X1 U13251 ( .A1(n20653), .A2(n20614), .ZN(n21207) );
  AND2_X1 U13252 ( .A1(n10419), .A2(n20648), .ZN(n21226) );
  INV_X1 U13253 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21251) );
  NAND2_X1 U13254 ( .A1(n20145), .A2(n20318), .ZN(n20313) );
  INV_X1 U13255 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20145) );
  OR2_X1 U13256 ( .A1(n15434), .A2(n12837), .ZN(n19549) );
  INV_X1 U13257 ( .A(n19549), .ZN(n19532) );
  INV_X1 U13258 ( .A(n12327), .ZN(n19553) );
  INV_X1 U13259 ( .A(n19551), .ZN(n19542) );
  INV_X1 U13260 ( .A(n19571), .ZN(n15883) );
  INV_X1 U13261 ( .A(n13220), .ZN(n13221) );
  INV_X1 U13262 ( .A(n19586), .ZN(n16010) );
  INV_X1 U13263 ( .A(n16013), .ZN(n19582) );
  INV_X1 U13264 ( .A(n13596), .ZN(n19626) );
  AND2_X1 U13265 ( .A1(n13563), .A2(n12004), .ZN(n19630) );
  INV_X1 U13266 ( .A(n16237), .ZN(n19634) );
  INV_X1 U13267 ( .A(n13261), .ZN(n13262) );
  CLKBUF_X1 U13268 ( .A(n16211), .Z(n16212) );
  NOR2_X1 U13269 ( .A1(n19840), .A2(n19942), .ZN(n19711) );
  NAND2_X1 U13270 ( .A1(n19723), .A2(n20152), .ZN(n19740) );
  OAI211_X1 U13271 ( .C1(n19754), .C2(n19753), .A(n20152), .B(n19752), .ZN(
        n19771) );
  NOR2_X1 U13272 ( .A1(n19881), .A2(n20304), .ZN(n19784) );
  INV_X1 U13273 ( .A(n19783), .ZN(n19833) );
  OAI21_X1 U13274 ( .B1(n19841), .B2(n19973), .A(n19839), .ZN(n19865) );
  OAI21_X1 U13275 ( .B1(n19981), .B2(n19980), .A(n20152), .ZN(n19998) );
  NOR2_X1 U13276 ( .A1(n20094), .A2(n20304), .ZN(n20019) );
  OAI211_X1 U13277 ( .C1(n20058), .C2(n20043), .A(n20042), .B(n20152), .ZN(
        n20060) );
  NOR2_X1 U13278 ( .A1(n20069), .A2(n20065), .ZN(n20088) );
  OAI22_X1 U13279 ( .A1(n20620), .A2(n16564), .B1(n18890), .B2(n16563), .ZN(
        n20123) );
  AND2_X1 U13280 ( .A1(n16566), .A2(n16565), .ZN(n20199) );
  INV_X1 U13281 ( .A(n17160), .ZN(n16626) );
  INV_X1 U13282 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20231) );
  NOR2_X1 U13283 ( .A1(n19293), .A2(n18188), .ZN(n19487) );
  NAND2_X1 U13284 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  NOR2_X1 U13285 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17308), .ZN(n17296) );
  NOR2_X1 U13286 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17329), .ZN(n17316) );
  NOR2_X1 U13287 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17350), .ZN(n17335) );
  NOR2_X1 U13288 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17368), .ZN(n17356) );
  NOR2_X1 U13289 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17456), .ZN(n17446) );
  NAND2_X1 U13290 ( .A1(n19338), .A2(n12928), .ZN(n17599) );
  OAI211_X1 U13291 ( .C1(n19349), .C2(n19350), .A(n12931), .B(n19486), .ZN(
        n17573) );
  INV_X1 U13292 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16657) );
  INV_X1 U13293 ( .A(n17573), .ZN(n17593) );
  AND3_X1 U13294 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17662), .ZN(n17651) );
  NOR2_X1 U13295 ( .A1(n17457), .A2(n17032), .ZN(n17844) );
  INV_X1 U13296 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17564) );
  INV_X1 U13297 ( .A(n17981), .ZN(n17984) );
  NOR2_X2 U13298 ( .A1(n11473), .A2(n11472), .ZN(n18896) );
  NOR2_X1 U13299 ( .A1(n18031), .A2(n18065), .ZN(n18059) );
  INV_X1 U13300 ( .A(n18094), .ZN(n18095) );
  NAND2_X1 U13301 ( .A1(n19294), .A2(n19469), .ZN(n18188) );
  AND2_X1 U13302 ( .A1(n18748), .A2(n18615), .ZN(n18622) );
  AND2_X1 U13303 ( .A1(n18663), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16835) );
  NOR2_X1 U13304 ( .A1(n16851), .A2(n18834), .ZN(n18742) );
  NOR2_X2 U13305 ( .A1(n16772), .A2(n16771), .ZN(n18760) );
  INV_X1 U13306 ( .A(n16772), .ZN(n18843) );
  INV_X1 U13307 ( .A(n18914), .ZN(n19216) );
  NOR2_X1 U13308 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19452), .ZN(
        n19342) );
  INV_X1 U13309 ( .A(n19037), .ZN(n19042) );
  INV_X1 U13310 ( .A(n19117), .ZN(n19131) );
  INV_X1 U13311 ( .A(n21311), .ZN(n19224) );
  INV_X1 U13312 ( .A(n18906), .ZN(n19188) );
  INV_X1 U13313 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n16879) );
  AND2_X1 U13314 ( .A1(n19434), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19379) );
  INV_X1 U13315 ( .A(n14866), .ZN(n14430) );
  NAND2_X1 U13316 ( .A1(n13241), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16533)
         );
  INV_X1 U13317 ( .A(U212), .ZN(n17203) );
  INV_X1 U13318 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20900) );
  OR2_X2 U13319 ( .A1(n14409), .A2(n13434), .ZN(n14772) );
  INV_X1 U13320 ( .A(n20411), .ZN(n20442) );
  INV_X2 U13321 ( .A(n20449), .ZN(n14838) );
  NAND2_X1 U13322 ( .A1(n13831), .A2(n14932), .ZN(n14931) );
  OR2_X1 U13323 ( .A1(n13792), .A2(n13791), .ZN(n20484) );
  NOR2_X1 U13324 ( .A1(n9667), .A2(n13943), .ZN(n13981) );
  OR2_X1 U13325 ( .A1(n17125), .A2(n21091), .ZN(n15122) );
  INV_X1 U13326 ( .A(n20544), .ZN(n20578) );
  OR2_X1 U13327 ( .A1(n20540), .A2(n14336), .ZN(n17123) );
  INV_X1 U13328 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20586) );
  INV_X1 U13329 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15392) );
  NAND2_X1 U13330 ( .A1(n20727), .A2(n9727), .ZN(n20690) );
  AOI22_X1 U13331 ( .A1(n20693), .A2(n20697), .B1(n20964), .B2(n10290), .ZN(
        n20718) );
  AOI22_X1 U13332 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20728), .B1(n20730), 
        .B2(n20726), .ZN(n20752) );
  NAND2_X1 U13333 ( .A1(n20753), .A2(n9727), .ZN(n20818) );
  AOI22_X1 U13334 ( .A1(n20827), .A2(n20824), .B1(n21129), .B2(n10290), .ZN(
        n20858) );
  OR2_X1 U13335 ( .A1(n20866), .A2(n20859), .ZN(n20904) );
  NAND2_X1 U13336 ( .A1(n20994), .A2(n9727), .ZN(n20959) );
  AOI22_X1 U13337 ( .A1(n20965), .A2(n20970), .B1(n20964), .B2(n21128), .ZN(
        n20992) );
  NAND2_X1 U13338 ( .A1(n20994), .A2(n20993), .ZN(n21043) );
  INV_X1 U13339 ( .A(n21177), .ZN(n21046) );
  INV_X1 U13340 ( .A(n21219), .ZN(n21069) );
  NAND2_X1 U13341 ( .A1(n21089), .A2(n21093), .ZN(n21124) );
  INV_X1 U13342 ( .A(n21104), .ZN(n21205) );
  NAND2_X1 U13343 ( .A1(n21180), .A2(n21126), .ZN(n21224) );
  INV_X1 U13344 ( .A(n21120), .ZN(n21242) );
  AND2_X1 U13345 ( .A1(n21251), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n14465) );
  INV_X1 U13346 ( .A(n12689), .ZN(n13539) );
  OR2_X1 U13347 ( .A1(n15434), .A2(n12830), .ZN(n19555) );
  INV_X1 U13348 ( .A(n19554), .ZN(n19546) );
  NAND2_X1 U13349 ( .A1(n12661), .A2(n12694), .ZN(n15903) );
  NAND2_X1 U13350 ( .A1(n19586), .A2(n13230), .ZN(n15981) );
  AND2_X1 U13351 ( .A1(n16013), .A2(n15981), .ZN(n16005) );
  NAND2_X1 U13352 ( .A1(n19586), .A2(n13229), .ZN(n16013) );
  OR2_X1 U13353 ( .A1(n19625), .A2(n13683), .ZN(n19588) );
  NAND2_X1 U13354 ( .A1(n13682), .A2(n20217), .ZN(n19625) );
  INV_X1 U13355 ( .A(n19630), .ZN(n13679) );
  NAND2_X1 U13356 ( .A1(n12944), .A2(n19672), .ZN(n12653) );
  INV_X1 U13357 ( .A(n19657), .ZN(n19668) );
  INV_X1 U13358 ( .A(n19711), .ZN(n19707) );
  INV_X1 U13359 ( .A(n19708), .ZN(n19743) );
  AOI21_X1 U13360 ( .B1(n19749), .B2(n19753), .A(n19748), .ZN(n19774) );
  INV_X1 U13361 ( .A(n19784), .ZN(n19807) );
  OR2_X1 U13362 ( .A1(n19881), .A2(n20072), .ZN(n19863) );
  AND2_X1 U13363 ( .A1(n19876), .A2(n19875), .ZN(n19886) );
  INV_X1 U13364 ( .A(n19882), .ZN(n19904) );
  OAI22_X1 U13365 ( .A1(n19909), .A2(n19928), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19912), .ZN(n19932) );
  AOI21_X1 U13366 ( .B1(n19937), .B2(n19940), .A(n19936), .ZN(n19970) );
  INV_X1 U13367 ( .A(n19974), .ZN(n20001) );
  INV_X1 U13368 ( .A(n20019), .ZN(n20032) );
  INV_X1 U13369 ( .A(n20039), .ZN(n20063) );
  INV_X1 U13370 ( .A(n20064), .ZN(n20092) );
  AOI211_X2 U13371 ( .C1(n20103), .C2(n20106), .A(n20101), .B(n20100), .ZN(
        n20142) );
  INV_X1 U13372 ( .A(n20123), .ZN(n20186) );
  NOR3_X1 U13373 ( .A1(n16625), .A2(n16624), .A3(n16623), .ZN(n17154) );
  INV_X1 U13374 ( .A(n20293), .ZN(n20210) );
  OR2_X1 U13375 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19492), .ZN(n20336) );
  INV_X1 U13376 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17254) );
  NOR2_X1 U13377 ( .A1(n12941), .A2(n12940), .ZN(n12942) );
  INV_X1 U13378 ( .A(n17518), .ZN(n17598) );
  INV_X1 U13379 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18495) );
  INV_X1 U13380 ( .A(n17584), .ZN(n17605) );
  INV_X1 U13381 ( .A(n17657), .ZN(n17662) );
  NOR2_X1 U13382 ( .A1(n17384), .A2(n17737), .ZN(n17756) );
  AND2_X1 U13383 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17927), .ZN(n17906) );
  INV_X1 U13384 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17962) );
  NOR2_X1 U13385 ( .A1(n18910), .A2(n13921), .ZN(n18100) );
  NOR2_X1 U13386 ( .A1(n11317), .A2(n11316), .ZN(n18114) );
  INV_X1 U13387 ( .A(n11587), .ZN(n18119) );
  NOR2_X1 U13388 ( .A1(n18184), .A2(n18171), .ZN(n18175) );
  INV_X1 U13389 ( .A(n18171), .ZN(n18186) );
  AOI211_X1 U13390 ( .C1(n19473), .C2(n19471), .A(n18189), .B(n18188), .ZN(
        n18220) );
  INV_X1 U13391 ( .A(n18436), .ZN(n18464) );
  NAND2_X1 U13392 ( .A1(n16835), .A2(n18742), .ZN(n18659) );
  INV_X1 U13393 ( .A(n18760), .ZN(n18753) );
  OR2_X1 U13394 ( .A1(n18813), .A2(n18846), .ZN(n18839) );
  INV_X1 U13395 ( .A(n18845), .ZN(n18833) );
  INV_X1 U13396 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19475) );
  INV_X1 U13397 ( .A(n19446), .ZN(n19443) );
  INV_X1 U13398 ( .A(n14430), .ZN(n14869) );
  NOR2_X1 U13399 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13452), .ZN(n17227)
         );
  INV_X1 U13400 ( .A(n17201), .ZN(n17206) );
  OAI21_X1 U13401 ( .B1(n15161), .B2(n15151), .A(n11248), .ZN(P1_U2970) );
  NAND2_X1 U13402 ( .A1(n12723), .A2(n12722), .ZN(P2_U2987) );
  OR4_X1 U13403 ( .A1(n13469), .A2(n13468), .A3(n13467), .A4(n13466), .ZN(
        P2_U3041) );
  OAI21_X1 U13404 ( .B1(n11641), .B2(n16828), .A(n10310), .ZN(P3_U2802) );
  INV_X1 U13405 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10314) );
  INV_X1 U13406 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10315) );
  AND2_X2 U13407 ( .A1(n10429), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10316) );
  NOR2_X4 U13408 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15361) );
  AND2_X4 U13409 ( .A1(n10316), .A2(n15361), .ZN(n10461) );
  AOI22_X1 U13410 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10321) );
  AND2_X2 U13411 ( .A1(n10317), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10322) );
  AOI22_X1 U13412 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13413 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10319) );
  AND2_X2 U13414 ( .A1(n15365), .A2(n14273), .ZN(n10448) );
  AOI22_X1 U13415 ( .A1(n10446), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13416 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10330) );
  AND2_X2 U13417 ( .A1(n10322), .A2(n14272), .ZN(n10453) );
  AOI22_X1 U13418 ( .A1(n10453), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10483), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10328) );
  AND2_X2 U13419 ( .A1(n15361), .A2(n14272), .ZN(n10402) );
  NAND4_X1 U13420 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10329) );
  AOI22_X1 U13421 ( .A1(n10453), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10532), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13422 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13423 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13424 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13426 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13427 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10402), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13428 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13429 ( .A1(n10532), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13430 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13431 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n9616), .ZN(n10342) );
  AOI22_X1 U13432 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13433 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13434 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10402), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13435 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10346) );
  NAND2_X2 U13436 ( .A1(n10350), .A2(n10349), .ZN(n10419) );
  INV_X2 U13437 ( .A(n10419), .ZN(n10437) );
  AOI22_X1 U13438 ( .A1(n10532), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13439 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13440 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13441 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13442 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13443 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13444 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10402), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13445 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13446 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13447 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13448 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10402), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13449 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13450 ( .A1(n10532), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13451 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13452 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13453 ( .A1(n10367), .A2(n10437), .A3(n14116), .A4(n20611), .ZN(
        n13711) );
  NAND2_X1 U13454 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13455 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10370) );
  NAND2_X1 U13456 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10369) );
  NAND2_X1 U13457 ( .A1(n9626), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10368) );
  NAND2_X1 U13458 ( .A1(n10446), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13459 ( .A1(n10402), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10373) );
  NAND2_X1 U13460 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10372) );
  NAND2_X1 U13461 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10378) );
  NAND2_X1 U13462 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U13463 ( .A1(n10532), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13464 ( .A1(n10453), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10383) );
  NAND2_X1 U13465 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13466 ( .A1(n9600), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10381) );
  NAND2_X1 U13467 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10380) );
  AOI22_X1 U13468 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13469 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13470 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10402), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13471 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10388) );
  NAND4_X1 U13472 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10397) );
  AOI22_X1 U13473 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13474 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13475 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10392) );
  NAND4_X1 U13476 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10396) );
  OR2_X2 U13477 ( .A1(n10397), .A2(n10396), .ZN(n10418) );
  AOI22_X1 U13478 ( .A1(n10530), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10466), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13479 ( .A1(n10555), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13480 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9626), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13481 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10398) );
  NAND4_X1 U13482 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10408) );
  AOI22_X1 U13483 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13484 ( .A1(n9600), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10403) );
  NAND4_X1 U13485 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10407) );
  XNOR2_X1 U13486 ( .A(n13525), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13385) );
  NAND2_X1 U13487 ( .A1(n10442), .A2(n10418), .ZN(n13830) );
  INV_X1 U13488 ( .A(n13830), .ZN(n13831) );
  NAND2_X1 U13489 ( .A1(n10497), .A2(n10419), .ZN(n10435) );
  NAND2_X1 U13490 ( .A1(n13831), .A2(n10292), .ZN(n10440) );
  INV_X1 U13491 ( .A(n10420), .ZN(n10409) );
  NAND3_X2 U13492 ( .A1(n10409), .A2(n10437), .A3(n10597), .ZN(n10441) );
  NOR2_X1 U13493 ( .A1(n20611), .A2(n20351), .ZN(n10410) );
  INV_X1 U13494 ( .A(n13266), .ZN(n10413) );
  NAND2_X1 U13495 ( .A1(n10413), .A2(n10412), .ZN(n14114) );
  NAND2_X1 U13496 ( .A1(n10476), .A2(n14187), .ZN(n13662) );
  NAND2_X1 U13497 ( .A1(n10436), .A2(n10414), .ZN(n10415) );
  NAND2_X1 U13498 ( .A1(n10432), .A2(n10431), .ZN(n13721) );
  NAND4_X1 U13499 ( .A1(n14114), .A2(n13662), .A3(n10415), .A4(n13721), .ZN(
        n10434) );
  NAND2_X1 U13500 ( .A1(n10434), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U13501 ( .A1(n10441), .A2(n20611), .ZN(n10422) );
  NAND2_X1 U13502 ( .A1(n10419), .A2(n10418), .ZN(n14429) );
  NAND2_X1 U13503 ( .A1(n13661), .A2(n14187), .ZN(n10424) );
  INV_X1 U13504 ( .A(n10553), .ZN(n10425) );
  NAND2_X1 U13505 ( .A1(n10433), .A2(n10425), .ZN(n10426) );
  NAND2_X1 U13506 ( .A1(n21278), .A2(n20351), .ZN(n11241) );
  NAND2_X1 U13507 ( .A1(n10433), .A2(n14770), .ZN(n14122) );
  INV_X1 U13508 ( .A(n10434), .ZN(n10444) );
  AND2_X1 U13509 ( .A1(n10435), .A2(n20649), .ZN(n10772) );
  INV_X1 U13510 ( .A(n21278), .ZN(n15422) );
  NOR2_X1 U13511 ( .A1(n15422), .A2(n20351), .ZN(n10438) );
  NAND2_X1 U13512 ( .A1(n15378), .A2(n10437), .ZN(n14124) );
  OAI211_X1 U13513 ( .C1(n10772), .C2(n21298), .A(n10438), .B(n14124), .ZN(
        n10439) );
  NAND2_X1 U13514 ( .A1(n10442), .A2(n20611), .ZN(n10443) );
  AOI22_X1 U13515 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13516 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13517 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10450) );
  INV_X1 U13518 ( .A(n10448), .ZN(n15363) );
  INV_X2 U13519 ( .A(n15363), .ZN(n13413) );
  AOI22_X1 U13520 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13521 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10460) );
  AOI22_X1 U13522 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13523 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13524 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13525 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U13526 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10459) );
  AOI22_X1 U13527 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13414), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13528 ( .A1(n10483), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13529 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13530 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10462) );
  NAND4_X1 U13531 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10473) );
  AOI22_X1 U13532 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13533 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13534 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13535 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10468) );
  NAND4_X1 U13536 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10472) );
  MUX2_X1 U13537 ( .A(n10482), .B(n10477), .S(n10609), .Z(n10474) );
  INV_X1 U13538 ( .A(n10474), .ZN(n10475) );
  INV_X1 U13539 ( .A(n10477), .ZN(n10494) );
  INV_X1 U13540 ( .A(n10479), .ZN(n10478) );
  NAND2_X1 U13541 ( .A1(n10494), .A2(n10478), .ZN(n10481) );
  NAND2_X1 U13542 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10480) );
  AOI22_X1 U13543 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10483), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13544 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13545 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13546 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13547 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10493) );
  AOI22_X1 U13548 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13549 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13550 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13551 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10488) );
  NAND4_X1 U13552 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10492) );
  NAND2_X1 U13553 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10495) );
  NOR2_X1 U13554 ( .A1(n13661), .A2(n10476), .ZN(n10496) );
  NAND2_X2 U13555 ( .A1(n13719), .A2(n13946), .ZN(n15394) );
  NOR2_X1 U13556 ( .A1(n13824), .A2(n14429), .ZN(n10498) );
  AOI21_X1 U13557 ( .B1(n13658), .B2(n13385), .A(n14130), .ZN(n10499) );
  NAND2_X1 U13558 ( .A1(n13658), .A2(n10431), .ZN(n14111) );
  NAND3_X1 U13559 ( .A1(n15394), .A2(n10499), .A3(n14111), .ZN(n10500) );
  NAND2_X1 U13560 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10520) );
  OAI21_X1 U13561 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10520), .ZN(n20963) );
  OR2_X1 U13562 ( .A1(n17084), .A2(n21033), .ZN(n10511) );
  OAI21_X1 U13563 ( .B1(n11241), .B2(n20963), .A(n10511), .ZN(n10501) );
  INV_X1 U13564 ( .A(n10504), .ZN(n10505) );
  OR2_X2 U13565 ( .A1(n20722), .A2(n10506), .ZN(n10516) );
  INV_X1 U13566 ( .A(n10511), .ZN(n10514) );
  INV_X1 U13567 ( .A(n10512), .ZN(n10513) );
  NOR2_X1 U13568 ( .A1(n17084), .A2(n10743), .ZN(n10518) );
  INV_X1 U13569 ( .A(n10544), .ZN(n10524) );
  INV_X1 U13570 ( .A(n11241), .ZN(n10522) );
  INV_X1 U13571 ( .A(n10520), .ZN(n10519) );
  NAND2_X1 U13572 ( .A1(n10519), .A2(n10743), .ZN(n20995) );
  NAND2_X1 U13573 ( .A1(n10520), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13574 ( .A1(n20995), .A2(n10521), .ZN(n14181) );
  NAND2_X1 U13575 ( .A1(n10522), .A2(n14181), .ZN(n10543) );
  INV_X1 U13576 ( .A(n10543), .ZN(n10523) );
  AOI21_X1 U13577 ( .B1(n10524), .B2(n20351), .A(n10523), .ZN(n10547) );
  AOI22_X1 U13578 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13579 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13580 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13581 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10526) );
  NAND4_X1 U13582 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10539) );
  AOI22_X1 U13583 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13584 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13585 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13586 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13587 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10538) );
  NAND2_X1 U13588 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10540) );
  OAI21_X1 U13589 ( .B1(n10605), .B2(n10553), .A(n10540), .ZN(n10542) );
  NOR2_X1 U13590 ( .A1(n10554), .A2(n10605), .ZN(n10541) );
  XNOR2_X1 U13591 ( .A(n10542), .B(n10541), .ZN(n10546) );
  NAND3_X1 U13592 ( .A1(n14167), .A2(n14168), .A3(n20351), .ZN(n10545) );
  OAI211_X1 U13593 ( .C1(n14167), .C2(n10547), .A(n10546), .B(n10545), .ZN(
        n10601) );
  NAND2_X1 U13594 ( .A1(n10517), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10552) );
  NOR3_X1 U13595 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10743), .A3(
        n21033), .ZN(n20869) );
  NAND2_X1 U13596 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20869), .ZN(
        n20874) );
  NAND2_X1 U13597 ( .A1(n17071), .A2(n20874), .ZN(n10549) );
  NAND3_X1 U13598 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21132) );
  INV_X1 U13599 ( .A(n21132), .ZN(n21185) );
  NAND2_X1 U13600 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21185), .ZN(
        n21198) );
  NAND2_X1 U13601 ( .A1(n10549), .A2(n21198), .ZN(n20896) );
  OAI22_X1 U13602 ( .A1(n11241), .A2(n20896), .B1(n17084), .B2(n17071), .ZN(
        n10550) );
  INV_X1 U13603 ( .A(n10550), .ZN(n10551) );
  AOI22_X1 U13604 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13605 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13606 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13607 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10557) );
  NAND4_X1 U13608 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10567) );
  AOI22_X1 U13609 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13610 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13611 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13612 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10562) );
  NAND4_X1 U13613 ( .A1(n10565), .A2(n10564), .A3(n10563), .A4(n10562), .ZN(
        n10566) );
  AOI22_X1 U13614 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10757), .B1(
        n10768), .B2(n10643), .ZN(n10568) );
  NAND2_X1 U13615 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10582) );
  AOI22_X1 U13616 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13617 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n9612), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13618 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13619 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13404), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10571) );
  NAND4_X1 U13620 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10580) );
  AOI22_X1 U13621 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11184), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13622 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10531), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13623 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10467), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13624 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10575) );
  NAND4_X1 U13625 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10579) );
  NAND2_X1 U13626 ( .A1(n10768), .A2(n10645), .ZN(n10581) );
  NAND2_X1 U13627 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10594) );
  AOI22_X1 U13628 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13629 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13630 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13631 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10583) );
  NAND4_X1 U13632 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10592) );
  AOI22_X1 U13633 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13634 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13635 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13636 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10587) );
  NAND4_X1 U13637 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10591) );
  NAND2_X1 U13638 ( .A1(n10768), .A2(n10670), .ZN(n10593) );
  NAND2_X1 U13639 ( .A1(n10642), .A2(n10595), .ZN(n10596) );
  NAND2_X1 U13640 ( .A1(n10668), .A2(n10596), .ZN(n10813) );
  INV_X1 U13641 ( .A(n13715), .ZN(n14068) );
  NAND2_X1 U13642 ( .A1(n10610), .A2(n10609), .ZN(n10608) );
  NAND2_X1 U13643 ( .A1(n10608), .A2(n10605), .ZN(n10644) );
  AND2_X1 U13644 ( .A1(n10645), .A2(n10643), .ZN(n10598) );
  NAND2_X1 U13645 ( .A1(n10644), .A2(n10598), .ZN(n10669) );
  XNOR2_X1 U13646 ( .A(n10669), .B(n10670), .ZN(n10599) );
  NAND2_X1 U13647 ( .A1(n10599), .A2(n14101), .ZN(n10600) );
  OAI21_X2 U13648 ( .B1(n10813), .B2(n14068), .A(n10600), .ZN(n14094) );
  INV_X1 U13649 ( .A(n10601), .ZN(n10602) );
  NAND2_X1 U13650 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  XNOR2_X1 U13651 ( .A(n10608), .B(n10605), .ZN(n10606) );
  AND2_X1 U13652 ( .A1(n10432), .A2(n20611), .ZN(n14065) );
  AOI21_X1 U13653 ( .B1(n10606), .B2(n14101), .A(n14065), .ZN(n10607) );
  OAI21_X1 U13654 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(n10611) );
  OAI21_X1 U13655 ( .B1(n10611), .B2(n21298), .A(n10312), .ZN(n10612) );
  INV_X1 U13656 ( .A(n10612), .ZN(n10613) );
  AND2_X1 U13657 ( .A1(n10614), .A2(n10613), .ZN(n14038) );
  INV_X1 U13658 ( .A(n10615), .ZN(n10620) );
  NAND2_X1 U13659 ( .A1(n14101), .A2(n10616), .ZN(n14066) );
  INV_X1 U13660 ( .A(n14065), .ZN(n10617) );
  NAND2_X1 U13661 ( .A1(n14066), .A2(n10617), .ZN(n10621) );
  NOR2_X1 U13662 ( .A1(n10780), .A2(n10621), .ZN(n10619) );
  OAI21_X1 U13663 ( .B1(n10621), .B2(n13715), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10618) );
  AOI21_X1 U13664 ( .B1(n10620), .B2(n10619), .A(n10618), .ZN(n10624) );
  OR2_X1 U13665 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  AND2_X1 U13666 ( .A1(n10624), .A2(n10623), .ZN(n10626) );
  NAND2_X1 U13667 ( .A1(n10626), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13668 ( .A1(n14038), .A2(n10625), .ZN(n10628) );
  INV_X1 U13669 ( .A(n10626), .ZN(n14070) );
  INV_X1 U13670 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20571) );
  NAND2_X1 U13671 ( .A1(n14070), .A2(n20571), .ZN(n10627) );
  NAND2_X1 U13672 ( .A1(n10628), .A2(n10627), .ZN(n10629) );
  XNOR2_X1 U13673 ( .A(n10629), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14078) );
  NAND2_X1 U13674 ( .A1(n14079), .A2(n14078), .ZN(n14077) );
  INV_X1 U13675 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20552) );
  OR2_X1 U13676 ( .A1(n10629), .A2(n20552), .ZN(n10630) );
  AND2_X1 U13677 ( .A1(n14077), .A2(n10630), .ZN(n14059) );
  INV_X1 U13678 ( .A(n10643), .ZN(n10632) );
  XNOR2_X1 U13679 ( .A(n10644), .B(n10632), .ZN(n10633) );
  NAND2_X1 U13680 ( .A1(n10633), .A2(n14101), .ZN(n10634) );
  NAND2_X1 U13681 ( .A1(n14059), .A2(n10635), .ZN(n10638) );
  INV_X1 U13682 ( .A(n14058), .ZN(n10636) );
  INV_X1 U13683 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20539) );
  NAND2_X1 U13684 ( .A1(n10636), .A2(n20539), .ZN(n10637) );
  NAND2_X1 U13685 ( .A1(n10640), .A2(n10639), .ZN(n10641) );
  NAND2_X1 U13686 ( .A1(n10644), .A2(n10643), .ZN(n10646) );
  XNOR2_X1 U13687 ( .A(n10646), .B(n10645), .ZN(n10647) );
  NAND2_X1 U13688 ( .A1(n10647), .A2(n14101), .ZN(n10648) );
  INV_X1 U13689 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14129) );
  AND2_X1 U13690 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13691 ( .A1(n10651), .A2(n14094), .B1(n10650), .B2(n20515), .ZN(
        n10652) );
  NAND2_X1 U13692 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10665) );
  AOI22_X1 U13693 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13694 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13695 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13696 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10654) );
  NAND4_X1 U13697 ( .A1(n10657), .A2(n10656), .A3(n10655), .A4(n10654), .ZN(
        n10663) );
  AOI22_X1 U13698 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13699 ( .A1(n13410), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13700 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13701 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10658) );
  NAND4_X1 U13702 ( .A1(n10661), .A2(n10660), .A3(n10659), .A4(n10658), .ZN(
        n10662) );
  NAND2_X1 U13703 ( .A1(n10768), .A2(n10682), .ZN(n10664) );
  INV_X1 U13704 ( .A(n10667), .ZN(n10666) );
  NAND2_X1 U13705 ( .A1(n10668), .A2(n10667), .ZN(n10825) );
  NAND3_X1 U13706 ( .A1(n10691), .A2(n13715), .A3(n10825), .ZN(n10674) );
  INV_X1 U13707 ( .A(n10669), .ZN(n10671) );
  NAND2_X1 U13708 ( .A1(n10671), .A2(n10670), .ZN(n10681) );
  XNOR2_X1 U13709 ( .A(n10681), .B(n10682), .ZN(n10672) );
  NAND2_X1 U13710 ( .A1(n10672), .A2(n14101), .ZN(n10673) );
  INV_X1 U13711 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U13712 ( .A1(n17101), .A2(n17100), .ZN(n10675) );
  INV_X1 U13713 ( .A(n17101), .ZN(n10676) );
  NAND2_X1 U13714 ( .A1(n10676), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10677) );
  NAND2_X1 U13715 ( .A1(n10757), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10679) );
  NAND2_X1 U13716 ( .A1(n10768), .A2(n10684), .ZN(n10678) );
  NAND2_X1 U13717 ( .A1(n10679), .A2(n10678), .ZN(n10680) );
  INV_X1 U13718 ( .A(n10681), .ZN(n10683) );
  NAND2_X1 U13719 ( .A1(n10683), .A2(n10682), .ZN(n10693) );
  XNOR2_X1 U13720 ( .A(n10693), .B(n10684), .ZN(n10685) );
  AND2_X1 U13721 ( .A1(n10685), .A2(n14101), .ZN(n10686) );
  AOI21_X2 U13722 ( .B1(n10831), .B2(n13715), .A(n10686), .ZN(n10687) );
  INV_X1 U13723 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17114) );
  NAND2_X1 U13724 ( .A1(n10687), .A2(n17114), .ZN(n17095) );
  INV_X1 U13725 ( .A(n10687), .ZN(n10688) );
  NAND2_X1 U13726 ( .A1(n10688), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17094) );
  NOR2_X1 U13727 ( .A1(n10689), .A2(n14068), .ZN(n10690) );
  OR3_X1 U13728 ( .A1(n10693), .A2(n21298), .A3(n10692), .ZN(n10694) );
  INV_X1 U13729 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U13730 ( .A1(n14209), .A2(n10695), .ZN(n10696) );
  INV_X1 U13731 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15352) );
  INV_X1 U13732 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15316) );
  NAND2_X1 U13733 ( .A1(n15098), .A2(n15316), .ZN(n10699) );
  INV_X1 U13734 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15132) );
  NAND2_X1 U13735 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U13736 ( .B1(n15132), .B2(n14338), .A(n15098), .ZN(n10700) );
  INV_X1 U13737 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U13738 ( .A1(n14964), .A2(n10705), .ZN(n15058) );
  NAND2_X1 U13739 ( .A1(n15098), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10701) );
  NAND2_X1 U13740 ( .A1(n15058), .A2(n10701), .ZN(n15065) );
  INV_X1 U13741 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15289) );
  NAND2_X1 U13742 ( .A1(n15098), .A2(n15289), .ZN(n15081) );
  NAND2_X1 U13743 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U13744 ( .A1(n15046), .A2(n10702), .ZN(n10703) );
  INV_X1 U13745 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15309) );
  NAND2_X1 U13746 ( .A1(n15046), .A2(n15309), .ZN(n15053) );
  NOR2_X1 U13747 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15099) );
  INV_X1 U13748 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15338) );
  NAND2_X1 U13749 ( .A1(n15099), .A2(n15338), .ZN(n15048) );
  INV_X1 U13750 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15283) );
  NAND3_X1 U13751 ( .A1(n15289), .A2(n10705), .A3(n15283), .ZN(n10706) );
  XNOR2_X1 U13752 ( .A(n15098), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15038) );
  AND2_X1 U13753 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15244) );
  NAND2_X1 U13754 ( .A1(n15244), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15227) );
  INV_X1 U13755 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15011) );
  INV_X1 U13756 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U13757 ( .A1(n15011), .A2(n15246), .ZN(n10710) );
  INV_X1 U13758 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14975) );
  INV_X1 U13759 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U13760 ( .A1(n14975), .A2(n15194), .ZN(n10711) );
  AND2_X1 U13761 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15180) );
  NAND2_X1 U13762 ( .A1(n15180), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15183) );
  INV_X1 U13763 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U13764 ( .A1(n10712), .A2(n9623), .ZN(n14973) );
  AND2_X1 U13765 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15154) );
  INV_X1 U13766 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14956) );
  INV_X1 U13767 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14945) );
  NAND2_X1 U13768 ( .A1(n14956), .A2(n14945), .ZN(n15162) );
  NAND2_X1 U13769 ( .A1(n14326), .A2(n14327), .ZN(n10715) );
  XNOR2_X1 U13770 ( .A(n10715), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15161) );
  NOR2_X1 U13771 ( .A1(n20629), .A2(n20351), .ZN(n10716) );
  NAND2_X1 U13772 ( .A1(n13946), .A2(n20629), .ZN(n10721) );
  XNOR2_X1 U13773 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10732) );
  XNOR2_X1 U13774 ( .A(n10732), .B(n10733), .ZN(n13368) );
  NAND2_X1 U13775 ( .A1(n10757), .A2(n13368), .ZN(n10717) );
  NAND2_X1 U13776 ( .A1(n10718), .A2(n10717), .ZN(n10727) );
  INV_X1 U13777 ( .A(n10727), .ZN(n10731) );
  AND2_X1 U13778 ( .A1(n10429), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10719) );
  NOR2_X1 U13779 ( .A1(n10733), .A2(n10719), .ZN(n10722) );
  NAND2_X1 U13780 ( .A1(n10768), .A2(n10722), .ZN(n10720) );
  NAND2_X1 U13781 ( .A1(n10764), .A2(n10720), .ZN(n10724) );
  OAI211_X1 U13782 ( .C1(n10432), .C2(n13661), .A(n10737), .B(n10722), .ZN(
        n10723) );
  INV_X1 U13783 ( .A(n10728), .ZN(n10730) );
  NAND2_X1 U13784 ( .A1(n10725), .A2(n10431), .ZN(n10755) );
  NAND2_X1 U13785 ( .A1(n10755), .A2(n13368), .ZN(n10726) );
  OAI21_X1 U13786 ( .B1(n10728), .B2(n10727), .A(n10726), .ZN(n10729) );
  NAND2_X1 U13787 ( .A1(n10733), .A2(n10732), .ZN(n10735) );
  NAND2_X1 U13788 ( .A1(n21033), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10734) );
  NAND2_X1 U13789 ( .A1(n10735), .A2(n10734), .ZN(n10742) );
  MUX2_X1 U13790 ( .A(n10743), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10741) );
  XNOR2_X1 U13791 ( .A(n10742), .B(n10741), .ZN(n13367) );
  INV_X1 U13792 ( .A(n13367), .ZN(n10736) );
  NAND2_X1 U13793 ( .A1(n10768), .A2(n10736), .ZN(n10738) );
  OAI211_X1 U13794 ( .C1(n10736), .C2(n10754), .A(n10738), .B(n10737), .ZN(
        n10740) );
  NOR2_X1 U13795 ( .A1(n10738), .A2(n10737), .ZN(n10739) );
  NAND2_X1 U13796 ( .A1(n10742), .A2(n10741), .ZN(n10745) );
  NAND2_X1 U13797 ( .A1(n10743), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10744) );
  NAND2_X1 U13798 ( .A1(n10745), .A2(n10744), .ZN(n10746) );
  MUX2_X1 U13799 ( .A(n17071), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10747) );
  INV_X1 U13800 ( .A(n10753), .ZN(n10751) );
  INV_X1 U13801 ( .A(n10746), .ZN(n10749) );
  INV_X1 U13802 ( .A(n10747), .ZN(n10748) );
  NAND2_X1 U13803 ( .A1(n10749), .A2(n10748), .ZN(n10750) );
  NAND2_X1 U13804 ( .A1(n10751), .A2(n10750), .ZN(n13369) );
  INV_X1 U13805 ( .A(n13369), .ZN(n10752) );
  NAND3_X1 U13806 ( .A1(n15392), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10763), .ZN(n13370) );
  INV_X1 U13807 ( .A(n13370), .ZN(n10756) );
  NAND2_X1 U13808 ( .A1(n10756), .A2(n10754), .ZN(n10761) );
  INV_X1 U13809 ( .A(n10755), .ZN(n10758) );
  NAND3_X1 U13810 ( .A1(n10758), .A2(n10757), .A3(n10756), .ZN(n10759) );
  OAI21_X1 U13811 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n15392), .A(n10759), 
        .ZN(n10760) );
  NOR2_X1 U13812 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20586), .ZN(
        n10762) );
  INV_X1 U13813 ( .A(n10764), .ZN(n10765) );
  NAND2_X1 U13814 ( .A1(n13372), .A2(n10768), .ZN(n10769) );
  NAND2_X1 U13815 ( .A1(n17084), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20348) );
  NAND2_X1 U13816 ( .A1(n10412), .A2(n10437), .ZN(n10771) );
  AND2_X1 U13817 ( .A1(n10772), .A2(n10771), .ZN(n14115) );
  NAND2_X1 U13818 ( .A1(n14116), .A2(n20611), .ZN(n10773) );
  AOI21_X1 U13819 ( .B1(n10441), .B2(n10432), .A(n10773), .ZN(n10774) );
  NAND2_X1 U13820 ( .A1(n13718), .A2(n10412), .ZN(n17079) );
  NAND2_X1 U13821 ( .A1(n20691), .A2(n10983), .ZN(n10779) );
  AOI22_X1 U13822 ( .A1(n14311), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21246), .ZN(n10777) );
  INV_X1 U13823 ( .A(n14429), .ZN(n14102) );
  AND2_X1 U13824 ( .A1(n14102), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10791) );
  NAND2_X1 U13825 ( .A1(n10791), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10776) );
  AND2_X1 U13826 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  NAND2_X1 U13827 ( .A1(n10779), .A2(n10778), .ZN(n13762) );
  NAND2_X1 U13828 ( .A1(n21093), .A2(n10437), .ZN(n10781) );
  NAND2_X1 U13829 ( .A1(n10781), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13779) );
  INV_X1 U13830 ( .A(n10791), .ZN(n10809) );
  NAND2_X1 U13831 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13832 ( .A1(n10783), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10784) );
  OAI211_X1 U13833 ( .C1(n10809), .C2(n10429), .A(n10785), .B(n10784), .ZN(
        n10786) );
  AOI21_X1 U13834 ( .B1(n10782), .B2(n10983), .A(n10786), .ZN(n10787) );
  OR2_X1 U13835 ( .A1(n13779), .A2(n10787), .ZN(n13780) );
  INV_X1 U13836 ( .A(n10787), .ZN(n13781) );
  OR2_X1 U13837 ( .A1(n13781), .A2(n13431), .ZN(n10788) );
  NAND2_X1 U13838 ( .A1(n13780), .A2(n10788), .ZN(n13761) );
  NAND2_X1 U13839 ( .A1(n13762), .A2(n13761), .ZN(n13760) );
  INV_X1 U13840 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10789) );
  XNOR2_X1 U13841 ( .A(n10789), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20427) );
  NAND2_X1 U13842 ( .A1(n21246), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10858) );
  OAI21_X1 U13843 ( .B1(n20427), .B2(n13431), .A(n10858), .ZN(n10790) );
  AOI21_X1 U13844 ( .B1(n14311), .B2(P1_EAX_REG_2__SCAN_IN), .A(n10790), .ZN(
        n10792) );
  NAND2_X1 U13845 ( .A1(n14310), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10795) );
  INV_X1 U13846 ( .A(n15413), .ZN(n10796) );
  INV_X1 U13847 ( .A(n10797), .ZN(n10799) );
  NOR2_X2 U13848 ( .A1(n10797), .A2(n14773), .ZN(n10806) );
  INV_X1 U13849 ( .A(n10806), .ZN(n10798) );
  OAI21_X1 U13850 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10799), .A(
        n10798), .ZN(n14783) );
  AOI22_X1 U13851 ( .A1(n13425), .A2(n14783), .B1(n14310), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13852 ( .A1(n14311), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10800) );
  OAI211_X1 U13853 ( .C1(n10809), .C2(n10317), .A(n10801), .B(n10800), .ZN(
        n10802) );
  INV_X1 U13854 ( .A(n10802), .ZN(n10803) );
  NAND2_X1 U13855 ( .A1(n10804), .A2(n10803), .ZN(n13884) );
  NAND2_X1 U13856 ( .A1(n13885), .A2(n13884), .ZN(n14055) );
  OAI21_X1 U13857 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10806), .A(
        n10814), .ZN(n20523) );
  OAI21_X1 U13858 ( .B1(n20900), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21246), .ZN(n10808) );
  NAND2_X1 U13859 ( .A1(n14311), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10807) );
  OAI211_X1 U13860 ( .C1(n10809), .C2(n15392), .A(n10808), .B(n10807), .ZN(
        n10810) );
  OAI21_X1 U13861 ( .B1(n13431), .B2(n20523), .A(n10810), .ZN(n10811) );
  INV_X1 U13862 ( .A(n10814), .ZN(n10816) );
  INV_X1 U13863 ( .A(n10821), .ZN(n10815) );
  OAI21_X1 U13864 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10816), .A(
        n10815), .ZN(n20401) );
  NAND2_X1 U13865 ( .A1(n20401), .A2(n13425), .ZN(n10817) );
  OAI21_X1 U13866 ( .B1(n20393), .B2(n10858), .A(n10817), .ZN(n10818) );
  AOI21_X1 U13867 ( .B1(n14311), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10818), .ZN(
        n10819) );
  INV_X1 U13868 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10823) );
  OAI21_X1 U13869 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10821), .A(
        n10826), .ZN(n20391) );
  AOI22_X1 U13870 ( .A1(n13425), .A2(n20391), .B1(n14310), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10822) );
  OAI21_X1 U13871 ( .B1(n11233), .B2(n10823), .A(n10822), .ZN(n10824) );
  INV_X1 U13872 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10829) );
  OAI21_X1 U13873 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10827), .A(
        n10856), .ZN(n20374) );
  AOI22_X1 U13874 ( .A1(n13425), .A2(n20374), .B1(n14310), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10828) );
  OAI21_X1 U13875 ( .B1(n11233), .B2(n10829), .A(n10828), .ZN(n10830) );
  AOI22_X1 U13876 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13877 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13878 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13879 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10833) );
  NAND4_X1 U13880 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10842) );
  AOI22_X1 U13881 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13882 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13414), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13883 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13884 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10837) );
  NAND4_X1 U13885 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10841) );
  OAI21_X1 U13886 ( .B1(n10842), .B2(n10841), .A(n10983), .ZN(n10845) );
  XNOR2_X1 U13887 ( .A(n10856), .B(n14761), .ZN(n14757) );
  AOI22_X1 U13888 ( .A1(n14757), .A2(n13425), .B1(n14310), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13889 ( .A1(n14311), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13890 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13404), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U13891 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13892 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13893 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10846) );
  NAND4_X1 U13894 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n10855) );
  AOI22_X1 U13895 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13896 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13897 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U13898 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10850) );
  NAND4_X1 U13899 ( .A1(n10853), .A2(n10852), .A3(n10851), .A4(n10850), .ZN(
        n10854) );
  NOR2_X1 U13900 ( .A1(n10855), .A2(n10854), .ZN(n10862) );
  INV_X1 U13901 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14746) );
  XNOR2_X1 U13902 ( .A(n10873), .B(n14746), .ZN(n15147) );
  NOR2_X1 U13903 ( .A1(n10858), .A2(n14746), .ZN(n10859) );
  AOI21_X1 U13904 ( .B1(n15147), .B2(n13425), .A(n10859), .ZN(n10861) );
  NAND2_X1 U13905 ( .A1(n14311), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10860) );
  OAI211_X1 U13906 ( .C1(n10973), .C2(n10862), .A(n10861), .B(n10860), .ZN(
        n14743) );
  INV_X1 U13907 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14933) );
  AOI22_X1 U13908 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13909 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13910 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13911 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10863) );
  NAND4_X1 U13912 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n10872) );
  AOI22_X1 U13913 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13914 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13915 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13916 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10867) );
  NAND4_X1 U13917 ( .A1(n10870), .A2(n10869), .A3(n10868), .A4(n10867), .ZN(
        n10871) );
  OAI21_X1 U13918 ( .B1(n10872), .B2(n10871), .A(n10983), .ZN(n10876) );
  INV_X1 U13919 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14733) );
  XNOR2_X1 U13920 ( .A(n10888), .B(n14733), .ZN(n15140) );
  AOI22_X1 U13921 ( .A1(n15140), .A2(n13425), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14310), .ZN(n10875) );
  OAI211_X1 U13922 ( .C1(n11233), .C2(n14933), .A(n10876), .B(n10875), .ZN(
        n14728) );
  AOI22_X1 U13923 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13924 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13925 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13926 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10877) );
  NAND4_X1 U13927 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n10886) );
  AOI22_X1 U13928 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13929 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U13930 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13931 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10881) );
  NAND4_X1 U13932 ( .A1(n10884), .A2(n10883), .A3(n10882), .A4(n10881), .ZN(
        n10885) );
  OR2_X1 U13933 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  NAND2_X1 U13934 ( .A1(n10983), .A2(n10887), .ZN(n14717) );
  NAND2_X1 U13935 ( .A1(n14311), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10895) );
  INV_X1 U13936 ( .A(n10890), .ZN(n10892) );
  INV_X1 U13937 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13938 ( .A1(n10892), .A2(n10891), .ZN(n10893) );
  NAND2_X1 U13939 ( .A1(n10940), .A2(n10893), .ZN(n15127) );
  AOI22_X1 U13940 ( .A1(n15127), .A2(n13425), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n14310), .ZN(n10894) );
  AOI22_X1 U13941 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13942 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13404), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13943 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13944 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10896) );
  NAND4_X1 U13945 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10905) );
  AOI22_X1 U13946 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13414), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13947 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13948 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10467), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13949 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10900) );
  NAND4_X1 U13950 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(
        n10904) );
  OAI21_X1 U13951 ( .B1(n10905), .B2(n10904), .A(n10983), .ZN(n10909) );
  NAND2_X1 U13952 ( .A1(n14311), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10908) );
  INV_X1 U13953 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15111) );
  XNOR2_X1 U13954 ( .A(n10940), .B(n15111), .ZN(n14711) );
  NAND2_X1 U13955 ( .A1(n14711), .A2(n13425), .ZN(n10907) );
  NAND2_X1 U13956 ( .A1(n14310), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10906) );
  NAND4_X1 U13957 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n14701) );
  AOI22_X1 U13958 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13959 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13960 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13961 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10910) );
  NAND4_X1 U13962 ( .A1(n10913), .A2(n10912), .A3(n10911), .A4(n10910), .ZN(
        n10919) );
  AOI22_X1 U13963 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11184), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13964 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13965 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13966 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10914) );
  NAND4_X1 U13967 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10918) );
  OAI21_X1 U13968 ( .B1(n10919), .B2(n10918), .A(n10983), .ZN(n10925) );
  NAND2_X1 U13969 ( .A1(n14311), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10924) );
  OR2_X1 U13970 ( .A1(n10940), .A2(n15111), .ZN(n10921) );
  INV_X1 U13971 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10920) );
  XNOR2_X1 U13972 ( .A(n10921), .B(n10920), .ZN(n15107) );
  NAND2_X1 U13973 ( .A1(n15107), .A2(n13425), .ZN(n10923) );
  NAND2_X1 U13974 ( .A1(n14310), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10922) );
  NAND4_X1 U13975 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n14689) );
  AOI22_X1 U13976 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13977 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13978 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13979 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U13980 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10935) );
  AOI22_X1 U13981 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13982 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13983 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13984 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10930) );
  NAND4_X1 U13985 ( .A1(n10933), .A2(n10932), .A3(n10931), .A4(n10930), .ZN(
        n10934) );
  NOR2_X1 U13986 ( .A1(n10935), .A2(n10934), .ZN(n10939) );
  OAI21_X1 U13987 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20900), .A(
        n21246), .ZN(n10936) );
  INV_X1 U13988 ( .A(n10936), .ZN(n10937) );
  AOI21_X1 U13989 ( .B1(n14311), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10937), .ZN(
        n10938) );
  OAI21_X1 U13990 ( .B1(n13428), .B2(n10939), .A(n10938), .ZN(n10946) );
  AND2_X1 U13991 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10941) );
  OR2_X2 U13992 ( .A1(n10943), .A2(n21437), .ZN(n10994) );
  NAND2_X1 U13993 ( .A1(n10943), .A2(n21437), .ZN(n10944) );
  AND2_X1 U13994 ( .A1(n10994), .A2(n10944), .ZN(n14646) );
  NAND2_X1 U13995 ( .A1(n14646), .A2(n13425), .ZN(n10945) );
  AOI22_X1 U13996 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13997 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13998 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13999 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10947) );
  NAND4_X1 U14000 ( .A1(n10950), .A2(n10949), .A3(n10948), .A4(n10947), .ZN(
        n10956) );
  AOI22_X1 U14001 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14002 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14003 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U14004 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10951) );
  NAND4_X1 U14005 ( .A1(n10954), .A2(n10953), .A3(n10952), .A4(n10951), .ZN(
        n10955) );
  NOR2_X1 U14006 ( .A1(n10956), .A2(n10955), .ZN(n10959) );
  INV_X1 U14007 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14634) );
  XNOR2_X1 U14008 ( .A(n10994), .B(n14634), .ZN(n15061) );
  NAND2_X1 U14009 ( .A1(n15061), .A2(n13425), .ZN(n10958) );
  AOI22_X1 U14010 ( .A1(n14311), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n14310), .ZN(n10957) );
  OAI211_X1 U14011 ( .C1(n13428), .C2(n10959), .A(n10958), .B(n10957), .ZN(
        n14628) );
  AOI22_X1 U14012 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U14013 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U14014 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U14015 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10960) );
  NAND4_X1 U14016 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(
        n10969) );
  AOI22_X1 U14017 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U14018 ( .A1(n13410), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U14019 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U14020 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10964) );
  NAND4_X1 U14021 ( .A1(n10967), .A2(n10966), .A3(n10965), .A4(n10964), .ZN(
        n10968) );
  NOR2_X1 U14022 ( .A1(n10969), .A2(n10968), .ZN(n10974) );
  XNOR2_X1 U14023 ( .A(n10970), .B(n14662), .ZN(n15085) );
  NAND2_X1 U14024 ( .A1(n15085), .A2(n13425), .ZN(n10972) );
  AOI22_X1 U14025 ( .A1(n14311), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n14310), .ZN(n10971) );
  OAI211_X1 U14026 ( .C1(n10974), .C2(n10973), .A(n10972), .B(n10971), .ZN(
        n14627) );
  AOI22_X1 U14027 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U14028 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14029 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U14030 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10975) );
  NAND4_X1 U14031 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        n10985) );
  AOI22_X1 U14032 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U14033 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U14034 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U14035 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10979) );
  NAND4_X1 U14036 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n10984) );
  OAI21_X1 U14037 ( .B1(n10985), .B2(n10984), .A(n10983), .ZN(n10992) );
  NAND2_X1 U14038 ( .A1(n14311), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10991) );
  INV_X1 U14039 ( .A(n10986), .ZN(n10988) );
  INV_X1 U14040 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10987) );
  XNOR2_X1 U14041 ( .A(n10988), .B(n10987), .ZN(n15094) );
  NAND2_X1 U14042 ( .A1(n15094), .A2(n13425), .ZN(n10990) );
  NAND2_X1 U14043 ( .A1(n14310), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10989) );
  NAND4_X1 U14044 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n14670) );
  NOR2_X2 U14045 ( .A1(n10994), .A2(n14634), .ZN(n11118) );
  AND2_X2 U14046 ( .A1(n10995), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11063) );
  AND2_X2 U14047 ( .A1(n10996), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11042) );
  XNOR2_X1 U14048 ( .A(n11157), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14513) );
  AOI22_X1 U14049 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13404), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14050 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14051 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14052 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10997) );
  NAND4_X1 U14053 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11006) );
  AOI22_X1 U14054 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14055 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14056 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14057 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11001) );
  NAND4_X1 U14058 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11005) );
  NOR2_X1 U14059 ( .A1(n11006), .A2(n11005), .ZN(n11054) );
  AOI22_X1 U14060 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14061 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14062 ( .A1(n13410), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14063 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11007) );
  NAND4_X1 U14064 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11016) );
  AOI22_X1 U14065 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14066 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14067 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U14068 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11011) );
  NAND4_X1 U14069 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11015) );
  NOR2_X1 U14070 ( .A1(n11016), .A2(n11015), .ZN(n11055) );
  NOR2_X1 U14071 ( .A1(n11054), .A2(n11055), .ZN(n11047) );
  AOI22_X1 U14072 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14073 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14074 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14075 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11017) );
  NAND4_X1 U14076 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11026) );
  AOI22_X1 U14077 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U14078 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11023) );
  INV_X1 U14079 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20606) );
  AOI22_X1 U14080 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14081 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11021) );
  NAND4_X1 U14082 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11025) );
  OR2_X1 U14083 ( .A1(n11026), .A2(n11025), .ZN(n11046) );
  NAND2_X1 U14084 ( .A1(n11047), .A2(n11046), .ZN(n11163) );
  AOI22_X1 U14085 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14086 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14087 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14088 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11027) );
  NAND4_X1 U14089 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11036) );
  AOI22_X1 U14090 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14091 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14092 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14093 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11031) );
  NAND4_X1 U14094 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11035) );
  NOR2_X1 U14095 ( .A1(n11036), .A2(n11035), .ZN(n11164) );
  XOR2_X1 U14096 ( .A(n11163), .B(n11164), .Z(n11040) );
  INV_X1 U14097 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U14098 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11037) );
  OAI211_X1 U14099 ( .C1(n11233), .C2(n11038), .A(n13431), .B(n11037), .ZN(
        n11039) );
  AOI21_X1 U14100 ( .B1(n11040), .B2(n11235), .A(n11039), .ZN(n11041) );
  AOI21_X1 U14101 ( .B1(n14513), .B2(n13425), .A(n11041), .ZN(n14510) );
  INV_X1 U14102 ( .A(n11042), .ZN(n11044) );
  INV_X1 U14103 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14104 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  NAND2_X1 U14105 ( .A1(n11157), .A2(n11045), .ZN(n14984) );
  OR2_X1 U14106 ( .A1(n14984), .A2(n13431), .ZN(n11053) );
  XNOR2_X1 U14107 ( .A(n11047), .B(n11046), .ZN(n11051) );
  NAND2_X1 U14108 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11048) );
  NAND2_X1 U14109 ( .A1(n13431), .A2(n11048), .ZN(n11049) );
  AOI21_X1 U14110 ( .B1(n14311), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11049), .ZN(
        n11050) );
  OAI21_X1 U14111 ( .B1(n11051), .B2(n13428), .A(n11050), .ZN(n11052) );
  INV_X1 U14112 ( .A(n14528), .ZN(n11082) );
  XNOR2_X1 U14113 ( .A(n11066), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14994) );
  NAND2_X1 U14114 ( .A1(n14994), .A2(n13425), .ZN(n11062) );
  XOR2_X1 U14115 ( .A(n11055), .B(n11054), .Z(n11056) );
  NAND2_X1 U14116 ( .A1(n11056), .A2(n11235), .ZN(n11060) );
  NAND2_X1 U14117 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11057) );
  NAND2_X1 U14118 ( .A1(n13431), .A2(n11057), .ZN(n11058) );
  AOI21_X1 U14119 ( .B1(n14311), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11058), .ZN(
        n11059) );
  NAND2_X1 U14120 ( .A1(n11060), .A2(n11059), .ZN(n11061) );
  NAND2_X1 U14121 ( .A1(n11062), .A2(n11061), .ZN(n14537) );
  INV_X1 U14122 ( .A(n11063), .ZN(n11064) );
  INV_X1 U14123 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14558) );
  NAND2_X1 U14124 ( .A1(n11064), .A2(n14558), .ZN(n11065) );
  NAND2_X1 U14125 ( .A1(n11066), .A2(n11065), .ZN(n15005) );
  OR2_X1 U14126 ( .A1(n15005), .A2(n13431), .ZN(n11081) );
  AOI22_X1 U14127 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14128 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14129 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14130 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11067) );
  NAND4_X1 U14131 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11076) );
  AOI22_X1 U14132 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14133 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14134 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14135 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U14136 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11075) );
  NOR2_X1 U14137 ( .A1(n11076), .A2(n11075), .ZN(n11079) );
  OAI21_X1 U14138 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20900), .A(
        n21246), .ZN(n11078) );
  NAND2_X1 U14139 ( .A1(n14311), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n11077) );
  OAI211_X1 U14140 ( .C1(n13428), .C2(n11079), .A(n11078), .B(n11077), .ZN(
        n11080) );
  NAND2_X1 U14141 ( .A1(n11081), .A2(n11080), .ZN(n14552) );
  NOR2_X1 U14142 ( .A1(n11082), .A2(n14525), .ZN(n14509) );
  AND2_X1 U14143 ( .A1(n14510), .A2(n14509), .ZN(n11155) );
  INV_X1 U14144 ( .A(n11083), .ZN(n11085) );
  INV_X1 U14145 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U14146 ( .A1(n11085), .A2(n11084), .ZN(n11086) );
  NAND2_X1 U14147 ( .A1(n11140), .A2(n11086), .ZN(n15025) );
  OR2_X1 U14148 ( .A1(n15025), .A2(n13431), .ZN(n11101) );
  AOI22_X1 U14149 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9613), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14150 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11184), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14151 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11220), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14152 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n13404), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11087) );
  NAND4_X1 U14153 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11096) );
  AOI22_X1 U14154 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9612), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14155 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14156 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U14157 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11091) );
  NAND4_X1 U14158 ( .A1(n11094), .A2(n11093), .A3(n11092), .A4(n11091), .ZN(
        n11095) );
  NOR2_X1 U14159 ( .A1(n11096), .A2(n11095), .ZN(n11099) );
  OAI21_X1 U14160 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20900), .A(
        n21246), .ZN(n11098) );
  NAND2_X1 U14161 ( .A1(n14311), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n11097) );
  OAI211_X1 U14162 ( .C1(n13428), .C2(n11099), .A(n11098), .B(n11097), .ZN(
        n11100) );
  NAND2_X1 U14163 ( .A1(n11101), .A2(n11100), .ZN(n14582) );
  INV_X1 U14164 ( .A(n11102), .ZN(n11122) );
  XNOR2_X1 U14165 ( .A(n11122), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14604) );
  NAND2_X1 U14166 ( .A1(n14604), .A2(n13425), .ZN(n11117) );
  AOI22_X1 U14167 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14168 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14169 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14170 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11103) );
  NAND4_X1 U14171 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11112) );
  AOI22_X1 U14172 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14173 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14174 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14175 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11107) );
  NAND4_X1 U14176 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n11111) );
  NOR2_X1 U14177 ( .A1(n11112), .A2(n11111), .ZN(n11115) );
  INV_X1 U14178 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14607) );
  AOI21_X1 U14179 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14607), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11113) );
  AOI21_X1 U14180 ( .B1(n14311), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11113), .ZN(
        n11114) );
  OAI21_X1 U14181 ( .B1(n13428), .B2(n11115), .A(n11114), .ZN(n11116) );
  NAND2_X1 U14182 ( .A1(n11117), .A2(n11116), .ZN(n14596) );
  INV_X1 U14183 ( .A(n11118), .ZN(n11120) );
  INV_X1 U14184 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U14185 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  NAND2_X1 U14186 ( .A1(n11122), .A2(n11121), .ZN(n15040) );
  OR2_X1 U14187 ( .A1(n15040), .A2(n13431), .ZN(n11139) );
  AOI22_X1 U14188 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14189 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14190 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14191 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11124) );
  NAND4_X1 U14192 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11133) );
  AOI22_X1 U14193 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10561), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14194 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14195 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14196 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11128) );
  NAND4_X1 U14197 ( .A1(n11131), .A2(n11130), .A3(n11129), .A4(n11128), .ZN(
        n11132) );
  NOR2_X1 U14198 ( .A1(n11133), .A2(n11132), .ZN(n11137) );
  NAND2_X1 U14199 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14200 ( .A1(n13431), .A2(n11134), .ZN(n11135) );
  AOI21_X1 U14201 ( .B1(n14311), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11135), .ZN(
        n11136) );
  OAI21_X1 U14202 ( .B1(n13428), .B2(n11137), .A(n11136), .ZN(n11138) );
  NAND2_X1 U14203 ( .A1(n11139), .A2(n11138), .ZN(n14566) );
  NOR3_X1 U14204 ( .A1(n14582), .A2(n14596), .A3(n14566), .ZN(n11154) );
  XNOR2_X1 U14205 ( .A(n11140), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15013) );
  INV_X1 U14206 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14571) );
  AOI21_X1 U14207 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14571), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11141) );
  AOI21_X1 U14208 ( .B1(n14311), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11141), .ZN(
        n11153) );
  AOI22_X1 U14209 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14210 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14211 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14212 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11142) );
  NAND4_X1 U14213 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11151) );
  AOI22_X1 U14214 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13414), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14215 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14216 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14217 ( .A1(n13405), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11146) );
  NAND4_X1 U14218 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11150) );
  OAI21_X1 U14219 ( .B1(n11151), .B2(n11150), .A(n11235), .ZN(n11152) );
  AOI22_X1 U14220 ( .A1(n15013), .A2(n13425), .B1(n11153), .B2(n11152), .ZN(
        n14568) );
  AND2_X2 U14221 ( .A1(n11158), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11159) );
  INV_X1 U14222 ( .A(n11159), .ZN(n11161) );
  INV_X1 U14223 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11160) );
  NAND2_X1 U14224 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  NAND2_X1 U14225 ( .A1(n11198), .A2(n11162), .ZN(n14969) );
  NOR2_X1 U14226 ( .A1(n11164), .A2(n11163), .ZN(n11183) );
  AOI22_X1 U14227 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14228 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14229 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14230 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11165) );
  NAND4_X1 U14231 ( .A1(n11168), .A2(n11167), .A3(n11166), .A4(n11165), .ZN(
        n11174) );
  AOI22_X1 U14232 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14233 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14234 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14235 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11169) );
  NAND4_X1 U14236 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11173) );
  OR2_X1 U14237 ( .A1(n11174), .A2(n11173), .ZN(n11182) );
  XNOR2_X1 U14238 ( .A(n11183), .B(n11182), .ZN(n11178) );
  NAND2_X1 U14239 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11175) );
  NAND2_X1 U14240 ( .A1(n13431), .A2(n11175), .ZN(n11176) );
  AOI21_X1 U14241 ( .B1(n14311), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11176), .ZN(
        n11177) );
  OAI21_X1 U14242 ( .B1(n11178), .B2(n13428), .A(n11177), .ZN(n11179) );
  NAND2_X1 U14243 ( .A1(n11180), .A2(n11179), .ZN(n14495) );
  XNOR2_X1 U14244 ( .A(n11198), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14484) );
  INV_X1 U14245 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14485) );
  NOR2_X1 U14246 ( .A1(n14485), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11181) );
  AOI211_X1 U14247 ( .C1(n14311), .C2(P1_EAX_REG_27__SCAN_IN), .A(n13425), .B(
        n11181), .ZN(n11197) );
  NAND2_X1 U14248 ( .A1(n11183), .A2(n11182), .ZN(n11202) );
  AOI22_X1 U14249 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11184), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14250 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9612), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14251 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14252 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11185) );
  NAND4_X1 U14253 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n11194) );
  AOI22_X1 U14254 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9613), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14255 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14256 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14257 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10467), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11189) );
  NAND4_X1 U14258 ( .A1(n11192), .A2(n11191), .A3(n11190), .A4(n11189), .ZN(
        n11193) );
  NOR2_X1 U14259 ( .A1(n11194), .A2(n11193), .ZN(n11203) );
  XOR2_X1 U14260 ( .A(n11202), .B(n11203), .Z(n11195) );
  NAND2_X1 U14261 ( .A1(n11195), .A2(n11235), .ZN(n11196) );
  AOI22_X1 U14262 ( .A1(n14484), .A2(n13425), .B1(n11197), .B2(n11196), .ZN(
        n14481) );
  OR2_X2 U14263 ( .A1(n11198), .A2(n14485), .ZN(n11200) );
  INV_X1 U14264 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11199) );
  OR2_X2 U14265 ( .A1(n11200), .A2(n11199), .ZN(n13378) );
  NAND2_X1 U14266 ( .A1(n11200), .A2(n11199), .ZN(n11201) );
  NAND2_X1 U14267 ( .A1(n13378), .A2(n11201), .ZN(n14948) );
  NOR2_X1 U14268 ( .A1(n11203), .A2(n11202), .ZN(n11219) );
  AOI22_X1 U14269 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10467), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14270 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14271 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14272 ( .A1(n13411), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11204) );
  NAND4_X1 U14273 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11213) );
  AOI22_X1 U14274 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14275 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10461), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14276 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14277 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11208) );
  NAND4_X1 U14278 ( .A1(n11211), .A2(n11210), .A3(n11209), .A4(n11208), .ZN(
        n11212) );
  OR2_X1 U14279 ( .A1(n11213), .A2(n11212), .ZN(n11218) );
  XNOR2_X1 U14280 ( .A(n11219), .B(n11218), .ZN(n11216) );
  AOI21_X1 U14281 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21246), .A(
        n13425), .ZN(n11215) );
  NAND2_X1 U14282 ( .A1(n14311), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11214) );
  OAI211_X1 U14283 ( .C1(n11216), .C2(n13428), .A(n11215), .B(n11214), .ZN(
        n11217) );
  OAI21_X1 U14284 ( .B1(n14948), .B2(n13431), .A(n11217), .ZN(n14468) );
  XNOR2_X1 U14285 ( .A(n13378), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14457) );
  NAND2_X1 U14286 ( .A1(n11219), .A2(n11218), .ZN(n13421) );
  AOI22_X1 U14287 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14288 ( .A1(n10531), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13410), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14289 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14290 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11221) );
  NAND4_X1 U14291 ( .A1(n11224), .A2(n11223), .A3(n11222), .A4(n11221), .ZN(
        n11230) );
  AOI22_X1 U14292 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14293 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14294 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14295 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11225) );
  NAND4_X1 U14296 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(
        n11229) );
  NOR2_X1 U14297 ( .A1(n11230), .A2(n11229), .ZN(n13422) );
  XOR2_X1 U14298 ( .A(n13421), .B(n13422), .Z(n11236) );
  INV_X1 U14299 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n11232) );
  NAND2_X1 U14300 ( .A1(n21246), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11231) );
  OAI211_X1 U14301 ( .C1(n11233), .C2(n11232), .A(n13431), .B(n11231), .ZN(
        n11234) );
  AOI21_X1 U14302 ( .B1(n11236), .B2(n11235), .A(n11234), .ZN(n11237) );
  AOI21_X1 U14303 ( .B1(n14457), .B2(n13425), .A(n11237), .ZN(n13432) );
  NAND2_X1 U14304 ( .A1(n20351), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17125) );
  NAND2_X1 U14305 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21186), .ZN(n21091) );
  NOR2_X1 U14306 ( .A1(n14443), .A2(n15122), .ZN(n11247) );
  NAND2_X1 U14307 ( .A1(n11241), .A2(n21184), .ZN(n21291) );
  NAND2_X1 U14308 ( .A1(n21291), .A2(n20351), .ZN(n11238) );
  NAND2_X1 U14309 ( .A1(n20351), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U14310 ( .A1(n20900), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14311 ( .A1(n11240), .A2(n11239), .ZN(n14071) );
  NAND2_X2 U14312 ( .A1(n15112), .A2(n14071), .ZN(n20524) );
  INV_X1 U14313 ( .A(n20524), .ZN(n15119) );
  NAND2_X1 U14314 ( .A1(n14457), .A2(n15119), .ZN(n11245) );
  INV_X1 U14315 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11242) );
  OR2_X2 U14316 ( .A1(n11241), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20416) );
  NAND2_X1 U14317 ( .A1(n20580), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15155) );
  OAI21_X1 U14318 ( .B1(n15112), .B2(n11242), .A(n15155), .ZN(n11243) );
  INV_X1 U14319 ( .A(n11243), .ZN(n11244) );
  NAND2_X4 U14320 ( .A1(n16930), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17950) );
  INV_X1 U14321 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n21374) );
  NAND2_X1 U14322 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11250) );
  NAND2_X1 U14323 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11249) );
  OAI211_X1 U14324 ( .C1(n17950), .C2(n21374), .A(n11250), .B(n11249), .ZN(
        n11251) );
  INV_X1 U14325 ( .A(n11251), .ZN(n11257) );
  AND2_X4 U14326 ( .A1(n16904), .A2(n11261), .ZN(n17931) );
  AOI22_X1 U14327 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11256) );
  AND2_X2 U14328 ( .A1(n11261), .A2(n17046), .ZN(n11411) );
  AOI22_X1 U14329 ( .A1(n17898), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U14330 ( .A1(n11465), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11254) );
  NAND4_X1 U14331 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11267) );
  AND2_X2 U14332 ( .A1(n11259), .A2(n17046), .ZN(n11447) );
  AOI22_X1 U14333 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11265) );
  AND2_X2 U14334 ( .A1(n11259), .A2(n16904), .ZN(n11467) );
  AOI22_X1 U14335 ( .A1(n11467), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17878), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11264) );
  INV_X4 U14336 ( .A(n17818), .ZN(n17933) );
  AOI22_X1 U14337 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11263) );
  AND2_X2 U14338 ( .A1(n16911), .A2(n11261), .ZN(n11509) );
  AOI22_X1 U14339 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11262) );
  NAND4_X1 U14340 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11266) );
  OR2_X2 U14341 ( .A1(n11267), .A2(n11266), .ZN(n16663) );
  INV_X1 U14342 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17909) );
  NAND2_X1 U14343 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11268) );
  AOI22_X1 U14344 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14345 ( .A1(n17793), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11270) );
  NAND2_X1 U14346 ( .A1(n11465), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11269) );
  AOI22_X1 U14347 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14348 ( .A1(n11467), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14349 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14350 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11272) );
  INV_X1 U14351 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17740) );
  NAND2_X1 U14352 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14353 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11276) );
  OAI211_X1 U14354 ( .C1(n17950), .C2(n17740), .A(n11277), .B(n11276), .ZN(
        n11278) );
  INV_X1 U14355 ( .A(n11278), .ZN(n11282) );
  AOI22_X1 U14356 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14357 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17793), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11280) );
  NAND2_X1 U14358 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11279) );
  NAND4_X1 U14359 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11288) );
  AOI22_X1 U14360 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14361 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14362 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14363 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14364 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11287) );
  INV_X1 U14365 ( .A(n11369), .ZN(n11304) );
  NAND2_X1 U14366 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14367 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11292) );
  NAND2_X1 U14368 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11291) );
  NAND2_X1 U14369 ( .A1(n17898), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11290) );
  AOI22_X1 U14370 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U14371 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11295) );
  NAND2_X1 U14372 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11294) );
  NAND4_X1 U14373 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n11303) );
  AOI22_X1 U14374 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14375 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14376 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14377 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14378 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11302) );
  NAND2_X1 U14379 ( .A1(n11304), .A2(n11587), .ZN(n11373) );
  INV_X1 U14380 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14381 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14382 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11305) );
  OAI211_X1 U14383 ( .C1(n17950), .C2(n11466), .A(n11306), .B(n11305), .ZN(
        n11307) );
  INV_X1 U14384 ( .A(n11307), .ZN(n11311) );
  AOI22_X1 U14385 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14386 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11322), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11309) );
  NAND2_X1 U14387 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11308) );
  NAND4_X1 U14388 ( .A1(n11311), .A2(n11310), .A3(n11309), .A4(n11308), .ZN(
        n11317) );
  AOI22_X1 U14389 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14390 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14391 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17793), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14392 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11312) );
  NAND4_X1 U14393 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n11316) );
  INV_X1 U14394 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14395 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11319) );
  NAND2_X1 U14396 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11318) );
  OAI211_X1 U14397 ( .C1(n17950), .C2(n11320), .A(n11319), .B(n11318), .ZN(
        n11321) );
  INV_X1 U14398 ( .A(n11321), .ZN(n11326) );
  AOI22_X1 U14399 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14400 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14401 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11323) );
  NAND4_X1 U14402 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11332) );
  AOI22_X1 U14403 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17912), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14404 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14405 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14406 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17793), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11327) );
  NAND4_X1 U14407 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11331) );
  INV_X1 U14408 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16996) );
  NAND2_X1 U14409 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14410 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11334) );
  OAI211_X1 U14411 ( .C1(n17950), .C2(n16996), .A(n11335), .B(n11334), .ZN(
        n11336) );
  INV_X1 U14412 ( .A(n11336), .ZN(n11340) );
  AOI22_X1 U14413 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14414 ( .A1(n17793), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U14415 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11337) );
  NAND4_X1 U14416 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11346) );
  AOI22_X1 U14417 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11344) );
  INV_X2 U14418 ( .A(n11434), .ZN(n17912) );
  AOI22_X1 U14419 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14420 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14421 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11341) );
  NAND4_X1 U14422 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11345) );
  OR2_X2 U14423 ( .A1(n16830), .A2(n16771), .ZN(n18369) );
  XNOR2_X1 U14424 ( .A(n11362), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18541) );
  INV_X1 U14425 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14426 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14427 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11347) );
  OAI211_X1 U14428 ( .C1(n17950), .C2(n11349), .A(n11348), .B(n11347), .ZN(
        n11350) );
  INV_X1 U14429 ( .A(n11350), .ZN(n11354) );
  AOI22_X1 U14430 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14431 ( .A1(n17793), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U14432 ( .A1(n11465), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11351) );
  NAND4_X1 U14433 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11360) );
  AOI22_X1 U14434 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14435 ( .A1(n11467), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17878), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14436 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14437 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14438 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  INV_X1 U14439 ( .A(n13923), .ZN(n11596) );
  NAND2_X1 U14440 ( .A1(n11596), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11361) );
  NAND2_X1 U14441 ( .A1(n18549), .A2(n11361), .ZN(n18540) );
  NAND2_X1 U14442 ( .A1(n18541), .A2(n18540), .ZN(n18539) );
  INV_X1 U14443 ( .A(n11362), .ZN(n11363) );
  NAND2_X1 U14444 ( .A1(n11363), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11364) );
  INV_X1 U14445 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18805) );
  XNOR2_X1 U14446 ( .A(n11367), .B(n18805), .ZN(n18524) );
  INV_X1 U14447 ( .A(n18126), .ZN(n11365) );
  NAND2_X1 U14448 ( .A1(n11593), .A2(n11365), .ZN(n11366) );
  AND2_X1 U14449 ( .A1(n11369), .A2(n11366), .ZN(n18523) );
  NAND2_X1 U14450 ( .A1(n18524), .A2(n18523), .ZN(n18526) );
  NAND2_X1 U14451 ( .A1(n11367), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11368) );
  NAND2_X1 U14452 ( .A1(n18526), .A2(n11368), .ZN(n18509) );
  XNOR2_X1 U14453 ( .A(n11369), .B(n18119), .ZN(n11370) );
  XNOR2_X1 U14454 ( .A(n11370), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18508) );
  NAND2_X1 U14455 ( .A1(n18509), .A2(n18508), .ZN(n18511) );
  INV_X1 U14456 ( .A(n11370), .ZN(n11371) );
  NAND2_X1 U14457 ( .A1(n11371), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11372) );
  NAND2_X2 U14458 ( .A1(n18511), .A2(n11372), .ZN(n11377) );
  NAND2_X1 U14459 ( .A1(n11373), .A2(n18114), .ZN(n11374) );
  NAND2_X1 U14460 ( .A1(n11380), .A2(n11374), .ZN(n11375) );
  INV_X1 U14461 ( .A(n11375), .ZN(n11376) );
  NAND2_X1 U14462 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  INV_X1 U14463 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11379) );
  XNOR2_X1 U14464 ( .A(n11605), .B(n11379), .ZN(n18482) );
  XNOR2_X1 U14465 ( .A(n11380), .B(n18482), .ZN(n18488) );
  XNOR2_X1 U14466 ( .A(n11380), .B(n11605), .ZN(n11381) );
  NAND2_X1 U14467 ( .A1(n11381), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U14468 ( .A1(n16830), .A2(n16771), .ZN(n11383) );
  NAND2_X1 U14469 ( .A1(n18369), .A2(n11383), .ZN(n11384) );
  NAND2_X1 U14470 ( .A1(n18473), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18472) );
  INV_X1 U14471 ( .A(n11384), .ZN(n11385) );
  NAND2_X1 U14472 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  INV_X1 U14473 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11388) );
  INV_X1 U14474 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18680) );
  NAND3_X1 U14475 ( .A1(n11388), .A2(n18680), .A3(n18374), .ZN(n11392) );
  NOR2_X1 U14476 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18445) );
  INV_X1 U14477 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11390) );
  INV_X1 U14478 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11389) );
  NAND3_X1 U14479 ( .A1(n18445), .A2(n11390), .A3(n11389), .ZN(n11391) );
  INV_X1 U14480 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18658) );
  NAND2_X1 U14481 ( .A1(n18367), .A2(n18658), .ZN(n11393) );
  NAND2_X1 U14482 ( .A1(n18348), .A2(n11393), .ZN(n18342) );
  NAND2_X2 U14483 ( .A1(n11394), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U14484 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18727) );
  NOR2_X1 U14485 ( .A1(n18727), .A2(n11390), .ZN(n18697) );
  NAND2_X1 U14486 ( .A1(n18697), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18677) );
  NOR2_X1 U14487 ( .A1(n18677), .A2(n11388), .ZN(n18386) );
  OR2_X2 U14488 ( .A1(n11633), .A2(n16850), .ZN(n18660) );
  AND2_X1 U14489 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18631) );
  INV_X1 U14490 ( .A(n18631), .ZN(n18627) );
  AND2_X1 U14491 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18606) );
  NAND2_X1 U14492 ( .A1(n18606), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18588) );
  NAND2_X1 U14493 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11395) );
  NOR2_X1 U14494 ( .A1(n18588), .A2(n11395), .ZN(n11396) );
  INV_X1 U14495 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18635) );
  NOR2_X1 U14496 ( .A1(n18627), .A2(n18635), .ZN(n18602) );
  INV_X1 U14497 ( .A(n18602), .ZN(n18600) );
  NOR2_X1 U14498 ( .A1(n18588), .A2(n18600), .ZN(n18273) );
  AND2_X1 U14499 ( .A1(n18273), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16852) );
  AND2_X1 U14500 ( .A1(n16852), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16750) );
  INV_X1 U14501 ( .A(n16750), .ZN(n11584) );
  INV_X1 U14502 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18620) );
  NAND2_X1 U14503 ( .A1(n18329), .A2(n18620), .ZN(n11397) );
  NOR2_X1 U14504 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11397), .ZN(
        n18285) );
  INV_X1 U14505 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18587) );
  INV_X1 U14506 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18591) );
  INV_X1 U14507 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18267) );
  NAND4_X1 U14508 ( .A1(n18285), .A2(n18587), .A3(n18591), .A4(n18267), .ZN(
        n11398) );
  OAI21_X1 U14509 ( .B1(n18660), .B2(n11584), .A(n11398), .ZN(n11399) );
  INV_X1 U14510 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16748) );
  NAND2_X1 U14511 ( .A1(n11401), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11400) );
  NAND2_X1 U14512 ( .A1(n16747), .A2(n18369), .ZN(n18251) );
  OAI211_X1 U14513 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18369), .A(
        n11400), .B(n18251), .ZN(n16734) );
  NAND2_X1 U14514 ( .A1(n11401), .A2(n18367), .ZN(n18252) );
  AND2_X1 U14515 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16844) );
  INV_X1 U14516 ( .A(n16844), .ZN(n11402) );
  NAND2_X1 U14517 ( .A1(n18367), .A2(n11402), .ZN(n11403) );
  INV_X1 U14518 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16854) );
  INV_X1 U14519 ( .A(n16724), .ZN(n16820) );
  INV_X1 U14520 ( .A(n16829), .ZN(n16723) );
  AOI21_X1 U14521 ( .B1(n16820), .B2(n18367), .A(n16723), .ZN(n11583) );
  INV_X1 U14522 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16808) );
  XNOR2_X1 U14523 ( .A(n18369), .B(n16808), .ZN(n11582) );
  NAND2_X1 U14524 ( .A1(n11583), .A2(n11582), .ZN(n11581) );
  AOI22_X1 U14525 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14526 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11447), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11409) );
  INV_X1 U14527 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17940) );
  INV_X1 U14528 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17942) );
  OAI22_X1 U14529 ( .A1(n17799), .A2(n17940), .B1(n17747), .B2(n17942), .ZN(
        n11406) );
  AOI21_X1 U14530 ( .B1(n17932), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n11406), .ZN(n11408) );
  NAND2_X1 U14531 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11407) );
  NAND4_X1 U14532 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11418) );
  AOI22_X1 U14533 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14534 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11415) );
  INV_X1 U14535 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17800) );
  OAI22_X1 U14536 ( .A1(n17709), .A2(n16980), .B1(n17939), .B2(n17800), .ZN(
        n11412) );
  AOI21_X1 U14537 ( .B1(n17020), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n11412), .ZN(n11414) );
  NAND2_X1 U14538 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11413) );
  NAND4_X1 U14539 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11417) );
  INV_X1 U14540 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11421) );
  NAND2_X1 U14541 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11420) );
  NAND2_X1 U14542 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11419) );
  OAI211_X1 U14543 ( .C1(n17950), .C2(n11421), .A(n11420), .B(n11419), .ZN(
        n11422) );
  INV_X1 U14544 ( .A(n11422), .ZN(n11426) );
  AOI22_X1 U14545 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14546 ( .A1(n17793), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U14547 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11423) );
  NAND4_X1 U14548 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11432) );
  AOI22_X1 U14549 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14550 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17878), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14551 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14552 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11427) );
  NAND4_X1 U14553 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n11431) );
  NAND2_X1 U14554 ( .A1(n13916), .A2(n18133), .ZN(n11524) );
  NAND2_X1 U14555 ( .A1(n11526), .A2(n11524), .ZN(n19485) );
  INV_X1 U14556 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U14557 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11322), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11433) );
  OAI21_X1 U14558 ( .B1(n11434), .B2(n17623), .A(n11433), .ZN(n11435) );
  AOI22_X1 U14559 ( .A1(n17898), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14560 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11437) );
  INV_X1 U14561 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17815) );
  INV_X1 U14562 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17816) );
  OAI22_X1 U14563 ( .A1(n17891), .A2(n17815), .B1(n9666), .B2(n17816), .ZN(
        n11439) );
  AOI21_X1 U14564 ( .B1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17867), .A(
        n11439), .ZN(n11443) );
  AOI22_X1 U14565 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14566 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17933), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14567 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11440) );
  NAND4_X1 U14568 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11444) );
  INV_X1 U14569 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U14570 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11322), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U14571 ( .A1(n17894), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11445) );
  OAI211_X1 U14572 ( .C1(n16961), .C2(n16942), .A(n11446), .B(n11445), .ZN(
        n11452) );
  INV_X1 U14573 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16960) );
  INV_X1 U14574 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11448) );
  OAI22_X1 U14575 ( .A1(n11436), .A2(n16960), .B1(n17709), .B2(n11448), .ZN(
        n11451) );
  INV_X1 U14576 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17870) );
  INV_X1 U14577 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11449) );
  OAI22_X1 U14578 ( .A1(n17943), .A2(n17870), .B1(n17918), .B2(n11449), .ZN(
        n11450) );
  INV_X1 U14579 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11453) );
  OAI22_X1 U14580 ( .A1(n17799), .A2(n11453), .B1(n17941), .B2(n17740), .ZN(
        n11454) );
  AOI21_X1 U14581 ( .B1(n17020), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n11454), .ZN(n11458) );
  AOI22_X1 U14582 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14583 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U14584 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11455) );
  NAND4_X1 U14585 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11459) );
  AOI22_X1 U14586 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14587 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14588 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14589 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U14590 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11473) );
  INV_X1 U14591 ( .A(n11465), .ZN(n11488) );
  INV_X1 U14592 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17708) );
  OAI22_X1 U14593 ( .A1(n9668), .A2(n17708), .B1(n17941), .B2(n11466), .ZN(
        n11469) );
  INV_X1 U14594 ( .A(n11467), .ZN(n17709) );
  INV_X1 U14595 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17706) );
  INV_X1 U14596 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16949) );
  OAI22_X1 U14597 ( .A1(n17709), .A2(n17706), .B1(n17747), .B2(n16949), .ZN(
        n11468) );
  AOI211_X1 U14598 ( .C1(n17872), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n11469), .B(n11468), .ZN(n11471) );
  AOI22_X1 U14599 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11470) );
  OAI211_X1 U14600 ( .C1(n17950), .C2(n17711), .A(n11471), .B(n11470), .ZN(
        n11472) );
  INV_X1 U14601 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U14602 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11475) );
  NAND2_X1 U14603 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11474) );
  OAI211_X1 U14604 ( .C1(n17950), .C2(n11476), .A(n11475), .B(n11474), .ZN(
        n11477) );
  INV_X1 U14605 ( .A(n11477), .ZN(n11481) );
  AOI22_X1 U14606 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14607 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U14608 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11478) );
  NAND4_X1 U14609 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n11487) );
  AOI22_X1 U14610 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14611 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11322), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14612 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14613 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14614 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11486) );
  NOR2_X1 U14615 ( .A1(n18896), .A2(n18880), .ZN(n13811) );
  INV_X1 U14616 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14617 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11489) );
  OAI21_X1 U14618 ( .B1(n17943), .B2(n11490), .A(n11489), .ZN(n11491) );
  AOI21_X1 U14619 ( .B1(n17894), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n11491), .ZN(n11494) );
  AOI22_X1 U14620 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17912), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14621 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11492) );
  NAND3_X1 U14622 ( .A1(n11494), .A2(n11493), .A3(n11492), .ZN(n11501) );
  INV_X1 U14623 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U14624 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11495) );
  OAI21_X1 U14625 ( .B1(n17918), .B2(n17017), .A(n11495), .ZN(n11496) );
  AOI21_X1 U14626 ( .B1(n17858), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n11496), .ZN(n11499) );
  AOI22_X1 U14627 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14628 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11497) );
  NAND3_X1 U14629 ( .A1(n11499), .A2(n11498), .A3(n11497), .ZN(n11500) );
  INV_X1 U14630 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17836) );
  NAND2_X1 U14631 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14632 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11502) );
  OAI211_X1 U14633 ( .C1(n17950), .C2(n17836), .A(n11503), .B(n11502), .ZN(
        n11504) );
  INV_X1 U14634 ( .A(n11504), .ZN(n11508) );
  AOI22_X1 U14635 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14636 ( .A1(n17793), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U14637 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11505) );
  NAND4_X1 U14638 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11515) );
  AOI22_X1 U14639 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14640 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17878), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14641 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14642 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11510) );
  NAND4_X1 U14643 ( .A1(n11513), .A2(n11512), .A3(n11511), .A4(n11510), .ZN(
        n11514) );
  NOR2_X1 U14644 ( .A1(n11517), .A2(n18899), .ZN(n16908) );
  NAND3_X1 U14645 ( .A1(n11544), .A2(n13811), .A3(n16908), .ZN(n13917) );
  NAND2_X1 U14646 ( .A1(n13809), .A2(n11531), .ZN(n11541) );
  NAND2_X1 U14647 ( .A1(n18896), .A2(n18899), .ZN(n13799) );
  INV_X1 U14648 ( .A(n11531), .ZN(n18885) );
  NAND2_X1 U14649 ( .A1(n11517), .A2(n17990), .ZN(n11533) );
  INV_X1 U14650 ( .A(n11544), .ZN(n11519) );
  AOI21_X1 U14651 ( .B1(n18133), .B2(n16886), .A(n18889), .ZN(n11518) );
  NAND2_X2 U14652 ( .A1(n11523), .A2(n13800), .ZN(n18189) );
  AOI21_X1 U14653 ( .B1(n18873), .B2(n13809), .A(n11520), .ZN(n11535) );
  INV_X1 U14654 ( .A(n11526), .ZN(n11522) );
  NOR2_X1 U14655 ( .A1(n11522), .A2(n11521), .ZN(n11530) );
  INV_X1 U14656 ( .A(n13811), .ZN(n13805) );
  INV_X1 U14657 ( .A(n11523), .ZN(n11525) );
  AOI21_X1 U14658 ( .B1(n18031), .B2(n16886), .A(n11524), .ZN(n13801) );
  AOI21_X1 U14659 ( .B1(n13805), .B2(n11525), .A(n13801), .ZN(n11528) );
  NAND2_X1 U14660 ( .A1(n13809), .A2(n11526), .ZN(n13803) );
  NAND2_X1 U14661 ( .A1(n11534), .A2(n13803), .ZN(n11527) );
  OAI21_X1 U14662 ( .B1(n11528), .B2(n11531), .A(n11527), .ZN(n11529) );
  AOI21_X1 U14663 ( .B1(n11531), .B2(n11530), .A(n11529), .ZN(n11532) );
  OAI221_X1 U14664 ( .B1(n11535), .B2(n11534), .C1(n11535), .C2(n11533), .A(
        n11532), .ZN(n11539) );
  NAND2_X1 U14665 ( .A1(n11540), .A2(n11543), .ZN(n12925) );
  NAND2_X2 U14666 ( .A1(n16914), .A2(n12925), .ZN(n18851) );
  INV_X1 U14667 ( .A(n11541), .ZN(n16907) );
  AOI21_X4 U14668 ( .B1(n16907), .B2(n16914), .A(n16906), .ZN(n18746) );
  MUX2_X1 U14669 ( .A(n19311), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11572) );
  INV_X1 U14670 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14671 ( .A1(n11572), .A2(n11554), .ZN(n11547) );
  NAND2_X1 U14672 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19311), .ZN(
        n11546) );
  NAND2_X1 U14673 ( .A1(n11547), .A2(n11546), .ZN(n11560) );
  MUX2_X1 U14674 ( .A(n18865), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11559) );
  NAND2_X1 U14675 ( .A1(n11560), .A2(n11559), .ZN(n11558) );
  NAND2_X1 U14676 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18865), .ZN(
        n11548) );
  NAND2_X1 U14677 ( .A1(n11558), .A2(n11548), .ZN(n11549) );
  NAND2_X1 U14678 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17054), .ZN(
        n11550) );
  OAI21_X1 U14679 ( .B1(n11549), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11550), .ZN(n11562) );
  NAND2_X1 U14680 ( .A1(n11562), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U14681 ( .A1(n11549), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11563) );
  INV_X1 U14682 ( .A(n11550), .ZN(n11551) );
  NAND2_X1 U14683 ( .A1(n11563), .A2(n11551), .ZN(n11552) );
  NAND2_X1 U14684 ( .A1(n11553), .A2(n11552), .ZN(n11561) );
  INV_X1 U14685 ( .A(n11554), .ZN(n11571) );
  NAND2_X1 U14686 ( .A1(n16909), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U14687 ( .A1(n11571), .A2(n11555), .ZN(n11556) );
  OR2_X1 U14688 ( .A1(n11561), .A2(n11556), .ZN(n11578) );
  INV_X1 U14689 ( .A(n11572), .ZN(n11557) );
  NOR2_X1 U14690 ( .A1(n11578), .A2(n11557), .ZN(n11568) );
  OAI21_X1 U14691 ( .B1(n11560), .B2(n11559), .A(n11558), .ZN(n11577) );
  INV_X1 U14692 ( .A(n11562), .ZN(n11566) );
  NAND2_X1 U14693 ( .A1(n11563), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11565) );
  NOR2_X1 U14694 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17054), .ZN(
        n11564) );
  AOI21_X1 U14695 ( .B1(n11566), .B2(n11565), .A(n11564), .ZN(n11575) );
  NAND2_X1 U14696 ( .A1(n11570), .A2(n11575), .ZN(n11567) );
  INV_X1 U14697 ( .A(n19299), .ZN(n11569) );
  AND2_X1 U14698 ( .A1(n13809), .A2(n19471), .ZN(n13807) );
  INV_X1 U14699 ( .A(n11570), .ZN(n11574) );
  XNOR2_X1 U14700 ( .A(n11572), .B(n11571), .ZN(n11573) );
  NAND2_X1 U14701 ( .A1(n11574), .A2(n11573), .ZN(n11576) );
  OR2_X1 U14702 ( .A1(n11578), .A2(n11577), .ZN(n11579) );
  AND2_X1 U14703 ( .A1(n19294), .A2(n11579), .ZN(n19296) );
  INV_X1 U14704 ( .A(n19296), .ZN(n11580) );
  NAND2_X1 U14705 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n16879), .ZN(n19349) );
  OR2_X2 U14706 ( .A1(n17257), .A2(n13916), .ZN(n18552) );
  NAND2_X1 U14707 ( .A1(n11581), .A2(n18436), .ZN(n11641) );
  NOR2_X1 U14708 ( .A1(n11583), .A2(n11582), .ZN(n16828) );
  NOR2_X4 U14709 ( .A1(n18552), .A2(n18104), .ZN(n18426) );
  NOR2_X1 U14710 ( .A1(n18660), .A2(n11584), .ZN(n16869) );
  AND2_X1 U14711 ( .A1(n16869), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18242) );
  INV_X1 U14712 ( .A(n16846), .ZN(n16679) );
  INV_X1 U14713 ( .A(n16663), .ZN(n11586) );
  NAND2_X1 U14714 ( .A1(n13923), .A2(n16667), .ZN(n11585) );
  NAND2_X1 U14715 ( .A1(n11586), .A2(n11585), .ZN(n11592) );
  NAND2_X1 U14716 ( .A1(n11590), .A2(n11587), .ZN(n11589) );
  NAND2_X1 U14717 ( .A1(n18481), .A2(n11605), .ZN(n11588) );
  NOR2_X1 U14718 ( .A1(n16771), .A2(n11588), .ZN(n11611) );
  XOR2_X1 U14719 ( .A(n16771), .B(n11588), .Z(n11607) );
  XOR2_X1 U14720 ( .A(n18114), .B(n11589), .Z(n11603) );
  AND2_X1 U14721 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11603), .ZN(
        n11604) );
  XNOR2_X1 U14722 ( .A(n18119), .B(n11590), .ZN(n11601) );
  AND2_X1 U14723 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11601), .ZN(
        n11602) );
  INV_X1 U14724 ( .A(n11590), .ZN(n11591) );
  OAI21_X1 U14725 ( .B1(n11592), .B2(n18126), .A(n11591), .ZN(n11600) );
  INV_X1 U14726 ( .A(n16667), .ZN(n11597) );
  OAI21_X1 U14727 ( .B1(n11593), .B2(n11597), .A(n11592), .ZN(n11594) );
  AND2_X1 U14728 ( .A1(n11594), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11599) );
  NOR2_X1 U14729 ( .A1(n11594), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11595) );
  OR2_X1 U14730 ( .A1(n11599), .A2(n11595), .ZN(n18538) );
  INV_X1 U14731 ( .A(n18550), .ZN(n18556) );
  NOR2_X1 U14732 ( .A1(n16667), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18555) );
  NAND2_X1 U14733 ( .A1(n18556), .A2(n18555), .ZN(n18554) );
  MUX2_X1 U14734 ( .A(n11597), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        n11596), .Z(n11598) );
  NAND2_X1 U14735 ( .A1(n18554), .A2(n11598), .ZN(n18537) );
  XNOR2_X1 U14736 ( .A(n18805), .B(n11600), .ZN(n18528) );
  XNOR2_X1 U14737 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11601), .ZN(
        n18517) );
  NOR2_X1 U14738 ( .A1(n18518), .A2(n18517), .ZN(n18516) );
  NOR2_X1 U14739 ( .A1(n11602), .A2(n18516), .ZN(n18499) );
  XNOR2_X1 U14740 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11603), .ZN(
        n18498) );
  INV_X1 U14741 ( .A(n11605), .ZN(n18110) );
  INV_X1 U14742 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18765) );
  NOR2_X1 U14743 ( .A1(n18469), .A2(n18765), .ZN(n11606) );
  NAND2_X1 U14744 ( .A1(n11611), .A2(n11606), .ZN(n11612) );
  INV_X1 U14745 ( .A(n11606), .ZN(n11610) );
  AND2_X1 U14746 ( .A1(n11608), .A2(n11607), .ZN(n18470) );
  AOI21_X1 U14747 ( .B1(n11611), .B2(n11610), .A(n18470), .ZN(n11609) );
  OAI21_X1 U14748 ( .B1(n11611), .B2(n11610), .A(n11609), .ZN(n16767) );
  NAND2_X1 U14749 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16767), .ZN(
        n16766) );
  NOR2_X1 U14750 ( .A1(n18267), .A2(n16748), .ZN(n18563) );
  NAND3_X1 U14751 ( .A1(n16852), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n18563), .ZN(n18241) );
  AOI22_X1 U14752 ( .A1(n16679), .A2(n18426), .B1(n16796), .B2(n18557), .ZN(
        n16735) );
  NAND2_X1 U14753 ( .A1(n16735), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16732) );
  OAI211_X1 U14754 ( .C1(n18426), .C2(n18557), .A(n16732), .B(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11640) );
  NOR2_X1 U14755 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U14756 ( .A1(n19472), .A2(n19452), .ZN(n17252) );
  AND2_X1 U14757 ( .A1(n16931), .A2(n17252), .ZN(n19468) );
  INV_X1 U14758 ( .A(n19468), .ZN(n11613) );
  NAND2_X1 U14759 ( .A1(n11613), .A2(n19475), .ZN(n11614) );
  NAND2_X1 U14760 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18519) );
  INV_X1 U14761 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11621) );
  INV_X1 U14762 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18243) );
  NAND2_X1 U14763 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18278) );
  NAND3_X1 U14764 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11618) );
  NAND2_X1 U14765 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18440) );
  INV_X1 U14766 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17504) );
  NAND3_X1 U14767 ( .A1(n11615), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18429) );
  INV_X1 U14768 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17484) );
  INV_X1 U14769 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18379) );
  NAND2_X1 U14770 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11620), .ZN(
        n12903) );
  NAND2_X1 U14771 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12910), .ZN(
        n12911) );
  NAND2_X1 U14772 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12914), .ZN(
        n12913) );
  NAND2_X1 U14773 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n12916), .ZN(
        n12915) );
  INV_X1 U14774 ( .A(n12915), .ZN(n12918) );
  NAND2_X1 U14775 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12918), .ZN(
        n12917) );
  INV_X1 U14776 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18561) );
  NAND2_X1 U14777 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18248) );
  NOR2_X1 U14778 ( .A1(n18561), .A2(n12899), .ZN(n16682) );
  AOI21_X1 U14779 ( .B1(n11621), .B2(n12917), .A(n16682), .ZN(n12919) );
  NOR2_X1 U14780 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n16931), .ZN(n19488) );
  NAND2_X2 U14781 ( .A1(n19488), .A2(n19475), .ZN(n18748) );
  INV_X2 U14782 ( .A(n18748), .ZN(n18846) );
  NAND2_X1 U14783 ( .A1(n18846), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n16837) );
  INV_X1 U14784 ( .A(n16837), .ZN(n11627) );
  NOR2_X1 U14785 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19472), .ZN(n18396) );
  NOR2_X1 U14786 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19478) );
  AOI21_X1 U14787 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n19478), .ZN(n19356) );
  NAND2_X2 U14788 ( .A1(n19216), .A2(n19159), .ZN(n18906) );
  NAND2_X1 U14789 ( .A1(n11622), .A2(n18906), .ZN(n18398) );
  NAND2_X1 U14790 ( .A1(n11623), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11629) );
  INV_X1 U14791 ( .A(n11629), .ZN(n11624) );
  NAND2_X1 U14792 ( .A1(n18398), .A2(n11624), .ZN(n11628) );
  INV_X1 U14793 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11625) );
  NOR3_X1 U14794 ( .A1(n11628), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        n11625), .ZN(n11626) );
  AOI211_X1 U14795 ( .C1(n18417), .C2(n12919), .A(n11627), .B(n11626), .ZN(
        n11639) );
  NOR2_X1 U14796 ( .A1(n11628), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16730) );
  INV_X1 U14797 ( .A(n18396), .ZN(n19360) );
  OAI21_X1 U14798 ( .B1(n12916), .B2(n19360), .A(n18547), .ZN(n11631) );
  INV_X1 U14799 ( .A(n18519), .ZN(n18859) );
  AND2_X1 U14800 ( .A1(n11629), .A2(n18859), .ZN(n11630) );
  NOR2_X1 U14801 ( .A1(n11631), .A2(n11630), .ZN(n16737) );
  OR2_X1 U14802 ( .A1(n18277), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11632) );
  NAND2_X1 U14803 ( .A1(n16737), .A2(n11632), .ZN(n16726) );
  OAI21_X1 U14804 ( .B1(n16730), .B2(n16726), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11638) );
  INV_X1 U14805 ( .A(n11633), .ZN(n18724) );
  NAND2_X1 U14806 ( .A1(n18426), .A2(n18724), .ZN(n11635) );
  NAND2_X1 U14807 ( .A1(n18557), .A2(n18373), .ZN(n11634) );
  INV_X1 U14808 ( .A(n16852), .ZN(n16873) );
  NAND2_X1 U14809 ( .A1(n18563), .A2(n16844), .ZN(n16853) );
  OR2_X1 U14810 ( .A1(n16853), .A2(n16854), .ZN(n16836) );
  INV_X1 U14811 ( .A(n16836), .ZN(n11636) );
  NAND3_X1 U14812 ( .A1(n18268), .A2(n11636), .A3(n16808), .ZN(n11637) );
  NOR2_X4 U14813 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16517) );
  AND2_X4 U14814 ( .A1(n13861), .A2(n13862), .ZN(n13083) );
  AND2_X4 U14815 ( .A1(n11643), .A2(n16519), .ZN(n13077) );
  NOR2_X2 U14816 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11644) );
  AND2_X4 U14817 ( .A1(n11644), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13078) );
  AOI22_X1 U14818 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11646) );
  AND2_X2 U14819 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11914) );
  AND2_X4 U14820 ( .A1(n11914), .A2(n11785), .ZN(n11909) );
  BUF_X4 U14821 ( .A(n11659), .Z(n11908) );
  AND2_X4 U14822 ( .A1(n16579), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13076) );
  AOI22_X1 U14823 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14824 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14825 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14826 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14827 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14828 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14829 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14830 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11654) );
  NAND4_X1 U14831 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11658) );
  INV_X2 U14832 ( .A(n11691), .ZN(n11737) );
  AOI22_X1 U14833 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14834 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11662) );
  BUF_X4 U14835 ( .A(n11659), .Z(n13081) );
  AOI22_X1 U14836 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14837 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U14838 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11664) );
  AOI22_X1 U14839 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14840 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n11909), .B1(
        n9620), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14841 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14842 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14843 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11669) );
  AOI22_X1 U14844 ( .A1(n11737), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14845 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11909), .B1(
        n9620), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14846 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14847 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11670) );
  NAND4_X1 U14848 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n11674) );
  NAND2_X4 U14849 ( .A1(n11676), .A2(n11675), .ZN(n16566) );
  NAND2_X1 U14850 ( .A1(n11962), .A2(n16566), .ZN(n11767) );
  NAND2_X1 U14851 ( .A1(n11677), .A2(n11767), .ZN(n11715) );
  AOI22_X1 U14852 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14853 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14854 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14855 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11680) );
  NAND3_X1 U14856 ( .A1(n10295), .A2(n11681), .A3(n11680), .ZN(n11688) );
  AOI22_X1 U14857 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14858 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14859 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11685) );
  NAND3_X1 U14860 ( .A1(n11686), .A2(n11685), .A3(n11684), .ZN(n11687) );
  AOI22_X1 U14861 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14862 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14863 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14864 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14865 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14866 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14867 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11697) );
  NAND3_X1 U14868 ( .A1(n11699), .A2(n11698), .A3(n11697), .ZN(n11700) );
  AOI22_X1 U14869 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14870 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14871 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U14872 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NAND2_X1 U14873 ( .A1(n11706), .A2(n13875), .ZN(n11713) );
  AOI22_X1 U14874 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14875 ( .A1(n13081), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14876 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11707) );
  NAND4_X1 U14877 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11711) );
  NAND2_X1 U14878 ( .A1(n11711), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11712) );
  OAI21_X1 U14879 ( .B1(n12065), .B2(n16546), .A(n11754), .ZN(n11714) );
  NAND3_X1 U14880 ( .A1(n11715), .A2(n16542), .A3(n11714), .ZN(n11731) );
  INV_X1 U14881 ( .A(n11759), .ZN(n12305) );
  AND4_X2 U14882 ( .A1(n11716), .A2(n12065), .A3(n16566), .A4(n12305), .ZN(
        n11717) );
  NAND2_X1 U14883 ( .A1(n11717), .A2(n11744), .ZN(n11761) );
  AOI22_X1 U14884 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14885 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14886 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11718) );
  NAND4_X1 U14887 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11722) );
  NAND2_X1 U14888 ( .A1(n11722), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11730) );
  AOI22_X1 U14889 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14890 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14891 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11724) );
  NAND4_X1 U14892 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11728) );
  NAND2_X1 U14893 ( .A1(n11728), .A2(n13875), .ZN(n11729) );
  NAND2_X2 U14894 ( .A1(n11730), .A2(n11729), .ZN(n11752) );
  INV_X2 U14895 ( .A(n11752), .ZN(n16535) );
  AND3_X2 U14896 ( .A1(n11731), .A2(n11761), .A3(n16535), .ZN(n12302) );
  NAND2_X1 U14897 ( .A1(n12302), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14898 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14899 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14900 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14901 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11732) );
  NAND4_X1 U14902 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11736) );
  AOI22_X1 U14903 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13076), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14904 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14905 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13083), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14906 ( .A1(n13077), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U14907 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11742) );
  AOI21_X2 U14908 ( .B1(n12308), .B2(n12309), .A(n17153), .ZN(n11806) );
  NAND2_X1 U14909 ( .A1(n11806), .A2(n16535), .ZN(n11750) );
  NAND2_X1 U14910 ( .A1(n11745), .A2(n11744), .ZN(n12003) );
  NAND3_X1 U14911 ( .A1(n12003), .A2(n16542), .A3(n12042), .ZN(n11748) );
  NAND2_X1 U14912 ( .A1(n12022), .A2(n16549), .ZN(n12030) );
  NAND2_X1 U14913 ( .A1(n12030), .A2(n16566), .ZN(n12298) );
  NAND2_X1 U14914 ( .A1(n12298), .A2(n16546), .ZN(n11757) );
  NAND2_X1 U14916 ( .A1(n12309), .A2(n11716), .ZN(n11755) );
  AOI21_X1 U14917 ( .B1(n17153), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11758) );
  INV_X1 U14918 ( .A(n13646), .ZN(n12979) );
  INV_X1 U14919 ( .A(n11761), .ZN(n11762) );
  NOR2_X1 U14920 ( .A1(n15806), .A2(n17153), .ZN(n11764) );
  INV_X1 U14921 ( .A(n11944), .ZN(n11765) );
  NAND3_X1 U14922 ( .A1(n11716), .A2(n16542), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11795) );
  NOR2_X1 U14923 ( .A1(n11795), .A2(n11767), .ZN(n11768) );
  AND2_X4 U14924 ( .A1(n11775), .A2(n11770), .ZN(n11902) );
  AOI22_X1 U14925 ( .A1(n11902), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11769) );
  INV_X1 U14926 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13775) );
  NAND2_X1 U14927 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  INV_X1 U14928 ( .A(n12397), .ZN(n11812) );
  NAND2_X1 U14929 ( .A1(n11784), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U14930 ( .A1(n17153), .A2(n16621), .ZN(n15432) );
  NAND2_X1 U14931 ( .A1(n11778), .A2(n11777), .ZN(n11782) );
  NAND2_X1 U14932 ( .A1(n11804), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11780) );
  INV_X1 U14933 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15761) );
  AOI22_X1 U14934 ( .A1(n11902), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11779) );
  INV_X1 U14935 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12343) );
  NAND3_X1 U14936 ( .A1(n11780), .A2(n11779), .A3(n9697), .ZN(n11781) );
  NAND2_X1 U14937 ( .A1(n11787), .A2(n12836), .ZN(n11794) );
  INV_X1 U14938 ( .A(n11788), .ZN(n11789) );
  INV_X1 U14939 ( .A(n11767), .ZN(n11791) );
  NAND2_X1 U14940 ( .A1(n11794), .A2(n16506), .ZN(n11797) );
  INV_X1 U14941 ( .A(n11795), .ZN(n11796) );
  INV_X1 U14942 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11800) );
  NAND2_X1 U14943 ( .A1(n11902), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14944 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U14945 ( .A1(n11804), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14946 ( .A1(n11807), .A2(n11806), .ZN(n11808) );
  INV_X1 U14947 ( .A(n12396), .ZN(n11817) );
  INV_X1 U14948 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12347) );
  NAND2_X1 U14949 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11816) );
  AOI22_X1 U14950 ( .A1(n11902), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U14951 ( .A1(n11817), .A2(n12393), .ZN(n16231) );
  INV_X1 U14952 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U14953 ( .A1(n11899), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U14954 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11818) );
  OAI211_X1 U14955 ( .C1(n11884), .C2(n11820), .A(n11819), .B(n11818), .ZN(
        n11821) );
  AOI21_X1 U14956 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11821), .ZN(n16230) );
  INV_X1 U14957 ( .A(n16230), .ZN(n11822) );
  INV_X1 U14958 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11827) );
  NAND2_X1 U14959 ( .A1(n11899), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11826) );
  NAND2_X1 U14960 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11825) );
  OAI211_X1 U14961 ( .C1(n11884), .C2(n11827), .A(n11826), .B(n11825), .ZN(
        n11828) );
  AOI21_X1 U14962 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11828), .ZN(n13454) );
  INV_X1 U14963 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U14964 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11830) );
  AOI22_X1 U14965 ( .A1(n11902), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11829) );
  OAI211_X1 U14966 ( .C1(n9619), .C2(n12352), .A(n11830), .B(n11829), .ZN(
        n13902) );
  INV_X1 U14967 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U14968 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11832) );
  AOI22_X1 U14969 ( .A1(n11902), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11831) );
  OAI211_X1 U14970 ( .C1(n9618), .C2(n12355), .A(n11832), .B(n11831), .ZN(
        n13880) );
  INV_X1 U14971 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20243) );
  NAND2_X1 U14972 ( .A1(n11899), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U14973 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11833) );
  OAI211_X1 U14974 ( .C1(n11884), .C2(n20243), .A(n11834), .B(n11833), .ZN(
        n11835) );
  AOI21_X1 U14975 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11835), .ZN(n15698) );
  INV_X1 U14976 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20245) );
  NAND2_X1 U14977 ( .A1(n11899), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U14978 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11838) );
  OAI211_X1 U14979 ( .C1(n11884), .C2(n20245), .A(n11839), .B(n11838), .ZN(
        n11840) );
  AOI21_X1 U14980 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11840), .ZN(n13995) );
  INV_X1 U14981 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20247) );
  NAND2_X1 U14982 ( .A1(n11899), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11842) );
  NAND2_X1 U14983 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11841) );
  OAI211_X1 U14984 ( .C1(n11884), .C2(n20247), .A(n11842), .B(n11841), .ZN(
        n11843) );
  AOI21_X1 U14985 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11843), .ZN(n13907) );
  NAND2_X1 U14986 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11845) );
  AOI22_X1 U14987 ( .A1(n11902), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11844) );
  OAI211_X1 U14988 ( .C1(n11904), .C2(n12356), .A(n11845), .B(n11844), .ZN(
        n13494) );
  INV_X1 U14989 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20250) );
  NAND2_X1 U14990 ( .A1(n11899), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U14991 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11846) );
  OAI211_X1 U14992 ( .C1(n11884), .C2(n20250), .A(n11847), .B(n11846), .ZN(
        n11848) );
  AOI21_X1 U14993 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11848), .ZN(n14044) );
  INV_X1 U14994 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16131) );
  NAND2_X1 U14995 ( .A1(n11899), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U14996 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11849) );
  OAI211_X1 U14997 ( .C1(n11884), .C2(n16131), .A(n11850), .B(n11849), .ZN(
        n11851) );
  AOI21_X1 U14998 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11851), .ZN(n13477) );
  INV_X1 U14999 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15664) );
  NAND2_X1 U15000 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11853) );
  AOI22_X1 U15001 ( .A1(n11902), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11852) );
  OAI211_X1 U15002 ( .C1(n15664), .C2(n11904), .A(n11853), .B(n11852), .ZN(
        n15654) );
  INV_X1 U15003 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U15004 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11855) );
  AOI22_X1 U15005 ( .A1(n11902), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11854) );
  OAI211_X1 U15006 ( .C1(n12528), .C2(n11904), .A(n11855), .B(n11854), .ZN(
        n15641) );
  INV_X1 U15007 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U15008 ( .A1(n11899), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U15009 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11856) );
  OAI211_X1 U15010 ( .C1(n11884), .C2(n16091), .A(n11857), .B(n11856), .ZN(
        n11858) );
  AOI21_X1 U15011 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11858), .ZN(n15622) );
  INV_X1 U15012 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20257) );
  NAND2_X1 U15013 ( .A1(n11899), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U15014 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11859) );
  OAI211_X1 U15015 ( .C1(n11884), .C2(n20257), .A(n11860), .B(n11859), .ZN(
        n11861) );
  AOI21_X1 U15016 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11861), .ZN(n14254) );
  INV_X1 U15017 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U15018 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11863) );
  AOI22_X1 U15019 ( .A1(n11902), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11862) );
  OAI211_X1 U15020 ( .C1(n11904), .C2(n15596), .A(n11863), .B(n11862), .ZN(
        n15604) );
  INV_X1 U15021 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n15586) );
  NAND2_X1 U15022 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11865) );
  AOI22_X1 U15023 ( .A1(n11902), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11864) );
  OAI211_X1 U15024 ( .C1(n11904), .C2(n15586), .A(n11865), .B(n11864), .ZN(
        n12869) );
  INV_X1 U15025 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15485) );
  NAND2_X1 U15026 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11867) );
  AOI22_X1 U15027 ( .A1(n11902), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11866) );
  OAI211_X1 U15028 ( .C1(n11904), .C2(n15485), .A(n11867), .B(n11866), .ZN(
        n14366) );
  INV_X1 U15029 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15818) );
  NAND2_X1 U15030 ( .A1(n11902), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U15031 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11868) );
  OAI211_X1 U15032 ( .C1(n15818), .C2(n11904), .A(n11869), .B(n11868), .ZN(
        n11870) );
  AOI21_X1 U15033 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11870), .ZN(n15496) );
  INV_X1 U15034 ( .A(n15496), .ZN(n11888) );
  INV_X1 U15035 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15828) );
  NAND2_X1 U15036 ( .A1(n11902), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11872) );
  NAND2_X1 U15037 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11871) );
  OAI211_X1 U15038 ( .C1(n15828), .C2(n11904), .A(n11872), .B(n11871), .ZN(
        n11873) );
  AOI21_X1 U15039 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11873), .ZN(n15512) );
  INV_X1 U15040 ( .A(n15512), .ZN(n11887) );
  INV_X1 U15041 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15529) );
  NAND2_X1 U15042 ( .A1(n11902), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U15043 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11874) );
  OAI211_X1 U15044 ( .C1(n15529), .C2(n11904), .A(n11875), .B(n11874), .ZN(
        n11876) );
  AOI21_X1 U15045 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11876), .ZN(n15527) );
  INV_X1 U15046 ( .A(n15527), .ZN(n11886) );
  INV_X1 U15047 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U15048 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11878) );
  AOI22_X1 U15049 ( .A1(n11902), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11877) );
  OAI211_X1 U15050 ( .C1(n15552), .C2(n11904), .A(n11878), .B(n11877), .ZN(
        n15540) );
  INV_X1 U15051 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20264) );
  NAND2_X1 U15052 ( .A1(n11899), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U15053 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11879) );
  OAI211_X1 U15054 ( .C1(n11884), .C2(n20264), .A(n11880), .B(n11879), .ZN(
        n11881) );
  AOI21_X1 U15055 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11881), .ZN(n12746) );
  INV_X1 U15056 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20262) );
  NAND2_X1 U15057 ( .A1(n11899), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U15058 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11882) );
  OAI211_X1 U15059 ( .C1(n11884), .C2(n20262), .A(n11883), .B(n11882), .ZN(
        n11885) );
  AOI21_X1 U15060 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11885), .ZN(n14294) );
  NOR2_X1 U15061 ( .A1(n12746), .A2(n14294), .ZN(n12745) );
  AND2_X1 U15062 ( .A1(n15540), .A2(n12745), .ZN(n15524) );
  INV_X1 U15063 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U15064 ( .A1(n11902), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U15065 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11890) );
  OAI211_X1 U15066 ( .C1(n11892), .C2(n11904), .A(n11891), .B(n11890), .ZN(
        n11893) );
  AOI21_X1 U15067 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11893), .ZN(n12713) );
  INV_X1 U15068 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U15069 ( .A1(n11902), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U15070 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11894) );
  OAI211_X1 U15071 ( .C1(n15459), .C2(n11904), .A(n11895), .B(n11894), .ZN(
        n11896) );
  AOI21_X1 U15072 ( .B1(n11906), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11896), .ZN(n15457) );
  INV_X1 U15073 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U15074 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11898) );
  AOI22_X1 U15075 ( .A1(n11902), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11897) );
  OAI211_X1 U15076 ( .C1(n15444), .C2(n11904), .A(n11898), .B(n11897), .ZN(
        n12665) );
  INV_X1 U15077 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15078 ( .A1(n11902), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11901) );
  NAND2_X1 U15079 ( .A1(n11899), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11900) );
  OAI211_X1 U15080 ( .C1(n11824), .C2(n12335), .A(n11901), .B(n11900), .ZN(
        n12675) );
  INV_X1 U15081 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U15082 ( .A1(n11902), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11903) );
  OAI21_X1 U15083 ( .B1(n11904), .B2(n12840), .A(n11903), .ZN(n11905) );
  AOI21_X1 U15084 ( .B1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11906), .A(
        n11905), .ZN(n11907) );
  INV_X1 U15085 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19492) );
  NOR2_X1 U15086 ( .A1(n19492), .A2(n20231), .ZN(n20223) );
  NAND2_X1 U15087 ( .A1(n19492), .A2(n20231), .ZN(n20226) );
  INV_X1 U15088 ( .A(n20226), .ZN(n20213) );
  NOR3_X1 U15089 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20223), .A3(n20213), 
        .ZN(n20217) );
  NAND2_X1 U15090 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n17147) );
  NAND2_X1 U15091 ( .A1(n20217), .A2(n17147), .ZN(n13632) );
  OR2_X1 U15092 ( .A1(n13632), .A2(n16542), .ZN(n11968) );
  AND2_X4 U15093 ( .A1(n13207), .A2(n13875), .ZN(n13060) );
  AOI22_X1 U15095 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11930), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11913) );
  AND2_X2 U15096 ( .A1(n11908), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11969) );
  AOI22_X1 U15097 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13866), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11912) );
  AND2_X2 U15098 ( .A1(n13083), .A2(n13875), .ZN(n12104) );
  AOI22_X1 U15099 ( .A1(n12104), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11911) );
  AND2_X2 U15100 ( .A1(n13083), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12105) );
  AOI22_X1 U15101 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11910) );
  NAND4_X1 U15102 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n11920) );
  AOI22_X1 U15103 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15105 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11917) );
  AND2_X2 U15106 ( .A1(n11723), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11989) );
  INV_X1 U15107 ( .A(n13864), .ZN(n13872) );
  NOR2_X1 U15108 ( .A1(n13872), .A2(n13875), .ZN(n12005) );
  AOI22_X1 U15109 ( .A1(n11989), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11916) );
  AND2_X2 U15110 ( .A1(n13077), .A2(n13875), .ZN(n13069) );
  AND2_X2 U15111 ( .A1(n13078), .A2(n13875), .ZN(n13068) );
  AOI22_X1 U15112 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11915) );
  NAND4_X1 U15113 ( .A1(n11918), .A2(n11917), .A3(n11916), .A4(n11915), .ZN(
        n11919) );
  NAND2_X1 U15114 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20335), .ZN(
        n11945) );
  NAND2_X1 U15115 ( .A1(n11983), .A2(n11947), .ZN(n11922) );
  NAND2_X1 U15116 ( .A1(n20034), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U15117 ( .A1(n11922), .A2(n11921), .ZN(n11943) );
  XNOR2_X1 U15118 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U15119 ( .A1(n11943), .A2(n11941), .ZN(n11924) );
  NAND2_X1 U15120 ( .A1(n20325), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11923) );
  INV_X1 U15121 ( .A(n11937), .ZN(n11925) );
  XNOR2_X1 U15122 ( .A(n11938), .B(n11925), .ZN(n12011) );
  AOI22_X1 U15123 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15124 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15125 ( .A1(n9673), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U15126 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12105), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11926) );
  NAND4_X1 U15127 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11936) );
  AOI22_X1 U15128 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15129 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13069), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15130 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U15131 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U15132 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11935) );
  NAND2_X1 U15133 ( .A1(n11938), .A2(n11937), .ZN(n11940) );
  NAND2_X1 U15134 ( .A1(n20317), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15135 ( .A1(n11940), .A2(n11939), .ZN(n11957) );
  NAND2_X1 U15136 ( .A1(n16605), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11958) );
  MUX2_X1 U15137 ( .A(n12451), .B(n12009), .S(n12609), .Z(n12348) );
  INV_X1 U15138 ( .A(n11941), .ZN(n11942) );
  XNOR2_X1 U15139 ( .A(n11943), .B(n11942), .ZN(n12010) );
  NAND2_X1 U15140 ( .A1(n11944), .A2(n12010), .ZN(n11950) );
  OAI21_X1 U15141 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20335), .A(
        n11945), .ZN(n12017) );
  INV_X1 U15142 ( .A(n12017), .ZN(n11982) );
  NAND2_X1 U15143 ( .A1(n11983), .A2(n11982), .ZN(n11946) );
  NAND2_X1 U15144 ( .A1(n12836), .A2(n11946), .ZN(n11949) );
  XNOR2_X1 U15145 ( .A(n11983), .B(n11945), .ZN(n12013) );
  OAI211_X1 U15146 ( .C1(n15806), .C2(n11982), .A(n16535), .B(n12013), .ZN(
        n11948) );
  NOR2_X1 U15147 ( .A1(n15425), .A2(n12004), .ZN(n11952) );
  MUX2_X1 U15148 ( .A(n11952), .B(n12836), .S(n12010), .Z(n11953) );
  OAI21_X1 U15149 ( .B1(n11954), .B2(n11953), .A(n12011), .ZN(n11955) );
  INV_X1 U15150 ( .A(n12009), .ZN(n11960) );
  NOR2_X1 U15151 ( .A1(n16605), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11956) );
  AOI21_X1 U15152 ( .B1(n12836), .B2(n11960), .A(n11964), .ZN(n11961) );
  NAND2_X1 U15153 ( .A1(n11966), .A2(n16535), .ZN(n11963) );
  NAND2_X1 U15154 ( .A1(n11963), .A2(n11962), .ZN(n11967) );
  NAND2_X1 U15155 ( .A1(n16592), .A2(n12042), .ZN(n13681) );
  MUX2_X1 U15156 ( .A(n11968), .B(n11967), .S(n13681), .Z(n12037) );
  AOI22_X1 U15157 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15158 ( .A1(n11989), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15159 ( .A1(n9673), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15160 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12105), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11970) );
  NAND4_X1 U15161 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n11981) );
  AOI22_X1 U15162 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15163 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15164 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15165 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11976) );
  NAND4_X1 U15166 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11980) );
  MUX2_X1 U15167 ( .A(n13732), .B(n11982), .S(n12609), .Z(n12436) );
  INV_X1 U15168 ( .A(n12436), .ZN(n11999) );
  INV_X1 U15169 ( .A(n11983), .ZN(n11998) );
  AOI22_X1 U15170 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11930), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15171 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13866), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15172 ( .A1(n12104), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15173 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11985) );
  NAND4_X1 U15174 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(
        n11995) );
  AOI22_X1 U15175 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15176 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15177 ( .A1(n11989), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15178 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U15179 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11994) );
  INV_X1 U15180 ( .A(n12010), .ZN(n11996) );
  NAND2_X1 U15181 ( .A1(n12609), .A2(n11996), .ZN(n11997) );
  OAI21_X1 U15182 ( .B1(n11999), .B2(n11998), .A(n12340), .ZN(n12001) );
  NAND2_X1 U15183 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  NAND2_X1 U15184 ( .A1(n12002), .A2(n12015), .ZN(n20342) );
  INV_X1 U15185 ( .A(n12003), .ZN(n16603) );
  AND2_X1 U15186 ( .A1(n12004), .A2(n11752), .ZN(n12021) );
  NAND2_X1 U15187 ( .A1(n16603), .A2(n12021), .ZN(n12650) );
  INV_X1 U15188 ( .A(n12005), .ZN(n12006) );
  AND2_X1 U15189 ( .A1(n12006), .A2(n16605), .ZN(n13641) );
  INV_X1 U15190 ( .A(n12058), .ZN(n12007) );
  NAND2_X1 U15191 ( .A1(n13641), .A2(n12007), .ZN(n12008) );
  INV_X1 U15192 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n16600) );
  NAND2_X1 U15193 ( .A1(n12008), .A2(n16600), .ZN(n20326) );
  NAND3_X1 U15194 ( .A1(n12011), .A2(n12010), .A3(n12009), .ZN(n12016) );
  INV_X1 U15195 ( .A(n12016), .ZN(n12012) );
  NAND2_X1 U15196 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  OAI21_X1 U15197 ( .B1(n12017), .B2(n12016), .A(n16591), .ZN(n12018) );
  INV_X1 U15198 ( .A(n12018), .ZN(n12019) );
  MUX2_X1 U15199 ( .A(n20326), .B(n12019), .S(n16621), .Z(n20338) );
  NAND3_X1 U15200 ( .A1(n16603), .A2(n15806), .A3(n20338), .ZN(n12020) );
  NAND2_X1 U15201 ( .A1(n16591), .A2(n17147), .ZN(n13223) );
  INV_X1 U15202 ( .A(n16566), .ZN(n13230) );
  OAI21_X1 U15203 ( .B1(n12022), .B2(n13230), .A(n12021), .ZN(n12300) );
  INV_X1 U15204 ( .A(n13632), .ZN(n13537) );
  NAND3_X1 U15205 ( .A1(n12023), .A2(n13537), .A3(n16591), .ZN(n12027) );
  NAND2_X1 U15206 ( .A1(n11752), .A2(n16566), .ZN(n12025) );
  OAI211_X1 U15207 ( .C1(n11767), .C2(n15806), .A(n16542), .B(n12025), .ZN(
        n12026) );
  NAND4_X1 U15208 ( .A1(n12300), .A2(n12027), .A3(n12303), .A4(n12026), .ZN(
        n12033) );
  NAND2_X1 U15209 ( .A1(n12296), .A2(n16542), .ZN(n12029) );
  NAND2_X1 U15210 ( .A1(n12028), .A2(n12029), .ZN(n12031) );
  NAND2_X1 U15211 ( .A1(n12031), .A2(n12030), .ZN(n12032) );
  NOR2_X1 U15212 ( .A1(n12033), .A2(n12032), .ZN(n13637) );
  OAI21_X1 U15213 ( .B1(n12034), .B2(n13223), .A(n13637), .ZN(n12035) );
  NAND3_X1 U15214 ( .A1(n16621), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17160) );
  NAND2_X1 U15215 ( .A1(n12038), .A2(n12004), .ZN(n12039) );
  INV_X1 U15216 ( .A(n16506), .ZN(n12292) );
  NAND2_X1 U15217 ( .A1(n12292), .A2(n12024), .ZN(n13870) );
  NAND2_X1 U15218 ( .A1(n12039), .A2(n13870), .ZN(n12040) );
  NOR2_X1 U15219 ( .A1(n14463), .A2(n17133), .ZN(n12339) );
  NAND2_X1 U15220 ( .A1(n12046), .A2(n12065), .ZN(n12116) );
  NAND2_X1 U15221 ( .A1(n13732), .A2(n12041), .ZN(n12044) );
  INV_X1 U15222 ( .A(n12066), .ZN(n13229) );
  NAND2_X1 U15223 ( .A1(n12042), .A2(n20318), .ZN(n12281) );
  NAND2_X1 U15224 ( .A1(n13229), .A2(n12282), .ZN(n12072) );
  MUX2_X1 U15225 ( .A(n16566), .B(n20335), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12043) );
  NAND3_X1 U15226 ( .A1(n12044), .A2(n12072), .A3(n12043), .ZN(n13733) );
  NAND2_X1 U15227 ( .A1(n12090), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12051) );
  INV_X1 U15228 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U15229 ( .A1(n15806), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12047) );
  OAI211_X1 U15230 ( .C1(n16566), .C2(n12048), .A(n12047), .B(n20318), .ZN(
        n12049) );
  INV_X1 U15231 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U15232 ( .A1(n12051), .A2(n12050), .ZN(n13735) );
  NAND2_X1 U15233 ( .A1(n13733), .A2(n13735), .ZN(n13734) );
  INV_X1 U15234 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20232) );
  NOR2_X1 U15235 ( .A1(n16566), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12052) );
  XNOR2_X1 U15236 ( .A(n13734), .B(n12069), .ZN(n13851) );
  AOI22_X1 U15237 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15238 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12105), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15239 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15240 ( .A1(n12104), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12054) );
  NAND4_X1 U15241 ( .A1(n12057), .A2(n12056), .A3(n12055), .A4(n12054), .ZN(
        n12064) );
  AOI22_X1 U15242 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15243 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15244 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15245 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U15246 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12063) );
  OR2_X2 U15247 ( .A1(n12064), .A2(n12063), .ZN(n12616) );
  INV_X1 U15248 ( .A(n12345), .ZN(n12067) );
  AOI22_X1 U15249 ( .A1(n12067), .A2(n12004), .B1(n12066), .B2(n16566), .ZN(
        n12068) );
  NAND2_X1 U15250 ( .A1(n13851), .A2(n13850), .ZN(n13849) );
  INV_X1 U15251 ( .A(n12069), .ZN(n12070) );
  NAND2_X1 U15252 ( .A1(n13734), .A2(n12070), .ZN(n12071) );
  NAND2_X1 U15253 ( .A1(n13849), .A2(n12071), .ZN(n12078) );
  NAND2_X1 U15254 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12073) );
  OAI211_X1 U15255 ( .C1(n12116), .C2(n12619), .A(n12073), .B(n12072), .ZN(
        n12076) );
  XNOR2_X1 U15256 ( .A(n12078), .B(n12076), .ZN(n13935) );
  NAND2_X1 U15257 ( .A1(n12285), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15258 ( .A1(n12288), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12074) );
  AND2_X1 U15259 ( .A1(n12075), .A2(n12074), .ZN(n13934) );
  INV_X1 U15260 ( .A(n12076), .ZN(n12077) );
  NAND2_X1 U15261 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  NAND2_X1 U15262 ( .A1(n13937), .A2(n12079), .ZN(n15741) );
  INV_X1 U15263 ( .A(n15741), .ZN(n12086) );
  INV_X1 U15264 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16476) );
  NOR2_X1 U15265 ( .A1(n12281), .A2(n16476), .ZN(n12080) );
  AOI21_X1 U15266 ( .B1(n12041), .B2(n12081), .A(n12080), .ZN(n12084) );
  AOI22_X1 U15267 ( .A1(n12288), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12083) );
  NAND2_X1 U15268 ( .A1(n12285), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U15269 ( .A1(n12086), .A2(n12085), .ZN(n15739) );
  NAND2_X1 U15270 ( .A1(n12285), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15271 ( .A1(n12288), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U15272 ( .A1(n12041), .A2(n12451), .ZN(n12087) );
  NAND2_X1 U15273 ( .A1(n12285), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15274 ( .A1(n12288), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15275 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15276 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15277 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15278 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12091) );
  NAND4_X1 U15279 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12100) );
  AOI22_X1 U15280 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15281 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15282 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15283 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15284 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12099) );
  NOR2_X1 U15285 ( .A1(n12100), .A2(n12099), .ZN(n12466) );
  INV_X1 U15286 ( .A(n12466), .ZN(n12349) );
  NAND2_X1 U15287 ( .A1(n12041), .A2(n12349), .ZN(n12101) );
  AOI22_X1 U15288 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11930), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15289 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15290 ( .A1(n12104), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15291 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12105), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12106) );
  NAND4_X1 U15292 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12115) );
  AOI22_X1 U15293 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15294 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15295 ( .A1(n11989), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15296 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12110) );
  NAND4_X1 U15297 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12114) );
  INV_X1 U15298 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20239) );
  AOI22_X1 U15299 ( .A1(n12288), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12117) );
  OAI21_X1 U15300 ( .B1(n12280), .B2(n20239), .A(n12117), .ZN(n13752) );
  NAND2_X1 U15301 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U15302 ( .A1(n11989), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12120) );
  NAND2_X1 U15303 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12119) );
  NAND2_X1 U15304 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12118) );
  INV_X1 U15305 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12125) );
  INV_X1 U15306 ( .A(n13060), .ZN(n12124) );
  INV_X1 U15307 ( .A(n13067), .ZN(n12123) );
  INV_X1 U15308 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12122) );
  OAI22_X1 U15309 ( .A1(n12125), .A2(n12124), .B1(n12123), .B2(n12122), .ZN(
        n12132) );
  INV_X1 U15310 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12130) );
  INV_X1 U15311 ( .A(n12126), .ZN(n12129) );
  INV_X1 U15312 ( .A(n13068), .ZN(n12128) );
  INV_X1 U15313 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12127) );
  OAI22_X1 U15314 ( .A1(n12130), .A2(n12129), .B1(n12128), .B2(n12127), .ZN(
        n12131) );
  NOR2_X1 U15315 ( .A1(n12132), .A2(n12131), .ZN(n12143) );
  NAND2_X1 U15316 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15317 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U15318 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12134) );
  NAND2_X1 U15319 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12133) );
  NAND2_X1 U15320 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U15321 ( .A1(n12104), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U15322 ( .A1(n9673), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12138) );
  NAND2_X1 U15323 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12137) );
  NAND2_X1 U15324 ( .A1(n12041), .A2(n12644), .ZN(n12145) );
  INV_X1 U15325 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20241) );
  AOI22_X1 U15326 ( .A1(n12288), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12146) );
  OAI21_X1 U15327 ( .B1(n12280), .B2(n20241), .A(n12146), .ZN(n13756) );
  NAND2_X1 U15328 ( .A1(n13757), .A2(n13756), .ZN(n13748) );
  INV_X1 U15329 ( .A(n13748), .ZN(n12161) );
  NAND2_X1 U15330 ( .A1(n12285), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15331 ( .A1(n12288), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15332 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15333 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13866), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15334 ( .A1(n12104), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15335 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15336 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12156) );
  AOI22_X1 U15337 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15338 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15339 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15340 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U15341 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12155) );
  NAND2_X1 U15342 ( .A1(n12041), .A2(n13991), .ZN(n12157) );
  NAND2_X1 U15343 ( .A1(n12161), .A2(n12160), .ZN(n13747) );
  NAND2_X1 U15344 ( .A1(n12285), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15345 ( .A1(n12288), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15346 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15347 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15348 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15349 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12162) );
  NAND4_X1 U15350 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n12171) );
  AOI22_X1 U15351 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15352 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15353 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15354 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15355 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12170) );
  OR2_X1 U15356 ( .A1(n12171), .A2(n12170), .ZN(n13993) );
  NAND2_X1 U15357 ( .A1(n12041), .A2(n13993), .ZN(n12172) );
  NAND2_X1 U15358 ( .A1(n12285), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15359 ( .A1(n12288), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15360 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15361 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15362 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15363 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U15364 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12184) );
  AOI22_X1 U15365 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15366 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15367 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15368 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15369 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  NAND2_X1 U15370 ( .A1(n12041), .A2(n13912), .ZN(n12185) );
  INV_X1 U15371 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20254) );
  AOI22_X1 U15372 ( .A1(n12288), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15373 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13060), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15374 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15375 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11984), .B1(
        n12105), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15376 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12104), .B1(
        n13866), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15377 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12197) );
  AOI22_X1 U15378 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12126), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15379 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15380 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15381 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U15382 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12196) );
  OR2_X1 U15383 ( .A1(n12197), .A2(n12196), .ZN(n15874) );
  NAND2_X1 U15384 ( .A1(n12041), .A2(n15874), .ZN(n12198) );
  OAI211_X1 U15385 ( .C1(n12280), .C2(n20254), .A(n12199), .B(n12198), .ZN(
        n14146) );
  INV_X1 U15386 ( .A(n14146), .ZN(n12239) );
  NAND2_X1 U15387 ( .A1(n12285), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15388 ( .A1(n12288), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15389 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15390 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15391 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15392 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U15393 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12209) );
  AOI22_X1 U15394 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15395 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15396 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15397 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15398 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  OR2_X1 U15399 ( .A1(n12209), .A2(n12208), .ZN(n15885) );
  NAND2_X1 U15400 ( .A1(n12041), .A2(n15885), .ZN(n12210) );
  AND3_X1 U15401 ( .A1(n12212), .A2(n12211), .A3(n12210), .ZN(n13481) );
  NAND2_X1 U15402 ( .A1(n12285), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15403 ( .A1(n12288), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15404 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15405 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15406 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15407 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12213) );
  NAND4_X1 U15408 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12222) );
  AOI22_X1 U15409 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15410 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15411 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15412 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15413 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12221) );
  OR2_X1 U15414 ( .A1(n12222), .A2(n12221), .ZN(n14050) );
  NAND2_X1 U15415 ( .A1(n12041), .A2(n14050), .ZN(n12223) );
  INV_X1 U15416 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n16119) );
  AOI22_X1 U15417 ( .A1(n12288), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15418 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15419 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12105), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15420 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15421 ( .A1(n9673), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12226) );
  NAND4_X1 U15422 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12235) );
  AOI22_X1 U15423 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15424 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15425 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15426 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12230) );
  NAND4_X1 U15427 ( .A1(n12233), .A2(n12232), .A3(n12231), .A4(n12230), .ZN(
        n12234) );
  OR2_X1 U15428 ( .A1(n12235), .A2(n12234), .ZN(n15879) );
  NAND2_X1 U15429 ( .A1(n12041), .A2(n15879), .ZN(n12236) );
  OAI211_X1 U15430 ( .C1(n12280), .C2(n16119), .A(n12237), .B(n12236), .ZN(
        n12238) );
  INV_X1 U15431 ( .A(n12238), .ZN(n14089) );
  NOR2_X1 U15432 ( .A1(n12239), .A2(n14086), .ZN(n12252) );
  INV_X1 U15433 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U15434 ( .A1(n12288), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15435 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15436 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15437 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15438 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15439 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12249) );
  AOI22_X1 U15440 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15441 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15442 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15443 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15444 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12248) );
  NAND2_X1 U15445 ( .A1(n12041), .A2(n14011), .ZN(n12250) );
  OAI211_X1 U15446 ( .C1(n12280), .C2(n13488), .A(n12251), .B(n12250), .ZN(
        n13491) );
  AND2_X1 U15447 ( .A1(n12252), .A2(n13491), .ZN(n12253) );
  NAND2_X1 U15448 ( .A1(n12285), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15449 ( .A1(n12288), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12254) );
  NAND2_X1 U15450 ( .A1(n12285), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12259) );
  INV_X2 U15451 ( .A(n12279), .ZN(n12288) );
  AOI22_X1 U15452 ( .A1(n12288), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12258) );
  INV_X1 U15453 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20260) );
  AOI22_X1 U15454 ( .A1(n12288), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12260) );
  OAI21_X1 U15455 ( .B1(n12280), .B2(n20260), .A(n12260), .ZN(n12876) );
  INV_X1 U15456 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U15457 ( .A1(n12288), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12261) );
  OAI21_X1 U15458 ( .B1(n12280), .B2(n16074), .A(n12261), .ZN(n15590) );
  AND2_X1 U15459 ( .A1(n12876), .A2(n15590), .ZN(n12262) );
  AOI22_X1 U15460 ( .A1(n12288), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12263) );
  OAI21_X1 U15461 ( .B1(n12280), .B2(n20262), .A(n12263), .ZN(n14295) );
  NAND2_X1 U15462 ( .A1(n12285), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15463 ( .A1(n12288), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12264) );
  AND2_X1 U15464 ( .A1(n12265), .A2(n12264), .ZN(n13253) );
  NAND2_X1 U15465 ( .A1(n12285), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15466 ( .A1(n12288), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12266) );
  AND2_X1 U15467 ( .A1(n12267), .A2(n12266), .ZN(n15542) );
  INV_X1 U15468 ( .A(n15542), .ZN(n12268) );
  NAND2_X1 U15469 ( .A1(n12285), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15470 ( .A1(n12288), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12269) );
  NAND2_X1 U15471 ( .A1(n12285), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15472 ( .A1(n12288), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U15473 ( .A1(n12272), .A2(n12271), .ZN(n15507) );
  NAND2_X1 U15474 ( .A1(n12285), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15475 ( .A1(n12288), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12273) );
  AND2_X1 U15476 ( .A1(n12274), .A2(n12273), .ZN(n15491) );
  NAND2_X1 U15477 ( .A1(n12285), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15478 ( .A1(n12288), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12275) );
  AND2_X1 U15479 ( .A1(n12276), .A2(n12275), .ZN(n14371) );
  NAND2_X1 U15480 ( .A1(n12285), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15481 ( .A1(n12288), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U15482 ( .A1(n12278), .A2(n12277), .ZN(n14416) );
  INV_X1 U15483 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12595) );
  INV_X1 U15484 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20279) );
  INV_X1 U15485 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13687) );
  OAI222_X1 U15486 ( .A1(n12595), .A2(n12281), .B1(n20279), .B2(n12280), .C1(
        n12279), .C2(n13687), .ZN(n12659) );
  NAND2_X1 U15487 ( .A1(n12285), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15488 ( .A1(n12288), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U15489 ( .A1(n12284), .A2(n12283), .ZN(n15452) );
  AND2_X1 U15490 ( .A1(n12659), .A2(n15452), .ZN(n12660) );
  AOI222_X1 U15491 ( .A1(n12285), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n12288), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n12282), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12695) );
  INV_X1 U15492 ( .A(n12695), .ZN(n12286) );
  AND2_X1 U15493 ( .A1(n12660), .A2(n12286), .ZN(n12287) );
  AOI222_X1 U15494 ( .A1(n12285), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12288), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12282), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12289) );
  INV_X1 U15495 ( .A(n12289), .ZN(n12290) );
  NAND2_X1 U15496 ( .A1(n9739), .A2(n12292), .ZN(n13859) );
  OAI21_X1 U15497 ( .B1(n12004), .B2(n12291), .A(n13859), .ZN(n12293) );
  NAND2_X1 U15498 ( .A1(n12651), .A2(n12293), .ZN(n19648) );
  INV_X1 U15499 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13456) );
  INV_X1 U15500 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19660) );
  NOR2_X1 U15501 ( .A1(n13456), .A2(n19660), .ZN(n13453) );
  INV_X1 U15502 ( .A(n13453), .ZN(n12321) );
  NAND3_X1 U15503 ( .A1(n12342), .A2(n12004), .A3(n16542), .ZN(n12294) );
  NAND2_X1 U15504 ( .A1(n12651), .A2(n16594), .ZN(n19683) );
  NAND2_X1 U15505 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19675) );
  INV_X1 U15506 ( .A(n19675), .ZN(n12295) );
  NAND2_X1 U15507 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12295), .ZN(
        n19682) );
  NOR2_X1 U15508 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12295), .ZN(
        n12320) );
  INV_X1 U15509 ( .A(n12296), .ZN(n12297) );
  OR2_X1 U15510 ( .A1(n12298), .A2(n12297), .ZN(n12299) );
  NAND2_X1 U15511 ( .A1(n12299), .A2(n15806), .ZN(n16507) );
  NAND2_X1 U15512 ( .A1(n16507), .A2(n12300), .ZN(n12301) );
  NAND2_X1 U15513 ( .A1(n12301), .A2(n16546), .ZN(n12317) );
  INV_X1 U15514 ( .A(n12302), .ZN(n12315) );
  NAND2_X1 U15515 ( .A1(n12303), .A2(n16549), .ZN(n12307) );
  INV_X1 U15516 ( .A(n15430), .ZN(n12306) );
  AOI22_X1 U15517 ( .A1(n12307), .A2(n12306), .B1(n11752), .B2(n12305), .ZN(
        n12314) );
  INV_X1 U15518 ( .A(n12308), .ZN(n12310) );
  NAND3_X1 U15519 ( .A1(n12310), .A2(n12024), .A3(n12309), .ZN(n12313) );
  NAND2_X1 U15520 ( .A1(n12311), .A2(n12312), .ZN(n13227) );
  AND4_X1 U15521 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n13227), .ZN(
        n12316) );
  NAND2_X1 U15522 ( .A1(n16571), .A2(n12309), .ZN(n12319) );
  NAND2_X1 U15523 ( .A1(n12651), .A2(n12319), .ZN(n14264) );
  NAND2_X1 U15524 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16464), .ZN(
        n17135) );
  INV_X1 U15525 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16457) );
  INV_X1 U15526 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16451) );
  NOR2_X1 U15527 ( .A1(n16457), .A2(n16451), .ZN(n16450) );
  INV_X1 U15528 ( .A(n16450), .ZN(n12322) );
  AND2_X1 U15529 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16375) );
  AND2_X1 U15530 ( .A1(n16375), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14257) );
  NAND2_X1 U15531 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14258) );
  AND3_X1 U15532 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U15533 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n14262), .ZN(
        n12323) );
  NOR2_X1 U15534 ( .A1(n14258), .A2(n12323), .ZN(n12324) );
  NAND2_X1 U15535 ( .A1(n14257), .A2(n12324), .ZN(n16334) );
  INV_X1 U15536 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16068) );
  INV_X1 U15537 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16306) );
  NAND2_X1 U15538 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16305) );
  NOR4_X1 U15539 ( .A1(n16334), .A2(n16068), .A3(n16306), .A4(n16305), .ZN(
        n13255) );
  INV_X1 U15540 ( .A(n13255), .ZN(n12325) );
  AND2_X1 U15541 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12332) );
  INV_X1 U15542 ( .A(n12332), .ZN(n16308) );
  AND2_X1 U15543 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12334) );
  NAND2_X1 U15544 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12376) );
  INV_X1 U15545 ( .A(n12376), .ZN(n12662) );
  NAND2_X1 U15546 ( .A1(n12662), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12696) );
  NOR3_X1 U15547 ( .A1(n12696), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12335), .ZN(n12337) );
  OR2_X1 U15548 ( .A1(n20313), .A2(n15432), .ZN(n12327) );
  INV_X2 U15549 ( .A(n19553), .ZN(n16032) );
  INV_X1 U15550 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12326) );
  NOR2_X1 U15551 ( .A1(n16032), .A2(n12326), .ZN(n12945) );
  INV_X1 U15552 ( .A(n14264), .ZN(n12328) );
  INV_X1 U15553 ( .A(n12327), .ZN(n19527) );
  NOR2_X1 U15554 ( .A1(n12651), .A2(n19527), .ZN(n16489) );
  AOI21_X1 U15555 ( .B1(n12328), .B2(n19675), .A(n16489), .ZN(n19662) );
  INV_X1 U15556 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12622) );
  NAND2_X1 U15557 ( .A1(n12328), .A2(n12622), .ZN(n19676) );
  INV_X1 U15558 ( .A(n19683), .ZN(n14261) );
  NAND3_X1 U15559 ( .A1(n14261), .A2(n12622), .A3(n19675), .ZN(n19680) );
  NAND3_X1 U15560 ( .A1(n19662), .A2(n19676), .A3(n19680), .ZN(n16477) );
  NOR2_X1 U15561 ( .A1(n16408), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12329) );
  NOR2_X1 U15562 ( .A1(n16477), .A2(n12329), .ZN(n19659) );
  OR2_X1 U15563 ( .A1(n16408), .A2(n13453), .ZN(n12330) );
  NAND2_X1 U15564 ( .A1(n19659), .A2(n12330), .ZN(n16463) );
  NOR2_X1 U15565 ( .A1(n16408), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12331) );
  NAND2_X1 U15566 ( .A1(n10023), .A2(n16408), .ZN(n12333) );
  INV_X1 U15567 ( .A(n12333), .ZN(n12336) );
  AND2_X1 U15568 ( .A1(n13255), .A2(n12332), .ZN(n12647) );
  OAI21_X1 U15569 ( .B1(n12334), .B2(n12336), .A(n16283), .ZN(n16270) );
  NAND2_X1 U15570 ( .A1(n12365), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12341) );
  NAND3_X1 U15571 ( .A1(n12365), .A2(n12343), .A3(n11800), .ZN(n12344) );
  INV_X1 U15572 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19574) );
  MUX2_X1 U15573 ( .A(n19574), .B(n12348), .S(n12342), .Z(n12442) );
  INV_X1 U15574 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12350) );
  MUX2_X1 U15575 ( .A(n12350), .B(n12349), .S(n12342), .Z(n12447) );
  INV_X1 U15576 ( .A(n12478), .ZN(n12351) );
  MUX2_X1 U15577 ( .A(n12352), .B(n12351), .S(n12342), .Z(n12479) );
  MUX2_X1 U15578 ( .A(n12355), .B(n12644), .S(n12342), .Z(n12483) );
  NAND2_X1 U15579 ( .A1(n16554), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12486) );
  INV_X1 U15580 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12356) );
  INV_X1 U15581 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12534) );
  NAND2_X1 U15582 ( .A1(n12356), .A2(n12534), .ZN(n12357) );
  NOR2_X1 U15583 ( .A1(n12357), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U15584 ( .A1(n16554), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12541) );
  INV_X1 U15585 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12360) );
  NOR2_X1 U15586 ( .A1(n12342), .A2(n12360), .ZN(n12544) );
  OAI21_X1 U15587 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n16554), .ZN(n12361) );
  NAND2_X1 U15588 ( .A1(n16554), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12362) );
  INV_X1 U15589 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12363) );
  NOR2_X1 U15590 ( .A1(n12342), .A2(n12363), .ZN(n12523) );
  NOR2_X1 U15591 ( .A1(n12342), .A2(n15596), .ZN(n12514) );
  NAND2_X1 U15592 ( .A1(n16554), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12511) );
  OR2_X1 U15593 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n12364) );
  AND2_X1 U15594 ( .A1(n16554), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U15595 ( .A1(n16554), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U15596 ( .A1(n16554), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12706) );
  AND2_X1 U15597 ( .A1(n16554), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12374) );
  NOR2_X2 U15598 ( .A1(n12373), .A2(n12374), .ZN(n12372) );
  NAND2_X1 U15599 ( .A1(n16554), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15600 ( .A1(n12372), .A2(n12593), .ZN(n12371) );
  INV_X1 U15601 ( .A(n12371), .ZN(n12367) );
  INV_X1 U15602 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12366) );
  NAND2_X1 U15603 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  INV_X1 U15604 ( .A(n12369), .ZN(n12858) );
  NAND2_X1 U15605 ( .A1(n12369), .A2(n12644), .ZN(n12601) );
  NAND2_X1 U15606 ( .A1(n16554), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12370) );
  XNOR2_X1 U15607 ( .A(n12371), .B(n12370), .ZN(n12834) );
  AOI21_X1 U15608 ( .B1(n12834), .B2(n12644), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12600) );
  INV_X1 U15609 ( .A(n12372), .ZN(n12594) );
  NAND2_X1 U15610 ( .A1(n12373), .A2(n12374), .ZN(n12375) );
  NAND2_X1 U15611 ( .A1(n16021), .A2(n12376), .ZN(n12391) );
  INV_X1 U15612 ( .A(n12377), .ZN(n15481) );
  NAND2_X1 U15613 ( .A1(n15481), .A2(n12644), .ZN(n12586) );
  XNOR2_X1 U15614 ( .A(n12586), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14363) );
  NAND2_X1 U15615 ( .A1(n16554), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12379) );
  MUX2_X1 U15616 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n12379), .S(n12386), .Z(
        n12380) );
  AND2_X1 U15617 ( .A1(n12380), .A2(n12492), .ZN(n15503) );
  NAND2_X1 U15618 ( .A1(n15503), .A2(n12644), .ZN(n12381) );
  INV_X1 U15619 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16286) );
  NAND2_X1 U15620 ( .A1(n12381), .A2(n16286), .ZN(n16028) );
  INV_X1 U15621 ( .A(n12382), .ZN(n12385) );
  AND2_X1 U15622 ( .A1(n16554), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12384) );
  INV_X1 U15623 ( .A(n12492), .ZN(n12383) );
  AOI21_X1 U15624 ( .B1(n12385), .B2(n12384), .A(n12383), .ZN(n12387) );
  INV_X1 U15625 ( .A(n12582), .ZN(n12389) );
  INV_X1 U15626 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U15627 ( .A1(n12389), .A2(n12388), .ZN(n16038) );
  AND2_X1 U15628 ( .A1(n16028), .A2(n16038), .ZN(n12390) );
  AND2_X1 U15629 ( .A1(n14363), .A2(n12390), .ZN(n12704) );
  AOI22_X1 U15630 ( .A1(n11784), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n12392), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15631 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n9606), .B1(
        n12453), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12410) );
  AND2_X2 U15632 ( .A1(n12411), .A2(n12406), .ZN(n12458) );
  INV_X1 U15633 ( .A(n13865), .ZN(n12405) );
  INV_X1 U15634 ( .A(n12403), .ZN(n12404) );
  AND2_X2 U15635 ( .A1(n12405), .A2(n12404), .ZN(n12412) );
  AND2_X2 U15636 ( .A1(n12412), .A2(n12415), .ZN(n12457) );
  AOI22_X1 U15637 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12458), .B1(
        n12457), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12409) );
  AND2_X2 U15638 ( .A1(n13865), .A2(n16572), .ZN(n12416) );
  AND2_X2 U15639 ( .A1(n12412), .A2(n12406), .ZN(n12459) );
  AOI22_X1 U15640 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12452), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15641 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n16529), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12407) );
  AND2_X2 U15642 ( .A1(n12412), .A2(n12413), .ZN(n19843) );
  AND2_X2 U15643 ( .A1(n12412), .A2(n12414), .ZN(n12454) );
  AOI22_X1 U15644 ( .A1(n12454), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12418) );
  AND2_X2 U15645 ( .A1(n12416), .A2(n12415), .ZN(n12460) );
  AOI22_X1 U15646 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19934), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15647 ( .A1(n12421), .A2(n12004), .ZN(n12422) );
  NAND2_X1 U15648 ( .A1(n19685), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12424) );
  NAND2_X1 U15649 ( .A1(n12459), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12423) );
  NAND3_X1 U15650 ( .A1(n12616), .A2(n13732), .A3(n12004), .ZN(n12620) );
  NAND2_X1 U15651 ( .A1(n12620), .A2(n12619), .ZN(n12425) );
  NAND2_X1 U15652 ( .A1(n12427), .A2(n12426), .ZN(n12428) );
  INV_X1 U15653 ( .A(n12429), .ZN(n12435) );
  INV_X1 U15654 ( .A(n12430), .ZN(n12431) );
  NAND2_X1 U15655 ( .A1(n12435), .A2(n12431), .ZN(n12432) );
  NAND2_X1 U15656 ( .A1(n12444), .A2(n12432), .ZN(n15738) );
  NAND2_X1 U15657 ( .A1(n12433), .A2(n12438), .ZN(n12434) );
  NAND2_X1 U15658 ( .A1(n12435), .A2(n12434), .ZN(n15754) );
  XNOR2_X1 U15659 ( .A(n15754), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14387) );
  MUX2_X1 U15660 ( .A(n12436), .B(P2_EBX_REG_0__SCAN_IN), .S(n16554), .Z(
        n15776) );
  NAND2_X1 U15661 ( .A1(n15776), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16262) );
  NAND3_X1 U15662 ( .A1(n16554), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12437) );
  AND2_X1 U15663 ( .A1(n12438), .A2(n12437), .ZN(n16260) );
  NAND2_X1 U15664 ( .A1(n16260), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12440) );
  INV_X1 U15665 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16514) );
  INV_X1 U15666 ( .A(n16260), .ZN(n12439) );
  AOI22_X1 U15667 ( .A1(n16262), .A2(n12440), .B1(n16514), .B2(n12439), .ZN(
        n14386) );
  NAND2_X1 U15668 ( .A1(n14387), .A2(n14386), .ZN(n19671) );
  OAI21_X1 U15669 ( .B1(n15754), .B2(n12622), .A(n19671), .ZN(n16245) );
  INV_X1 U15670 ( .A(n12442), .ZN(n12443) );
  NAND2_X1 U15671 ( .A1(n12444), .A2(n12443), .ZN(n12445) );
  NAND2_X1 U15672 ( .A1(n12441), .A2(n12445), .ZN(n19550) );
  XNOR2_X1 U15673 ( .A(n19550), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16229) );
  INV_X1 U15674 ( .A(n19550), .ZN(n12446) );
  XNOR2_X1 U15675 ( .A(n12441), .B(n12447), .ZN(n12448) );
  NAND2_X1 U15676 ( .A1(n12448), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12450) );
  INV_X1 U15677 ( .A(n12448), .ZN(n15725) );
  NAND2_X1 U15678 ( .A1(n15725), .A2(n13456), .ZN(n12449) );
  AND2_X1 U15679 ( .A1(n12450), .A2(n12449), .ZN(n13464) );
  NAND2_X1 U15680 ( .A1(n13463), .A2(n13464), .ZN(n12469) );
  INV_X1 U15681 ( .A(n12451), .ZN(n12627) );
  AOI22_X1 U15682 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n12452), .B1(
        n20104), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15683 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12454), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15684 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12459), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15685 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19977), .B1(
        n19934), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15686 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19718), .B1(
        n19843), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U15687 ( .A1(n12466), .A2(n12004), .ZN(n12467) );
  AOI22_X1 U15688 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12452), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15689 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20104), .B1(
        n12453), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15690 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16529), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15691 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19934), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15692 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19977), .B1(
        n12454), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15693 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19843), .B1(
        n19685), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15694 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19718), .B1(
        n20037), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12474) );
  XNOR2_X1 U15695 ( .A(n12480), .B(n12479), .ZN(n19531) );
  INV_X1 U15696 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16469) );
  INV_X1 U15697 ( .A(n12482), .ZN(n12484) );
  XNOR2_X1 U15698 ( .A(n12484), .B(n12483), .ZN(n15714) );
  NAND2_X1 U15699 ( .A1(n15714), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16202) );
  NAND2_X1 U15700 ( .A1(n12485), .A2(n12486), .ZN(n12497) );
  INV_X1 U15701 ( .A(n12485), .ZN(n12488) );
  INV_X1 U15702 ( .A(n12486), .ZN(n12487) );
  NAND2_X1 U15703 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  NAND2_X1 U15704 ( .A1(n12497), .A2(n12489), .ZN(n15701) );
  NOR2_X1 U15705 ( .A1(n15701), .A2(n12354), .ZN(n12494) );
  NAND2_X1 U15706 ( .A1(n12494), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16189) );
  NAND2_X1 U15707 ( .A1(n16554), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12491) );
  MUX2_X1 U15708 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n12491), .S(n12533), .Z(
        n12493) );
  NAND2_X1 U15709 ( .A1(n12493), .A2(n12492), .ZN(n15672) );
  INV_X1 U15710 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16431) );
  OAI21_X1 U15711 ( .B1(n15672), .B2(n12354), .A(n16431), .ZN(n16164) );
  INV_X1 U15712 ( .A(n12494), .ZN(n12495) );
  NAND2_X1 U15713 ( .A1(n12495), .A2(n16457), .ZN(n16188) );
  INV_X1 U15714 ( .A(n15714), .ZN(n12496) );
  NAND2_X1 U15715 ( .A1(n12496), .A2(n16451), .ZN(n16205) );
  AND2_X1 U15716 ( .A1(n16188), .A2(n16205), .ZN(n16161) );
  NAND2_X1 U15717 ( .A1(n16554), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12498) );
  MUX2_X1 U15718 ( .A(n16554), .B(n12498), .S(n12497), .Z(n12499) );
  NAND2_X1 U15719 ( .A1(n12499), .A2(n12533), .ZN(n15689) );
  OR2_X1 U15720 ( .A1(n15689), .A2(n12354), .ZN(n12500) );
  INV_X1 U15721 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16444) );
  NAND2_X1 U15722 ( .A1(n12500), .A2(n16444), .ZN(n16176) );
  NAND3_X1 U15723 ( .A1(n16164), .A2(n16161), .A3(n16176), .ZN(n12501) );
  INV_X1 U15724 ( .A(n12501), .ZN(n12502) );
  NAND2_X1 U15725 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12504) );
  NOR2_X1 U15726 ( .A1(n15672), .A2(n12504), .ZN(n16163) );
  INV_X1 U15727 ( .A(n15689), .ZN(n12506) );
  AND2_X1 U15728 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12505) );
  OR2_X1 U15729 ( .A1(n12551), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12552) );
  NAND3_X1 U15730 ( .A1(n12552), .A2(n16554), .A3(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n12508) );
  NAND2_X1 U15731 ( .A1(n9704), .A2(n12508), .ZN(n15563) );
  NOR2_X1 U15732 ( .A1(n15563), .A2(n12354), .ZN(n12557) );
  INV_X1 U15733 ( .A(n12557), .ZN(n12509) );
  NAND2_X1 U15734 ( .A1(n12509), .A2(n10099), .ZN(n12732) );
  INV_X1 U15735 ( .A(n12510), .ZN(n12512) );
  XNOR2_X1 U15736 ( .A(n12512), .B(n12511), .ZN(n15582) );
  INV_X1 U15737 ( .A(n12558), .ZN(n12513) );
  NAND2_X1 U15738 ( .A1(n12513), .A2(n16306), .ZN(n12864) );
  INV_X1 U15739 ( .A(n12514), .ZN(n12515) );
  XNOR2_X1 U15740 ( .A(n12526), .B(n12515), .ZN(n15603) );
  NAND2_X1 U15741 ( .A1(n15603), .A2(n12644), .ZN(n12516) );
  NAND2_X1 U15742 ( .A1(n12516), .A2(n16068), .ZN(n16071) );
  NAND3_X1 U15743 ( .A1(n12517), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n16554), 
        .ZN(n12518) );
  OAI211_X1 U15744 ( .C1(n12517), .C2(P2_EBX_REG_16__SCAN_IN), .A(n12518), .B(
        n12492), .ZN(n15624) );
  OR2_X1 U15745 ( .A1(n15624), .A2(n12354), .ZN(n12519) );
  XNOR2_X1 U15746 ( .A(n12519), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16090) );
  NAND2_X1 U15747 ( .A1(n16554), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12521) );
  MUX2_X1 U15748 ( .A(n16554), .B(n12521), .S(n12546), .Z(n12522) );
  NAND2_X1 U15749 ( .A1(n12520), .A2(n15664), .ZN(n12530) );
  AOI21_X1 U15750 ( .B1(n15660), .B2(n12644), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16102) );
  INV_X1 U15751 ( .A(n16102), .ZN(n16117) );
  NAND2_X1 U15752 ( .A1(n12524), .A2(n12523), .ZN(n12525) );
  NAND2_X1 U15753 ( .A1(n12526), .A2(n12525), .ZN(n15611) );
  NOR2_X1 U15754 ( .A1(n15611), .A2(n12354), .ZN(n12560) );
  INV_X1 U15755 ( .A(n12560), .ZN(n12527) );
  INV_X1 U15756 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U15757 ( .A1(n12527), .A2(n16081), .ZN(n12729) );
  NOR2_X1 U15758 ( .A1(n12342), .A2(n12528), .ZN(n12529) );
  NAND2_X1 U15759 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  NAND2_X1 U15760 ( .A1(n12531), .A2(n12517), .ZN(n15651) );
  OR2_X1 U15761 ( .A1(n15651), .A2(n12354), .ZN(n12532) );
  INV_X1 U15762 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16364) );
  NAND2_X1 U15763 ( .A1(n12532), .A2(n16364), .ZN(n16104) );
  INV_X1 U15764 ( .A(n12533), .ZN(n12535) );
  NAND2_X1 U15765 ( .A1(n12535), .A2(n12534), .ZN(n12536) );
  AND3_X1 U15766 ( .A1(n12536), .A2(n16554), .A3(P2_EBX_REG_11__SCAN_IN), .ZN(
        n12537) );
  OR2_X1 U15767 ( .A1(n12538), .A2(n12537), .ZN(n13492) );
  NOR2_X1 U15768 ( .A1(n13492), .A2(n12354), .ZN(n12556) );
  INV_X1 U15769 ( .A(n12556), .ZN(n12539) );
  INV_X1 U15770 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16410) );
  NAND2_X1 U15771 ( .A1(n12539), .A2(n16410), .ZN(n16149) );
  NAND2_X1 U15772 ( .A1(n12542), .A2(n10171), .ZN(n12543) );
  NAND2_X1 U15773 ( .A1(n12540), .A2(n12543), .ZN(n19514) );
  INV_X1 U15774 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16384) );
  NAND2_X1 U15775 ( .A1(n12555), .A2(n16384), .ZN(n12725) );
  NAND2_X1 U15776 ( .A1(n12540), .A2(n12544), .ZN(n12545) );
  NAND2_X1 U15777 ( .A1(n12546), .A2(n12545), .ZN(n13476) );
  NOR2_X1 U15778 ( .A1(n13476), .A2(n12354), .ZN(n12562) );
  INV_X1 U15779 ( .A(n12562), .ZN(n12547) );
  INV_X1 U15780 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16383) );
  NAND2_X1 U15781 ( .A1(n12547), .A2(n16383), .ZN(n16101) );
  AND4_X1 U15782 ( .A1(n16104), .A2(n16149), .A3(n12725), .A4(n16101), .ZN(
        n12548) );
  AND4_X1 U15783 ( .A1(n16090), .A2(n16117), .A3(n12729), .A4(n12548), .ZN(
        n12549) );
  AND2_X1 U15784 ( .A1(n14283), .A2(n12549), .ZN(n12554) );
  NAND2_X1 U15785 ( .A1(n12551), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12550) );
  MUX2_X1 U15786 ( .A(n12551), .B(n12550), .S(n16554), .Z(n12553) );
  INV_X1 U15787 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14290) );
  AND3_X1 U15788 ( .A1(n12732), .A2(n12554), .A3(n14285), .ZN(n12570) );
  XNOR2_X1 U15789 ( .A(n12555), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16139) );
  AND2_X1 U15790 ( .A1(n12556), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12724) );
  INV_X1 U15791 ( .A(n12724), .ZN(n16150) );
  NAND2_X1 U15792 ( .A1(n16139), .A2(n16150), .ZN(n12569) );
  NAND2_X1 U15793 ( .A1(n12557), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12733) );
  NAND2_X1 U15794 ( .A1(n12558), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12865) );
  AND2_X1 U15795 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12559) );
  NAND2_X1 U15796 ( .A1(n15603), .A2(n12559), .ZN(n16070) );
  NAND2_X1 U15797 ( .A1(n12865), .A2(n16070), .ZN(n12731) );
  NAND2_X1 U15798 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12730) );
  AND2_X1 U15799 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12561) );
  NAND2_X1 U15800 ( .A1(n15660), .A2(n12561), .ZN(n16116) );
  NAND2_X1 U15801 ( .A1(n12562), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16128) );
  OR3_X1 U15802 ( .A1(n15651), .A2(n12354), .A3(n16364), .ZN(n16103) );
  AND3_X1 U15803 ( .A1(n16116), .A2(n16128), .A3(n16103), .ZN(n12727) );
  NAND2_X1 U15804 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12563) );
  NOR2_X1 U15805 ( .A1(n15624), .A2(n12563), .ZN(n12728) );
  INV_X1 U15806 ( .A(n12728), .ZN(n12564) );
  NAND3_X1 U15807 ( .A1(n12730), .A2(n12727), .A3(n12564), .ZN(n12565) );
  NOR2_X1 U15808 ( .A1(n12731), .A2(n12565), .ZN(n12567) );
  NAND2_X1 U15809 ( .A1(n12566), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14286) );
  NAND3_X1 U15810 ( .A1(n12733), .A2(n12567), .A3(n14286), .ZN(n12568) );
  AOI21_X1 U15811 ( .B1(n12570), .B2(n12569), .A(n12568), .ZN(n16056) );
  INV_X1 U15812 ( .A(n12571), .ZN(n12580) );
  INV_X1 U15813 ( .A(n12572), .ZN(n12574) );
  NAND2_X1 U15814 ( .A1(n12574), .A2(n12573), .ZN(n12575) );
  NAND2_X1 U15815 ( .A1(n12580), .A2(n12575), .ZN(n15546) );
  INV_X1 U15816 ( .A(n12578), .ZN(n12576) );
  NAND2_X1 U15817 ( .A1(n12576), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16055) );
  AND2_X1 U15818 ( .A1(n16056), .A2(n16055), .ZN(n12577) );
  INV_X1 U15819 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16324) );
  NAND2_X1 U15820 ( .A1(n12578), .A2(n16324), .ZN(n16054) );
  XNOR2_X1 U15821 ( .A(n12580), .B(n12579), .ZN(n15536) );
  NAND2_X1 U15822 ( .A1(n15536), .A2(n12644), .ZN(n12584) );
  XNOR2_X1 U15823 ( .A(n12584), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16050) );
  AND2_X1 U15824 ( .A1(n16054), .A2(n16050), .ZN(n12581) );
  NAND2_X1 U15825 ( .A1(n12582), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16039) );
  INV_X1 U15826 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12583) );
  OR2_X1 U15827 ( .A1(n12584), .A2(n12583), .ZN(n14360) );
  AND2_X1 U15828 ( .A1(n16039), .A2(n14360), .ZN(n12585) );
  INV_X1 U15829 ( .A(n16021), .ZN(n12591) );
  INV_X1 U15830 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21443) );
  INV_X1 U15831 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16019) );
  NAND2_X1 U15832 ( .A1(n21443), .A2(n16019), .ZN(n12590) );
  INV_X1 U15833 ( .A(n12586), .ZN(n12587) );
  NAND2_X1 U15834 ( .A1(n12587), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12589) );
  AND2_X1 U15835 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12588) );
  NAND2_X1 U15836 ( .A1(n15503), .A2(n12588), .ZN(n16027) );
  NAND2_X1 U15837 ( .A1(n12589), .A2(n16027), .ZN(n16017) );
  AOI21_X1 U15838 ( .B1(n12591), .B2(n12590), .A(n16017), .ZN(n12592) );
  XNOR2_X1 U15839 ( .A(n12594), .B(n12593), .ZN(n15442) );
  NAND2_X1 U15840 ( .A1(n15442), .A2(n12644), .ZN(n12596) );
  NAND2_X1 U15841 ( .A1(n12596), .A2(n12595), .ZN(n12656) );
  INV_X1 U15842 ( .A(n12687), .ZN(n12607) );
  AND2_X1 U15843 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12597) );
  NAND2_X1 U15844 ( .A1(n12834), .A2(n12597), .ZN(n12684) );
  AND2_X1 U15845 ( .A1(n12644), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12598) );
  NAND2_X1 U15846 ( .A1(n15442), .A2(n12598), .ZN(n12686) );
  NOR2_X1 U15847 ( .A1(n9691), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12603) );
  INV_X1 U15848 ( .A(n12600), .ZN(n12685) );
  NOR2_X1 U15849 ( .A1(n12685), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12602) );
  INV_X1 U15850 ( .A(n12604), .ZN(n12605) );
  OAI21_X1 U15851 ( .B1(n12607), .B2(n12606), .A(n12605), .ZN(n12608) );
  NOR2_X1 U15852 ( .A1(n12003), .A2(n12609), .ZN(n20339) );
  NAND2_X1 U15853 ( .A1(n12640), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12612) );
  NAND2_X1 U15854 ( .A1(n12632), .A2(n13456), .ZN(n12611) );
  MUX2_X1 U15855 ( .A(n12612), .B(n12611), .S(n12634), .Z(n12636) );
  INV_X1 U15856 ( .A(n12616), .ZN(n12614) );
  INV_X1 U15857 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12613) );
  NOR3_X1 U15858 ( .A1(n12614), .A2(n13732), .A3(n12613), .ZN(n12618) );
  NOR2_X1 U15859 ( .A1(n13732), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12615) );
  XNOR2_X1 U15860 ( .A(n12616), .B(n12615), .ZN(n16259) );
  AND2_X1 U15861 ( .A1(n16259), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12617) );
  NOR2_X1 U15862 ( .A1(n12618), .A2(n12617), .ZN(n12623) );
  XNOR2_X1 U15863 ( .A(n12622), .B(n12623), .ZN(n14390) );
  INV_X1 U15864 ( .A(n14390), .ZN(n12621) );
  XNOR2_X1 U15865 ( .A(n12620), .B(n12619), .ZN(n14388) );
  NAND2_X1 U15866 ( .A1(n12621), .A2(n14388), .ZN(n14392) );
  OR2_X1 U15867 ( .A1(n12623), .A2(n12622), .ZN(n12624) );
  NAND2_X1 U15868 ( .A1(n14392), .A2(n12624), .ZN(n12625) );
  XNOR2_X1 U15869 ( .A(n12625), .B(n16476), .ZN(n16250) );
  NAND2_X1 U15870 ( .A1(n12625), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12626) );
  NAND2_X1 U15871 ( .A1(n12628), .A2(n12627), .ZN(n12629) );
  INV_X1 U15872 ( .A(n12638), .ZN(n12633) );
  NAND2_X1 U15873 ( .A1(n12634), .A2(n13456), .ZN(n13460) );
  INV_X1 U15874 ( .A(n12634), .ZN(n12635) );
  NAND2_X1 U15875 ( .A1(n13459), .A2(n13460), .ZN(n13458) );
  NAND2_X1 U15876 ( .A1(n13458), .A2(n12637), .ZN(n12639) );
  NAND3_X1 U15877 ( .A1(n12645), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n12644), .ZN(n12646) );
  INV_X1 U15878 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14374) );
  NOR2_X1 U15879 ( .A1(n14374), .A2(n12696), .ZN(n12648) );
  INV_X1 U15880 ( .A(n12650), .ZN(n20341) );
  NAND2_X1 U15881 ( .A1(n9695), .A2(n19657), .ZN(n12652) );
  NAND3_X1 U15882 ( .A1(n12654), .A2(n12653), .A3(n12652), .ZN(P2_U3015) );
  NOR2_X4 U15883 ( .A1(n14369), .A2(n16019), .ZN(n16015) );
  AOI21_X1 U15884 ( .B1(n16015), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12655) );
  NOR2_X1 U15885 ( .A1(n12655), .A2(n12674), .ZN(n12889) );
  NAND2_X1 U15886 ( .A1(n12889), .A2(n19657), .ZN(n12671) );
  NAND2_X1 U15887 ( .A1(n12656), .A2(n12686), .ZN(n12657) );
  XNOR2_X1 U15888 ( .A(n12658), .B(n12657), .ZN(n12893) );
  NAND2_X1 U15889 ( .A1(n12893), .A2(n19672), .ZN(n12670) );
  NOR2_X1 U15890 ( .A1(n16032), .A2(n20279), .ZN(n12891) );
  AOI21_X1 U15891 ( .B1(n16270), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12891), .ZN(n12664) );
  OAI211_X1 U15892 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n12662), .A(
        n16272), .B(n12696), .ZN(n12663) );
  OAI211_X1 U15893 ( .C1(n15903), .C2(n19648), .A(n12664), .B(n12663), .ZN(
        n12668) );
  NOR2_X1 U15894 ( .A1(n15456), .A2(n12665), .ZN(n12666) );
  NOR2_X1 U15895 ( .A1(n15791), .A2(n17133), .ZN(n12667) );
  NAND3_X1 U15896 ( .A1(n12671), .A2(n12670), .A3(n12669), .ZN(P2_U3017) );
  AND2_X1 U15897 ( .A1(n11752), .A2(n16626), .ZN(n12672) );
  NOR2_X1 U15898 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20305) );
  INV_X1 U15899 ( .A(n20305), .ZN(n20297) );
  NAND2_X1 U15900 ( .A1(n20313), .A2(n20297), .ZN(n20306) );
  NAND2_X1 U15901 ( .A1(n20306), .A2(n17153), .ZN(n12679) );
  AND2_X1 U15902 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12680) );
  NAND2_X1 U15903 ( .A1(n12770), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12772) );
  INV_X1 U15904 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12783) );
  INV_X1 U15905 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16075) );
  INV_X1 U15906 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12868) );
  INV_X1 U15907 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12801) );
  INV_X1 U15908 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12804) );
  INV_X1 U15909 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12808) );
  INV_X1 U15910 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12816) );
  INV_X1 U15911 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12714) );
  XNOR2_X1 U15912 ( .A(n12754), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12826) );
  NAND2_X1 U15913 ( .A1(n17153), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15428) );
  INV_X1 U15914 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n16495) );
  NAND2_X1 U15915 ( .A1(n16495), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U15916 ( .A1(n15428), .A2(n12825), .ZN(n19633) );
  NAND2_X1 U15917 ( .A1(n19553), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12698) );
  OAI21_X1 U15918 ( .B1(n16237), .B2(n10186), .A(n12698), .ZN(n12681) );
  AOI21_X1 U15919 ( .B1(n12826), .B2(n16234), .A(n12681), .ZN(n12682) );
  OAI21_X1 U15920 ( .B1(n14382), .B2(n16222), .A(n12682), .ZN(n12683) );
  AOI21_X1 U15921 ( .B1(n19636), .B2(n12701), .A(n12683), .ZN(n12692) );
  NAND2_X1 U15922 ( .A1(n12685), .A2(n12684), .ZN(n12688) );
  INV_X1 U15923 ( .A(n12702), .ZN(n12690) );
  NAND2_X1 U15924 ( .A1(n12690), .A2(n16263), .ZN(n12691) );
  NAND2_X1 U15925 ( .A1(n12692), .A2(n12691), .ZN(P2_U2984) );
  AOI21_X1 U15926 ( .B1(n12695), .B2(n12694), .A(n12693), .ZN(n13248) );
  INV_X1 U15927 ( .A(n12696), .ZN(n12697) );
  AOI21_X1 U15928 ( .B1(n16272), .B2(n12697), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15929 ( .A1(n12703), .A2(n10297), .ZN(P2_U3016) );
  INV_X1 U15930 ( .A(n12706), .ZN(n12707) );
  NAND2_X1 U15931 ( .A1(n12708), .A2(n12707), .ZN(n12709) );
  NAND2_X1 U15932 ( .A1(n12373), .A2(n12709), .ZN(n15470) );
  NOR2_X1 U15933 ( .A1(n15470), .A2(n12354), .ZN(n16016) );
  NAND3_X1 U15934 ( .A1(n14414), .A2(n14415), .A3(n16263), .ZN(n12723) );
  NAND2_X1 U15935 ( .A1(n14369), .A2(n16019), .ZN(n14413) );
  NAND2_X1 U15936 ( .A1(n14413), .A2(n19636), .ZN(n12720) );
  INV_X1 U15937 ( .A(n9662), .ZN(n12712) );
  AOI21_X1 U15938 ( .B1(n12713), .B2(n9632), .A(n12712), .ZN(n15801) );
  AND2_X1 U15939 ( .A1(n9663), .A2(n12714), .ZN(n12716) );
  OR2_X1 U15940 ( .A1(n12716), .A2(n12715), .ZN(n15471) );
  INV_X1 U15941 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20276) );
  NOR2_X1 U15942 ( .A1(n16032), .A2(n20276), .ZN(n14418) );
  AOI21_X1 U15943 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14418), .ZN(n12717) );
  OAI21_X1 U15944 ( .B1(n15471), .B2(n16264), .A(n12717), .ZN(n12718) );
  AOI21_X1 U15945 ( .B1(n15801), .B2(n19642), .A(n12718), .ZN(n12719) );
  NAND2_X1 U15946 ( .A1(n16117), .A2(n10296), .ZN(n12726) );
  AOI21_X2 U15947 ( .B1(n16100), .B2(n12727), .A(n12726), .ZN(n16089) );
  NAND2_X1 U15948 ( .A1(n12730), .A2(n12729), .ZN(n14251) );
  NAND2_X1 U15949 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  XNOR2_X1 U15950 ( .A(n12735), .B(n12734), .ZN(n13250) );
  NAND2_X1 U15951 ( .A1(n13250), .A2(n16263), .ZN(n12753) );
  OR2_X1 U15952 ( .A1(n16410), .A2(n16431), .ZN(n16141) );
  OR2_X1 U15953 ( .A1(n16141), .A2(n16384), .ZN(n12736) );
  NOR2_X1 U15954 ( .A1(n16444), .A2(n12736), .ZN(n12737) );
  INV_X1 U15955 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12738) );
  NOR2_X1 U15956 ( .A1(n16383), .A2(n12738), .ZN(n14256) );
  INV_X1 U15957 ( .A(n14258), .ZN(n12739) );
  AND2_X1 U15958 ( .A1(n14256), .A2(n12739), .ZN(n12740) );
  NAND2_X1 U15959 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12741) );
  INV_X1 U15960 ( .A(n13251), .ZN(n12743) );
  INV_X1 U15961 ( .A(n12744), .ZN(n14293) );
  INV_X1 U15962 ( .A(n12798), .ZN(n12747) );
  INV_X1 U15963 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21452) );
  NAND2_X1 U15964 ( .A1(n12747), .A2(n21452), .ZN(n12748) );
  NAND2_X1 U15965 ( .A1(n12802), .A2(n12748), .ZN(n15559) );
  NOR2_X1 U15966 ( .A1(n15559), .A2(n16264), .ZN(n12750) );
  NAND2_X1 U15967 ( .A1(n19553), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n13256) );
  OAI21_X1 U15968 ( .B1(n16237), .B2(n21452), .A(n13256), .ZN(n12749) );
  AOI211_X1 U15969 ( .C1(n15845), .C2(n19642), .A(n12750), .B(n12749), .ZN(
        n12751) );
  NAND3_X1 U15970 ( .A1(n12753), .A2(n12752), .A3(n12751), .ZN(P2_U2993) );
  MUX2_X1 U15971 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16504) );
  MUX2_X1 U15972 ( .A(n15761), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15765) );
  INV_X1 U15973 ( .A(n12760), .ZN(n12758) );
  INV_X1 U15974 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U15975 ( .A1(n15761), .A2(n12756), .ZN(n12757) );
  NAND2_X1 U15976 ( .A1(n12758), .A2(n12757), .ZN(n15748) );
  AND2_X1 U15977 ( .A1(n15767), .A2(n15748), .ZN(n15731) );
  OAI21_X1 U15978 ( .B1(n12760), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n12759), .ZN(n16248) );
  NAND2_X1 U15979 ( .A1(n15731), .A2(n16248), .ZN(n19558) );
  AND2_X1 U15980 ( .A1(n12759), .A2(n16236), .ZN(n12762) );
  NOR2_X1 U15981 ( .A1(n12761), .A2(n12762), .ZN(n19561) );
  OR2_X1 U15982 ( .A1(n19558), .A2(n19561), .ZN(n19562) );
  OR2_X1 U15983 ( .A1(n12761), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12764) );
  AND2_X1 U15984 ( .A1(n12763), .A2(n12764), .ZN(n16219) );
  NAND2_X1 U15985 ( .A1(n12763), .A2(n12766), .ZN(n12767) );
  NAND2_X1 U15986 ( .A1(n12765), .A2(n12767), .ZN(n19536) );
  NAND2_X1 U15987 ( .A1(n19534), .A2(n19536), .ZN(n15711) );
  AND2_X1 U15988 ( .A1(n12765), .A2(n16201), .ZN(n12769) );
  NOR2_X1 U15989 ( .A1(n12768), .A2(n12769), .ZN(n16199) );
  OR2_X1 U15990 ( .A1(n15711), .A2(n16199), .ZN(n15694) );
  NOR2_X1 U15991 ( .A1(n12768), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12771) );
  OR2_X1 U15992 ( .A1(n12770), .A2(n12771), .ZN(n16193) );
  INV_X1 U15993 ( .A(n16193), .ZN(n15695) );
  NOR2_X1 U15994 ( .A1(n15694), .A2(n15695), .ZN(n15682) );
  OR2_X1 U15995 ( .A1(n12770), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12773) );
  NAND2_X1 U15996 ( .A1(n12772), .A2(n12773), .ZN(n16182) );
  AND2_X1 U15997 ( .A1(n15682), .A2(n16182), .ZN(n15669) );
  OR2_X1 U15998 ( .A1(n12772), .A2(n15675), .ZN(n12775) );
  NAND2_X1 U15999 ( .A1(n12772), .A2(n15675), .ZN(n12774) );
  NAND2_X1 U16000 ( .A1(n12775), .A2(n12774), .ZN(n16169) );
  NAND2_X1 U16001 ( .A1(n15669), .A2(n16169), .ZN(n13487) );
  NAND2_X1 U16002 ( .A1(n12775), .A2(n16152), .ZN(n12776) );
  AND2_X1 U16003 ( .A1(n12777), .A2(n12776), .ZN(n16154) );
  AND2_X1 U16004 ( .A1(n12777), .A2(n16142), .ZN(n12778) );
  NOR2_X1 U16005 ( .A1(n12780), .A2(n12778), .ZN(n19518) );
  OR2_X1 U16006 ( .A1(n12780), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12781) );
  NAND2_X1 U16007 ( .A1(n12779), .A2(n12781), .ZN(n16134) );
  INV_X1 U16008 ( .A(n12782), .ZN(n12785) );
  NAND2_X1 U16009 ( .A1(n12779), .A2(n12783), .ZN(n12784) );
  NAND2_X1 U16010 ( .A1(n12785), .A2(n12784), .ZN(n16120) );
  NAND2_X1 U16011 ( .A1(n15657), .A2(n16120), .ZN(n15643) );
  AND2_X1 U16012 ( .A1(n12785), .A2(n16107), .ZN(n12786) );
  NOR2_X1 U16013 ( .A1(n12788), .A2(n12786), .ZN(n16109) );
  OR2_X1 U16014 ( .A1(n15643), .A2(n16109), .ZN(n15628) );
  NOR2_X1 U16015 ( .A1(n12788), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12789) );
  OR2_X1 U16016 ( .A1(n12787), .A2(n12789), .ZN(n16093) );
  INV_X1 U16017 ( .A(n16093), .ZN(n12790) );
  OR2_X1 U16018 ( .A1(n12787), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12792) );
  NAND2_X1 U16019 ( .A1(n12791), .A2(n12792), .ZN(n16084) );
  NAND2_X1 U16020 ( .A1(n15609), .A2(n16084), .ZN(n15598) );
  NAND2_X1 U16021 ( .A1(n12791), .A2(n16075), .ZN(n12793) );
  AND2_X1 U16022 ( .A1(n12794), .A2(n12793), .ZN(n16077) );
  OR2_X1 U16023 ( .A1(n15598), .A2(n16077), .ZN(n15578) );
  AND2_X1 U16024 ( .A1(n12794), .A2(n12868), .ZN(n12795) );
  NOR2_X1 U16025 ( .A1(n12796), .A2(n12795), .ZN(n15579) );
  NOR2_X1 U16026 ( .A1(n12796), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12797) );
  OR2_X1 U16027 ( .A1(n12798), .A2(n12797), .ZN(n15571) );
  NAND2_X1 U16028 ( .A1(n15567), .A2(n15571), .ZN(n12799) );
  NAND2_X1 U16029 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U16030 ( .A1(n12805), .A2(n12803), .ZN(n16064) );
  NAND2_X1 U16031 ( .A1(n15530), .A2(n19559), .ZN(n12807) );
  NAND2_X1 U16032 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  NAND2_X1 U16033 ( .A1(n12809), .A2(n12806), .ZN(n16047) );
  NAND2_X1 U16034 ( .A1(n15514), .A2(n19559), .ZN(n12811) );
  AND2_X1 U16035 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  OR2_X1 U16036 ( .A1(n12810), .A2(n12813), .ZN(n16043) );
  NAND2_X1 U16037 ( .A1(n15498), .A2(n19559), .ZN(n12815) );
  OR2_X1 U16038 ( .A1(n12813), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12814) );
  NAND2_X1 U16039 ( .A1(n12812), .A2(n12814), .ZN(n16035) );
  NAND2_X1 U16040 ( .A1(n15478), .A2(n19559), .ZN(n12818) );
  NAND2_X1 U16041 ( .A1(n12812), .A2(n12816), .ZN(n12817) );
  NAND2_X1 U16042 ( .A1(n9663), .A2(n12817), .ZN(n15479) );
  NOR2_X1 U16043 ( .A1(n12715), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12820) );
  OR2_X1 U16044 ( .A1(n12819), .A2(n12820), .ZN(n16025) );
  NAND2_X1 U16045 ( .A1(n15439), .A2(n19559), .ZN(n12823) );
  OR2_X1 U16046 ( .A1(n12819), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12822) );
  NAND2_X1 U16047 ( .A1(n12754), .A2(n12822), .ZN(n15440) );
  NAND2_X1 U16048 ( .A1(n17153), .A2(n20145), .ZN(n12824) );
  OR2_X1 U16049 ( .A1(n12825), .A2(n12824), .ZN(n19537) );
  AOI21_X1 U16050 ( .B1(n12827), .B2(n19559), .A(n12826), .ZN(n12853) );
  INV_X1 U16051 ( .A(n12291), .ZN(n16597) );
  NAND2_X1 U16052 ( .A1(n16597), .A2(n12832), .ZN(n15434) );
  NAND2_X1 U16053 ( .A1(n17147), .A2(n16495), .ZN(n12835) );
  INV_X1 U16054 ( .A(n12835), .ZN(n12829) );
  NAND2_X1 U16055 ( .A1(n12836), .A2(n12829), .ZN(n12830) );
  NOR2_X1 U16056 ( .A1(n13632), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12843) );
  NAND2_X1 U16057 ( .A1(n19630), .A2(n12843), .ZN(n19551) );
  INV_X1 U16058 ( .A(n12834), .ZN(n12847) );
  NAND3_X1 U16059 ( .A1(n12836), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12835), 
        .ZN(n12837) );
  NAND2_X1 U16060 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20145), .ZN(n19684) );
  NOR2_X1 U16061 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19684), .ZN(n12838) );
  NAND2_X1 U16062 ( .A1(n12838), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17148) );
  AND3_X1 U16063 ( .A1(n16032), .A2(n19537), .A3(n17148), .ZN(n12839) );
  AOI22_X1 U16064 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19554), .ZN(n12846) );
  INV_X1 U16065 ( .A(n13563), .ZN(n13531) );
  INV_X1 U16066 ( .A(n17147), .ZN(n20224) );
  OAI21_X1 U16067 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20224), .A(n12840), 
        .ZN(n12841) );
  OR2_X1 U16068 ( .A1(n13531), .A2(n12841), .ZN(n12842) );
  NAND2_X1 U16069 ( .A1(n13679), .A2(n12842), .ZN(n12844) );
  INV_X1 U16070 ( .A(n12843), .ZN(n16622) );
  NAND2_X1 U16071 ( .A1(n19547), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12845) );
  OAI211_X1 U16072 ( .C1(n12847), .C2(n19549), .A(n12846), .B(n12845), .ZN(
        n12848) );
  NAND2_X1 U16073 ( .A1(n12852), .A2(n12851), .ZN(P2_U2825) );
  AOI22_X1 U16074 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19554), .ZN(n12857) );
  NAND2_X1 U16075 ( .A1(n19547), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12856) );
  OAI211_X1 U16076 ( .C1(n12858), .C2(n19549), .A(n12857), .B(n12856), .ZN(
        n12859) );
  INV_X1 U16077 ( .A(n12859), .ZN(n12860) );
  OAI211_X1 U16078 ( .C1(n12828), .C2(n15784), .A(n12863), .B(n12862), .ZN(
        P2_U2824) );
  AND2_X1 U16079 ( .A1(n12865), .A2(n12864), .ZN(n12866) );
  XNOR2_X1 U16080 ( .A(n12867), .B(n12866), .ZN(n12875) );
  NAND2_X1 U16081 ( .A1(n12875), .A2(n16263), .ZN(n12874) );
  NAND2_X1 U16082 ( .A1(n19553), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12882) );
  OAI21_X1 U16083 ( .B1(n16237), .B2(n12868), .A(n12882), .ZN(n12871) );
  OAI21_X1 U16084 ( .B1(n9640), .B2(n12869), .A(n14293), .ZN(n15858) );
  NOR2_X1 U16085 ( .A1(n15858), .A2(n16222), .ZN(n12870) );
  AOI211_X1 U16086 ( .C1(n16234), .C2(n15579), .A(n12871), .B(n12870), .ZN(
        n12872) );
  NAND2_X1 U16087 ( .A1(n12874), .A2(n12873), .ZN(P2_U2995) );
  NAND2_X1 U16088 ( .A1(n12875), .A2(n19672), .ZN(n12888) );
  INV_X1 U16089 ( .A(n12876), .ZN(n12879) );
  AND2_X1 U16090 ( .A1(n15591), .A2(n15590), .ZN(n15593) );
  INV_X1 U16091 ( .A(n15593), .ZN(n12878) );
  AOI21_X1 U16092 ( .B1(n12879), .B2(n12878), .A(n12877), .ZN(n15972) );
  NOR2_X1 U16093 ( .A1(n16334), .A2(n16068), .ZN(n12880) );
  NAND2_X1 U16094 ( .A1(n16411), .A2(n12880), .ZN(n16307) );
  OR2_X1 U16095 ( .A1(n16408), .A2(n12880), .ZN(n12881) );
  NAND2_X1 U16096 ( .A1(n9631), .A2(n12881), .ZN(n16337) );
  NAND2_X1 U16097 ( .A1(n16337), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12883) );
  OAI211_X1 U16098 ( .C1(n16307), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12883), .B(n12882), .ZN(n12885) );
  NOR2_X1 U16099 ( .A1(n15858), .A2(n17133), .ZN(n12884) );
  AOI211_X1 U16100 ( .C1(n19665), .C2(n15972), .A(n12885), .B(n12884), .ZN(
        n12886) );
  NAND2_X1 U16101 ( .A1(n12888), .A2(n12887), .ZN(P2_U3027) );
  NAND2_X1 U16102 ( .A1(n12889), .A2(n19636), .ZN(n12898) );
  NOR2_X1 U16103 ( .A1(n15440), .A2(n16264), .ZN(n12890) );
  AOI211_X1 U16104 ( .C1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19634), .A(
        n12891), .B(n12890), .ZN(n12892) );
  OAI21_X1 U16105 ( .B1(n15791), .B2(n16222), .A(n12892), .ZN(n12896) );
  INV_X1 U16106 ( .A(n12893), .ZN(n12894) );
  NOR2_X1 U16107 ( .A1(n12896), .A2(n12895), .ZN(n12897) );
  NAND2_X1 U16108 ( .A1(n12898), .A2(n12897), .ZN(P2_U2985) );
  INV_X1 U16109 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17285) );
  NOR2_X1 U16110 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18561), .ZN(
        n17579) );
  NAND2_X1 U16111 ( .A1(n9734), .A2(n17579), .ZN(n17430) );
  INV_X1 U16112 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18363) );
  NAND2_X1 U16113 ( .A1(n17508), .A2(n10301), .ZN(n17424) );
  INV_X1 U16114 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18400) );
  INV_X1 U16115 ( .A(n18394), .ZN(n12901) );
  INV_X1 U16116 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18494) );
  NAND2_X1 U16117 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n12900), .ZN(
        n17551) );
  NOR2_X1 U16118 ( .A1(n18494), .A2(n17551), .ZN(n17543) );
  NAND2_X1 U16119 ( .A1(n12901), .A2(n17543), .ZN(n18395) );
  NOR2_X1 U16120 ( .A1(n18400), .A2(n18395), .ZN(n17470) );
  NAND2_X1 U16121 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17470), .ZN(
        n17454) );
  NOR2_X1 U16122 ( .A1(n18379), .A2(n17454), .ZN(n17442) );
  INV_X1 U16123 ( .A(n17442), .ZN(n18354) );
  NOR2_X1 U16124 ( .A1(n18363), .A2(n18354), .ZN(n17429) );
  NAND3_X1 U16125 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17442), .ZN(n12904) );
  OAI21_X1 U16126 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17429), .A(
        n12904), .ZN(n18353) );
  NAND2_X1 U16127 ( .A1(n17424), .A2(n18353), .ZN(n17425) );
  INV_X1 U16128 ( .A(n12903), .ZN(n18314) );
  AOI21_X1 U16129 ( .B1(n18339), .B2(n12904), .A(n18314), .ZN(n18341) );
  INV_X1 U16130 ( .A(n18341), .ZN(n17411) );
  NAND2_X1 U16131 ( .A1(n17410), .A2(n17411), .ZN(n17409) );
  NAND2_X1 U16132 ( .A1(n17508), .A2(n17409), .ZN(n17402) );
  INV_X1 U16133 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21318) );
  AOI22_X1 U16134 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n12903), .B1(
        n18314), .B2(n21318), .ZN(n18325) );
  NAND2_X1 U16135 ( .A1(n17508), .A2(n17403), .ZN(n17391) );
  NOR2_X1 U16136 ( .A1(n21318), .A2(n12903), .ZN(n12906) );
  NAND3_X1 U16137 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18304) );
  NOR2_X1 U16138 ( .A1(n12904), .A2(n18304), .ZN(n18275) );
  INV_X1 U16139 ( .A(n18275), .ZN(n12905) );
  OAI21_X1 U16140 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12906), .A(
        n12905), .ZN(n18320) );
  OAI21_X1 U16141 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18275), .A(
        n12907), .ZN(n18305) );
  NAND2_X1 U16142 ( .A1(n17508), .A2(n17379), .ZN(n17369) );
  INV_X1 U16143 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18292) );
  NOR2_X1 U16144 ( .A1(n18292), .A2(n12907), .ZN(n12909) );
  AOI21_X1 U16145 ( .B1(n18292), .B2(n12907), .A(n12909), .ZN(n12908) );
  INV_X1 U16146 ( .A(n12908), .ZN(n18289) );
  NAND2_X1 U16147 ( .A1(n17508), .A2(n17370), .ZN(n17358) );
  INV_X1 U16148 ( .A(n12910), .ZN(n16753) );
  OAI21_X1 U16149 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12909), .A(
        n16753), .ZN(n18281) );
  OAI21_X1 U16150 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12910), .A(
        n12911), .ZN(n18263) );
  NAND2_X1 U16151 ( .A1(n17508), .A2(n17351), .ZN(n17340) );
  AOI21_X1 U16152 ( .B1(n18243), .B2(n12911), .A(n12914), .ZN(n12912) );
  INV_X1 U16153 ( .A(n12912), .ZN(n17342) );
  NAND2_X1 U16154 ( .A1(n17508), .A2(n17341), .ZN(n17330) );
  OAI21_X1 U16155 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12914), .A(
        n12913), .ZN(n18244) );
  OAI21_X1 U16156 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n12916), .A(
        n12915), .ZN(n17321) );
  NAND2_X1 U16157 ( .A1(n17508), .A2(n17319), .ZN(n17310) );
  OAI21_X1 U16158 ( .B1(n12918), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n12917), .ZN(n17312) );
  NAND2_X1 U16159 ( .A1(n17508), .A2(n17311), .ZN(n17298) );
  INV_X1 U16160 ( .A(n12919), .ZN(n17300) );
  INV_X1 U16161 ( .A(n12920), .ZN(n12921) );
  OAI21_X1 U16162 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16682), .A(
        n12921), .ZN(n17290) );
  NAND2_X1 U16163 ( .A1(n17508), .A2(n17289), .ZN(n17280) );
  OAI21_X1 U16164 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12920), .A(
        n12922), .ZN(n17281) );
  INV_X2 U16165 ( .A(n19355), .ZN(n17558) );
  INV_X2 U16166 ( .A(n19482), .ZN(n19434) );
  NOR2_X1 U16167 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19361) );
  NOR3_X1 U16168 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19379), .A3(n19361), 
        .ZN(n19470) );
  INV_X1 U16169 ( .A(n19470), .ZN(n19366) );
  NAND2_X1 U16170 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19466) );
  INV_X1 U16171 ( .A(n19466), .ZN(n19473) );
  AOI211_X1 U16172 ( .C1(n13916), .C2(n19366), .A(n19473), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19338) );
  INV_X1 U16173 ( .A(n12925), .ZN(n12926) );
  INV_X1 U16174 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19423) );
  INV_X1 U16175 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19419) );
  INV_X1 U16176 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19408) );
  INV_X1 U16177 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19402) );
  INV_X1 U16178 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19400) );
  INV_X1 U16179 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19396) );
  INV_X1 U16180 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19382) );
  NAND3_X1 U16181 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16639) );
  NOR2_X1 U16182 ( .A1(n19382), .A2(n16639), .ZN(n17568) );
  NAND2_X1 U16183 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17568), .ZN(n17492) );
  INV_X1 U16184 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19391) );
  NAND2_X1 U16185 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17516) );
  NOR2_X1 U16186 ( .A1(n19391), .A2(n17516), .ZN(n17496) );
  NAND3_X1 U16187 ( .A1(n17496), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n17477) );
  NOR3_X1 U16188 ( .A1(n19396), .A2(n17492), .A3(n17477), .ZN(n17469) );
  NAND2_X1 U16189 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17469), .ZN(n17440) );
  NOR3_X1 U16190 ( .A1(n19402), .A2(n19400), .A3(n17440), .ZN(n17428) );
  NAND3_X1 U16191 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n17428), .ZN(n17408) );
  NOR2_X1 U16192 ( .A1(n19408), .A2(n17408), .ZN(n17406) );
  NAND4_X1 U16193 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n17406), .ZN(n17360) );
  NAND2_X1 U16194 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n17361) );
  OR3_X1 U16195 ( .A1(n19419), .A2(n17360), .A3(n17361), .ZN(n17337) );
  NOR2_X1 U16196 ( .A1(n19423), .A2(n17337), .ZN(n12932) );
  NAND3_X1 U16197 ( .A1(n17328), .A2(P3_REIP_REG_25__SCAN_IN), .A3(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17301) );
  NAND2_X1 U16198 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n12934) );
  NOR2_X1 U16199 ( .A1(n17301), .A2(n12934), .ZN(n17288) );
  NAND2_X1 U16200 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17288), .ZN(n17273) );
  NOR2_X1 U16201 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17273), .ZN(n17279) );
  INV_X1 U16202 ( .A(n12928), .ZN(n12936) );
  NAND2_X1 U16203 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19471), .ZN(n12929) );
  AOI211_X4 U16204 ( .C1(n17254), .C2(n19466), .A(n12936), .B(n12929), .ZN(
        n17584) );
  NOR3_X2 U16205 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17582) );
  NAND2_X1 U16206 ( .A1(n17582), .A2(n16657), .ZN(n16656) );
  NAND2_X1 U16207 ( .A1(n17562), .A2(n17564), .ZN(n17561) );
  NOR2_X2 U16208 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17561), .ZN(n17542) );
  NAND2_X1 U16209 ( .A1(n17542), .A2(n17962), .ZN(n17538) );
  NOR2_X2 U16210 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17538), .ZN(n17522) );
  INV_X1 U16211 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17928) );
  NAND2_X1 U16212 ( .A1(n17522), .A2(n17928), .ZN(n17509) );
  NOR2_X2 U16213 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17509), .ZN(n17490) );
  INV_X1 U16214 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17489) );
  NAND2_X1 U16215 ( .A1(n17490), .A2(n17489), .ZN(n17481) );
  NOR2_X2 U16216 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17481), .ZN(n17466) );
  INV_X1 U16217 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17457) );
  NAND2_X1 U16218 ( .A1(n17466), .A2(n17457), .ZN(n17456) );
  INV_X1 U16219 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17437) );
  NAND2_X1 U16220 ( .A1(n17446), .A2(n17437), .ZN(n17436) );
  NOR2_X2 U16221 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17436), .ZN(n17420) );
  INV_X1 U16222 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17415) );
  NAND2_X1 U16223 ( .A1(n17420), .A2(n17415), .ZN(n17412) );
  NOR2_X2 U16224 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17412), .ZN(n17397) );
  INV_X1 U16225 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U16226 ( .A1(n17397), .A2(n17384), .ZN(n17387) );
  NOR2_X2 U16227 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17387), .ZN(n17374) );
  INV_X1 U16228 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17717) );
  NAND2_X1 U16229 ( .A1(n17374), .A2(n17717), .ZN(n17368) );
  INV_X1 U16230 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17607) );
  NAND2_X1 U16231 ( .A1(n17356), .A2(n17607), .ZN(n17350) );
  INV_X1 U16232 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17610) );
  NAND2_X1 U16233 ( .A1(n17335), .A2(n17610), .ZN(n17329) );
  INV_X1 U16234 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17309) );
  NAND2_X1 U16235 ( .A1(n17316), .A2(n17309), .ZN(n17308) );
  INV_X1 U16236 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17650) );
  NAND2_X1 U16237 ( .A1(n17296), .A2(n17650), .ZN(n12937) );
  NAND2_X1 U16238 ( .A1(n17584), .A2(n12937), .ZN(n17294) );
  NAND2_X1 U16239 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19472), .ZN(n19350) );
  NOR2_X1 U16240 ( .A1(n18846), .A2(n17558), .ZN(n12931) );
  NOR2_X1 U16241 ( .A1(n17581), .A2(n17593), .ZN(n17493) );
  INV_X1 U16242 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19431) );
  INV_X1 U16243 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21348) );
  INV_X1 U16244 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19426) );
  NOR2_X1 U16245 ( .A1(n21348), .A2(n19426), .ZN(n12933) );
  OAI221_X1 U16246 ( .B1(n17599), .B2(n12933), .C1(n17599), .C2(n12932), .A(
        n17573), .ZN(n17318) );
  AOI221_X1 U16247 ( .B1(n12934), .B2(n17450), .C1(n19431), .C2(n17450), .A(
        n17318), .ZN(n17278) );
  INV_X1 U16248 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19436) );
  INV_X1 U16249 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16696) );
  OAI22_X1 U16250 ( .A1(n17278), .A2(n19436), .B1(n16696), .B2(n17595), .ZN(
        n12935) );
  INV_X1 U16251 ( .A(n12935), .ZN(n12939) );
  AOI211_X4 U16252 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19471), .A(n19338), .B(
        n12936), .ZN(n17518) );
  NOR2_X1 U16253 ( .A1(n17605), .A2(n12937), .ZN(n17277) );
  OAI21_X1 U16254 ( .B1(n17518), .B2(n17277), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n12938) );
  NAND2_X1 U16255 ( .A1(n12943), .A2(n12942), .ZN(P3_U2641) );
  NAND2_X1 U16256 ( .A1(n12944), .A2(n16263), .ZN(n12952) );
  AOI21_X1 U16257 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12945), .ZN(n12948) );
  NAND2_X1 U16258 ( .A1(n12946), .A2(n16234), .ZN(n12947) );
  OAI211_X1 U16259 ( .C1(n14463), .C2(n16222), .A(n12948), .B(n12947), .ZN(
        n12949) );
  NAND2_X1 U16260 ( .A1(n9695), .A2(n19636), .ZN(n12950) );
  NAND3_X1 U16261 ( .A1(n12952), .A2(n12951), .A3(n12950), .ZN(P2_U2983) );
  NAND2_X1 U16262 ( .A1(n12979), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U16263 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19747) );
  NAND2_X1 U16264 ( .A1(n19747), .A2(n20325), .ZN(n12954) );
  NAND2_X1 U16265 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20097) );
  INV_X1 U16266 ( .A(n20097), .ZN(n20146) );
  NAND2_X1 U16267 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20146), .ZN(
        n16527) );
  NAND2_X1 U16268 ( .A1(n12954), .A2(n16527), .ZN(n19781) );
  NOR2_X1 U16269 ( .A1(n19781), .A2(n20313), .ZN(n19775) );
  AOI21_X1 U16270 ( .B1(n12972), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19775), .ZN(n12955) );
  OAI21_X2 U16271 ( .B1(n16572), .B2(n15428), .A(n12955), .ZN(n12966) );
  NAND2_X1 U16272 ( .A1(n13846), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12964) );
  INV_X1 U16273 ( .A(n20313), .ZN(n20099) );
  NAND2_X1 U16274 ( .A1(n20335), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19971) );
  NOR2_X1 U16275 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20335), .ZN(
        n19935) );
  INV_X1 U16276 ( .A(n19935), .ZN(n19808) );
  NAND2_X1 U16277 ( .A1(n19971), .A2(n19808), .ZN(n19780) );
  AND2_X1 U16278 ( .A1(n20099), .A2(n19780), .ZN(n19838) );
  AOI21_X1 U16279 ( .B1(n12972), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19838), .ZN(n12957) );
  INV_X1 U16280 ( .A(n15428), .ZN(n12968) );
  NOR2_X1 U16281 ( .A1(n20313), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12958) );
  AOI21_X1 U16282 ( .B1(n12972), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12958), .ZN(n12959) );
  NAND2_X1 U16283 ( .A1(n13846), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12961) );
  INV_X1 U16284 ( .A(n12961), .ZN(n12962) );
  NOR2_X1 U16285 ( .A1(n13644), .A2(n12962), .ZN(n12963) );
  INV_X1 U16286 ( .A(n12964), .ZN(n12965) );
  NAND2_X1 U16287 ( .A1(n12966), .A2(n12965), .ZN(n12967) );
  NAND2_X1 U16288 ( .A1(n13865), .A2(n12968), .ZN(n12974) );
  INV_X1 U16289 ( .A(n19747), .ZN(n20003) );
  NAND2_X1 U16290 ( .A1(n20317), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19841) );
  INV_X1 U16291 ( .A(n19841), .ZN(n12969) );
  NAND2_X1 U16292 ( .A1(n20003), .A2(n12969), .ZN(n19911) );
  NAND2_X1 U16293 ( .A1(n16527), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12970) );
  NAND2_X1 U16294 ( .A1(n19911), .A2(n12970), .ZN(n12971) );
  AND2_X1 U16295 ( .A1(n12971), .A2(n20099), .ZN(n20033) );
  AOI21_X1 U16296 ( .B1(n12972), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20033), .ZN(n12973) );
  NAND2_X1 U16297 ( .A1(n12974), .A2(n12973), .ZN(n12977) );
  INV_X1 U16298 ( .A(n13846), .ZN(n13163) );
  INV_X1 U16299 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12975) );
  NAND2_X1 U16300 ( .A1(n12977), .A2(n12976), .ZN(n12981) );
  OR2_X1 U16301 ( .A1(n12977), .A2(n12976), .ZN(n12978) );
  NAND2_X1 U16302 ( .A1(n13784), .A2(n13783), .ZN(n12983) );
  NAND2_X1 U16303 ( .A1(n12979), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12980) );
  AND2_X1 U16304 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  AND2_X1 U16305 ( .A1(n13991), .A2(n13993), .ZN(n13911) );
  NAND2_X1 U16306 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13878) );
  NAND2_X1 U16307 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12984) );
  NOR2_X1 U16308 ( .A1(n13878), .A2(n12984), .ZN(n13910) );
  AND4_X1 U16309 ( .A1(n13846), .A2(n13911), .A3(n13910), .A4(n13912), .ZN(
        n12985) );
  AOI22_X1 U16310 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U16311 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16312 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16313 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12986) );
  NAND4_X1 U16314 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        n12995) );
  AOI22_X1 U16315 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16316 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16317 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16318 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12990) );
  NAND4_X1 U16319 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n12990), .ZN(
        n12994) );
  OR2_X1 U16320 ( .A1(n12995), .A2(n12994), .ZN(n15869) );
  AND2_X1 U16321 ( .A1(n15874), .A2(n15869), .ZN(n12996) );
  NAND4_X1 U16322 ( .A1(n12996), .A2(n15879), .A3(n15885), .A4(n14050), .ZN(
        n12997) );
  AOI22_X1 U16323 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16324 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16325 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16326 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12998) );
  NAND4_X1 U16327 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13007) );
  AOI22_X1 U16328 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16329 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16330 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16331 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13002) );
  NAND4_X1 U16332 ( .A1(n13005), .A2(n13004), .A3(n13003), .A4(n13002), .ZN(
        n13006) );
  OR2_X1 U16333 ( .A1(n13007), .A2(n13006), .ZN(n14155) );
  INV_X2 U16334 ( .A(n14154), .ZN(n13019) );
  AOI22_X1 U16335 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U16336 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U16337 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13009) );
  AOI22_X1 U16338 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13008) );
  NAND4_X1 U16339 ( .A1(n13011), .A2(n13010), .A3(n13009), .A4(n13008), .ZN(
        n13017) );
  AOI22_X1 U16340 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U16341 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16342 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16343 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13012) );
  NAND4_X1 U16344 ( .A1(n13015), .A2(n13014), .A3(n13013), .A4(n13012), .ZN(
        n13016) );
  NOR2_X1 U16345 ( .A1(n13017), .A2(n13016), .ZN(n15862) );
  INV_X1 U16346 ( .A(n15862), .ZN(n13018) );
  AOI22_X1 U16347 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U16348 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16349 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16350 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13020) );
  NAND4_X1 U16351 ( .A1(n13023), .A2(n13022), .A3(n13021), .A4(n13020), .ZN(
        n13029) );
  AOI22_X1 U16352 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U16353 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16354 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16355 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13024) );
  NAND4_X1 U16356 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        n13028) );
  NOR2_X1 U16357 ( .A1(n13029), .A2(n13028), .ZN(n15854) );
  AOI22_X1 U16358 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U16359 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16360 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U16361 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13030) );
  NAND4_X1 U16362 ( .A1(n13033), .A2(n13032), .A3(n13031), .A4(n13030), .ZN(
        n13039) );
  AOI22_X1 U16363 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16364 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16365 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U16366 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13034) );
  NAND4_X1 U16367 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n13038) );
  OR2_X1 U16368 ( .A1(n13039), .A2(n13038), .ZN(n15849) );
  AOI22_X1 U16369 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16370 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16371 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16372 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13040) );
  NAND4_X1 U16373 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13040), .ZN(
        n13049) );
  AOI22_X1 U16374 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16375 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16376 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16377 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13044) );
  NAND4_X1 U16378 ( .A1(n13047), .A2(n13046), .A3(n13045), .A4(n13044), .ZN(
        n13048) );
  OR2_X1 U16379 ( .A1(n13049), .A2(n13048), .ZN(n15844) );
  AOI22_X1 U16380 ( .A1(n13060), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16381 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16382 ( .A1(n12105), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U16383 ( .A1(n13866), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13050) );
  NAND4_X1 U16384 ( .A1(n13053), .A2(n13052), .A3(n13051), .A4(n13050), .ZN(
        n13059) );
  AOI22_X1 U16385 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16386 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16387 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16388 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13054) );
  NAND4_X1 U16389 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        n13058) );
  NOR2_X1 U16390 ( .A1(n13059), .A2(n13058), .ZN(n15840) );
  OR2_X2 U16391 ( .A1(n15837), .A2(n15840), .ZN(n15821) );
  AOI22_X1 U16392 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11989), .B1(
        n13060), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16393 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16394 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n12105), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16395 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12104), .B1(
        n13866), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13061) );
  NAND4_X1 U16396 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13075) );
  AOI22_X1 U16397 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16398 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U16399 ( .A1(n11930), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13067), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16400 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13068), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13070) );
  NAND4_X1 U16401 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13074) );
  OR2_X1 U16402 ( .A1(n13075), .A2(n13074), .ZN(n13110) );
  AOI22_X1 U16403 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16404 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13079) );
  AND2_X1 U16405 ( .A1(n13080), .A2(n13079), .ZN(n13086) );
  AOI22_X1 U16406 ( .A1(n16574), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13084) );
  XNOR2_X1 U16407 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13203) );
  NAND4_X1 U16408 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13203), .ZN(
        n13093) );
  AOI22_X1 U16409 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16410 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13087) );
  AND2_X1 U16411 ( .A1(n13088), .A2(n13087), .ZN(n13091) );
  INV_X1 U16412 ( .A(n13203), .ZN(n13213) );
  AOI22_X1 U16413 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13090) );
  NAND4_X1 U16414 ( .A1(n13091), .A2(n13213), .A3(n13090), .A4(n13089), .ZN(
        n13092) );
  AND2_X1 U16415 ( .A1(n13093), .A2(n13092), .ZN(n15822) );
  AND2_X1 U16416 ( .A1(n13110), .A2(n15822), .ZN(n13106) );
  AOI22_X1 U16417 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16418 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13094) );
  AND2_X1 U16419 ( .A1(n13095), .A2(n13094), .ZN(n13098) );
  AOI22_X1 U16420 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13097) );
  NAND4_X1 U16421 ( .A1(n13098), .A2(n13097), .A3(n13096), .A4(n13203), .ZN(
        n13105) );
  AOI22_X1 U16422 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16423 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13099) );
  AND2_X1 U16424 ( .A1(n13100), .A2(n13099), .ZN(n13103) );
  AOI22_X1 U16425 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13102) );
  NAND4_X1 U16426 ( .A1(n13103), .A2(n13213), .A3(n13102), .A4(n13101), .ZN(
        n13104) );
  AND2_X1 U16427 ( .A1(n13105), .A2(n13104), .ZN(n13107) );
  NAND2_X1 U16428 ( .A1(n13106), .A2(n13107), .ZN(n13115) );
  INV_X1 U16429 ( .A(n13106), .ZN(n13108) );
  INV_X1 U16430 ( .A(n13107), .ZN(n13112) );
  NAND2_X1 U16431 ( .A1(n13108), .A2(n13112), .ZN(n13109) );
  AND3_X1 U16432 ( .A1(n13115), .A2(n13846), .A3(n13109), .ZN(n15825) );
  NAND2_X1 U16433 ( .A1(n15822), .A2(n15806), .ZN(n13111) );
  XNOR2_X1 U16434 ( .A(n13111), .B(n13110), .ZN(n15823) );
  NAND2_X1 U16435 ( .A1(n15825), .A2(n15823), .ZN(n13114) );
  NOR2_X1 U16436 ( .A1(n15806), .A2(n13112), .ZN(n15824) );
  NAND3_X1 U16437 ( .A1(n15823), .A2(n15822), .A3(n15824), .ZN(n13113) );
  OAI21_X2 U16438 ( .B1(n15821), .B2(n13114), .A(n13113), .ZN(n13145) );
  INV_X1 U16439 ( .A(n13115), .ZN(n13128) );
  AOI22_X1 U16440 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16441 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13116) );
  AND2_X1 U16442 ( .A1(n13117), .A2(n13116), .ZN(n13120) );
  AOI22_X1 U16443 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13119) );
  NAND4_X1 U16444 ( .A1(n13120), .A2(n13119), .A3(n13118), .A4(n13203), .ZN(
        n13127) );
  AOI22_X1 U16445 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16446 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13121) );
  AND2_X1 U16447 ( .A1(n13122), .A2(n13121), .ZN(n13125) );
  AOI22_X1 U16448 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13124) );
  NAND4_X1 U16449 ( .A1(n13125), .A2(n13213), .A3(n13124), .A4(n13123), .ZN(
        n13126) );
  AND2_X1 U16450 ( .A1(n13127), .A2(n13126), .ZN(n13129) );
  NAND2_X1 U16451 ( .A1(n13128), .A2(n13129), .ZN(n13147) );
  OAI211_X1 U16452 ( .C1(n13128), .C2(n13129), .A(n13147), .B(n13846), .ZN(
        n13143) );
  XNOR2_X1 U16453 ( .A(n13145), .B(n13143), .ZN(n15804) );
  INV_X1 U16454 ( .A(n13129), .ZN(n13130) );
  NOR2_X1 U16455 ( .A1(n15806), .A2(n13130), .ZN(n15817) );
  AOI22_X1 U16456 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16457 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13131) );
  AND2_X1 U16458 ( .A1(n13132), .A2(n13131), .ZN(n13135) );
  AOI22_X1 U16459 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13134) );
  NAND4_X1 U16460 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13203), .ZN(
        n13142) );
  AOI22_X1 U16461 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16462 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13136) );
  AND2_X1 U16463 ( .A1(n13137), .A2(n13136), .ZN(n13140) );
  AOI22_X1 U16464 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13139) );
  NAND4_X1 U16465 ( .A1(n13140), .A2(n13213), .A3(n13139), .A4(n13138), .ZN(
        n13141) );
  AND2_X1 U16466 ( .A1(n13142), .A2(n13141), .ZN(n13146) );
  AND2_X1 U16467 ( .A1(n15817), .A2(n13146), .ZN(n13150) );
  INV_X1 U16468 ( .A(n13143), .ZN(n13144) );
  INV_X1 U16469 ( .A(n13146), .ZN(n15807) );
  AOI21_X1 U16470 ( .B1(n13147), .B2(n15807), .A(n13163), .ZN(n13148) );
  OR2_X1 U16471 ( .A1(n13147), .A2(n15807), .ZN(n13164) );
  AND2_X1 U16472 ( .A1(n13148), .A2(n13164), .ZN(n15809) );
  AOI22_X1 U16473 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U16474 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13151) );
  AND2_X1 U16475 ( .A1(n13152), .A2(n13151), .ZN(n13155) );
  AOI22_X1 U16476 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13154) );
  NAND4_X1 U16477 ( .A1(n13155), .A2(n13154), .A3(n13153), .A4(n13203), .ZN(
        n13162) );
  AOI22_X1 U16478 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16479 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13156) );
  AND2_X1 U16480 ( .A1(n13157), .A2(n13156), .ZN(n13160) );
  AOI22_X1 U16481 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13159) );
  NAND4_X1 U16482 ( .A1(n13160), .A2(n13213), .A3(n13159), .A4(n13158), .ZN(
        n13161) );
  NAND2_X1 U16483 ( .A1(n13162), .A2(n13161), .ZN(n13168) );
  AOI21_X1 U16484 ( .B1(n13164), .B2(n13168), .A(n13163), .ZN(n13165) );
  OR2_X1 U16485 ( .A1(n13164), .A2(n13168), .ZN(n13194) );
  NAND2_X1 U16486 ( .A1(n13165), .A2(n13194), .ZN(n13166) );
  NOR2_X1 U16487 ( .A1(n15806), .A2(n13168), .ZN(n15800) );
  AOI22_X1 U16488 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U16489 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13169) );
  AND2_X1 U16490 ( .A1(n13170), .A2(n13169), .ZN(n13173) );
  AOI22_X1 U16491 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13172) );
  NAND4_X1 U16492 ( .A1(n13173), .A2(n13172), .A3(n13171), .A4(n13203), .ZN(
        n13180) );
  AOI22_X1 U16493 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16494 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13174) );
  AND2_X1 U16495 ( .A1(n13175), .A2(n13174), .ZN(n13178) );
  AOI22_X1 U16496 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13177) );
  NAND4_X1 U16497 ( .A1(n13178), .A2(n13213), .A3(n13177), .A4(n13176), .ZN(
        n13179) );
  NAND2_X1 U16498 ( .A1(n13180), .A2(n13179), .ZN(n15794) );
  AOI22_X1 U16499 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16500 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13181) );
  AND2_X1 U16501 ( .A1(n13182), .A2(n13181), .ZN(n13185) );
  AOI22_X1 U16502 ( .A1(n16574), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13183) );
  NAND4_X1 U16503 ( .A1(n13185), .A2(n13184), .A3(n13183), .A4(n13203), .ZN(
        n13193) );
  AOI22_X1 U16504 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U16505 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13186) );
  AND2_X1 U16506 ( .A1(n13187), .A2(n13186), .ZN(n13191) );
  AOI22_X1 U16507 ( .A1(n16574), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13189) );
  NAND4_X1 U16508 ( .A1(n13191), .A2(n13213), .A3(n13190), .A4(n13189), .ZN(
        n13192) );
  NAND2_X1 U16509 ( .A1(n13193), .A2(n13192), .ZN(n13198) );
  INV_X1 U16510 ( .A(n13194), .ZN(n15792) );
  INV_X1 U16511 ( .A(n15794), .ZN(n13195) );
  AND2_X1 U16512 ( .A1(n15806), .A2(n13195), .ZN(n13196) );
  NAND2_X1 U16513 ( .A1(n15792), .A2(n13196), .ZN(n13197) );
  NOR2_X1 U16514 ( .A1(n13197), .A2(n13198), .ZN(n13199) );
  AOI21_X1 U16515 ( .B1(n13198), .B2(n13197), .A(n13199), .ZN(n15786) );
  NAND2_X1 U16516 ( .A1(n15787), .A2(n15786), .ZN(n15788) );
  INV_X1 U16517 ( .A(n13199), .ZN(n13200) );
  NAND2_X1 U16518 ( .A1(n15788), .A2(n13200), .ZN(n13222) );
  AOI22_X1 U16519 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16574), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13201) );
  NAND2_X1 U16520 ( .A1(n13202), .A2(n13201), .ZN(n13219) );
  AOI22_X1 U16521 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16522 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13204) );
  NAND3_X1 U16523 ( .A1(n13205), .A2(n13204), .A3(n13203), .ZN(n13218) );
  AOI22_X1 U16524 ( .A1(n13207), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13206), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16525 ( .A1(n13209), .A2(n13208), .ZN(n13217) );
  AOI22_X1 U16526 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13210), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U16527 ( .A1(n13212), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13211), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13214) );
  NAND3_X1 U16528 ( .A1(n13215), .A2(n13214), .A3(n13213), .ZN(n13216) );
  OAI22_X1 U16529 ( .A1(n13219), .A2(n13218), .B1(n13217), .B2(n13216), .ZN(
        n13220) );
  XNOR2_X1 U16530 ( .A(n13222), .B(n13221), .ZN(n14385) );
  INV_X1 U16531 ( .A(n13223), .ZN(n13224) );
  NAND2_X1 U16532 ( .A1(n13224), .A2(n15430), .ZN(n13225) );
  NOR2_X1 U16533 ( .A1(n12291), .A2(n13225), .ZN(n13226) );
  AOI21_X1 U16534 ( .B1(n16592), .B2(n16594), .A(n13226), .ZN(n13636) );
  NAND2_X1 U16535 ( .A1(n13636), .A2(n13227), .ZN(n13228) );
  AND2_X1 U16536 ( .A1(n16558), .A2(n16566), .ZN(n13231) );
  NOR4_X1 U16537 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13235) );
  NOR4_X1 U16538 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13234) );
  NOR4_X1 U16539 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13233) );
  NOR4_X1 U16540 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13232) );
  AND4_X1 U16541 ( .A1(n13235), .A2(n13234), .A3(n13233), .A4(n13232), .ZN(
        n13240) );
  NOR4_X1 U16542 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_1__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n13238) );
  NOR4_X1 U16543 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13237) );
  NOR4_X1 U16544 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13236) );
  INV_X1 U16545 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20237) );
  AND4_X1 U16546 ( .A1(n13238), .A2(n13237), .A3(n13236), .A4(n20237), .ZN(
        n13239) );
  NAND2_X1 U16547 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  NAND2_X1 U16548 ( .A1(n15983), .A2(BUF1_REG_30__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U16549 ( .A1(n15984), .A2(BUF2_REG_30__SCAN_IN), .ZN(n13245) );
  INV_X1 U16550 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13243) );
  INV_X2 U16551 ( .A(n16533), .ZN(n13618) );
  NAND2_X1 U16552 ( .A1(n13618), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13242) );
  OAI21_X1 U16553 ( .B1(n13618), .B2(n13243), .A(n13242), .ZN(n19627) );
  AOI22_X1 U16554 ( .A1(n15985), .A2(n19627), .B1(n16010), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n13244) );
  NAND3_X1 U16555 ( .A1(n13246), .A2(n13245), .A3(n13244), .ZN(n13247) );
  AOI21_X1 U16556 ( .B1(n13248), .B2(n19578), .A(n13247), .ZN(n13249) );
  OAI21_X1 U16557 ( .B1(n14385), .B2(n16013), .A(n13249), .ZN(P2_U2889) );
  NAND2_X1 U16558 ( .A1(n13250), .A2(n19672), .ZN(n13265) );
  NAND2_X1 U16559 ( .A1(n9690), .A2(n13253), .ZN(n13254) );
  NAND2_X1 U16560 ( .A1(n15543), .A2(n13254), .ZN(n15557) );
  OAI21_X1 U16561 ( .B1(n13255), .B2(n16408), .A(n9631), .ZN(n16320) );
  INV_X1 U16562 ( .A(n13256), .ZN(n13258) );
  NAND2_X1 U16563 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14297) );
  NOR3_X1 U16564 ( .A1(n16307), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n14297), .ZN(n13257) );
  AOI211_X1 U16565 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n16320), .A(
        n13258), .B(n13257), .ZN(n13259) );
  OAI21_X1 U16566 ( .B1(n19648), .B2(n15557), .A(n13259), .ZN(n13260) );
  AOI21_X1 U16567 ( .B1(n15845), .B2(n19669), .A(n13260), .ZN(n13261) );
  NOR2_X1 U16568 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  NAND2_X1 U16569 ( .A1(n13265), .A2(n13264), .ZN(P2_U3025) );
  OR2_X2 U16570 ( .A1(n20611), .A2(n10432), .ZN(n13274) );
  INV_X1 U16571 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13267) );
  OAI22_X1 U16572 ( .A1(n13274), .A2(n13267), .B1(n14305), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13777) );
  NAND2_X1 U16573 ( .A1(n13269), .A2(n10304), .ZN(n13270) );
  XNOR2_X1 U16574 ( .A(n13777), .B(n13270), .ZN(n13768) );
  INV_X1 U16575 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n20443) );
  NAND2_X1 U16576 ( .A1(n13347), .A2(n20443), .ZN(n13273) );
  INV_X2 U16577 ( .A(n10302), .ZN(n13376) );
  NAND2_X1 U16578 ( .A1(n14305), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13271) );
  OAI211_X1 U16579 ( .C1(n13376), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13274), .B(
        n13271), .ZN(n13272) );
  MUX2_X1 U16580 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13278) );
  INV_X1 U16581 ( .A(n13274), .ZN(n13275) );
  NAND2_X1 U16582 ( .A1(n13275), .A2(n13376), .ZN(n13296) );
  NAND2_X1 U16583 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13376), .ZN(
        n13276) );
  AND2_X1 U16584 ( .A1(n13296), .A2(n13276), .ZN(n13277) );
  NAND2_X1 U16585 ( .A1(n13278), .A2(n13277), .ZN(n13887) );
  NAND2_X1 U16586 ( .A1(n13839), .A2(n13887), .ZN(n13886) );
  INV_X1 U16587 ( .A(n13886), .ZN(n13282) );
  NAND2_X1 U16588 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13279) );
  OAI211_X1 U16589 ( .C1(n13376), .C2(P1_EBX_REG_4__SCAN_IN), .A(n13274), .B(
        n13279), .ZN(n13280) );
  OAI21_X1 U16590 ( .B1(n13337), .B2(P1_EBX_REG_4__SCAN_IN), .A(n13280), .ZN(
        n20410) );
  NAND2_X1 U16591 ( .A1(n13282), .A2(n13281), .ZN(n14005) );
  MUX2_X1 U16592 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n13285) );
  NAND2_X1 U16593 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13376), .ZN(
        n13283) );
  AND2_X1 U16594 ( .A1(n13296), .A2(n13283), .ZN(n13284) );
  NAND2_X1 U16595 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13287) );
  OAI211_X1 U16596 ( .C1(n13376), .C2(P1_EBX_REG_6__SCAN_IN), .A(n13274), .B(
        n13287), .ZN(n13288) );
  OAI21_X1 U16597 ( .B1(n13337), .B2(P1_EBX_REG_6__SCAN_IN), .A(n13288), .ZN(
        n17117) );
  MUX2_X1 U16598 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13291) );
  NAND2_X1 U16599 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n13376), .ZN(
        n13289) );
  AND2_X1 U16600 ( .A1(n13296), .A2(n13289), .ZN(n13290) );
  NAND2_X1 U16601 ( .A1(n13291), .A2(n13290), .ZN(n14203) );
  INV_X1 U16602 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13292) );
  MUX2_X1 U16603 ( .A(n13360), .B(n13347), .S(n13292), .Z(n13294) );
  NOR2_X1 U16604 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13293) );
  NOR2_X1 U16605 ( .A1(n13294), .A2(n13293), .ZN(n14217) );
  MUX2_X1 U16606 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13298) );
  NAND2_X1 U16607 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n13376), .ZN(
        n13295) );
  AND2_X1 U16608 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  NAND2_X1 U16609 ( .A1(n13298), .A2(n13297), .ZN(n14234) );
  MUX2_X1 U16610 ( .A(n13347), .B(n13360), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13299) );
  INV_X1 U16611 ( .A(n13299), .ZN(n13300) );
  NAND2_X1 U16612 ( .A1(n13300), .A2(n10300), .ZN(n14735) );
  INV_X1 U16613 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21357) );
  NAND2_X1 U16614 ( .A1(n13347), .A2(n21357), .ZN(n13303) );
  NAND2_X1 U16615 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13301) );
  OAI211_X1 U16616 ( .C1(n13376), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13274), .B(
        n13301), .ZN(n13302) );
  INV_X1 U16617 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15346) );
  NAND2_X1 U16618 ( .A1(n13274), .A2(n15346), .ZN(n13304) );
  OAI211_X1 U16619 ( .C1(n13376), .C2(P1_EBX_REG_11__SCAN_IN), .A(n13361), .B(
        n13304), .ZN(n13305) );
  OAI21_X1 U16620 ( .B1(n13338), .B2(P1_EBX_REG_11__SCAN_IN), .A(n13305), .ZN(
        n14718) );
  MUX2_X1 U16621 ( .A(n13347), .B(n13360), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13307) );
  NOR2_X1 U16622 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13306) );
  NOR2_X1 U16623 ( .A1(n13307), .A2(n13306), .ZN(n14675) );
  MUX2_X1 U16624 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13309) );
  NAND2_X1 U16625 ( .A1(n13376), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13308) );
  NAND2_X1 U16626 ( .A1(n13309), .A2(n13308), .ZN(n14687) );
  NAND2_X1 U16627 ( .A1(n14704), .A2(n13310), .ZN(n14657) );
  MUX2_X1 U16628 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13312) );
  NAND2_X1 U16629 ( .A1(n13376), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13311) );
  NAND2_X1 U16630 ( .A1(n13312), .A2(n13311), .ZN(n14659) );
  INV_X1 U16631 ( .A(n14659), .ZN(n13313) );
  NOR2_X2 U16632 ( .A1(n14657), .A2(n13313), .ZN(n14644) );
  NAND2_X1 U16633 ( .A1(n14305), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13314) );
  OAI211_X1 U16634 ( .C1(n13376), .C2(P1_EBX_REG_16__SCAN_IN), .A(n13274), .B(
        n13314), .ZN(n13315) );
  OAI21_X1 U16635 ( .B1(n13337), .B2(P1_EBX_REG_16__SCAN_IN), .A(n13315), .ZN(
        n14645) );
  INV_X1 U16636 ( .A(n14645), .ZN(n13316) );
  NAND2_X1 U16637 ( .A1(n13274), .A2(n15283), .ZN(n13317) );
  OAI211_X1 U16638 ( .C1(n13376), .C2(P1_EBX_REG_17__SCAN_IN), .A(n13361), .B(
        n13317), .ZN(n13318) );
  OAI21_X1 U16639 ( .B1(n13338), .B2(P1_EBX_REG_17__SCAN_IN), .A(n13318), .ZN(
        n14632) );
  NAND2_X1 U16640 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13319) );
  OAI211_X1 U16641 ( .C1(n13376), .C2(P1_EBX_REG_18__SCAN_IN), .A(n13274), .B(
        n13319), .ZN(n13320) );
  OAI21_X1 U16642 ( .B1(n13337), .B2(P1_EBX_REG_18__SCAN_IN), .A(n13320), .ZN(
        n14617) );
  INV_X1 U16643 ( .A(n13338), .ZN(n13357) );
  INV_X1 U16644 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U16645 ( .A1(n13357), .A2(n13321), .ZN(n13324) );
  NAND2_X1 U16646 ( .A1(n13274), .A2(n10709), .ZN(n13322) );
  OAI211_X1 U16647 ( .C1(n13376), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13361), .B(
        n13322), .ZN(n13323) );
  INV_X1 U16648 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14819) );
  NAND2_X1 U16649 ( .A1(n13347), .A2(n14819), .ZN(n13327) );
  NAND2_X1 U16650 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13325) );
  OAI211_X1 U16651 ( .C1(n13376), .C2(P1_EBX_REG_20__SCAN_IN), .A(n13274), .B(
        n13325), .ZN(n13326) );
  NAND2_X1 U16652 ( .A1(n13274), .A2(n15011), .ZN(n13328) );
  OAI211_X1 U16653 ( .C1(n13376), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14305), .B(
        n13328), .ZN(n13329) );
  OAI21_X1 U16654 ( .B1(n13338), .B2(P1_EBX_REG_21__SCAN_IN), .A(n13329), .ZN(
        n14565) );
  NAND2_X1 U16655 ( .A1(n14564), .A2(n14565), .ZN(n14553) );
  NAND2_X1 U16656 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13330) );
  OAI211_X1 U16657 ( .C1(n13376), .C2(P1_EBX_REG_22__SCAN_IN), .A(n13274), .B(
        n13330), .ZN(n13331) );
  OAI21_X1 U16658 ( .B1(n13337), .B2(P1_EBX_REG_22__SCAN_IN), .A(n13331), .ZN(
        n14555) );
  MUX2_X1 U16659 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13333) );
  NAND2_X1 U16660 ( .A1(n13376), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13332) );
  AND2_X1 U16661 ( .A1(n13333), .A2(n13332), .ZN(n14543) );
  NAND2_X1 U16662 ( .A1(n13361), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13335) );
  OAI211_X1 U16663 ( .C1(n13376), .C2(P1_EBX_REG_24__SCAN_IN), .A(n13274), .B(
        n13335), .ZN(n13336) );
  OAI21_X1 U16664 ( .B1(n13337), .B2(P1_EBX_REG_24__SCAN_IN), .A(n13336), .ZN(
        n14523) );
  MUX2_X1 U16665 ( .A(n13338), .B(n13274), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13340) );
  NAND2_X1 U16666 ( .A1(n13376), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13339) );
  NAND2_X1 U16667 ( .A1(n13340), .A2(n13339), .ZN(n14512) );
  MUX2_X1 U16668 ( .A(n13347), .B(n13360), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13341) );
  INV_X1 U16669 ( .A(n13341), .ZN(n13344) );
  INV_X1 U16670 ( .A(n14307), .ZN(n13342) );
  NAND2_X1 U16671 ( .A1(n13342), .A2(n15182), .ZN(n13343) );
  NAND2_X1 U16672 ( .A1(n13344), .A2(n13343), .ZN(n14497) );
  INV_X1 U16673 ( .A(n14497), .ZN(n13345) );
  NAND2_X1 U16674 ( .A1(n13346), .A2(n13345), .ZN(n14469) );
  MUX2_X1 U16675 ( .A(n13347), .B(n13360), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13349) );
  NOR2_X1 U16676 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13348) );
  NOR2_X1 U16677 ( .A1(n13349), .A2(n13348), .ZN(n14470) );
  INV_X1 U16678 ( .A(n14470), .ZN(n13354) );
  INV_X1 U16679 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U16680 ( .A1(n13357), .A2(n13350), .ZN(n13353) );
  NAND2_X1 U16681 ( .A1(n13274), .A2(n14956), .ZN(n13351) );
  OAI211_X1 U16682 ( .C1(n13376), .C2(P1_EBX_REG_27__SCAN_IN), .A(n14305), .B(
        n13351), .ZN(n13352) );
  AND2_X1 U16683 ( .A1(n13353), .A2(n13352), .ZN(n14483) );
  OR2_X1 U16684 ( .A1(n13376), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U16685 ( .B1(n14307), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13356), .ZN(n13363) );
  OR2_X1 U16686 ( .A1(n13363), .A2(n13360), .ZN(n13359) );
  INV_X1 U16687 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U16688 ( .A1(n13357), .A2(n14459), .ZN(n13358) );
  NAND2_X1 U16689 ( .A1(n13359), .A2(n13358), .ZN(n14454) );
  NAND2_X1 U16690 ( .A1(n14472), .A2(n14454), .ZN(n14304) );
  NAND2_X1 U16691 ( .A1(n14304), .A2(n13360), .ZN(n13364) );
  INV_X1 U16692 ( .A(n14472), .ZN(n13362) );
  AOI22_X1 U16693 ( .A1(n14307), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13376), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14306) );
  INV_X1 U16694 ( .A(n14306), .ZN(n13365) );
  XNOR2_X1 U16695 ( .A(n13366), .B(n13365), .ZN(n14323) );
  INV_X1 U16696 ( .A(n14323), .ZN(n14357) );
  NOR3_X1 U16697 ( .A1(n13369), .A2(n13368), .A3(n13367), .ZN(n13371) );
  OAI21_X1 U16698 ( .B1(n13372), .B2(n13371), .A(n13370), .ZN(n13714) );
  AND2_X1 U16699 ( .A1(n13714), .A2(n13719), .ZN(n13657) );
  INV_X1 U16700 ( .A(n20348), .ZN(n13828) );
  NAND2_X1 U16701 ( .A1(n13657), .A2(n13828), .ZN(n21294) );
  NOR2_X1 U16702 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21296) );
  NAND2_X1 U16703 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21296), .ZN(n17127) );
  OR2_X1 U16704 ( .A1(n17125), .A2(n13431), .ZN(n13434) );
  OAI211_X1 U16705 ( .C1(n17127), .C2(n20351), .A(n20416), .B(n13434), .ZN(
        n13373) );
  INV_X1 U16706 ( .A(n13373), .ZN(n13374) );
  INV_X1 U16707 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14315) );
  OR2_X1 U16708 ( .A1(n13376), .A2(n14315), .ZN(n13399) );
  NAND2_X1 U16709 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21293) );
  NAND2_X1 U16710 ( .A1(n21293), .A2(n20900), .ZN(n17057) );
  INV_X1 U16711 ( .A(n17057), .ZN(n13386) );
  NOR2_X1 U16712 ( .A1(n13399), .A2(n13386), .ZN(n13377) );
  INV_X1 U16713 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14314) );
  INV_X1 U16714 ( .A(n13434), .ZN(n13382) );
  INV_X2 U16715 ( .A(n20426), .ZN(n20402) );
  INV_X1 U16716 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13383) );
  XNOR2_X1 U16717 ( .A(n13384), .B(n13383), .ZN(n14331) );
  AND2_X1 U16718 ( .A1(n13385), .A2(n21251), .ZN(n13787) );
  OAI21_X1 U16719 ( .B1(n10431), .B2(n13787), .A(n13386), .ZN(n13398) );
  NOR2_X1 U16720 ( .A1(n13398), .A2(n10432), .ZN(n13387) );
  AND2_X1 U16721 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14499) );
  INV_X1 U16722 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21264) );
  INV_X1 U16723 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21260) );
  INV_X1 U16724 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20381) );
  INV_X1 U16725 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20400) );
  NAND4_X1 U16726 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20398)
         );
  NOR2_X1 U16727 ( .A1(n20400), .A2(n20398), .ZN(n20383) );
  NAND2_X1 U16728 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20383), .ZN(n20372) );
  NOR3_X1 U16729 ( .A1(n21260), .A2(n20381), .A3(n20372), .ZN(n14750) );
  NAND2_X1 U16730 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n14750), .ZN(n14738) );
  INV_X1 U16731 ( .A(n14738), .ZN(n13388) );
  NAND2_X1 U16732 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n13388), .ZN(n14720) );
  NAND2_X1 U16733 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n13389) );
  NOR2_X1 U16734 ( .A1(n14720), .A2(n13389), .ZN(n14598) );
  NAND2_X1 U16735 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14605) );
  INV_X1 U16736 ( .A(n14605), .ZN(n13390) );
  NAND2_X1 U16737 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n13390), .ZN(n14601) );
  NAND2_X1 U16738 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n13391) );
  NOR2_X1 U16739 ( .A1(n14601), .A2(n13391), .ZN(n13392) );
  NAND2_X1 U16740 ( .A1(n14598), .A2(n13392), .ZN(n14586) );
  INV_X1 U16741 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15023) );
  INV_X1 U16742 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15092) );
  INV_X1 U16743 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15105) );
  NOR2_X1 U16744 ( .A1(n15092), .A2(n15105), .ZN(n14600) );
  INV_X1 U16745 ( .A(n14600), .ZN(n14585) );
  OR3_X1 U16746 ( .A1(n14586), .A2(n15023), .A3(n14585), .ZN(n14572) );
  INV_X1 U16747 ( .A(n14572), .ZN(n13393) );
  NAND2_X1 U16748 ( .A1(n13393), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14556) );
  NOR2_X1 U16749 ( .A1(n21264), .A2(n14556), .ZN(n14538) );
  AND2_X1 U16750 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14538), .ZN(n14514) );
  AND3_X1 U16751 ( .A1(n14499), .A2(n14514), .A3(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14489) );
  AND2_X1 U16752 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n13394) );
  NAND2_X1 U16753 ( .A1(n14489), .A2(n13394), .ZN(n13396) );
  INV_X1 U16754 ( .A(n13396), .ZN(n13395) );
  NAND2_X1 U16755 ( .A1(n20433), .A2(n13395), .ZN(n14453) );
  INV_X1 U16756 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n13544) );
  NOR2_X1 U16757 ( .A1(n14453), .A2(n13544), .ZN(n13397) );
  AND2_X1 U16758 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14316) );
  NOR2_X1 U16759 ( .A1(n20399), .A2(n13396), .ZN(n14450) );
  INV_X1 U16760 ( .A(n20399), .ZN(n20428) );
  AOI21_X1 U16761 ( .B1(n14316), .B2(n14450), .A(n14798), .ZN(n14320) );
  OAI21_X1 U16762 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n13397), .A(n14320), 
        .ZN(n13402) );
  AND3_X1 U16763 ( .A1(n13399), .A2(n10476), .A3(n13398), .ZN(n13400) );
  AND2_X2 U16764 ( .A1(n14779), .A2(n13400), .ZN(n20411) );
  NOR2_X2 U16765 ( .A1(n20399), .A2(n21041), .ZN(n20430) );
  AOI22_X1 U16766 ( .A1(n20411), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20430), .ZN(n13401) );
  OAI211_X1 U16767 ( .C1(n20402), .C2(n14331), .A(n13402), .B(n13401), .ZN(
        n13403) );
  AOI21_X1 U16768 ( .B1(n14357), .B2(n20425), .A(n13403), .ZN(n13437) );
  AOI22_X1 U16769 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10531), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U16770 ( .A1(n13404), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11123), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U16771 ( .A1(n10467), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13405), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U16772 ( .A1(n9613), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13406) );
  NAND4_X1 U16773 ( .A1(n13409), .A2(n13408), .A3(n13407), .A4(n13406), .ZN(
        n13420) );
  AOI22_X1 U16774 ( .A1(n13410), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U16775 ( .A1(n10561), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13411), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16776 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U16777 ( .A1(n13414), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13415) );
  NAND4_X1 U16778 ( .A1(n13418), .A2(n13417), .A3(n13416), .A4(n13415), .ZN(
        n13419) );
  NOR2_X1 U16779 ( .A1(n13420), .A2(n13419), .ZN(n13424) );
  NOR2_X1 U16780 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  XOR2_X1 U16781 ( .A(n13424), .B(n13423), .Z(n13429) );
  AOI21_X1 U16782 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21246), .A(
        n13425), .ZN(n13427) );
  NAND2_X1 U16783 ( .A1(n14311), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13426) );
  OAI211_X1 U16784 ( .C1(n13429), .C2(n13428), .A(n13427), .B(n13426), .ZN(
        n13430) );
  OAI21_X1 U16785 ( .B1(n14331), .B2(n13431), .A(n13430), .ZN(n13433) );
  INV_X1 U16786 ( .A(n14839), .ZN(n14325) );
  NAND2_X1 U16787 ( .A1(n14839), .A2(n13435), .ZN(n13436) );
  NAND2_X1 U16788 ( .A1(n13437), .A2(n13436), .ZN(P1_U2810) );
  NOR2_X1 U16789 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13439) );
  NOR4_X1 U16790 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13438) );
  NAND4_X1 U16791 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13439), .A4(n13438), .ZN(n13452) );
  NOR2_X1 U16792 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21449) );
  NOR3_X1 U16793 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(
        P1_ADDRESS_REG_2__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13442) );
  NOR4_X1 U16794 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13441) );
  NOR4_X1 U16795 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n13440) );
  AND4_X1 U16796 ( .A1(n21449), .A2(n13442), .A3(n13441), .A4(n13440), .ZN(
        n13448) );
  NOR4_X1 U16797 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13446) );
  NOR4_X1 U16798 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13445) );
  NOR4_X1 U16799 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13444) );
  NOR4_X1 U16800 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13443) );
  AND4_X1 U16801 ( .A1(n13446), .A2(n13445), .A3(n13444), .A4(n13443), .ZN(
        n13447) );
  NAND2_X1 U16802 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  INV_X1 U16803 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n13521) );
  NOR3_X1 U16804 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n13521), .ZN(n13451) );
  NOR4_X1 U16805 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13450) );
  NAND4_X1 U16806 ( .A1(n14869), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13451), .A4(
        n13450), .ZN(U214) );
  NOR2_X1 U16807 ( .A1(n16533), .A2(n13452), .ZN(n17164) );
  NAND2_X1 U16808 ( .A1(n17164), .A2(U214), .ZN(U212) );
  AOI211_X1 U16809 ( .C1(n13456), .C2(n19660), .A(n13453), .B(n19661), .ZN(
        n13469) );
  AND2_X1 U16810 ( .A1(n16233), .A2(n13454), .ZN(n13455) );
  OR2_X1 U16811 ( .A1(n13455), .A2(n9753), .ZN(n16223) );
  OAI22_X1 U16812 ( .A1(n19659), .A2(n13456), .B1(n17133), .B2(n16223), .ZN(
        n13468) );
  XOR2_X1 U16813 ( .A(n15997), .B(n13457), .Z(n15728) );
  INV_X1 U16814 ( .A(n15728), .ZN(n16006) );
  OAI22_X1 U16815 ( .A1(n16006), .A2(n19648), .B1(n11827), .B2(n16032), .ZN(
        n13467) );
  INV_X1 U16816 ( .A(n13458), .ZN(n13462) );
  AOI21_X1 U16817 ( .B1(n12637), .B2(n13460), .A(n13459), .ZN(n13461) );
  AOI21_X1 U16818 ( .B1(n13462), .B2(n12637), .A(n13461), .ZN(n16225) );
  INV_X1 U16819 ( .A(n16225), .ZN(n13465) );
  XNOR2_X1 U16820 ( .A(n13463), .B(n13464), .ZN(n16227) );
  OAI22_X1 U16821 ( .A1(n13465), .A2(n19668), .B1(n16227), .B2(n19653), .ZN(
        n13466) );
  INV_X1 U16822 ( .A(n16134), .ZN(n13473) );
  INV_X1 U16823 ( .A(n13470), .ZN(n13472) );
  INV_X1 U16824 ( .A(n15657), .ZN(n13471) );
  NAND2_X1 U16825 ( .A1(n15733), .A2(n13471), .ZN(n15658) );
  AOI21_X1 U16826 ( .B1(n13473), .B2(n13472), .A(n15658), .ZN(n13485) );
  OAI21_X1 U16827 ( .B1(n19546), .B2(n16131), .A(n16032), .ZN(n13474) );
  AOI21_X1 U16828 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19548), .A(
        n13474), .ZN(n13475) );
  OAI21_X1 U16829 ( .B1(n12360), .B2(n19529), .A(n13475), .ZN(n13484) );
  OAI22_X1 U16830 ( .A1(n15772), .A2(n16134), .B1(n13476), .B2(n19549), .ZN(
        n13483) );
  AND2_X1 U16831 ( .A1(n14046), .A2(n13477), .ZN(n13478) );
  NOR2_X1 U16832 ( .A1(n15655), .A2(n13478), .ZN(n16130) );
  INV_X1 U16833 ( .A(n16130), .ZN(n16391) );
  NAND2_X1 U16834 ( .A1(n13893), .A2(n13491), .ZN(n14087) );
  OR2_X1 U16835 ( .A1(n14087), .A2(n13986), .ZN(n13480) );
  NOR2_X1 U16836 ( .A1(n14087), .A2(n13479), .ZN(n14085) );
  AOI21_X1 U16837 ( .B1(n13481), .B2(n13480), .A(n14085), .ZN(n16388) );
  INV_X1 U16838 ( .A(n16388), .ZN(n14153) );
  OAI22_X1 U16839 ( .A1(n16391), .A2(n19555), .B1(n14153), .B2(n19551), .ZN(
        n13482) );
  OR4_X1 U16840 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        P2_U2842) );
  INV_X1 U16841 ( .A(n19517), .ZN(n13486) );
  AOI211_X1 U16842 ( .C1(n16154), .C2(n13487), .A(n13486), .B(n15784), .ZN(
        n13500) );
  OAI21_X1 U16843 ( .B1(n19546), .B2(n13488), .A(n16032), .ZN(n13489) );
  AOI21_X1 U16844 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19548), .A(
        n13489), .ZN(n13490) );
  OAI21_X1 U16845 ( .B1(n12356), .B2(n19529), .A(n13490), .ZN(n13499) );
  OAI21_X1 U16846 ( .B1(n13893), .B2(n13491), .A(n14087), .ZN(n16412) );
  OAI22_X1 U16847 ( .A1(n16412), .A2(n19551), .B1(n13492), .B2(n19549), .ZN(
        n13498) );
  INV_X1 U16848 ( .A(n16154), .ZN(n13496) );
  OR2_X1 U16849 ( .A1(n13908), .A2(n13494), .ZN(n13495) );
  NAND2_X1 U16850 ( .A1(n13493), .A2(n13495), .ZN(n16418) );
  OAI22_X1 U16851 ( .A1(n15772), .A2(n13496), .B1(n19555), .B2(n16418), .ZN(
        n13497) );
  OR4_X1 U16852 ( .A1(n13500), .A2(n13499), .A3(n13498), .A4(n13497), .ZN(
        P2_U2844) );
  MUX2_X1 U16853 ( .A(n17147), .B(P2_STATEBS16_REG_SCAN_IN), .S(n17153), .Z(
        n13501) );
  AOI21_X1 U16854 ( .B1(n13501), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U16855 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20327) );
  INV_X1 U16856 ( .A(n20327), .ZN(n13502) );
  AND2_X1 U16857 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13502), .ZN(n17151) );
  NOR2_X1 U16858 ( .A1(n13503), .A2(n17151), .ZN(P2_U3178) );
  AOI22_X1 U16859 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n13506) );
  INV_X1 U16860 ( .A(HOLD), .ZN(n21254) );
  NOR2_X1 U16861 ( .A1(n21254), .A2(n13525), .ZN(n13505) );
  INV_X1 U16862 ( .A(n13787), .ZN(n14100) );
  INV_X1 U16863 ( .A(n21293), .ZN(n17126) );
  NAND2_X1 U16864 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n17126), .ZN(n13504) );
  OAI211_X1 U16865 ( .C1(n13506), .C2(n13505), .A(n14100), .B(n13504), .ZN(
        P1_U3195) );
  INV_X1 U16866 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20370) );
  INV_X1 U16867 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n13507) );
  OR2_X1 U16868 ( .A1(n14465), .A2(n13507), .ZN(n13508) );
  OAI21_X1 U16869 ( .B1(n21265), .B2(n20370), .A(n13508), .ZN(P1_U3458) );
  INV_X1 U16870 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21287) );
  INV_X1 U16871 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n13509) );
  OR2_X1 U16872 ( .A1(n14465), .A2(n13509), .ZN(n13510) );
  OAI21_X1 U16873 ( .B1(n21265), .B2(n21287), .A(n13510), .ZN(P1_U3459) );
  INV_X1 U16874 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21289) );
  INV_X1 U16875 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n13511) );
  OR2_X1 U16876 ( .A1(n14465), .A2(n13511), .ZN(n13512) );
  OAI21_X1 U16877 ( .B1(n21265), .B2(n21289), .A(n13512), .ZN(P1_U3461) );
  INV_X1 U16878 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20367) );
  INV_X1 U16879 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n13513) );
  OR2_X1 U16880 ( .A1(n14465), .A2(n13513), .ZN(n13514) );
  OAI21_X1 U16881 ( .B1(n21265), .B2(n20367), .A(n13514), .ZN(P1_U3460) );
  NOR2_X1 U16882 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20353) );
  OAI21_X1 U16883 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n20353), .A(n21265), .ZN(
        n13515) );
  OAI21_X1 U16884 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21265), .A(n13515), 
        .ZN(P1_U2804) );
  INV_X1 U16885 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21302) );
  INV_X1 U16886 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n13518) );
  AOI21_X1 U16887 ( .B1(n13518), .B2(n13525), .A(n21254), .ZN(n13516) );
  AOI211_X1 U16888 ( .C1(n21251), .C2(NA), .A(n21302), .B(n13516), .ZN(n13517)
         );
  AOI21_X1 U16889 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n17126), .A(n21251), 
        .ZN(n21256) );
  OAI22_X1 U16890 ( .A1(n13517), .A2(n13559), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21256), .ZN(P1_U3194) );
  INV_X1 U16891 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n13520) );
  OAI21_X1 U16892 ( .B1(n13518), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n13519) );
  OAI21_X1 U16893 ( .B1(n13559), .B2(n13520), .A(n21271), .ZN(P1_U2802) );
  OR2_X1 U16894 ( .A1(n13521), .A2(n13559), .ZN(n13522) );
  OAI21_X1 U16895 ( .B1(n21265), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13522), 
        .ZN(P1_U3483) );
  INV_X1 U16896 ( .A(n15434), .ZN(n13523) );
  INV_X1 U16897 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19493) );
  NAND2_X1 U16898 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20145), .ZN(n17146) );
  OAI22_X1 U16899 ( .A1(n13523), .A2(n19493), .B1(n20297), .B2(n17146), .ZN(
        P2_U2816) );
  NOR2_X1 U16900 ( .A1(n12028), .A2(n17160), .ZN(n13678) );
  NAND2_X1 U16901 ( .A1(n13678), .A2(n16591), .ZN(n19556) );
  INV_X1 U16902 ( .A(n19556), .ZN(n15781) );
  INV_X1 U16903 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13524) );
  OR2_X1 U16904 ( .A1(n20313), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13529) );
  OAI211_X1 U16905 ( .C1(n15781), .C2(n13524), .A(n13531), .B(n13529), .ZN(
        P2_U2814) );
  NAND2_X1 U16906 ( .A1(n13559), .A2(n13525), .ZN(n13561) );
  INV_X1 U16907 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21258) );
  INV_X1 U16908 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20432) );
  INV_X1 U16909 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21343) );
  OAI222_X1 U16910 ( .A1(n13561), .A2(n21258), .B1(n21268), .B2(n20432), .C1(
        n13559), .C2(n21343), .ZN(P1_U3198) );
  INV_X1 U16911 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13527) );
  INV_X1 U16912 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13526) );
  OAI222_X1 U16913 ( .A1(n13527), .A2(n21268), .B1(n13526), .B2(n13559), .C1(
        n13561), .C2(n20400), .ZN(P1_U3200) );
  INV_X1 U16914 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14946) );
  INV_X1 U16915 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13528) );
  OAI222_X1 U16916 ( .A1(n21268), .A2(n14946), .B1(n13528), .B2(n13559), .C1(
        n13544), .C2(n13561), .ZN(P1_U3224) );
  INV_X1 U16917 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n13530) );
  NAND4_X1 U16918 ( .A1(n13531), .A2(n19556), .A3(n13530), .A4(n13529), .ZN(
        n13532) );
  OAI21_X1 U16919 ( .B1(n15434), .B2(n15430), .A(n13532), .ZN(n13533) );
  INV_X1 U16920 ( .A(n13533), .ZN(P2_U3612) );
  INV_X1 U16921 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21262) );
  INV_X1 U16922 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13534) );
  INV_X1 U16923 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15059) );
  OAI222_X1 U16924 ( .A1(n13561), .A2(n21262), .B1(n14465), .B2(n13534), .C1(
        n15059), .C2(n21268), .ZN(P1_U3213) );
  INV_X1 U16925 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15125) );
  INV_X1 U16926 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n13535) );
  INV_X1 U16927 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15138) );
  OAI222_X1 U16928 ( .A1(n13561), .A2(n15125), .B1(n14465), .B2(n13535), .C1(
        n15138), .C2(n21268), .ZN(P1_U3206) );
  INV_X1 U16929 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13536) );
  INV_X1 U16930 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15031) );
  OAI222_X1 U16931 ( .A1(n13561), .A2(n15023), .B1(n13536), .B2(n13559), .C1(
        n15031), .C2(n21268), .ZN(P1_U3215) );
  AOI21_X1 U16932 ( .B1(n17147), .B2(n15430), .A(n13537), .ZN(n13538) );
  NAND3_X1 U16933 ( .A1(n16597), .A2(n16591), .A3(n13538), .ZN(n16598) );
  AND2_X1 U16934 ( .A1(n16598), .A2(n16626), .ZN(n20345) );
  OAI21_X1 U16935 ( .B1(n16600), .B2(n20345), .A(n13539), .ZN(P2_U2819) );
  INV_X1 U16936 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21404) );
  INV_X1 U16937 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13540) );
  INV_X1 U16938 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14983) );
  OAI222_X1 U16939 ( .A1(n13561), .A2(n21404), .B1(n14465), .B2(n13540), .C1(
        n14983), .C2(n21268), .ZN(P1_U3220) );
  INV_X1 U16940 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n13541) );
  INV_X1 U16941 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14995) );
  OAI222_X1 U16942 ( .A1(n13561), .A2(n14983), .B1(n13541), .B2(n13559), .C1(
        n14995), .C2(n21268), .ZN(P1_U3219) );
  INV_X1 U16943 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20386) );
  INV_X1 U16944 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n13542) );
  OAI222_X1 U16945 ( .A1(n13561), .A2(n20381), .B1(n21268), .B2(n20386), .C1(
        n13559), .C2(n13542), .ZN(P1_U3202) );
  INV_X1 U16946 ( .A(n13561), .ZN(n21266) );
  AOI22_X1 U16947 ( .A1(n21266), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21265), .ZN(n13543) );
  OAI21_X1 U16948 ( .B1(n13544), .B2(n21268), .A(n13543), .ZN(P1_U3225) );
  INV_X1 U16949 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13546) );
  AOI22_X1 U16950 ( .A1(n21266), .A2(P1_REIP_REG_31__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21265), .ZN(n13545) );
  OAI21_X1 U16951 ( .B1(n13546), .B2(n21268), .A(n13545), .ZN(P1_U3226) );
  INV_X1 U16952 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13547) );
  INV_X1 U16953 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15083) );
  OAI222_X1 U16954 ( .A1(n21268), .A2(n15092), .B1(n14465), .B2(n13547), .C1(
        n15083), .C2(n13561), .ZN(P1_U3210) );
  INV_X1 U16955 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n13548) );
  OAI222_X1 U16956 ( .A1(n21268), .A2(n20381), .B1(n13561), .B2(n21260), .C1(
        n13548), .C2(n13559), .ZN(P1_U3203) );
  INV_X1 U16957 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14706) );
  INV_X1 U16958 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13549) );
  OAI222_X1 U16959 ( .A1(n21268), .A2(n14706), .B1(n14465), .B2(n13549), .C1(
        n15105), .C2(n13561), .ZN(P1_U3208) );
  INV_X1 U16960 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n13550) );
  INV_X1 U16961 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15070) );
  OAI222_X1 U16962 ( .A1(n21268), .A2(n15083), .B1(n14465), .B2(n13550), .C1(
        n15070), .C2(n13561), .ZN(P1_U3211) );
  INV_X1 U16963 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21284) );
  INV_X1 U16964 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13551) );
  OAI222_X1 U16965 ( .A1(n21268), .A2(n21284), .B1(n13561), .B2(n20432), .C1(
        n13559), .C2(n13551), .ZN(P1_U3197) );
  INV_X1 U16966 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21390) );
  INV_X1 U16967 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15014) );
  OAI222_X1 U16968 ( .A1(n21268), .A2(n15023), .B1(n14465), .B2(n21390), .C1(
        n15014), .C2(n13561), .ZN(P1_U3216) );
  INV_X1 U16969 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14235) );
  INV_X1 U16970 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13552) );
  OAI222_X1 U16971 ( .A1(n21268), .A2(n14235), .B1(n13552), .B2(n13559), .C1(
        n15138), .C2(n13561), .ZN(P1_U3205) );
  INV_X1 U16972 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13553) );
  INV_X1 U16973 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14967) );
  OAI222_X1 U16974 ( .A1(n21268), .A2(n21404), .B1(n14465), .B2(n13553), .C1(
        n14967), .C2(n13561), .ZN(P1_U3221) );
  INV_X1 U16975 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n13554) );
  INV_X1 U16976 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21269) );
  OAI222_X1 U16977 ( .A1(n21268), .A2(n14967), .B1(n13559), .B2(n13554), .C1(
        n21269), .C2(n13561), .ZN(P1_U3222) );
  INV_X1 U16978 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n13555) );
  OAI222_X1 U16979 ( .A1(n21268), .A2(n15125), .B1(n14465), .B2(n13555), .C1(
        n14706), .C2(n13561), .ZN(P1_U3207) );
  INV_X1 U16980 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13556) );
  OAI222_X1 U16981 ( .A1(n21268), .A2(n15014), .B1(n13559), .B2(n13556), .C1(
        n21264), .C2(n13561), .ZN(P1_U3217) );
  INV_X1 U16982 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13557) );
  OAI222_X1 U16983 ( .A1(n21268), .A2(n15070), .B1(n13559), .B2(n13557), .C1(
        n15059), .C2(n13561), .ZN(P1_U3212) );
  INV_X1 U16984 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13558) );
  OAI222_X1 U16985 ( .A1(n13561), .A2(n20386), .B1(n21268), .B2(n20400), .C1(
        n13559), .C2(n13558), .ZN(P1_U3201) );
  INV_X1 U16986 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13560) );
  OAI222_X1 U16987 ( .A1(n13561), .A2(n15092), .B1(n14465), .B2(n13560), .C1(
        n15105), .C2(n21268), .ZN(P1_U3209) );
  INV_X1 U16988 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13695) );
  NAND3_X1 U16989 ( .A1(n13563), .A2(n17147), .A3(n15806), .ZN(n13593) );
  INV_X1 U16990 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18891) );
  NAND2_X1 U16991 ( .A1(n13618), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13562) );
  OAI21_X1 U16992 ( .B1(n13618), .B2(n18891), .A(n13562), .ZN(n19576) );
  NAND2_X1 U16993 ( .A1(n19628), .A2(n19576), .ZN(n13600) );
  OAI21_X1 U16994 ( .B1(n12004), .B2(n17147), .A(n13563), .ZN(n13574) );
  NAND2_X1 U16995 ( .A1(n13574), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13564) );
  OAI211_X1 U16996 ( .C1(n13679), .C2(n13695), .A(n13600), .B(n13564), .ZN(
        P2_U2956) );
  INV_X1 U16997 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13710) );
  INV_X1 U16998 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18902) );
  NAND2_X1 U16999 ( .A1(n13618), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13565) );
  OAI21_X1 U17000 ( .B1(n13618), .B2(n18902), .A(n13565), .ZN(n16557) );
  NAND2_X1 U17001 ( .A1(n19628), .A2(n16557), .ZN(n13607) );
  INV_X1 U17002 ( .A(n13574), .ZN(n13596) );
  NAND2_X1 U17003 ( .A1(n13574), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13566) );
  OAI211_X1 U17004 ( .C1(n13679), .C2(n13710), .A(n13607), .B(n13566), .ZN(
        P2_U2958) );
  INV_X1 U17005 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13689) );
  INV_X1 U17006 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18871) );
  NAND2_X1 U17007 ( .A1(n13618), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13567) );
  OAI21_X1 U17008 ( .B1(n13618), .B2(n18871), .A(n13567), .ZN(n16525) );
  NAND2_X1 U17009 ( .A1(n19628), .A2(n16525), .ZN(n13572) );
  NAND2_X1 U17010 ( .A1(n13574), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13568) );
  OAI211_X1 U17011 ( .C1(n13679), .C2(n13689), .A(n13572), .B(n13568), .ZN(
        P2_U2952) );
  INV_X1 U17012 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19607) );
  INV_X1 U17013 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18222) );
  NAND2_X1 U17014 ( .A1(n13618), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13569) );
  OAI21_X1 U17015 ( .B1(n13618), .B2(n18222), .A(n13569), .ZN(n15934) );
  NAND2_X1 U17016 ( .A1(n19628), .A2(n15934), .ZN(n13598) );
  NAND2_X1 U17017 ( .A1(n19626), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13570) );
  OAI211_X1 U17018 ( .C1(n13679), .C2(n19607), .A(n13598), .B(n13570), .ZN(
        P2_U2975) );
  NAND2_X1 U17019 ( .A1(n19626), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13571) );
  OAI211_X1 U17020 ( .C1(n13679), .C2(n12048), .A(n13572), .B(n13571), .ZN(
        P2_U2967) );
  INV_X1 U17021 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19599) );
  INV_X1 U17022 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18231) );
  NAND2_X1 U17023 ( .A1(n13618), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13573) );
  OAI21_X1 U17024 ( .B1(n13618), .B2(n18231), .A(n13573), .ZN(n15904) );
  NAND2_X1 U17025 ( .A1(n19628), .A2(n15904), .ZN(n13602) );
  NAND2_X1 U17026 ( .A1(n13574), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13575) );
  OAI211_X1 U17027 ( .C1(n13679), .C2(n19599), .A(n13602), .B(n13575), .ZN(
        P2_U2979) );
  INV_X1 U17028 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19603) );
  INV_X1 U17029 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18225) );
  NAND2_X1 U17030 ( .A1(n13618), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13576) );
  OAI21_X1 U17031 ( .B1(n13618), .B2(n18225), .A(n13576), .ZN(n15919) );
  NAND2_X1 U17032 ( .A1(n19628), .A2(n15919), .ZN(n13606) );
  NAND2_X1 U17033 ( .A1(n19626), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13577) );
  OAI211_X1 U17034 ( .C1(n13679), .C2(n19603), .A(n13606), .B(n13577), .ZN(
        P2_U2977) );
  AOI22_X1 U17035 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n19630), .B1(n13574), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13580) );
  INV_X1 U17036 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13579) );
  NAND2_X1 U17037 ( .A1(n13618), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13578) );
  OAI21_X1 U17038 ( .B1(n13618), .B2(n13579), .A(n13578), .ZN(n15927) );
  NAND2_X1 U17039 ( .A1(n19628), .A2(n15927), .ZN(n13614) );
  NAND2_X1 U17040 ( .A1(n13580), .A2(n13614), .ZN(P2_U2961) );
  AOI22_X1 U17041 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(n19630), .B1(n13574), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13583) );
  INV_X1 U17042 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n13582) );
  NAND2_X1 U17043 ( .A1(n13618), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13581) );
  OAI21_X1 U17044 ( .B1(n13618), .B2(n13582), .A(n13581), .ZN(n16552) );
  NAND2_X1 U17045 ( .A1(n19628), .A2(n16552), .ZN(n13616) );
  NAND2_X1 U17046 ( .A1(n13583), .A2(n13616), .ZN(P2_U2957) );
  AOI22_X1 U17047 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(n19630), .B1(n13574), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13586) );
  INV_X1 U17048 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n13585) );
  NAND2_X1 U17049 ( .A1(n13618), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13584) );
  OAI21_X1 U17050 ( .B1(n13618), .B2(n13585), .A(n13584), .ZN(n16545) );
  NAND2_X1 U17051 ( .A1(n19628), .A2(n16545), .ZN(n13628) );
  NAND2_X1 U17052 ( .A1(n13586), .A2(n13628), .ZN(P2_U2955) );
  AOI22_X1 U17053 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(n19630), .B1(n13574), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13589) );
  INV_X1 U17054 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U17055 ( .A1(n13618), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13587) );
  OAI21_X1 U17056 ( .B1(n13618), .B2(n13588), .A(n13587), .ZN(n16561) );
  NAND2_X1 U17057 ( .A1(n19628), .A2(n16561), .ZN(n13630) );
  NAND2_X1 U17058 ( .A1(n13589), .A2(n13630), .ZN(P2_U2959) );
  AOI22_X1 U17059 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n19630), .B1(n13574), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13591) );
  INV_X1 U17060 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U17061 ( .A1(n13618), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13590) );
  OAI21_X1 U17062 ( .B1(n13618), .B2(n13926), .A(n13590), .ZN(n16538) );
  NAND2_X1 U17063 ( .A1(n19628), .A2(n16538), .ZN(n13622) );
  NAND2_X1 U17064 ( .A1(n13591), .A2(n13622), .ZN(P2_U2953) );
  INV_X1 U17065 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13595) );
  INV_X1 U17066 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13594) );
  INV_X1 U17067 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13978) );
  NOR2_X1 U17068 ( .A1(n16533), .A2(n13978), .ZN(n13592) );
  AOI21_X1 U17069 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n16533), .A(n13592), .ZN(
        n14149) );
  OAI222_X1 U17070 ( .A1(n13679), .A2(n13595), .B1(n13594), .B2(n13596), .C1(
        n13593), .C2(n14149), .ZN(P2_U2982) );
  INV_X1 U17071 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13702) );
  NAND2_X1 U17072 ( .A1(n19626), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13597) );
  OAI211_X1 U17073 ( .C1(n13679), .C2(n13702), .A(n13598), .B(n13597), .ZN(
        P2_U2960) );
  INV_X1 U17074 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19615) );
  NAND2_X1 U17075 ( .A1(n19626), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n13599) );
  OAI211_X1 U17076 ( .C1(n13679), .C2(n19615), .A(n13600), .B(n13599), .ZN(
        P2_U2971) );
  INV_X1 U17077 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21386) );
  NAND2_X1 U17078 ( .A1(n19626), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13601) );
  OAI211_X1 U17079 ( .C1(n13679), .C2(n21386), .A(n13602), .B(n13601), .ZN(
        P2_U2964) );
  INV_X1 U17080 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13685) );
  INV_X1 U17081 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18881) );
  NAND2_X1 U17082 ( .A1(n13618), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13603) );
  OAI21_X1 U17083 ( .B1(n13618), .B2(n18881), .A(n13603), .ZN(n16541) );
  NAND2_X1 U17084 ( .A1(n19628), .A2(n16541), .ZN(n13612) );
  NAND2_X1 U17085 ( .A1(n19626), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13604) );
  OAI211_X1 U17086 ( .C1(n13679), .C2(n13685), .A(n13612), .B(n13604), .ZN(
        P2_U2954) );
  INV_X1 U17087 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U17088 ( .A1(n19626), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13605) );
  OAI211_X1 U17089 ( .C1(n13679), .C2(n13706), .A(n13606), .B(n13605), .ZN(
        P2_U2962) );
  AOI22_X1 U17090 ( .A1(P2_EAX_REG_6__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U17091 ( .A1(n13608), .A2(n13607), .ZN(P2_U2973) );
  AOI22_X1 U17092 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n19630), .B1(n19626), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13611) );
  INV_X1 U17093 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n13610) );
  NAND2_X1 U17094 ( .A1(n13618), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13609) );
  OAI21_X1 U17095 ( .B1(n13618), .B2(n13610), .A(n13609), .ZN(n15897) );
  NAND2_X1 U17096 ( .A1(n19628), .A2(n15897), .ZN(n13626) );
  NAND2_X1 U17097 ( .A1(n13611), .A2(n13626), .ZN(P2_U2980) );
  AOI22_X1 U17098 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U17099 ( .A1(n13613), .A2(n13612), .ZN(P2_U2969) );
  AOI22_X1 U17100 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U17101 ( .A1(n13615), .A2(n13614), .ZN(P2_U2976) );
  AOI22_X1 U17102 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U17103 ( .A1(n13617), .A2(n13616), .ZN(P2_U2972) );
  AOI22_X1 U17104 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n19630), .B1(n19626), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13621) );
  INV_X1 U17105 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13620) );
  NAND2_X1 U17106 ( .A1(n13618), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13619) );
  OAI21_X1 U17107 ( .B1(n13618), .B2(n13620), .A(n13619), .ZN(n15911) );
  NAND2_X1 U17108 ( .A1(n19628), .A2(n15911), .ZN(n13624) );
  NAND2_X1 U17109 ( .A1(n13621), .A2(n13624), .ZN(P2_U2963) );
  AOI22_X1 U17110 ( .A1(P2_EAX_REG_1__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U17111 ( .A1(n13623), .A2(n13622), .ZN(P2_U2968) );
  AOI22_X1 U17112 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n19630), .B1(n19626), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U17113 ( .A1(n13625), .A2(n13624), .ZN(P2_U2978) );
  AOI22_X1 U17114 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n19630), .B1(n19626), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U17115 ( .A1(n13627), .A2(n13626), .ZN(P2_U2965) );
  AOI22_X1 U17116 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U17117 ( .A1(n13629), .A2(n13628), .ZN(P2_U2970) );
  AOI22_X1 U17118 ( .A1(P2_EAX_REG_7__SCAN_IN), .A2(n19630), .B1(n19626), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13631) );
  NAND2_X1 U17119 ( .A1(n13631), .A2(n13630), .ZN(P2_U2974) );
  INV_X1 U17120 ( .A(n13681), .ZN(n13634) );
  NOR2_X1 U17121 ( .A1(n12028), .A2(n13632), .ZN(n13633) );
  NAND2_X1 U17122 ( .A1(n13634), .A2(n13633), .ZN(n13638) );
  INV_X1 U17123 ( .A(n16592), .ZN(n13635) );
  INV_X1 U17124 ( .A(n13859), .ZN(n16593) );
  NAND2_X1 U17125 ( .A1(n13635), .A2(n16593), .ZN(n13648) );
  NAND4_X1 U17126 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13648), .ZN(
        n16610) );
  NAND2_X1 U17127 ( .A1(n16610), .A2(n16626), .ZN(n13640) );
  AOI22_X1 U17128 ( .A1(n17151), .A2(P2_FLUSH_REG_SCAN_IN), .B1(n17153), .B2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13639) );
  INV_X1 U17129 ( .A(n20301), .ZN(n13643) );
  NOR3_X1 U17130 ( .A1(n12028), .A2(n13641), .A3(n15806), .ZN(n16602) );
  NAND3_X1 U17131 ( .A1(n13643), .A2(n16602), .A3(n20305), .ZN(n13642) );
  OAI21_X1 U17132 ( .B1(n13643), .B2(n16605), .A(n13642), .ZN(P2_U3595) );
  NAND2_X1 U17133 ( .A1(n15806), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13645) );
  NAND4_X1 U17134 ( .A1(n13646), .A2(n13645), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20318), .ZN(n13647) );
  NAND2_X1 U17135 ( .A1(n16571), .A2(n12311), .ZN(n13871) );
  NAND2_X1 U17136 ( .A1(n13648), .A2(n13871), .ZN(n13649) );
  NAND2_X1 U17137 ( .A1(n19575), .A2(n16566), .ZN(n19571) );
  MUX2_X1 U17138 ( .A(n11800), .B(n15779), .S(n19575), .Z(n13650) );
  OAI21_X1 U17139 ( .B1(n20330), .B2(n19571), .A(n13650), .ZN(P2_U2887) );
  OR2_X1 U17140 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21184), .ZN(n20352) );
  NAND2_X1 U17141 ( .A1(n9667), .A2(n20352), .ZN(n13655) );
  NOR2_X1 U17142 ( .A1(n13655), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13654)
         );
  INV_X1 U17143 ( .A(n13652), .ZN(n13651) );
  AOI21_X1 U17144 ( .B1(n9667), .B2(n21294), .A(n13651), .ZN(n13653) );
  OAI22_X1 U17145 ( .A1(n13654), .A2(n13653), .B1(n13652), .B2(n21294), .ZN(
        P1_U3487) );
  AOI21_X1 U17146 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(n21294), .A(n13655), 
        .ZN(n13656) );
  INV_X1 U17147 ( .A(n13656), .ZN(P1_U2801) );
  INV_X1 U17148 ( .A(n14173), .ZN(n13659) );
  OAI22_X1 U17149 ( .A1(n13659), .A2(n14770), .B1(n13658), .B2(n13657), .ZN(
        n20349) );
  NOR3_X1 U17150 ( .A1(n10302), .A2(n14770), .A3(n13787), .ZN(n13660) );
  NOR2_X1 U17151 ( .A1(n13660), .A2(n17126), .ZN(n21297) );
  NOR2_X1 U17152 ( .A1(n20349), .A2(n21297), .ZN(n17076) );
  NOR2_X1 U17153 ( .A1(n17076), .A2(n20348), .ZN(n20355) );
  INV_X1 U17154 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13673) );
  INV_X1 U17155 ( .A(n13721), .ZN(n14778) );
  NAND2_X1 U17156 ( .A1(n14778), .A2(n13661), .ZN(n13663) );
  AND3_X1 U17157 ( .A1(n13663), .A2(n13662), .A3(n13274), .ZN(n14120) );
  NOR2_X1 U17158 ( .A1(n10441), .A2(n13946), .ZN(n14108) );
  NAND2_X1 U17159 ( .A1(n13718), .A2(n14770), .ZN(n15368) );
  AND2_X1 U17160 ( .A1(n17079), .A2(n15368), .ZN(n14112) );
  INV_X1 U17161 ( .A(n13664), .ZN(n13665) );
  NAND2_X1 U17162 ( .A1(n14112), .A2(n13665), .ZN(n13666) );
  MUX2_X1 U17163 ( .A(n15367), .B(n13666), .S(n14173), .Z(n13669) );
  INV_X1 U17164 ( .A(n13719), .ZN(n13667) );
  NOR2_X1 U17165 ( .A1(n13714), .A2(n13667), .ZN(n13668) );
  OR2_X1 U17166 ( .A1(n13669), .A2(n13668), .ZN(n13670) );
  NAND2_X1 U17167 ( .A1(n13670), .A2(n20649), .ZN(n17078) );
  INV_X1 U17168 ( .A(n17078), .ZN(n13671) );
  NAND2_X1 U17169 ( .A1(n20355), .A2(n13671), .ZN(n13672) );
  OAI21_X1 U17170 ( .B1(n20355), .B2(n13673), .A(n13672), .ZN(P1_U3484) );
  MUX2_X1 U17171 ( .A(n12343), .B(n16486), .S(n19575), .Z(n13677) );
  OAI21_X1 U17172 ( .B1(n19782), .B2(n19571), .A(n13677), .ZN(P2_U2886) );
  INV_X1 U17173 ( .A(n13678), .ZN(n13680) );
  INV_X1 U17174 ( .A(n15425), .ZN(n13683) );
  OR2_X1 U17175 ( .A1(n20327), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15435) );
  INV_X2 U17176 ( .A(n15435), .ZN(n19623) );
  AOI22_X1 U17177 ( .A1(n19623), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13684) );
  OAI21_X1 U17178 ( .B1(n13685), .B2(n19588), .A(n13684), .ZN(P2_U2933) );
  AOI22_X1 U17179 ( .A1(n19623), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13686) );
  OAI21_X1 U17180 ( .B1(n13687), .B2(n19588), .A(n13686), .ZN(P2_U2922) );
  AOI22_X1 U17181 ( .A1(n19623), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13688) );
  OAI21_X1 U17182 ( .B1(n13689), .B2(n19588), .A(n13688), .ZN(P2_U2935) );
  INV_X1 U17183 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13691) );
  AOI22_X1 U17184 ( .A1(n19623), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13690) );
  OAI21_X1 U17185 ( .B1(n13691), .B2(n19588), .A(n13690), .ZN(P2_U2928) );
  INV_X1 U17186 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U17187 ( .A1(n19623), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U17188 ( .B1(n13693), .B2(n19588), .A(n13692), .ZN(P2_U2934) );
  AOI22_X1 U17189 ( .A1(n19623), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13694) );
  OAI21_X1 U17190 ( .B1(n13695), .B2(n19588), .A(n13694), .ZN(P2_U2931) );
  INV_X1 U17191 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17192 ( .A1(n19623), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13696) );
  OAI21_X1 U17193 ( .B1(n13697), .B2(n19588), .A(n13696), .ZN(P2_U2930) );
  INV_X1 U17194 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U17195 ( .A1(n19623), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13698) );
  OAI21_X1 U17196 ( .B1(n13699), .B2(n19588), .A(n13698), .ZN(P2_U2924) );
  AOI22_X1 U17197 ( .A1(n19623), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13700) );
  OAI21_X1 U17198 ( .B1(n21386), .B2(n19588), .A(n13700), .ZN(P2_U2923) );
  AOI22_X1 U17199 ( .A1(n19623), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13701) );
  OAI21_X1 U17200 ( .B1(n13702), .B2(n19588), .A(n13701), .ZN(P2_U2927) );
  INV_X1 U17201 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U17202 ( .A1(n19623), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13703) );
  OAI21_X1 U17203 ( .B1(n13704), .B2(n19588), .A(n13703), .ZN(P2_U2926) );
  AOI22_X1 U17204 ( .A1(n19623), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13705) );
  OAI21_X1 U17205 ( .B1(n13706), .B2(n19588), .A(n13705), .ZN(P2_U2925) );
  INV_X1 U17206 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13708) );
  AOI22_X1 U17207 ( .A1(n19623), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13707) );
  OAI21_X1 U17208 ( .B1(n13708), .B2(n19588), .A(n13707), .ZN(P2_U2932) );
  AOI22_X1 U17209 ( .A1(n19623), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U17210 ( .B1(n13710), .B2(n19588), .A(n13709), .ZN(P2_U2929) );
  NAND2_X1 U17211 ( .A1(n17060), .A2(n13787), .ZN(n13790) );
  INV_X1 U17212 ( .A(n20649), .ZN(n14444) );
  OR2_X1 U17213 ( .A1(n13711), .A2(n14444), .ZN(n14268) );
  INV_X1 U17214 ( .A(n14268), .ZN(n13789) );
  OAI21_X1 U17215 ( .B1(n13787), .B2(n10302), .A(n13789), .ZN(n13712) );
  AOI21_X1 U17216 ( .B1(n13790), .B2(n13712), .A(n17126), .ZN(n13713) );
  MUX2_X1 U17217 ( .A(n13713), .B(n15367), .S(n14173), .Z(n13724) );
  NAND2_X1 U17218 ( .A1(n21293), .A2(n13714), .ZN(n14097) );
  OAI22_X1 U17219 ( .A1(n14173), .A2(n15368), .B1(n14097), .B2(n15394), .ZN(
        n13827) );
  AOI21_X1 U17220 ( .B1(n13715), .B2(n10437), .A(n10432), .ZN(n13716) );
  NAND2_X1 U17221 ( .A1(n10440), .A2(n13716), .ZN(n14119) );
  AND2_X1 U17222 ( .A1(n13718), .A2(n14119), .ZN(n13720) );
  NOR2_X1 U17223 ( .A1(n13720), .A2(n13719), .ZN(n14107) );
  NOR2_X1 U17224 ( .A1(n13721), .A2(n14187), .ZN(n13722) );
  OR2_X1 U17225 ( .A1(n14107), .A2(n13722), .ZN(n13723) );
  NAND2_X1 U17226 ( .A1(n17063), .A2(n13828), .ZN(n13727) );
  NOR2_X1 U17227 ( .A1(n21246), .A2(n15388), .ZN(n17131) );
  NAND2_X1 U17228 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17131), .ZN(n17132) );
  INV_X1 U17229 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20354) );
  OAI22_X1 U17230 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21041), .B1(n17132), 
        .B2(n20354), .ZN(n13725) );
  INV_X1 U17231 ( .A(n13725), .ZN(n13726) );
  INV_X1 U17232 ( .A(n21281), .ZN(n14282) );
  INV_X1 U17233 ( .A(n15394), .ZN(n13728) );
  NAND3_X1 U17234 ( .A1(n14282), .A2(n13728), .A3(n21278), .ZN(n13731) );
  INV_X1 U17235 ( .A(n21030), .ZN(n20754) );
  NOR2_X1 U17236 ( .A1(n13729), .A2(n20754), .ZN(n13730) );
  XNOR2_X1 U17237 ( .A(n13730), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20412) );
  OAI22_X1 U17238 ( .A1(n13731), .A2(n20412), .B1(n14282), .B2(n15392), .ZN(
        P1_U3468) );
  XNOR2_X1 U17239 ( .A(n13732), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19635) );
  OAI21_X1 U17240 ( .B1(n13733), .B2(n13735), .A(n13734), .ZN(n15774) );
  NAND2_X1 U17241 ( .A1(n19553), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19638) );
  OAI21_X1 U17242 ( .B1(n19648), .B2(n15774), .A(n19638), .ZN(n13737) );
  OAI21_X1 U17243 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15776), .A(
        n16262), .ZN(n19639) );
  OAI22_X1 U17244 ( .A1(n15779), .A2(n17133), .B1(n19653), .B2(n19639), .ZN(
        n13736) );
  AOI211_X1 U17245 ( .C1(n19657), .C2(n19635), .A(n13737), .B(n13736), .ZN(
        n13740) );
  INV_X1 U17246 ( .A(n16489), .ZN(n13738) );
  MUX2_X1 U17247 ( .A(n16408), .B(n13738), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13739) );
  NAND2_X1 U17248 ( .A1(n13740), .A2(n13739), .ZN(P2_U3046) );
  INV_X1 U17249 ( .A(n16525), .ZN(n13746) );
  INV_X1 U17250 ( .A(n15774), .ZN(n13743) );
  NOR2_X1 U17251 ( .A1(n20330), .A2(n15774), .ZN(n13853) );
  INV_X1 U17252 ( .A(n13853), .ZN(n13742) );
  OAI211_X1 U17253 ( .C1(n19691), .C2(n13743), .A(n13742), .B(n19582), .ZN(
        n13745) );
  AOI22_X1 U17254 ( .A1(n19578), .A2(n13743), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n16010), .ZN(n13744) );
  OAI211_X1 U17255 ( .C1(n13746), .C2(n14151), .A(n13745), .B(n13744), .ZN(
        P2_U2919) );
  NAND2_X1 U17256 ( .A1(n13748), .A2(n13749), .ZN(n13750) );
  NAND2_X1 U17257 ( .A1(n13747), .A2(n13750), .ZN(n16453) );
  AOI22_X1 U17258 ( .A1(n19577), .A2(n15934), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n16010), .ZN(n13751) );
  OAI21_X1 U17259 ( .B1(n16453), .B2(n16005), .A(n13751), .ZN(P2_U2911) );
  XNOR2_X1 U17260 ( .A(n13753), .B(n10229), .ZN(n19543) );
  INV_X1 U17261 ( .A(n19543), .ZN(n13755) );
  INV_X1 U17262 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19611) );
  INV_X1 U17263 ( .A(n16557), .ZN(n13754) );
  OAI222_X1 U17264 ( .A1(n13755), .A2(n16005), .B1(n19611), .B2(n19586), .C1(
        n14151), .C2(n13754), .ZN(P2_U2913) );
  OR2_X1 U17265 ( .A1(n13757), .A2(n13756), .ZN(n13758) );
  NAND2_X1 U17266 ( .A1(n13748), .A2(n13758), .ZN(n17138) );
  INV_X1 U17267 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19609) );
  INV_X1 U17268 ( .A(n16561), .ZN(n13759) );
  OAI222_X1 U17269 ( .A1(n17138), .A2(n16005), .B1(n19609), .B2(n19586), .C1(
        n14151), .C2(n13759), .ZN(P2_U2912) );
  OR2_X1 U17270 ( .A1(n13762), .A2(n13761), .ZN(n13763) );
  NAND2_X1 U17271 ( .A1(n13760), .A2(n13763), .ZN(n14794) );
  NAND2_X1 U17272 ( .A1(n14173), .A2(n15367), .ZN(n13766) );
  INV_X1 U17273 ( .A(n10435), .ZN(n13764) );
  NAND4_X1 U17274 ( .A1(n13764), .A2(n10445), .A3(n14444), .A4(n15378), .ZN(
        n13823) );
  OR2_X1 U17275 ( .A1(n13823), .A2(n13376), .ZN(n13765) );
  NAND2_X1 U17276 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  AND2_X1 U17277 ( .A1(n20452), .A2(n20649), .ZN(n20449) );
  XNOR2_X1 U17278 ( .A(n13768), .B(n13376), .ZN(n20561) );
  OAI222_X1 U17279 ( .A1(n14794), .A2(n14838), .B1(n13268), .B2(n20452), .C1(
        n14835), .C2(n20561), .ZN(P1_U2871) );
  INV_X1 U17280 ( .A(n13769), .ZN(n13772) );
  INV_X1 U17281 ( .A(n13770), .ZN(n13771) );
  NAND2_X1 U17282 ( .A1(n13772), .A2(n13771), .ZN(n13774) );
  INV_X1 U17283 ( .A(n20323), .ZN(n20299) );
  MUX2_X1 U17284 ( .A(n16572), .B(n13775), .S(n19570), .Z(n13776) );
  OAI21_X1 U17285 ( .B1(n20299), .B2(n19571), .A(n13776), .ZN(P2_U2885) );
  NOR2_X1 U17286 ( .A1(n14307), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13778) );
  OR2_X1 U17287 ( .A1(n13778), .A2(n13777), .ZN(n20577) );
  INV_X1 U17288 ( .A(n13779), .ZN(n13782) );
  OAI21_X1 U17289 ( .B1(n13782), .B2(n13781), .A(n13780), .ZN(n14802) );
  OAI222_X1 U17290 ( .A1(n20577), .A2(n14835), .B1(n13267), .B2(n20452), .C1(
        n14802), .C2(n14838), .ZN(P1_U2872) );
  CLKBUF_X1 U17291 ( .A(n13785), .Z(n16481) );
  MUX2_X1 U17292 ( .A(n12347), .B(n16481), .S(n19575), .Z(n13786) );
  OAI21_X1 U17293 ( .B1(n19692), .B2(n19571), .A(n13786), .ZN(P2_U2884) );
  INV_X1 U17294 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13794) );
  AND2_X1 U17295 ( .A1(n14101), .A2(n13787), .ZN(n13788) );
  NAND2_X1 U17296 ( .A1(n13789), .A2(n13788), .ZN(n17058) );
  NAND2_X1 U17297 ( .A1(n20453), .A2(n10476), .ZN(n14036) );
  NAND2_X1 U17298 ( .A1(n20351), .A2(n17131), .ZN(n20455) );
  INV_X2 U17299 ( .A(n20455), .ZN(n21292) );
  NOR2_X4 U17300 ( .A1(n20453), .A2(n21292), .ZN(n20471) );
  AOI22_X1 U17301 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13793) );
  OAI21_X1 U17302 ( .B1(n13794), .B2(n14036), .A(n13793), .ZN(P1_U2910) );
  AOI22_X1 U17303 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13795) );
  OAI21_X1 U17304 ( .B1(n11232), .B2(n14036), .A(n13795), .ZN(P1_U2907) );
  AOI22_X1 U17305 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13796) );
  OAI21_X1 U17306 ( .B1(n11038), .B2(n14036), .A(n13796), .ZN(P1_U2911) );
  INV_X1 U17307 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17308 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13797) );
  OAI21_X1 U17309 ( .B1(n13798), .B2(n14036), .A(n13797), .ZN(P1_U2908) );
  NOR2_X1 U17310 ( .A1(n18555), .A2(n10308), .ZN(n14002) );
  NAND2_X1 U17311 ( .A1(n13800), .A2(n13799), .ZN(n13802) );
  AOI221_X1 U17312 ( .B1(n13803), .B2(n17249), .C1(n13802), .C2(n17249), .A(
        n13801), .ZN(n16880) );
  NAND3_X1 U17313 ( .A1(n13807), .A2(n19296), .A3(n18899), .ZN(n13804) );
  OAI21_X1 U17314 ( .B1(n13805), .B2(n19299), .A(n13804), .ZN(n13806) );
  INV_X1 U17315 ( .A(n13806), .ZN(n13813) );
  INV_X1 U17316 ( .A(n19294), .ZN(n17248) );
  INV_X1 U17317 ( .A(n13807), .ZN(n13808) );
  OAI21_X1 U17318 ( .B1(n13809), .B2(n19471), .A(n13808), .ZN(n13810) );
  OAI21_X1 U17319 ( .B1(n19470), .B2(n13810), .A(n19466), .ZN(n17255) );
  OR3_X1 U17320 ( .A1(n13811), .A2(n17248), .A3(n17255), .ZN(n13812) );
  NAND3_X1 U17321 ( .A1(n16880), .A2(n13813), .A3(n13812), .ZN(n13814) );
  INV_X1 U17322 ( .A(n18746), .ZN(n16903) );
  NOR2_X1 U17323 ( .A1(n19300), .A2(n16903), .ZN(n18681) );
  NOR3_X1 U17324 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18681), .A3(
        n18834), .ZN(n18847) );
  INV_X1 U17325 ( .A(n18847), .ZN(n13818) );
  INV_X1 U17326 ( .A(n18851), .ZN(n18585) );
  INV_X1 U17327 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16842) );
  AOI21_X1 U17328 ( .B1(n18585), .B2(n18813), .A(n16842), .ZN(n13815) );
  MUX2_X1 U17329 ( .A(n13815), .B(P3_REIP_REG_0__SCAN_IN), .S(n18846), .Z(
        n13816) );
  AOI21_X1 U17330 ( .B1(n18843), .B2(n14002), .A(n13816), .ZN(n13817) );
  OAI211_X1 U17331 ( .C1(n14002), .C2(n18833), .A(n13818), .B(n13817), .ZN(
        P3_U2862) );
  INV_X1 U17332 ( .A(n13891), .ZN(n13819) );
  AOI21_X1 U17333 ( .B1(n13820), .B2(n13747), .A(n13819), .ZN(n16440) );
  INV_X1 U17334 ( .A(n16440), .ZN(n13822) );
  INV_X1 U17335 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19605) );
  INV_X1 U17336 ( .A(n15927), .ZN(n13821) );
  OAI222_X1 U17337 ( .A1(n13822), .A2(n16005), .B1(n19586), .B2(n19605), .C1(
        n14151), .C2(n13821), .ZN(P2_U2910) );
  OR2_X1 U17338 ( .A1(n14111), .A2(n17126), .ZN(n13825) );
  OAI22_X1 U17339 ( .A1(n14173), .A2(n13825), .B1(n13824), .B2(n13823), .ZN(
        n13826) );
  AND2_X1 U17340 ( .A1(n14932), .A2(n13830), .ZN(n14917) );
  INV_X1 U17341 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20482) );
  INV_X1 U17342 ( .A(DATAI_1_), .ZN(n13833) );
  NAND2_X1 U17343 ( .A1(n14866), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13832) );
  OAI21_X1 U17344 ( .B1(n14869), .B2(n13833), .A(n13832), .ZN(n20600) );
  INV_X1 U17345 ( .A(n20600), .ZN(n13834) );
  OAI222_X1 U17346 ( .A1(n14938), .A2(n14794), .B1(n14932), .B2(n20482), .C1(
        n14931), .C2(n13834), .ZN(P1_U2903) );
  INV_X1 U17347 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20485) );
  INV_X1 U17348 ( .A(DATAI_0_), .ZN(n13836) );
  NAND2_X1 U17349 ( .A1(n14866), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13835) );
  OAI21_X1 U17350 ( .B1(n14869), .B2(n13836), .A(n13835), .ZN(n20591) );
  INV_X1 U17351 ( .A(n20591), .ZN(n13837) );
  OAI222_X1 U17352 ( .A1(n14938), .A2(n14802), .B1(n14932), .B2(n20485), .C1(
        n14931), .C2(n13837), .ZN(P1_U2904) );
  OAI21_X1 U17353 ( .B1(n10289), .B2(n10794), .A(n13838), .ZN(n20437) );
  NOR2_X1 U17354 ( .A1(n13840), .A2(n13841), .ZN(n13842) );
  OR2_X1 U17355 ( .A1(n13839), .A2(n13842), .ZN(n20424) );
  OAI22_X1 U17356 ( .A1(n14835), .A2(n20424), .B1(n20443), .B2(n20452), .ZN(
        n13843) );
  INV_X1 U17357 ( .A(n13843), .ZN(n13844) );
  OAI21_X1 U17358 ( .B1(n20437), .B2(n14838), .A(n13844), .ZN(P1_U2870) );
  AND2_X1 U17359 ( .A1(n13846), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n15999) );
  NAND2_X1 U17360 ( .A1(n13845), .A2(n15999), .ZN(n16001) );
  XOR2_X1 U17361 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n16001), .Z(n13848)
         );
  MUX2_X1 U17362 ( .A(n16223), .B(n12350), .S(n19570), .Z(n13847) );
  OAI21_X1 U17363 ( .B1(n13848), .B2(n19571), .A(n13847), .ZN(P2_U2882) );
  OAI21_X1 U17364 ( .B1(n13851), .B2(n13850), .A(n13849), .ZN(n15763) );
  INV_X1 U17365 ( .A(n15763), .ZN(n16498) );
  NAND2_X1 U17366 ( .A1(n19782), .A2(n16498), .ZN(n13931) );
  OAI21_X1 U17367 ( .B1(n19782), .B2(n16498), .A(n13931), .ZN(n13852) );
  NOR2_X1 U17368 ( .A1(n13852), .A2(n13853), .ZN(n13933) );
  AOI21_X1 U17369 ( .B1(n13853), .B2(n13852), .A(n13933), .ZN(n13856) );
  INV_X1 U17370 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19621) );
  OAI22_X1 U17371 ( .A1(n15981), .A2(n16498), .B1(n19586), .B2(n19621), .ZN(
        n13854) );
  AOI21_X1 U17372 ( .B1(n19577), .B2(n16538), .A(n13854), .ZN(n13855) );
  OAI21_X1 U17373 ( .B1(n13856), .B2(n16013), .A(n13855), .ZN(P2_U2918) );
  INV_X1 U17374 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20480) );
  INV_X1 U17375 ( .A(DATAI_2_), .ZN(n21388) );
  NAND2_X1 U17376 ( .A1(n14869), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13857) );
  OAI21_X1 U17377 ( .B1(n14869), .B2(n21388), .A(n13857), .ZN(n14900) );
  INV_X1 U17378 ( .A(n14900), .ZN(n13858) );
  OAI222_X1 U17379 ( .A1(n20437), .A2(n14938), .B1(n14932), .B2(n20480), .C1(
        n14931), .C2(n13858), .ZN(P1_U2902) );
  INV_X1 U17380 ( .A(n16594), .ZN(n13860) );
  NAND2_X1 U17381 ( .A1(n13860), .A2(n13859), .ZN(n16576) );
  INV_X1 U17382 ( .A(n16518), .ZN(n13863) );
  NAND2_X1 U17383 ( .A1(n13863), .A2(n13862), .ZN(n16573) );
  AOI22_X1 U17384 ( .A1(n16576), .A2(n16573), .B1(n13864), .B2(n12038), .ZN(
        n13869) );
  INV_X1 U17385 ( .A(n16571), .ZN(n16515) );
  NAND2_X1 U17386 ( .A1(n16257), .A2(n16515), .ZN(n13868) );
  INV_X1 U17387 ( .A(n13866), .ZN(n13867) );
  OAI211_X1 U17388 ( .C1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n13869), .A(
        n13868), .B(n13867), .ZN(n16586) );
  AOI22_X1 U17389 ( .A1(n20309), .A2(n17152), .B1(n16586), .B2(n20305), .ZN(
        n13877) );
  NAND2_X1 U17390 ( .A1(n13871), .A2(n13870), .ZN(n16582) );
  NAND2_X1 U17391 ( .A1(n12038), .A2(n13872), .ZN(n16578) );
  NAND2_X1 U17392 ( .A1(n16578), .A2(n16573), .ZN(n13873) );
  AOI21_X1 U17393 ( .B1(n16582), .B2(n9609), .A(n13873), .ZN(n16587) );
  INV_X1 U17394 ( .A(n16587), .ZN(n13874) );
  AOI21_X1 U17395 ( .B1(n13874), .B2(n20305), .A(n20301), .ZN(n13876) );
  OAI22_X1 U17396 ( .A1(n13877), .A2(n20301), .B1(n13876), .B2(n13875), .ZN(
        P2_U3596) );
  NOR2_X1 U17397 ( .A1(n16001), .A2(n13878), .ZN(n13990) );
  XNOR2_X1 U17398 ( .A(n13990), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13883) );
  OR2_X1 U17399 ( .A1(n9731), .A2(n13880), .ZN(n13881) );
  AND2_X1 U17400 ( .A1(n13879), .A2(n13881), .ZN(n16209) );
  INV_X1 U17401 ( .A(n16209), .ZN(n17134) );
  MUX2_X1 U17402 ( .A(n17134), .B(n12355), .S(n19570), .Z(n13882) );
  OAI21_X1 U17403 ( .B1(n13883), .B2(n19571), .A(n13882), .ZN(P2_U2880) );
  OAI21_X1 U17404 ( .B1(n13885), .B2(n13884), .A(n14055), .ZN(n14061) );
  INV_X1 U17405 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13889) );
  OR2_X1 U17406 ( .A1(n13839), .A2(n13887), .ZN(n13888) );
  NAND2_X1 U17407 ( .A1(n13886), .A2(n13888), .ZN(n20535) );
  OAI222_X1 U17408 ( .A1(n14061), .A2(n14838), .B1(n20452), .B2(n13889), .C1(
        n20535), .C2(n14835), .ZN(P1_U2869) );
  AND2_X1 U17409 ( .A1(n13891), .A2(n13890), .ZN(n13892) );
  NOR2_X1 U17410 ( .A1(n13893), .A2(n13892), .ZN(n16426) );
  INV_X1 U17411 ( .A(n16426), .ZN(n13895) );
  AOI22_X1 U17412 ( .A1(n19577), .A2(n15919), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n16010), .ZN(n13894) );
  OAI21_X1 U17413 ( .B1(n13895), .B2(n16005), .A(n13894), .ZN(P2_U2909) );
  INV_X1 U17414 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20478) );
  INV_X1 U17415 ( .A(DATAI_3_), .ZN(n13897) );
  NAND2_X1 U17416 ( .A1(n14866), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13896) );
  OAI21_X1 U17417 ( .B1(n14866), .B2(n13897), .A(n13896), .ZN(n20614) );
  INV_X1 U17418 ( .A(n20614), .ZN(n13898) );
  OAI222_X1 U17419 ( .A1(n14938), .A2(n14061), .B1(n14932), .B2(n20478), .C1(
        n14931), .C2(n13898), .ZN(P1_U2901) );
  INV_X1 U17420 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13899) );
  NOR2_X1 U17421 ( .A1(n16001), .A2(n13899), .ZN(n13901) );
  INV_X1 U17422 ( .A(n13990), .ZN(n13900) );
  OAI211_X1 U17423 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13901), .A(
        n13900), .B(n15883), .ZN(n13906) );
  NOR2_X1 U17424 ( .A1(n9753), .A2(n13902), .ZN(n13903) );
  OR2_X1 U17425 ( .A1(n9731), .A2(n13903), .ZN(n19533) );
  INV_X1 U17426 ( .A(n19533), .ZN(n13904) );
  NAND2_X1 U17427 ( .A1(n13904), .A2(n19575), .ZN(n13905) );
  OAI211_X1 U17428 ( .C1(n19575), .C2(n12352), .A(n13906), .B(n13905), .ZN(
        P2_U2881) );
  AND2_X1 U17429 ( .A1(n13994), .A2(n13907), .ZN(n13909) );
  OR2_X1 U17430 ( .A1(n13909), .A2(n13908), .ZN(n16427) );
  NAND3_X1 U17431 ( .A1(n13845), .A2(n13911), .A3(n13910), .ZN(n13992) );
  INV_X1 U17432 ( .A(n13992), .ZN(n13913) );
  OAI211_X1 U17433 ( .C1(n13913), .C2(n13912), .A(n15883), .B(n14010), .ZN(
        n13915) );
  NAND2_X1 U17434 ( .A1(n19570), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13914) );
  OAI211_X1 U17435 ( .C1(n16427), .C2(n19570), .A(n13915), .B(n13914), .ZN(
        P2_U2877) );
  NAND2_X1 U17436 ( .A1(n19294), .A2(n19466), .ZN(n16881) );
  AOI21_X2 U17437 ( .B1(n17051), .B2(n10309), .A(n16881), .ZN(n16884) );
  NOR2_X1 U17438 ( .A1(n18031), .A2(n18889), .ZN(n13918) );
  NOR3_X1 U17439 ( .A1(n16937), .A2(n18133), .A3(n19471), .ZN(n13920) );
  OAI21_X2 U17440 ( .B1(n16884), .B2(n13920), .A(n19469), .ZN(n13921) );
  NAND2_X1 U17441 ( .A1(n16886), .A2(n18100), .ZN(n18123) );
  INV_X1 U17442 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18187) );
  NOR2_X1 U17443 ( .A1(n13921), .A2(n18187), .ZN(n16662) );
  INV_X1 U17444 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21450) );
  INV_X1 U17445 ( .A(n16662), .ZN(n13922) );
  OAI221_X1 U17446 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n16662), .C1(n21450), 
        .C2(n13922), .A(n18118), .ZN(n13925) );
  NAND2_X1 U17447 ( .A1(n13923), .A2(n18127), .ZN(n13924) );
  OAI211_X1 U17448 ( .C1(n18123), .C2(n13926), .A(n13925), .B(n13924), .ZN(
        P3_U2734) );
  OAI21_X1 U17449 ( .B1(n17518), .B2(n17584), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n13930) );
  NOR2_X1 U17450 ( .A1(n18133), .A2(n19486), .ZN(n19489) );
  INV_X1 U17451 ( .A(n19489), .ZN(n16660) );
  NAND3_X1 U17452 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16931), .A3(
        n17573), .ZN(n13927) );
  OAI21_X1 U17453 ( .B1(n16660), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13927), .ZN(n13928) );
  AOI21_X1 U17454 ( .B1(n17450), .B2(P3_REIP_REG_0__SCAN_IN), .A(n13928), .ZN(
        n13929) );
  NAND2_X1 U17455 ( .A1(n13930), .A2(n13929), .ZN(P3_U2671) );
  INV_X1 U17456 ( .A(n13931), .ZN(n13932) );
  NOR2_X1 U17457 ( .A1(n13933), .A2(n13932), .ZN(n13939) );
  OR2_X1 U17458 ( .A1(n13935), .A2(n13934), .ZN(n13936) );
  NAND2_X1 U17459 ( .A1(n13937), .A2(n13936), .ZN(n19664) );
  INV_X1 U17460 ( .A(n19664), .ZN(n20319) );
  NAND2_X1 U17461 ( .A1(n20299), .A2(n20319), .ZN(n15992) );
  OAI21_X1 U17462 ( .B1(n20299), .B2(n20319), .A(n15992), .ZN(n13938) );
  NOR2_X1 U17463 ( .A1(n13938), .A2(n13939), .ZN(n15994) );
  AOI21_X1 U17464 ( .B1(n13939), .B2(n13938), .A(n15994), .ZN(n13942) );
  INV_X1 U17465 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19619) );
  OAI22_X1 U17466 ( .A1(n15981), .A2(n20319), .B1(n19586), .B2(n19619), .ZN(
        n13940) );
  AOI21_X1 U17467 ( .B1(n16541), .B2(n19577), .A(n13940), .ZN(n13941) );
  OAI21_X1 U17468 ( .B1(n13942), .B2(n16013), .A(n13941), .ZN(P2_U2917) );
  NOR2_X1 U17469 ( .A1(n14101), .A2(n21293), .ZN(n13943) );
  NOR2_X2 U17470 ( .A1(n20512), .A2(n13946), .ZN(n20497) );
  INV_X1 U17471 ( .A(DATAI_5_), .ZN(n13945) );
  NAND2_X1 U17472 ( .A1(n14866), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13944) );
  OAI21_X1 U17473 ( .B1(n14869), .B2(n13945), .A(n13944), .ZN(n20631) );
  NAND2_X1 U17474 ( .A1(n20497), .A2(n20631), .ZN(n13968) );
  AND2_X2 U17475 ( .A1(n13981), .A2(n13946), .ZN(n20509) );
  AOI22_X1 U17476 ( .A1(n20509), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13947) );
  NAND2_X1 U17477 ( .A1(n13968), .A2(n13947), .ZN(P1_U2957) );
  INV_X1 U17478 ( .A(DATAI_7_), .ZN(n13949) );
  NAND2_X1 U17479 ( .A1(n14866), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13948) );
  OAI21_X1 U17480 ( .B1(n14869), .B2(n13949), .A(n13948), .ZN(n20652) );
  NAND2_X1 U17481 ( .A1(n20497), .A2(n20652), .ZN(n13957) );
  AOI22_X1 U17482 ( .A1(n20509), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U17483 ( .A1(n13957), .A2(n13950), .ZN(P1_U2959) );
  INV_X1 U17484 ( .A(DATAI_6_), .ZN(n13952) );
  NAND2_X1 U17485 ( .A1(n14866), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13951) );
  OAI21_X1 U17486 ( .B1(n14869), .B2(n13952), .A(n13951), .ZN(n20639) );
  NAND2_X1 U17487 ( .A1(n20497), .A2(n20639), .ZN(n13955) );
  AOI22_X1 U17488 ( .A1(n20509), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13953) );
  NAND2_X1 U17489 ( .A1(n13955), .A2(n13953), .ZN(P1_U2958) );
  AOI22_X1 U17490 ( .A1(n20509), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13954) );
  NAND2_X1 U17491 ( .A1(n13955), .A2(n13954), .ZN(P1_U2943) );
  AOI22_X1 U17492 ( .A1(n20509), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U17493 ( .A1(n13957), .A2(n13956), .ZN(P1_U2944) );
  NAND2_X1 U17494 ( .A1(n20497), .A2(n14900), .ZN(n13970) );
  AOI22_X1 U17495 ( .A1(n20509), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13958) );
  NAND2_X1 U17496 ( .A1(n13970), .A2(n13958), .ZN(P1_U2954) );
  NAND2_X1 U17497 ( .A1(n20497), .A2(n20591), .ZN(n13961) );
  AOI22_X1 U17498 ( .A1(n20509), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13959) );
  NAND2_X1 U17499 ( .A1(n13961), .A2(n13959), .ZN(P1_U2952) );
  AOI22_X1 U17500 ( .A1(n20509), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13960) );
  NAND2_X1 U17501 ( .A1(n13961), .A2(n13960), .ZN(P1_U2937) );
  NAND2_X1 U17502 ( .A1(n20497), .A2(n20600), .ZN(n13972) );
  AOI22_X1 U17503 ( .A1(n20509), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U17504 ( .A1(n13972), .A2(n13962), .ZN(P1_U2953) );
  NAND2_X1 U17505 ( .A1(n20497), .A2(n20614), .ZN(n13976) );
  AOI22_X1 U17506 ( .A1(n20509), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13963) );
  NAND2_X1 U17507 ( .A1(n13976), .A2(n13963), .ZN(P1_U2955) );
  INV_X1 U17508 ( .A(DATAI_4_), .ZN(n13965) );
  NAND2_X1 U17509 ( .A1(n14866), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13964) );
  OAI21_X1 U17510 ( .B1(n14866), .B2(n13965), .A(n13964), .ZN(n20622) );
  NAND2_X1 U17511 ( .A1(n20497), .A2(n20622), .ZN(n13974) );
  AOI22_X1 U17512 ( .A1(n20509), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U17513 ( .A1(n13974), .A2(n13966), .ZN(P1_U2956) );
  AOI22_X1 U17514 ( .A1(n20509), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13967) );
  NAND2_X1 U17515 ( .A1(n13968), .A2(n13967), .ZN(P1_U2942) );
  AOI22_X1 U17516 ( .A1(n20509), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13969) );
  NAND2_X1 U17517 ( .A1(n13970), .A2(n13969), .ZN(P1_U2939) );
  AOI22_X1 U17518 ( .A1(n20509), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13971) );
  NAND2_X1 U17519 ( .A1(n13972), .A2(n13971), .ZN(P1_U2938) );
  AOI22_X1 U17520 ( .A1(n20509), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13973) );
  NAND2_X1 U17521 ( .A1(n13974), .A2(n13973), .ZN(P1_U2941) );
  AOI22_X1 U17522 ( .A1(n20509), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13975) );
  NAND2_X1 U17523 ( .A1(n13976), .A2(n13975), .ZN(P1_U2940) );
  INV_X1 U17524 ( .A(n15911), .ZN(n13977) );
  INV_X1 U17525 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19601) );
  OAI222_X1 U17526 ( .A1(n16412), .A2(n16005), .B1(n13977), .B2(n14151), .C1(
        n19601), .C2(n19586), .ZN(P2_U2908) );
  INV_X1 U17527 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14919) );
  INV_X1 U17528 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20456) );
  INV_X1 U17529 ( .A(n20497), .ZN(n13980) );
  INV_X1 U17530 ( .A(DATAI_15_), .ZN(n13979) );
  MUX2_X1 U17531 ( .A(n13979), .B(n13978), .S(n14869), .Z(n14920) );
  OAI222_X1 U17532 ( .A1(n13985), .A2(n14919), .B1(n13981), .B2(n20456), .C1(
        n13980), .C2(n14920), .ZN(P1_U2967) );
  INV_X1 U17533 ( .A(DATAI_13_), .ZN(n13983) );
  NAND2_X1 U17534 ( .A1(n14866), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13982) );
  OAI21_X1 U17535 ( .B1(n14866), .B2(n13983), .A(n13982), .ZN(n14924) );
  NAND2_X1 U17536 ( .A1(n20497), .A2(n14924), .ZN(n20510) );
  NAND2_X1 U17537 ( .A1(n20512), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13984) );
  OAI211_X1 U17538 ( .C1(n11232), .C2(n13985), .A(n20510), .B(n13984), .ZN(
        P1_U2950) );
  INV_X1 U17539 ( .A(n13986), .ZN(n13987) );
  XNOR2_X1 U17540 ( .A(n14087), .B(n13987), .ZN(n19520) );
  INV_X1 U17541 ( .A(n19520), .ZN(n13989) );
  AOI22_X1 U17542 ( .A1(n19577), .A2(n15904), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n16010), .ZN(n13988) );
  OAI21_X1 U17543 ( .B1(n13989), .B2(n16005), .A(n13988), .ZN(P2_U2907) );
  INV_X1 U17544 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13998) );
  NAND2_X1 U17545 ( .A1(n13990), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n15891) );
  INV_X1 U17546 ( .A(n13991), .ZN(n15892) );
  NOR2_X1 U17547 ( .A1(n15891), .A2(n15892), .ZN(n15890) );
  OAI211_X1 U17548 ( .C1(n15890), .C2(n13993), .A(n15883), .B(n13992), .ZN(
        n13997) );
  AOI21_X1 U17549 ( .B1(n13995), .B2(n15700), .A(n10224), .ZN(n16441) );
  NAND2_X1 U17550 ( .A1(n16441), .A2(n19575), .ZN(n13996) );
  OAI211_X1 U17551 ( .C1(n19575), .C2(n13998), .A(n13997), .B(n13996), .ZN(
        P2_U2878) );
  INV_X1 U17552 ( .A(n18552), .ZN(n18515) );
  NAND2_X1 U17553 ( .A1(n18515), .A2(n14002), .ZN(n14001) );
  NAND3_X1 U17554 ( .A1(n16879), .A2(n19360), .A3(n18547), .ZN(n13999) );
  AOI22_X1 U17555 ( .A1(n18846), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13999), .ZN(n14000) );
  OAI211_X1 U17556 ( .C1(n14002), .C2(n18484), .A(n14001), .B(n14000), .ZN(
        P3_U2830) );
  OAI21_X1 U17557 ( .B1(n14004), .B2(n14003), .A(n14193), .ZN(n17106) );
  INV_X1 U17558 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14008) );
  NAND2_X1 U17559 ( .A1(n14005), .A2(n14006), .ZN(n14007) );
  NAND2_X1 U17560 ( .A1(n17116), .A2(n14007), .ZN(n20407) );
  OAI222_X1 U17561 ( .A1(n17106), .A2(n14838), .B1(n14008), .B2(n20452), .C1(
        n14835), .C2(n20407), .ZN(P1_U2867) );
  INV_X1 U17562 ( .A(n16418), .ZN(n14009) );
  NAND2_X1 U17563 ( .A1(n14009), .A2(n19575), .ZN(n14013) );
  OAI211_X1 U17564 ( .C1(n10204), .C2(n14011), .A(n15883), .B(n14048), .ZN(
        n14012) );
  OAI211_X1 U17565 ( .C1(n19575), .C2(n12356), .A(n14013), .B(n14012), .ZN(
        P2_U2876) );
  INV_X1 U17566 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20474) );
  INV_X1 U17567 ( .A(n20631), .ZN(n14014) );
  OAI222_X1 U17568 ( .A1(n14938), .A2(n17106), .B1(n14932), .B2(n20474), .C1(
        n14931), .C2(n14014), .ZN(P1_U2899) );
  INV_X1 U17569 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14016) );
  AOI22_X1 U17570 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14015) );
  OAI21_X1 U17571 ( .B1(n14016), .B2(n14036), .A(n14015), .ZN(P1_U2906) );
  INV_X1 U17572 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14018) );
  AOI22_X1 U17573 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14017) );
  OAI21_X1 U17574 ( .B1(n14018), .B2(n14036), .A(n14017), .ZN(P1_U2913) );
  INV_X1 U17575 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U17576 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14019) );
  OAI21_X1 U17577 ( .B1(n14020), .B2(n14036), .A(n14019), .ZN(P1_U2917) );
  INV_X1 U17578 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17579 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14021) );
  OAI21_X1 U17580 ( .B1(n14022), .B2(n14036), .A(n14021), .ZN(P1_U2920) );
  INV_X1 U17581 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14024) );
  AOI22_X1 U17582 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14023) );
  OAI21_X1 U17583 ( .B1(n14024), .B2(n14036), .A(n14023), .ZN(P1_U2909) );
  INV_X1 U17584 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U17585 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14025) );
  OAI21_X1 U17586 ( .B1(n14026), .B2(n14036), .A(n14025), .ZN(P1_U2914) );
  INV_X1 U17587 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14028) );
  AOI22_X1 U17588 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14027) );
  OAI21_X1 U17589 ( .B1(n14028), .B2(n14036), .A(n14027), .ZN(P1_U2915) );
  INV_X1 U17590 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17591 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14029) );
  OAI21_X1 U17592 ( .B1(n14030), .B2(n14036), .A(n14029), .ZN(P1_U2916) );
  INV_X1 U17593 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17594 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14031) );
  OAI21_X1 U17595 ( .B1(n14032), .B2(n14036), .A(n14031), .ZN(P1_U2912) );
  INV_X1 U17596 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14034) );
  AOI22_X1 U17597 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14033) );
  OAI21_X1 U17598 ( .B1(n14034), .B2(n14036), .A(n14033), .ZN(P1_U2918) );
  INV_X1 U17599 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n21451) );
  AOI22_X1 U17600 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14035) );
  OAI21_X1 U17601 ( .B1(n21451), .B2(n14036), .A(n14035), .ZN(P1_U2919) );
  INV_X1 U17602 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14792) );
  NAND2_X1 U17603 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14037) );
  NAND2_X1 U17604 ( .A1(n20580), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20560) );
  NAND2_X1 U17605 ( .A1(n14037), .A2(n20560), .ZN(n14042) );
  XNOR2_X1 U17606 ( .A(n14038), .B(n14070), .ZN(n14039) );
  NOR2_X1 U17607 ( .A1(n14039), .A2(n20571), .ZN(n20564) );
  INV_X1 U17608 ( .A(n14039), .ZN(n14040) );
  NOR2_X1 U17609 ( .A1(n14040), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20563) );
  INV_X2 U17610 ( .A(n20518), .ZN(n15151) );
  NOR3_X1 U17611 ( .A1(n20564), .A2(n20563), .A3(n15151), .ZN(n14041) );
  AOI211_X1 U17612 ( .C1(n15119), .C2(n14792), .A(n14042), .B(n14041), .ZN(
        n14043) );
  OAI21_X1 U17613 ( .B1(n15122), .B2(n14794), .A(n14043), .ZN(P1_U2998) );
  NAND2_X1 U17614 ( .A1(n13493), .A2(n14044), .ZN(n14045) );
  NAND2_X1 U17615 ( .A1(n14046), .A2(n14045), .ZN(n19521) );
  INV_X1 U17616 ( .A(n14048), .ZN(n14051) );
  INV_X1 U17617 ( .A(n14050), .ZN(n14047) );
  NOR2_X1 U17618 ( .A1(n14048), .A2(n14047), .ZN(n15886) );
  INV_X1 U17619 ( .A(n15886), .ZN(n14049) );
  OAI211_X1 U17620 ( .C1(n14051), .C2(n14050), .A(n14049), .B(n15883), .ZN(
        n14053) );
  NAND2_X1 U17621 ( .A1(n19570), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14052) );
  OAI211_X1 U17622 ( .C1(n19521), .C2(n19570), .A(n14053), .B(n14052), .ZN(
        P2_U2875) );
  INV_X1 U17623 ( .A(n20622), .ZN(n14057) );
  XOR2_X1 U17624 ( .A(n14055), .B(n14054), .Z(n20520) );
  INV_X1 U17625 ( .A(n20520), .ZN(n14056) );
  INV_X1 U17626 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20476) );
  OAI222_X1 U17627 ( .A1(n14931), .A2(n14057), .B1(n14938), .B2(n14056), .C1(
        n20476), .C2(n14932), .ZN(P1_U2900) );
  XNOR2_X1 U17628 ( .A(n14058), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14060) );
  XNOR2_X1 U17629 ( .A(n14060), .B(n14059), .ZN(n20534) );
  INV_X1 U17630 ( .A(n14061), .ZN(n14785) );
  AOI22_X1 U17631 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20580), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14062) );
  OAI21_X1 U17632 ( .B1(n20524), .B2(n14783), .A(n14062), .ZN(n14063) );
  AOI21_X1 U17633 ( .B1(n14785), .B2(n20519), .A(n14063), .ZN(n14064) );
  OAI21_X1 U17634 ( .B1(n15151), .B2(n20534), .A(n14064), .ZN(P1_U2996) );
  NOR2_X1 U17635 ( .A1(n14065), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14067) );
  OAI211_X1 U17636 ( .C1(n21093), .C2(n14068), .A(n14067), .B(n14066), .ZN(
        n14069) );
  NAND2_X1 U17637 ( .A1(n14070), .A2(n14069), .ZN(n20575) );
  INV_X1 U17638 ( .A(n20575), .ZN(n14075) );
  INV_X1 U17639 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14073) );
  OAI21_X1 U17640 ( .B1(n17105), .B2(n14071), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14072) );
  OAI21_X1 U17641 ( .B1(n14073), .B2(n20416), .A(n14072), .ZN(n14074) );
  AOI21_X1 U17642 ( .B1(n20518), .B2(n14075), .A(n14074), .ZN(n14076) );
  OAI21_X1 U17643 ( .B1(n15122), .B2(n14802), .A(n14076), .ZN(P1_U2999) );
  OAI21_X1 U17644 ( .B1(n14079), .B2(n14078), .A(n14077), .ZN(n14080) );
  INV_X1 U17645 ( .A(n14080), .ZN(n20551) );
  INV_X1 U17646 ( .A(n20427), .ZN(n14082) );
  AOI22_X1 U17647 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20580), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14081) );
  OAI21_X1 U17648 ( .B1(n20524), .B2(n14082), .A(n14081), .ZN(n14083) );
  AOI21_X1 U17649 ( .B1(n20551), .B2(n20518), .A(n14083), .ZN(n14084) );
  OAI21_X1 U17650 ( .B1(n20437), .B2(n15122), .A(n14084), .ZN(P1_U2997) );
  INV_X1 U17651 ( .A(n14085), .ZN(n14088) );
  NOR2_X1 U17652 ( .A1(n14087), .A2(n14086), .ZN(n14147) );
  AOI21_X1 U17653 ( .B1(n14089), .B2(n14088), .A(n14147), .ZN(n16372) );
  INV_X1 U17654 ( .A(n16372), .ZN(n14091) );
  AOI22_X1 U17655 ( .A1(n19577), .A2(n19627), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n16010), .ZN(n14090) );
  OAI21_X1 U17656 ( .B1(n14091), .B2(n16005), .A(n14090), .ZN(P2_U2905) );
  INV_X1 U17657 ( .A(n20517), .ZN(n14092) );
  INV_X1 U17658 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20533) );
  NOR2_X1 U17659 ( .A1(n14092), .A2(n20533), .ZN(n14093) );
  OAI22_X1 U17660 ( .A1(n14093), .A2(n20515), .B1(n20517), .B2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14096) );
  XNOR2_X1 U17661 ( .A(n14094), .B(n14129), .ZN(n14095) );
  XNOR2_X1 U17662 ( .A(n14096), .B(n14095), .ZN(n17107) );
  NAND2_X1 U17663 ( .A1(n10431), .A2(n14100), .ZN(n14099) );
  INV_X1 U17664 ( .A(n14097), .ZN(n14098) );
  NAND2_X1 U17665 ( .A1(n14099), .A2(n14098), .ZN(n14106) );
  OAI21_X1 U17666 ( .B1(n14268), .B2(n17126), .A(n10476), .ZN(n14104) );
  NAND2_X1 U17667 ( .A1(n14101), .A2(n14100), .ZN(n14103) );
  AOI21_X1 U17668 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(n14105) );
  AOI21_X1 U17669 ( .B1(n14173), .B2(n14108), .A(n14107), .ZN(n14109) );
  NAND2_X1 U17670 ( .A1(n14130), .A2(n10414), .ZN(n14110) );
  NAND4_X1 U17671 ( .A1(n14112), .A2(n15394), .A3(n14111), .A4(n14110), .ZN(
        n14113) );
  NAND2_X2 U17672 ( .A1(n14134), .A2(n14113), .ZN(n20576) );
  NAND2_X1 U17673 ( .A1(n14134), .A2(n17060), .ZN(n20582) );
  OR2_X1 U17674 ( .A1(n14115), .A2(n13361), .ZN(n14121) );
  OAI21_X1 U17675 ( .B1(n14116), .B2(n10419), .A(n20649), .ZN(n14117) );
  OAI21_X1 U17676 ( .B1(n14117), .B2(n15378), .A(n10431), .ZN(n14118) );
  AND4_X1 U17677 ( .A1(n14121), .A2(n14120), .A3(n14119), .A4(n14118), .ZN(
        n14123) );
  AND2_X1 U17678 ( .A1(n14123), .A2(n14122), .ZN(n14270) );
  OAI211_X1 U17679 ( .C1(n14114), .C2(n10476), .A(n14270), .B(n14124), .ZN(
        n14125) );
  NAND2_X1 U17680 ( .A1(n14134), .A2(n14125), .ZN(n20572) );
  INV_X1 U17681 ( .A(n20582), .ZN(n14126) );
  NOR2_X1 U17682 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14126), .ZN(
        n20565) );
  INV_X1 U17683 ( .A(n20565), .ZN(n14127) );
  NAND2_X1 U17684 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14226) );
  INV_X1 U17685 ( .A(n14226), .ZN(n14337) );
  NAND2_X1 U17686 ( .A1(n20553), .A2(n14337), .ZN(n14212) );
  INV_X1 U17687 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20559) );
  OAI21_X1 U17688 ( .B1(n20559), .B2(n20571), .A(n20552), .ZN(n20541) );
  NAND2_X1 U17689 ( .A1(n20573), .A2(n20541), .ZN(n14128) );
  NOR2_X1 U17690 ( .A1(n20533), .A2(n20539), .ZN(n20528) );
  NAND2_X1 U17691 ( .A1(n20528), .A2(n14129), .ZN(n14211) );
  NAND2_X1 U17692 ( .A1(n14130), .A2(n10445), .ZN(n14131) );
  OAI21_X1 U17693 ( .B1(n14268), .B2(n21298), .A(n14131), .ZN(n14132) );
  INV_X1 U17694 ( .A(n20407), .ZN(n14133) );
  AOI22_X1 U17695 ( .A1(n20544), .A2(n14133), .B1(n20580), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n14142) );
  OR2_X1 U17696 ( .A1(n20572), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14136) );
  NAND2_X1 U17697 ( .A1(n14136), .A2(n14135), .ZN(n20558) );
  NAND2_X1 U17698 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20528), .ZN(
        n14336) );
  INV_X1 U17699 ( .A(n14336), .ZN(n14137) );
  NAND2_X1 U17700 ( .A1(n14137), .A2(n20541), .ZN(n14228) );
  NAND2_X1 U17701 ( .A1(n20573), .A2(n14228), .ZN(n14138) );
  NAND2_X1 U17702 ( .A1(n20547), .A2(n14138), .ZN(n15330) );
  NAND2_X1 U17703 ( .A1(n14337), .A2(n20528), .ZN(n14139) );
  AND2_X1 U17704 ( .A1(n20546), .A2(n14139), .ZN(n14140) );
  OR2_X1 U17705 ( .A1(n15330), .A2(n14140), .ZN(n14214) );
  NAND2_X1 U17706 ( .A1(n14214), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14141) );
  OAI211_X1 U17707 ( .C1(n20540), .C2(n14211), .A(n14142), .B(n14141), .ZN(
        n14143) );
  AOI21_X1 U17708 ( .B1(n17107), .B2(n20550), .A(n14143), .ZN(n14144) );
  INV_X1 U17709 ( .A(n14144), .ZN(P1_U3026) );
  OR2_X1 U17710 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  AND2_X1 U17711 ( .A1(n14145), .A2(n14148), .ZN(n16358) );
  INV_X1 U17712 ( .A(n16358), .ZN(n14150) );
  OAI222_X1 U17713 ( .A1(n14150), .A2(n16005), .B1(n19586), .B2(n13595), .C1(
        n14149), .C2(n14151), .ZN(P2_U2904) );
  INV_X1 U17714 ( .A(n15897), .ZN(n14152) );
  INV_X1 U17715 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19597) );
  OAI222_X1 U17716 ( .A1(n14153), .A2(n16005), .B1(n14152), .B2(n14151), .C1(
        n19597), .C2(n19586), .ZN(P2_U2906) );
  OAI21_X1 U17717 ( .B1(n15870), .B2(n14155), .A(n15861), .ZN(n15867) );
  AOI21_X1 U17718 ( .B1(n14156), .B2(n15635), .A(n15591), .ZN(n14255) );
  NAND2_X1 U17719 ( .A1(n15983), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U17720 ( .A1(n15984), .A2(BUF2_REG_17__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U17721 ( .A1(n15985), .A2(n16538), .B1(n16010), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14157) );
  NAND3_X1 U17722 ( .A1(n14159), .A2(n14158), .A3(n14157), .ZN(n14160) );
  AOI21_X1 U17723 ( .B1(n14255), .B2(n19578), .A(n14160), .ZN(n14161) );
  OAI21_X1 U17724 ( .B1(n16013), .B2(n15867), .A(n14161), .ZN(P2_U2902) );
  INV_X1 U17725 ( .A(n21093), .ZN(n14163) );
  NAND2_X1 U17726 ( .A1(n20690), .A2(n21241), .ZN(n14164) );
  NAND2_X1 U17727 ( .A1(n14164), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14165) );
  NAND2_X1 U17728 ( .A1(n14165), .A2(n21186), .ZN(n14180) );
  INV_X1 U17729 ( .A(n14167), .ZN(n14169) );
  NAND2_X1 U17730 ( .A1(n14169), .A2(n14168), .ZN(n14170) );
  OR2_X1 U17731 ( .A1(n20893), .A2(n21031), .ZN(n20721) );
  INV_X1 U17732 ( .A(n14172), .ZN(n21133) );
  NOR2_X1 U17733 ( .A1(n20721), .A2(n21133), .ZN(n14178) );
  OR2_X1 U17734 ( .A1(n14180), .A2(n14178), .ZN(n14177) );
  NAND2_X1 U17735 ( .A1(n20896), .A2(n20963), .ZN(n20756) );
  NAND3_X1 U17736 ( .A1(n17071), .A2(n10743), .A3(n21033), .ZN(n20659) );
  NOR2_X1 U17737 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20659), .ZN(
        n20590) );
  INV_X1 U17738 ( .A(n20590), .ZN(n20650) );
  NAND2_X1 U17739 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20650), .ZN(n14174) );
  NAND2_X1 U17740 ( .A1(n14181), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20821) );
  NAND2_X1 U17741 ( .A1(n20653), .A2(n20821), .ZN(n20694) );
  NAND2_X1 U17742 ( .A1(n14174), .A2(n20967), .ZN(n14175) );
  AOI21_X1 U17743 ( .B1(n20756), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n14175), 
        .ZN(n14176) );
  INV_X1 U17744 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14192) );
  NAND2_X1 U17745 ( .A1(n20653), .A2(n14900), .ZN(n21200) );
  INV_X1 U17746 ( .A(n21200), .ZN(n14190) );
  INV_X1 U17747 ( .A(n14178), .ZN(n14179) );
  NOR2_X1 U17748 ( .A1(n14181), .A2(n21246), .ZN(n20964) );
  INV_X1 U17749 ( .A(n20756), .ZN(n14182) );
  NAND2_X1 U17750 ( .A1(n20964), .A2(n14182), .ZN(n14183) );
  INV_X1 U17751 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17178) );
  INV_X1 U17752 ( .A(DATAI_18_), .ZN(n14185) );
  OAI22_X1 U17753 ( .A1(n17178), .A2(n20644), .B1(n14185), .B2(n20646), .ZN(
        n21104) );
  INV_X1 U17754 ( .A(n21241), .ZN(n21221) );
  INV_X1 U17755 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21377) );
  INV_X1 U17756 ( .A(DATAI_26_), .ZN(n14186) );
  OAI22_X2 U17757 ( .A1(n21377), .A2(n20644), .B1(n14186), .B2(n20646), .ZN(
        n21202) );
  NAND2_X1 U17758 ( .A1(n14187), .A2(n20648), .ZN(n21197) );
  INV_X1 U17759 ( .A(n21197), .ZN(n20976) );
  AOI22_X1 U17760 ( .A1(n21221), .A2(n21202), .B1(n20976), .B2(n20590), .ZN(
        n14188) );
  OAI21_X1 U17761 ( .B1(n20690), .B2(n21205), .A(n14188), .ZN(n14189) );
  AOI21_X1 U17762 ( .B1(n14190), .B2(n20654), .A(n14189), .ZN(n14191) );
  OAI21_X1 U17763 ( .B1(n20613), .B2(n14192), .A(n14191), .ZN(P1_U3035) );
  INV_X1 U17764 ( .A(n20639), .ZN(n14196) );
  XOR2_X1 U17765 ( .A(n14194), .B(n14193), .Z(n20445) );
  INV_X1 U17766 ( .A(n20445), .ZN(n14195) );
  OAI222_X1 U17767 ( .A1(n14931), .A2(n14196), .B1(n14938), .B2(n14195), .C1(
        n10823), .C2(n14932), .ZN(P1_U2898) );
  INV_X1 U17768 ( .A(n14198), .ZN(n14200) );
  NAND2_X1 U17769 ( .A1(n14200), .A2(n14199), .ZN(n14201) );
  AND2_X1 U17770 ( .A1(n14197), .A2(n14201), .ZN(n20376) );
  INV_X1 U17771 ( .A(n20376), .ZN(n14207) );
  INV_X1 U17772 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14205) );
  NOR2_X1 U17773 ( .A1(n9722), .A2(n14203), .ZN(n14204) );
  OR2_X1 U17774 ( .A1(n14202), .A2(n14204), .ZN(n20373) );
  OAI222_X1 U17775 ( .A1(n14207), .A2(n14838), .B1(n14205), .B2(n20452), .C1(
        n14835), .C2(n20373), .ZN(P1_U2865) );
  INV_X1 U17776 ( .A(n20652), .ZN(n14206) );
  OAI222_X1 U17777 ( .A1(n14938), .A2(n14207), .B1(n14932), .B2(n10829), .C1(
        n14931), .C2(n14206), .ZN(P1_U2897) );
  XNOR2_X1 U17778 ( .A(n14209), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14210) );
  XNOR2_X1 U17779 ( .A(n14208), .B(n14210), .ZN(n14246) );
  NOR2_X1 U17780 ( .A1(n14212), .A2(n14211), .ZN(n14213) );
  NOR2_X1 U17781 ( .A1(n14214), .A2(n14213), .ZN(n17118) );
  NAND2_X1 U17782 ( .A1(n15293), .A2(n17100), .ZN(n14215) );
  AND2_X1 U17783 ( .A1(n17118), .A2(n14215), .ZN(n17113) );
  INV_X1 U17784 ( .A(n17113), .ZN(n14222) );
  OAI21_X1 U17785 ( .B1(n14202), .B2(n14217), .A(n14216), .ZN(n14760) );
  NAND2_X1 U17786 ( .A1(n20580), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n14241) );
  OAI21_X1 U17787 ( .B1(n14760), .B2(n20578), .A(n14241), .ZN(n14221) );
  INV_X1 U17788 ( .A(n17123), .ZN(n14218) );
  NAND2_X1 U17789 ( .A1(n14218), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17115) );
  XNOR2_X1 U17790 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14219) );
  NOR2_X1 U17791 ( .A1(n17115), .A2(n14219), .ZN(n14220) );
  AOI211_X1 U17792 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n14222), .A(
        n14221), .B(n14220), .ZN(n14223) );
  OAI21_X1 U17793 ( .B1(n14246), .B2(n20576), .A(n14223), .ZN(P1_U3023) );
  INV_X1 U17794 ( .A(n15098), .ZN(n14964) );
  XNOR2_X1 U17795 ( .A(n9623), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14225) );
  XNOR2_X1 U17796 ( .A(n14224), .B(n14225), .ZN(n15152) );
  NAND2_X1 U17797 ( .A1(n20546), .A2(n14226), .ZN(n14227) );
  NAND2_X1 U17798 ( .A1(n20547), .A2(n14227), .ZN(n20525) );
  INV_X1 U17799 ( .A(n14228), .ZN(n14229) );
  AND3_X1 U17800 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14335) );
  NAND2_X1 U17801 ( .A1(n14229), .A2(n14335), .ZN(n14230) );
  OR2_X1 U17802 ( .A1(n20525), .A2(n14230), .ZN(n14232) );
  INV_X1 U17803 ( .A(n15293), .ZN(n20566) );
  NAND2_X1 U17804 ( .A1(n20566), .A2(n20547), .ZN(n14231) );
  AND2_X1 U17805 ( .A1(n14232), .A2(n14231), .ZN(n15356) );
  OAI21_X1 U17806 ( .B1(n10134), .B2(n14234), .A(n14233), .ZN(n14836) );
  OR2_X1 U17807 ( .A1(n20416), .A2(n14235), .ZN(n15144) );
  OAI21_X1 U17808 ( .B1(n14836), .B2(n20578), .A(n15144), .ZN(n14236) );
  INV_X1 U17809 ( .A(n14335), .ZN(n15351) );
  NOR3_X1 U17810 ( .A1(n17123), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n15351), .ZN(n15357) );
  AOI211_X1 U17811 ( .C1(n15356), .C2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14236), .B(n15357), .ZN(n14237) );
  OAI21_X1 U17812 ( .B1(n15152), .B2(n20576), .A(n14237), .ZN(P1_U3022) );
  AOI21_X1 U17813 ( .B1(n14240), .B2(n14197), .A(n14239), .ZN(n14247) );
  INV_X1 U17814 ( .A(n14241), .ZN(n14242) );
  AOI21_X1 U17815 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n14242), .ZN(n14243) );
  OAI21_X1 U17816 ( .B1(n20524), .B2(n14757), .A(n14243), .ZN(n14244) );
  AOI21_X1 U17817 ( .B1(n14247), .B2(n20519), .A(n14244), .ZN(n14245) );
  OAI21_X1 U17818 ( .B1(n15151), .B2(n14246), .A(n14245), .ZN(P1_U2991) );
  INV_X1 U17819 ( .A(n14247), .ZN(n14769) );
  INV_X1 U17820 ( .A(DATAI_8_), .ZN(n14249) );
  NAND2_X1 U17821 ( .A1(n14866), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U17822 ( .B1(n14869), .B2(n14249), .A(n14248), .ZN(n20486) );
  AOI22_X1 U17823 ( .A1(n14936), .A2(n20486), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14935), .ZN(n14250) );
  OAI21_X1 U17824 ( .B1(n14769), .B2(n14938), .A(n14250), .ZN(P1_U2896) );
  OAI222_X1 U17825 ( .A1(n14769), .A2(n14838), .B1(n20452), .B2(n13292), .C1(
        n14760), .C2(n14835), .ZN(P1_U2864) );
  AOI21_X1 U17826 ( .B1(n14254), .B2(n9628), .A(n14253), .ZN(n16087) );
  INV_X1 U17827 ( .A(n14255), .ZN(n15620) );
  NAND2_X1 U17828 ( .A1(n19553), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16083) );
  OAI21_X1 U17829 ( .B1(n15620), .B2(n19648), .A(n16083), .ZN(n14259) );
  NAND2_X1 U17830 ( .A1(n16411), .A2(n14262), .ZN(n16400) );
  INV_X1 U17831 ( .A(n14257), .ZN(n14263) );
  NOR2_X1 U17832 ( .A1(n16400), .A2(n14263), .ZN(n16365) );
  OAI21_X1 U17833 ( .B1(n16408), .B2(n14262), .A(n9631), .ZN(n16403) );
  AOI21_X1 U17834 ( .B1(n14263), .B2(n9986), .A(n16403), .ZN(n16361) );
  NOR2_X1 U17835 ( .A1(n16408), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14265) );
  INV_X1 U17836 ( .A(n14266), .ZN(n14267) );
  AND3_X1 U17837 ( .A1(n14114), .A2(n14268), .A3(n14267), .ZN(n14269) );
  AND2_X1 U17838 ( .A1(n15394), .A2(n14269), .ZN(n14271) );
  NAND2_X1 U17839 ( .A1(n14271), .A2(n14270), .ZN(n15386) );
  INV_X1 U17840 ( .A(n15386), .ZN(n14275) );
  NOR2_X1 U17841 ( .A1(n14272), .A2(n14273), .ZN(n14276) );
  AOI22_X1 U17842 ( .A1(n17060), .A2(n15379), .B1(n14276), .B2(n14425), .ZN(
        n14274) );
  OAI21_X1 U17843 ( .B1(n14172), .B2(n14275), .A(n14274), .ZN(n17064) );
  AND2_X1 U17844 ( .A1(n17064), .A2(n21278), .ZN(n14280) );
  INV_X1 U17845 ( .A(n14276), .ZN(n14278) );
  NAND2_X1 U17846 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15417) );
  INV_X1 U17847 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14277) );
  AOI22_X1 U17848 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20571), .B2(n14277), .ZN(
        n15419) );
  OAI22_X1 U17849 ( .A1(n17056), .A2(n14278), .B1(n15417), .B2(n15419), .ZN(
        n14279) );
  OAI21_X1 U17850 ( .B1(n14280), .B2(n14279), .A(n14282), .ZN(n14281) );
  OAI21_X1 U17851 ( .B1(n14282), .B2(n15379), .A(n14281), .ZN(P1_U3473) );
  INV_X1 U17852 ( .A(n14283), .ZN(n14284) );
  NOR2_X1 U17853 ( .A1(n9692), .A2(n14284), .ZN(n14287) );
  XNOR2_X1 U17854 ( .A(n14287), .B(n10293), .ZN(n14442) );
  AOI21_X1 U17855 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14440) );
  NAND2_X1 U17856 ( .A1(n14440), .A2(n19657), .ZN(n14303) );
  INV_X1 U17857 ( .A(n14291), .ZN(n14292) );
  AOI21_X1 U17858 ( .B1(n14294), .B2(n14293), .A(n14292), .ZN(n15851) );
  OR2_X1 U17859 ( .A1(n12877), .A2(n14295), .ZN(n14296) );
  NAND2_X1 U17860 ( .A1(n9690), .A2(n14296), .ZN(n15962) );
  NOR2_X1 U17861 ( .A1(n15962), .A2(n19648), .ZN(n14301) );
  OAI21_X1 U17862 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n14297), .ZN(n14299) );
  NOR2_X1 U17863 ( .A1(n16032), .A2(n20262), .ZN(n14436) );
  AOI21_X1 U17864 ( .B1(n16337), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14436), .ZN(n14298) );
  OAI21_X1 U17865 ( .B1(n16307), .B2(n14299), .A(n14298), .ZN(n14300) );
  AOI211_X1 U17866 ( .C1(n15851), .C2(n19669), .A(n14301), .B(n14300), .ZN(
        n14302) );
  OAI211_X1 U17867 ( .C1(n14442), .C2(n19653), .A(n14303), .B(n14302), .ZN(
        P2_U3026) );
  MUX2_X2 U17868 ( .A(n14306), .B(n14305), .S(n14304), .Z(n14309) );
  AOI22_X1 U17869 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n14307), .B1(n13376), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14308) );
  OAI22_X1 U17870 ( .A1(n14404), .A2(n14835), .B1(n20452), .B2(n14315), .ZN(
        P1_U2841) );
  AOI22_X1 U17871 ( .A1(n14311), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14310), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17872 ( .A1(n14432), .A2(n13435), .ZN(n14322) );
  OAI22_X1 U17873 ( .A1(n20442), .A2(n14315), .B1(n14314), .B2(n20394), .ZN(
        n14319) );
  INV_X1 U17874 ( .A(n14316), .ZN(n14317) );
  NOR3_X1 U17875 ( .A1(n14453), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14317), 
        .ZN(n14318) );
  AOI211_X1 U17876 ( .C1(n14320), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14319), 
        .B(n14318), .ZN(n14321) );
  OAI211_X1 U17877 ( .C1(n14404), .C2(n20408), .A(n14322), .B(n14321), .ZN(
        P1_U2809) );
  INV_X1 U17878 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14324) );
  OAI222_X1 U17879 ( .A1(n14838), .A2(n14325), .B1(n14324), .B2(n20452), .C1(
        n14835), .C2(n14323), .ZN(P1_U2842) );
  INV_X1 U17880 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14353) );
  NAND2_X1 U17881 ( .A1(n20580), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14354) );
  NAND2_X1 U17882 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14330) );
  OAI211_X1 U17883 ( .C1(n14331), .C2(n20524), .A(n14354), .B(n14330), .ZN(
        n14332) );
  AOI21_X1 U17884 ( .B1(n14839), .B2(n20519), .A(n14332), .ZN(n14333) );
  OAI21_X1 U17885 ( .B1(n14359), .B2(n15151), .A(n14333), .ZN(P1_U2969) );
  AND2_X1 U17886 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U17887 ( .A1(n14335), .A2(n14334), .ZN(n15327) );
  NOR2_X1 U17888 ( .A1(n15327), .A2(n14336), .ZN(n14340) );
  AND2_X1 U17889 ( .A1(n14340), .A2(n14337), .ZN(n15326) );
  INV_X1 U17890 ( .A(n14338), .ZN(n15310) );
  AND2_X1 U17891 ( .A1(n15326), .A2(n15310), .ZN(n15219) );
  INV_X1 U17892 ( .A(n15219), .ZN(n15223) );
  NOR2_X1 U17893 ( .A1(n15223), .A2(n15316), .ZN(n15267) );
  NAND2_X1 U17894 ( .A1(n20553), .A2(n15267), .ZN(n15202) );
  INV_X1 U17895 ( .A(n20541), .ZN(n20526) );
  NOR2_X1 U17896 ( .A1(n14338), .A2(n20526), .ZN(n14339) );
  NAND2_X1 U17897 ( .A1(n14340), .A2(n14339), .ZN(n14346) );
  INV_X1 U17898 ( .A(n14346), .ZN(n15270) );
  NAND3_X1 U17899 ( .A1(n20573), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15270), .ZN(n14341) );
  NAND2_X1 U17900 ( .A1(n15202), .A2(n14341), .ZN(n15280) );
  NAND2_X1 U17901 ( .A1(n9991), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14343) );
  NAND4_X1 U17902 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15272) );
  INV_X1 U17903 ( .A(n15272), .ZN(n14342) );
  NAND2_X1 U17904 ( .A1(n14342), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14345) );
  NOR2_X1 U17905 ( .A1(n14343), .A2(n14345), .ZN(n14344) );
  NAND2_X1 U17906 ( .A1(n15280), .A2(n14344), .ZN(n15210) );
  INV_X1 U17907 ( .A(n15154), .ZN(n15163) );
  NOR3_X1 U17908 ( .A1(n15171), .A2(n14353), .A3(n15163), .ZN(n14401) );
  INV_X1 U17909 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15203) );
  NOR2_X1 U17910 ( .A1(n15316), .A2(n14345), .ZN(n15225) );
  NAND2_X1 U17911 ( .A1(n15219), .A2(n15225), .ZN(n14348) );
  OR3_X1 U17912 ( .A1(n14346), .A2(n14345), .A3(n15316), .ZN(n14347) );
  AOI22_X1 U17913 ( .A1(n20546), .A2(n14348), .B1(n20573), .B2(n14347), .ZN(
        n14349) );
  INV_X1 U17914 ( .A(n15244), .ZN(n15226) );
  NAND2_X1 U17915 ( .A1(n15293), .A2(n15226), .ZN(n14350) );
  NAND2_X1 U17916 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14351) );
  NOR3_X1 U17917 ( .A1(n15179), .A2(n15194), .A3(n15182), .ZN(n14352) );
  NOR2_X1 U17918 ( .A1(n15213), .A2(n15293), .ZN(n14399) );
  NAND2_X1 U17919 ( .A1(n14355), .A2(n14354), .ZN(n14356) );
  OAI21_X1 U17920 ( .B1(n14359), .B2(n20576), .A(n14358), .ZN(P1_U3001) );
  NAND2_X1 U17921 ( .A1(n16314), .A2(n14360), .ZN(n16040) );
  INV_X1 U17922 ( .A(n16039), .ZN(n14361) );
  OAI21_X1 U17923 ( .B1(n16040), .B2(n14361), .A(n16038), .ZN(n16030) );
  INV_X1 U17924 ( .A(n16028), .ZN(n14362) );
  AOI21_X1 U17925 ( .B1(n16030), .B2(n16027), .A(n14362), .ZN(n14364) );
  XNOR2_X1 U17926 ( .A(n14364), .B(n14363), .ZN(n14381) );
  AND2_X1 U17927 ( .A1(n12744), .A2(n14365), .ZN(n15495) );
  OR2_X1 U17928 ( .A1(n15495), .A2(n14366), .ZN(n14367) );
  NAND2_X1 U17929 ( .A1(n19553), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n14373) );
  NAND2_X1 U17930 ( .A1(n19634), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14368) );
  OAI211_X1 U17931 ( .C1(n15479), .C2(n16264), .A(n14373), .B(n14368), .ZN(
        n14370) );
  AOI21_X1 U17932 ( .B1(n14371), .B2(n15493), .A(n9710), .ZN(n15924) );
  INV_X1 U17933 ( .A(n15924), .ZN(n14378) );
  INV_X1 U17934 ( .A(n14372), .ZN(n16287) );
  XNOR2_X1 U17935 ( .A(n16286), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14376) );
  OAI21_X1 U17936 ( .B1(n16283), .B2(n14374), .A(n14373), .ZN(n14375) );
  AOI21_X1 U17937 ( .B1(n16287), .B2(n14376), .A(n14375), .ZN(n14377) );
  OAI21_X1 U17938 ( .B1(n14378), .B2(n19648), .A(n14377), .ZN(n14380) );
  NOR2_X1 U17939 ( .A1(n14382), .A2(n19570), .ZN(n14383) );
  AOI21_X1 U17940 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19570), .A(n14383), .ZN(
        n14384) );
  OAI21_X1 U17941 ( .B1(n14385), .B2(n19571), .A(n14384), .ZN(P2_U2857) );
  INV_X1 U17942 ( .A(n15748), .ZN(n14396) );
  OR2_X1 U17943 ( .A1(n14387), .A2(n14386), .ZN(n19670) );
  AND3_X1 U17944 ( .A1(n19670), .A2(n16263), .A3(n19671), .ZN(n14395) );
  INV_X1 U17945 ( .A(n14388), .ZN(n14389) );
  NAND2_X1 U17946 ( .A1(n14390), .A2(n14389), .ZN(n14391) );
  NAND2_X1 U17947 ( .A1(n14392), .A2(n14391), .ZN(n19667) );
  INV_X1 U17948 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20234) );
  NOR2_X1 U17949 ( .A1(n16032), .A2(n20234), .ZN(n19663) );
  AOI21_X1 U17950 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19663), .ZN(n14393) );
  OAI21_X1 U17951 ( .B1(n19667), .B2(n16253), .A(n14393), .ZN(n14394) );
  AOI211_X1 U17952 ( .C1(n14396), .C2(n16234), .A(n14395), .B(n14394), .ZN(
        n14397) );
  OAI21_X1 U17953 ( .B1(n16572), .B2(n16222), .A(n14397), .ZN(P2_U3012) );
  NAND3_X1 U17954 ( .A1(n14400), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n9946), .ZN(n14403) );
  NAND2_X1 U17955 ( .A1(n20580), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14408) );
  NAND3_X1 U17956 ( .A1(n14401), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14277), .ZN(n14402) );
  OAI21_X1 U17957 ( .B1(n14404), .B2(n20578), .A(n10299), .ZN(n14405) );
  INV_X1 U17958 ( .A(n14405), .ZN(n14406) );
  OAI21_X1 U17959 ( .B1(n14412), .B2(n20576), .A(n14406), .ZN(P1_U3000) );
  NAND2_X1 U17960 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14407) );
  OAI211_X1 U17961 ( .C1(n14409), .C2(n20524), .A(n14408), .B(n14407), .ZN(
        n14410) );
  AOI21_X1 U17962 ( .B1(n14432), .B2(n20519), .A(n14410), .ZN(n14411) );
  OAI21_X1 U17963 ( .B1(n14412), .B2(n15151), .A(n14411), .ZN(P1_U2968) );
  NAND2_X1 U17964 ( .A1(n14413), .A2(n19657), .ZN(n14424) );
  NAND3_X1 U17965 ( .A1(n14415), .A2(n14414), .A3(n19672), .ZN(n14423) );
  NOR2_X1 U17966 ( .A1(n9710), .A2(n14416), .ZN(n14417) );
  OR2_X1 U17967 ( .A1(n15453), .A2(n14417), .ZN(n15467) );
  AOI21_X1 U17968 ( .B1(n16270), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14418), .ZN(n14420) );
  NAND2_X1 U17969 ( .A1(n16272), .A2(n16019), .ZN(n14419) );
  OAI211_X1 U17970 ( .C1(n15467), .C2(n19648), .A(n14420), .B(n14419), .ZN(
        n14421) );
  AOI21_X1 U17971 ( .B1(n15801), .B2(n19669), .A(n14421), .ZN(n14422) );
  OAI211_X1 U17972 ( .C1(n16015), .C2(n14424), .A(n14423), .B(n14422), .ZN(
        P2_U3019) );
  AOI21_X1 U17973 ( .B1(n17060), .B2(n21278), .A(n21281), .ZN(n14428) );
  INV_X1 U17974 ( .A(n17056), .ZN(n21276) );
  AOI22_X1 U17975 ( .A1(n10782), .A2(n15386), .B1(n14425), .B2(n10429), .ZN(
        n17061) );
  OAI21_X1 U17976 ( .B1(n17061), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n15388), 
        .ZN(n14426) );
  AOI22_X1 U17977 ( .A1(n21276), .A2(n10429), .B1(n14426), .B2(n15417), .ZN(
        n14427) );
  OAI22_X1 U17978 ( .A1(n14428), .A2(n10429), .B1(n21281), .B2(n14427), .ZN(
        P1_U3474) );
  OR2_X1 U17979 ( .A1(n14935), .A2(n14429), .ZN(n14433) );
  INV_X1 U17980 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20645) );
  AOI22_X1 U17981 ( .A1(n14912), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14935), .ZN(n14434) );
  OAI211_X1 U17982 ( .C1(n14915), .C2(n20645), .A(n14435), .B(n14434), .ZN(
        P1_U2873) );
  NAND2_X1 U17983 ( .A1(n15851), .A2(n19642), .ZN(n14438) );
  AOI21_X1 U17984 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14436), .ZN(n14437) );
  OAI211_X1 U17985 ( .C1(n16264), .C2(n15571), .A(n14438), .B(n14437), .ZN(
        n14439) );
  AOI21_X1 U17986 ( .B1(n14440), .B2(n19636), .A(n14439), .ZN(n14441) );
  OAI21_X1 U17987 ( .B1(n19640), .B2(n14442), .A(n14441), .ZN(P2_U2994) );
  INV_X1 U17988 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20628) );
  NOR2_X1 U17989 ( .A1(n14444), .A2(n20629), .ZN(n14445) );
  AOI22_X1 U17990 ( .A1(n14911), .A2(n14924), .B1(n14935), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U17991 ( .A1(n14912), .A2(DATAI_29_), .ZN(n14446) );
  OAI211_X1 U17992 ( .C1(n14915), .C2(n20628), .A(n14447), .B(n14446), .ZN(
        n14448) );
  INV_X1 U17993 ( .A(n14448), .ZN(n14449) );
  OAI21_X1 U17994 ( .B1(n14443), .B2(n14938), .A(n14449), .ZN(P1_U2875) );
  NOR2_X1 U17995 ( .A1(n14798), .A2(n14450), .ZN(n14473) );
  NAND2_X1 U17996 ( .A1(n14473), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U17997 ( .A1(n20411), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20430), .ZN(n14451) );
  OAI211_X1 U17998 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14453), .A(n14452), 
        .B(n14451), .ZN(n14456) );
  XNOR2_X1 U17999 ( .A(n14472), .B(n14454), .ZN(n15153) );
  NOR2_X1 U18000 ( .A1(n15153), .A2(n20408), .ZN(n14455) );
  AOI211_X1 U18001 ( .C1(n14457), .C2(n20426), .A(n14456), .B(n14455), .ZN(
        n14458) );
  OAI21_X1 U18002 ( .B1(n14443), .B2(n14772), .A(n14458), .ZN(P1_U2811) );
  OAI222_X1 U18003 ( .A1(n14443), .A2(n14838), .B1(n14459), .B2(n20452), .C1(
        n14835), .C2(n15153), .ZN(P1_U2843) );
  AOI22_X1 U18004 ( .A1(n15984), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n16010), .ZN(n14461) );
  NAND2_X1 U18005 ( .A1(n15983), .A2(BUF1_REG_31__SCAN_IN), .ZN(n14460) );
  OAI211_X1 U18006 ( .C1(n14462), .C2(n15981), .A(n14461), .B(n14460), .ZN(
        P2_U2888) );
  NAND2_X1 U18007 ( .A1(n19570), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14464) );
  OAI21_X1 U18008 ( .B1(n14463), .B2(n19570), .A(n14464), .ZN(P2_U2856) );
  MUX2_X1 U18009 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n14465), .Z(P1_U3486) );
  AOI21_X1 U18010 ( .B1(n14468), .B2(n14480), .A(n14467), .ZN(n14950) );
  INV_X1 U18011 ( .A(n14950), .ZN(n14805) );
  NOR2_X1 U18012 ( .A1(n14469), .A2(n14483), .ZN(n14482) );
  NOR2_X1 U18013 ( .A1(n14482), .A2(n14470), .ZN(n14471) );
  OR2_X1 U18014 ( .A1(n14472), .A2(n14471), .ZN(n14803) );
  INV_X1 U18015 ( .A(n14803), .ZN(n15167) );
  AOI22_X1 U18016 ( .A1(n20411), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20430), .ZN(n14476) );
  INV_X1 U18017 ( .A(n14489), .ZN(n14486) );
  NOR3_X1 U18018 ( .A1(n20392), .A2(n21269), .A3(n14486), .ZN(n14474) );
  OAI21_X1 U18019 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14474), .A(n14473), 
        .ZN(n14475) );
  OAI211_X1 U18020 ( .C1(n20402), .C2(n14948), .A(n14476), .B(n14475), .ZN(
        n14477) );
  AOI21_X1 U18021 ( .B1(n15167), .B2(n20425), .A(n14477), .ZN(n14478) );
  OAI21_X1 U18022 ( .B1(n14805), .B2(n14772), .A(n14478), .ZN(P1_U2812) );
  OAI21_X1 U18023 ( .B1(n14479), .B2(n14481), .A(n14480), .ZN(n14852) );
  AOI21_X1 U18024 ( .B1(n14483), .B2(n14469), .A(n14482), .ZN(n15175) );
  INV_X1 U18025 ( .A(n14484), .ZN(n14958) );
  NOR2_X1 U18026 ( .A1(n20394), .A2(n14485), .ZN(n14488) );
  NOR3_X1 U18027 ( .A1(n20392), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14486), 
        .ZN(n14487) );
  AOI211_X1 U18028 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20411), .A(n14488), .B(
        n14487), .ZN(n14491) );
  OAI21_X1 U18029 ( .B1(n20392), .B2(n14489), .A(n20428), .ZN(n14501) );
  NAND2_X1 U18030 ( .A1(n14501), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14490) );
  OAI211_X1 U18031 ( .C1(n20402), .C2(n14958), .A(n14491), .B(n14490), .ZN(
        n14492) );
  AOI21_X1 U18032 ( .B1(n15175), .B2(n20425), .A(n14492), .ZN(n14493) );
  OAI21_X1 U18033 ( .B1(n14852), .B2(n14772), .A(n14493), .ZN(P1_U2813) );
  AOI21_X1 U18034 ( .B1(n14495), .B2(n14494), .A(n14479), .ZN(n14971) );
  INV_X1 U18035 ( .A(n14971), .ZN(n14809) );
  NAND2_X1 U18036 ( .A1(n14496), .A2(n14497), .ZN(n14498) );
  NAND2_X1 U18037 ( .A1(n14469), .A2(n14498), .ZN(n14807) );
  INV_X1 U18038 ( .A(n14807), .ZN(n15187) );
  AOI22_X1 U18039 ( .A1(n20411), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20430), .ZN(n14504) );
  NAND2_X1 U18040 ( .A1(n20433), .A2(n14514), .ZN(n14530) );
  INV_X1 U18041 ( .A(n14499), .ZN(n14500) );
  NOR2_X1 U18042 ( .A1(n14530), .A2(n14500), .ZN(n14502) );
  OAI21_X1 U18043 ( .B1(n14502), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14501), 
        .ZN(n14503) );
  OAI211_X1 U18044 ( .C1(n20402), .C2(n14969), .A(n14504), .B(n14503), .ZN(
        n14505) );
  AOI21_X1 U18045 ( .B1(n15187), .B2(n20425), .A(n14505), .ZN(n14506) );
  OAI21_X1 U18046 ( .B1(n14809), .B2(n14772), .A(n14506), .ZN(P1_U2814) );
  OAI21_X1 U18047 ( .B1(n14526), .B2(n14510), .A(n14494), .ZN(n14865) );
  OAI21_X1 U18048 ( .B1(n14511), .B2(n14512), .A(n14496), .ZN(n14811) );
  INV_X1 U18049 ( .A(n14811), .ZN(n15197) );
  INV_X1 U18050 ( .A(n14513), .ZN(n14979) );
  INV_X1 U18051 ( .A(n14514), .ZN(n14515) );
  OAI21_X1 U18052 ( .B1(n20399), .B2(n14515), .A(n20397), .ZN(n14541) );
  OAI21_X1 U18053 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20392), .A(n14541), 
        .ZN(n14519) );
  INV_X1 U18054 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14810) );
  INV_X1 U18055 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14516) );
  OAI22_X1 U18056 ( .A1(n20442), .A2(n14810), .B1(n14516), .B2(n20394), .ZN(
        n14518) );
  NOR3_X1 U18057 ( .A1(n14530), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14983), 
        .ZN(n14517) );
  AOI211_X1 U18058 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14519), .A(n14518), 
        .B(n14517), .ZN(n14520) );
  OAI21_X1 U18059 ( .B1(n14979), .B2(n20402), .A(n14520), .ZN(n14521) );
  AOI21_X1 U18060 ( .B1(n15197), .B2(n20425), .A(n14521), .ZN(n14522) );
  OAI21_X1 U18061 ( .B1(n14865), .B2(n14772), .A(n14522), .ZN(P1_U2815) );
  AND2_X1 U18062 ( .A1(n14545), .A2(n14523), .ZN(n14524) );
  OR2_X1 U18063 ( .A1(n14524), .A2(n14511), .ZN(n15209) );
  NOR2_X1 U18064 ( .A1(n14551), .A2(n14525), .ZN(n14536) );
  INV_X1 U18065 ( .A(n14526), .ZN(n14527) );
  OAI21_X1 U18066 ( .B1(n14528), .B2(n14536), .A(n14527), .ZN(n14991) );
  INV_X1 U18067 ( .A(n14991), .ZN(n14877) );
  NAND2_X1 U18068 ( .A1(n14877), .A2(n13435), .ZN(n14535) );
  INV_X1 U18069 ( .A(n14541), .ZN(n14533) );
  AOI22_X1 U18070 ( .A1(n20411), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20430), .ZN(n14529) );
  OAI21_X1 U18071 ( .B1(n14530), .B2(P1_REIP_REG_24__SCAN_IN), .A(n14529), 
        .ZN(n14532) );
  NOR2_X1 U18072 ( .A1(n20402), .A2(n14984), .ZN(n14531) );
  AOI211_X1 U18073 ( .C1(n14533), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14532), 
        .B(n14531), .ZN(n14534) );
  OAI211_X1 U18074 ( .C1(n15209), .C2(n20408), .A(n14535), .B(n14534), .ZN(
        P1_U2816) );
  AOI21_X1 U18075 ( .B1(n14537), .B2(n14549), .A(n14536), .ZN(n14999) );
  INV_X1 U18076 ( .A(n14999), .ZN(n14814) );
  AOI21_X1 U18077 ( .B1(n20433), .B2(n14538), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14540) );
  AOI22_X1 U18078 ( .A1(n20411), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20430), .ZN(n14539) );
  OAI21_X1 U18079 ( .B1(n14541), .B2(n14540), .A(n14539), .ZN(n14547) );
  NAND2_X1 U18080 ( .A1(n14554), .A2(n14543), .ZN(n14544) );
  NAND2_X1 U18081 ( .A1(n14545), .A2(n14544), .ZN(n15214) );
  NOR2_X1 U18082 ( .A1(n15214), .A2(n20408), .ZN(n14546) );
  AOI211_X1 U18083 ( .C1(n20426), .C2(n14994), .A(n14547), .B(n14546), .ZN(
        n14548) );
  OAI21_X1 U18084 ( .B1(n14814), .B2(n14772), .A(n14548), .ZN(P1_U2817) );
  INV_X1 U18085 ( .A(n14549), .ZN(n14550) );
  AOI21_X1 U18086 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n15007) );
  INV_X1 U18087 ( .A(n15007), .ZN(n14816) );
  AOI21_X1 U18088 ( .B1(n14555), .B2(n14553), .A(n14542), .ZN(n15231) );
  MUX2_X1 U18089 ( .A(n14556), .B(P1_REIP_REG_21__SCAN_IN), .S(
        P1_REIP_REG_22__SCAN_IN), .Z(n14557) );
  OAI22_X1 U18090 ( .A1(n14558), .A2(n20394), .B1(n20392), .B2(n14557), .ZN(
        n14560) );
  AOI21_X1 U18091 ( .B1(n20433), .B2(n14572), .A(n20399), .ZN(n14587) );
  NOR2_X1 U18092 ( .A1(n14587), .A2(n21264), .ZN(n14559) );
  AOI211_X1 U18093 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n20411), .A(n14560), .B(
        n14559), .ZN(n14561) );
  OAI21_X1 U18094 ( .B1(n15005), .B2(n20402), .A(n14561), .ZN(n14562) );
  AOI21_X1 U18095 ( .B1(n15231), .B2(n20425), .A(n14562), .ZN(n14563) );
  OAI21_X1 U18096 ( .B1(n14816), .B2(n14772), .A(n14563), .ZN(P1_U2818) );
  OAI21_X1 U18097 ( .B1(n14564), .B2(n14565), .A(n14553), .ZN(n15238) );
  INV_X1 U18098 ( .A(n14566), .ZN(n14615) );
  INV_X1 U18099 ( .A(n14582), .ZN(n14567) );
  NAND2_X1 U18100 ( .A1(n14595), .A2(n14567), .ZN(n14579) );
  INV_X1 U18101 ( .A(n14568), .ZN(n14570) );
  NAND2_X1 U18102 ( .A1(n15018), .A2(n13435), .ZN(n14578) );
  NOR2_X1 U18103 ( .A1(n20394), .A2(n14571), .ZN(n14574) );
  NOR3_X1 U18104 ( .A1(n20392), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14572), 
        .ZN(n14573) );
  AOI211_X1 U18105 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n20411), .A(n14574), .B(
        n14573), .ZN(n14575) );
  OAI21_X1 U18106 ( .B1(n14587), .B2(n15014), .A(n14575), .ZN(n14576) );
  AOI21_X1 U18107 ( .B1(n15013), .B2(n20426), .A(n14576), .ZN(n14577) );
  OAI211_X1 U18108 ( .C1(n15238), .C2(n20408), .A(n14578), .B(n14577), .ZN(
        P1_U2819) );
  INV_X1 U18109 ( .A(n14595), .ZN(n14581) );
  INV_X1 U18110 ( .A(n14579), .ZN(n14580) );
  AOI21_X1 U18111 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n15027) );
  INV_X1 U18112 ( .A(n15027), .ZN(n14820) );
  NOR2_X1 U18113 ( .A1(n9723), .A2(n14583), .ZN(n14584) );
  OR2_X1 U18114 ( .A1(n14564), .A2(n14584), .ZN(n15252) );
  INV_X1 U18115 ( .A(n15252), .ZN(n14593) );
  AOI22_X1 U18116 ( .A1(n20411), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20430), .ZN(n14591) );
  NOR3_X1 U18117 ( .A1(n20392), .A2(n14586), .A3(n14585), .ZN(n14589) );
  INV_X1 U18118 ( .A(n14587), .ZN(n14588) );
  OAI21_X1 U18119 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n14589), .A(n14588), 
        .ZN(n14590) );
  OAI211_X1 U18120 ( .C1(n20402), .C2(n15025), .A(n14591), .B(n14590), .ZN(
        n14592) );
  AOI21_X1 U18121 ( .B1(n14593), .B2(n20425), .A(n14592), .ZN(n14594) );
  OAI21_X1 U18122 ( .B1(n14820), .B2(n14772), .A(n14594), .ZN(P1_U2820) );
  AOI21_X1 U18123 ( .B1(n14596), .B2(n14614), .A(n14595), .ZN(n15035) );
  INV_X1 U18124 ( .A(n15035), .ZN(n14822) );
  AOI21_X1 U18125 ( .B1(n14597), .B2(n14618), .A(n9723), .ZN(n15261) );
  INV_X1 U18126 ( .A(n14598), .ZN(n14693) );
  NOR2_X1 U18127 ( .A1(n20399), .A2(n14693), .ZN(n14599) );
  OR2_X1 U18128 ( .A1(n14798), .A2(n14599), .ZN(n14692) );
  OAI21_X1 U18129 ( .B1(n14798), .B2(n14600), .A(n14692), .ZN(n14681) );
  AOI21_X1 U18130 ( .B1(n20397), .B2(n14601), .A(n14681), .ZN(n14639) );
  OR3_X1 U18131 ( .A1(n20392), .A2(n15105), .A3(n14693), .ZN(n14680) );
  NAND2_X1 U18132 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n14602) );
  NOR2_X1 U18133 ( .A1(n14680), .A2(n14602), .ZN(n14650) );
  NOR2_X1 U18134 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14605), .ZN(n14603) );
  NAND2_X1 U18135 ( .A1(n14650), .A2(n14603), .ZN(n14621) );
  AOI21_X1 U18136 ( .B1(n14639), .B2(n14621), .A(n15031), .ZN(n14612) );
  INV_X1 U18137 ( .A(n14604), .ZN(n15033) );
  NOR3_X1 U18138 ( .A1(n21262), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n14605), 
        .ZN(n14609) );
  NAND2_X1 U18139 ( .A1(n20411), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14606) );
  OAI211_X1 U18140 ( .C1(n20394), .C2(n14607), .A(n14606), .B(n20416), .ZN(
        n14608) );
  AOI21_X1 U18141 ( .B1(n14650), .B2(n14609), .A(n14608), .ZN(n14610) );
  OAI21_X1 U18142 ( .B1(n20402), .B2(n15033), .A(n14610), .ZN(n14611) );
  AOI211_X1 U18143 ( .C1(n15261), .C2(n20425), .A(n14612), .B(n14611), .ZN(
        n14613) );
  OAI21_X1 U18144 ( .B1(n14822), .B2(n14772), .A(n14613), .ZN(P1_U2821) );
  OAI21_X1 U18145 ( .B1(n14629), .B2(n14615), .A(n14614), .ZN(n15044) );
  INV_X1 U18146 ( .A(n14616), .ZN(n14619) );
  OAI21_X1 U18147 ( .B1(n14619), .B2(n10130), .A(n14618), .ZN(n15279) );
  INV_X1 U18148 ( .A(n15279), .ZN(n14625) );
  NOR2_X1 U18149 ( .A1(n14639), .A2(n21262), .ZN(n14624) );
  INV_X1 U18150 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21444) );
  NOR2_X1 U18151 ( .A1(n20442), .A2(n21444), .ZN(n14620) );
  AOI211_X1 U18152 ( .C1(n20430), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20580), .B(n14620), .ZN(n14622) );
  OAI211_X1 U18153 ( .C1(n20402), .C2(n15040), .A(n14622), .B(n14621), .ZN(
        n14623) );
  AOI211_X1 U18154 ( .C1(n14625), .C2(n20425), .A(n14624), .B(n14623), .ZN(
        n14626) );
  OAI21_X1 U18155 ( .B1(n15044), .B2(n14772), .A(n14626), .ZN(P1_U2822) );
  NAND2_X1 U18156 ( .A1(n14690), .A2(n14670), .ZN(n14671) );
  INV_X1 U18157 ( .A(n14627), .ZN(n14656) );
  NAND2_X1 U18158 ( .A1(n14655), .A2(n14643), .ZN(n14642) );
  INV_X1 U18159 ( .A(n14628), .ZN(n14630) );
  AOI21_X1 U18160 ( .B1(n14642), .B2(n14630), .A(n14629), .ZN(n15063) );
  INV_X1 U18161 ( .A(n15063), .ZN(n14825) );
  OAI21_X1 U18162 ( .B1(n14631), .B2(n14632), .A(n14616), .ZN(n14823) );
  INV_X1 U18163 ( .A(n14823), .ZN(n15286) );
  AOI21_X1 U18164 ( .B1(n14650), .B2(P1_REIP_REG_16__SCAN_IN), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14638) );
  INV_X1 U18165 ( .A(n15061), .ZN(n14636) );
  NAND2_X1 U18166 ( .A1(n20411), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14633) );
  OAI211_X1 U18167 ( .C1(n20394), .C2(n14634), .A(n14633), .B(n20416), .ZN(
        n14635) );
  AOI21_X1 U18168 ( .B1(n20426), .B2(n14636), .A(n14635), .ZN(n14637) );
  OAI21_X1 U18169 ( .B1(n14639), .B2(n14638), .A(n14637), .ZN(n14640) );
  AOI21_X1 U18170 ( .B1(n15286), .B2(n20425), .A(n14640), .ZN(n14641) );
  OAI21_X1 U18171 ( .B1(n14825), .B2(n14772), .A(n14641), .ZN(P1_U2823) );
  OAI21_X1 U18172 ( .B1(n14655), .B2(n14643), .A(n14642), .ZN(n14910) );
  INV_X1 U18173 ( .A(n14644), .ZN(n14658) );
  AOI21_X1 U18174 ( .B1(n14645), .B2(n14658), .A(n14631), .ZN(n15292) );
  INV_X1 U18175 ( .A(n14646), .ZN(n15072) );
  NAND2_X1 U18176 ( .A1(n15083), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14647) );
  NOR2_X1 U18177 ( .A1(n14680), .A2(n14647), .ZN(n14663) );
  OAI21_X1 U18178 ( .B1(n14681), .B2(n14663), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14652) );
  NAND2_X1 U18179 ( .A1(n20411), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n14648) );
  OAI211_X1 U18180 ( .C1(n20394), .C2(n21437), .A(n14648), .B(n20416), .ZN(
        n14649) );
  AOI21_X1 U18181 ( .B1(n14650), .B2(n15070), .A(n14649), .ZN(n14651) );
  OAI211_X1 U18182 ( .C1(n20402), .C2(n15072), .A(n14652), .B(n14651), .ZN(
        n14653) );
  AOI21_X1 U18183 ( .B1(n15292), .B2(n20425), .A(n14653), .ZN(n14654) );
  OAI21_X1 U18184 ( .B1(n14910), .B2(n14772), .A(n14654), .ZN(P1_U2824) );
  AOI21_X1 U18185 ( .B1(n14656), .B2(n14671), .A(n14655), .ZN(n15087) );
  INV_X1 U18186 ( .A(n15087), .ZN(n14921) );
  INV_X1 U18187 ( .A(n14657), .ZN(n14660) );
  OAI21_X1 U18188 ( .B1(n14660), .B2(n14659), .A(n14658), .ZN(n14827) );
  INV_X1 U18189 ( .A(n14827), .ZN(n15300) );
  INV_X1 U18190 ( .A(n14681), .ZN(n14667) );
  INV_X1 U18191 ( .A(n15085), .ZN(n14665) );
  NAND2_X1 U18192 ( .A1(n20411), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n14661) );
  OAI211_X1 U18193 ( .C1(n20394), .C2(n14662), .A(n14661), .B(n20416), .ZN(
        n14664) );
  AOI211_X1 U18194 ( .C1(n20426), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14666) );
  OAI21_X1 U18195 ( .B1(n14667), .B2(n15083), .A(n14666), .ZN(n14668) );
  AOI21_X1 U18196 ( .B1(n15300), .B2(n20425), .A(n14668), .ZN(n14669) );
  OAI21_X1 U18197 ( .B1(n14921), .B2(n14772), .A(n14669), .ZN(P1_U2825) );
  INV_X1 U18198 ( .A(n14670), .ZN(n14674) );
  INV_X1 U18199 ( .A(n14690), .ZN(n14673) );
  INV_X1 U18200 ( .A(n14671), .ZN(n14672) );
  AOI21_X1 U18201 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(n15096) );
  INV_X1 U18202 ( .A(n15096), .ZN(n14923) );
  NAND2_X1 U18203 ( .A1(n14704), .A2(n14687), .ZN(n14677) );
  INV_X1 U18204 ( .A(n14675), .ZN(n14676) );
  NAND2_X1 U18205 ( .A1(n14677), .A2(n14676), .ZN(n14678) );
  NAND2_X1 U18206 ( .A1(n14678), .A2(n14657), .ZN(n14829) );
  INV_X1 U18207 ( .A(n14829), .ZN(n15308) );
  INV_X1 U18208 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14830) );
  NOR2_X1 U18209 ( .A1(n20442), .A2(n14830), .ZN(n14679) );
  AOI211_X1 U18210 ( .C1(n20430), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20580), .B(n14679), .ZN(n14684) );
  INV_X1 U18211 ( .A(n14680), .ZN(n14682) );
  OAI21_X1 U18212 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14682), .A(n14681), 
        .ZN(n14683) );
  OAI211_X1 U18213 ( .C1(n20402), .C2(n15094), .A(n14684), .B(n14683), .ZN(
        n14685) );
  AOI21_X1 U18214 ( .B1(n20425), .B2(n15308), .A(n14685), .ZN(n14686) );
  OAI21_X1 U18215 ( .B1(n14923), .B2(n14772), .A(n14686), .ZN(P1_U2826) );
  XNOR2_X1 U18216 ( .A(n14704), .B(n14687), .ZN(n15321) );
  OAI21_X1 U18217 ( .B1(n9670), .B2(n10303), .A(n14688), .ZN(n14716) );
  OAI21_X1 U18218 ( .B1(n14716), .B2(n14717), .A(n14688), .ZN(n14702) );
  NAND2_X1 U18219 ( .A1(n14702), .A2(n14701), .ZN(n14700) );
  INV_X1 U18220 ( .A(n14689), .ZN(n14691) );
  AOI21_X1 U18221 ( .B1(n14700), .B2(n14691), .A(n14690), .ZN(n15109) );
  NAND2_X1 U18222 ( .A1(n15109), .A2(n13435), .ZN(n14699) );
  INV_X1 U18223 ( .A(n14692), .ZN(n14710) );
  NOR2_X1 U18224 ( .A1(n20402), .A2(n15107), .ZN(n14697) );
  INV_X1 U18225 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14831) );
  NOR3_X1 U18226 ( .A1(n20392), .A2(P1_REIP_REG_13__SCAN_IN), .A3(n14693), 
        .ZN(n14694) );
  AOI211_X1 U18227 ( .C1(n20430), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20580), .B(n14694), .ZN(n14695) );
  OAI21_X1 U18228 ( .B1(n20442), .B2(n14831), .A(n14695), .ZN(n14696) );
  AOI211_X1 U18229 ( .C1(n14710), .C2(P1_REIP_REG_13__SCAN_IN), .A(n14697), 
        .B(n14696), .ZN(n14698) );
  OAI211_X1 U18230 ( .C1(n15321), .C2(n20408), .A(n14699), .B(n14698), .ZN(
        P1_U2827) );
  OAI21_X1 U18231 ( .B1(n14702), .B2(n14701), .A(n14700), .ZN(n15121) );
  INV_X1 U18232 ( .A(n14719), .ZN(n14734) );
  AOI21_X1 U18233 ( .B1(n14734), .B2(n14718), .A(n14703), .ZN(n14705) );
  OR2_X1 U18234 ( .A1(n14705), .A2(n14704), .ZN(n15335) );
  OR2_X1 U18235 ( .A1(n20392), .A2(n14720), .ZN(n14723) );
  OAI21_X1 U18236 ( .B1(n14723), .B2(n15125), .A(n14706), .ZN(n14709) );
  NAND2_X1 U18237 ( .A1(n20411), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n14707) );
  OAI211_X1 U18238 ( .C1(n20394), .C2(n15111), .A(n14707), .B(n20416), .ZN(
        n14708) );
  AOI21_X1 U18239 ( .B1(n14710), .B2(n14709), .A(n14708), .ZN(n14713) );
  INV_X1 U18240 ( .A(n14711), .ZN(n15118) );
  NAND2_X1 U18241 ( .A1(n20426), .A2(n15118), .ZN(n14712) );
  OAI211_X1 U18242 ( .C1(n15335), .C2(n20408), .A(n14713), .B(n14712), .ZN(
        n14714) );
  INV_X1 U18243 ( .A(n14714), .ZN(n14715) );
  OAI21_X1 U18244 ( .B1(n15121), .B2(n14772), .A(n14715), .ZN(P1_U2828) );
  XOR2_X1 U18245 ( .A(n14717), .B(n14716), .Z(n15129) );
  INV_X1 U18246 ( .A(n15129), .ZN(n14929) );
  XNOR2_X1 U18247 ( .A(n14719), .B(n14718), .ZN(n15345) );
  NAND2_X1 U18248 ( .A1(n20433), .A2(n14720), .ZN(n14737) );
  NAND2_X1 U18249 ( .A1(n14737), .A2(n20428), .ZN(n14731) );
  AOI21_X1 U18250 ( .B1(n20430), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20580), .ZN(n14722) );
  NAND2_X1 U18251 ( .A1(n20411), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n14721) );
  OAI211_X1 U18252 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n14723), .A(n14722), 
        .B(n14721), .ZN(n14724) );
  AOI21_X1 U18253 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n14731), .A(n14724), 
        .ZN(n14725) );
  OAI21_X1 U18254 ( .B1(n15127), .B2(n20402), .A(n14725), .ZN(n14726) );
  AOI21_X1 U18255 ( .B1(n20425), .B2(n15345), .A(n14726), .ZN(n14727) );
  OAI21_X1 U18256 ( .B1(n14929), .B2(n14772), .A(n14727), .ZN(P1_U2829) );
  INV_X1 U18257 ( .A(n14729), .ZN(n14730) );
  AOI21_X1 U18258 ( .B1(n10119), .B2(n14730), .A(n9670), .ZN(n15142) );
  INV_X1 U18259 ( .A(n15142), .ZN(n14934) );
  INV_X1 U18260 ( .A(n15140), .ZN(n14741) );
  NAND2_X1 U18261 ( .A1(n14731), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n14732) );
  OAI211_X1 U18262 ( .C1(n20394), .C2(n14733), .A(n14732), .B(n20416), .ZN(
        n14740) );
  AOI21_X1 U18263 ( .B1(n14735), .B2(n14233), .A(n14734), .ZN(n15355) );
  AOI22_X1 U18264 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n20411), .B1(n20425), 
        .B2(n15355), .ZN(n14736) );
  OAI21_X1 U18265 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14739) );
  AOI211_X1 U18266 ( .C1(n20426), .C2(n14741), .A(n14740), .B(n14739), .ZN(
        n14742) );
  OAI21_X1 U18267 ( .B1(n14934), .B2(n14772), .A(n14742), .ZN(P1_U2830) );
  INV_X1 U18268 ( .A(n14743), .ZN(n14745) );
  INV_X1 U18269 ( .A(n14239), .ZN(n14744) );
  AOI21_X1 U18270 ( .B1(n14745), .B2(n14744), .A(n14729), .ZN(n15149) );
  INV_X1 U18271 ( .A(n15149), .ZN(n14939) );
  INV_X1 U18272 ( .A(n15147), .ZN(n14755) );
  OAI21_X1 U18273 ( .B1(n20394), .B2(n14746), .A(n20416), .ZN(n14749) );
  NAND2_X1 U18274 ( .A1(n20433), .A2(n14750), .ZN(n14747) );
  OAI22_X1 U18275 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n14747), .B1(n20408), 
        .B2(n14836), .ZN(n14748) );
  AOI211_X1 U18276 ( .C1(n20411), .C2(P1_EBX_REG_9__SCAN_IN), .A(n14749), .B(
        n14748), .ZN(n14753) );
  OR2_X1 U18277 ( .A1(n20392), .A2(n14750), .ZN(n14751) );
  NAND2_X1 U18278 ( .A1(n14751), .A2(n20428), .ZN(n14759) );
  NAND2_X1 U18279 ( .A1(n14759), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14752) );
  NAND2_X1 U18280 ( .A1(n14753), .A2(n14752), .ZN(n14754) );
  AOI21_X1 U18281 ( .B1(n14755), .B2(n20426), .A(n14754), .ZN(n14756) );
  OAI21_X1 U18282 ( .B1(n14939), .B2(n14772), .A(n14756), .ZN(P1_U2831) );
  INV_X1 U18283 ( .A(n14757), .ZN(n14767) );
  NAND3_X1 U18284 ( .A1(n20433), .A2(n20383), .A3(P1_REIP_REG_6__SCAN_IN), 
        .ZN(n20382) );
  OAI21_X1 U18285 ( .B1(n20381), .B2(n20382), .A(n21260), .ZN(n14758) );
  NAND2_X1 U18286 ( .A1(n14759), .A2(n14758), .ZN(n14765) );
  NAND2_X1 U18287 ( .A1(n20411), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n14764) );
  INV_X1 U18288 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14761) );
  OAI22_X1 U18289 ( .A1(n14761), .A2(n20394), .B1(n20408), .B2(n14760), .ZN(
        n14762) );
  INV_X1 U18290 ( .A(n14762), .ZN(n14763) );
  NAND4_X1 U18291 ( .A1(n14765), .A2(n20416), .A3(n14764), .A4(n14763), .ZN(
        n14766) );
  AOI21_X1 U18292 ( .B1(n14767), .B2(n20426), .A(n14766), .ZN(n14768) );
  OAI21_X1 U18293 ( .B1(n14769), .B2(n14772), .A(n14768), .ZN(P1_U2832) );
  NAND2_X1 U18294 ( .A1(n14779), .A2(n14770), .ZN(n14771) );
  NAND2_X1 U18295 ( .A1(n14772), .A2(n14771), .ZN(n20419) );
  OAI22_X1 U18296 ( .A1(n14773), .A2(n20394), .B1(n20408), .B2(n20535), .ZN(
        n14775) );
  NAND2_X1 U18297 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14776) );
  NOR3_X1 U18298 ( .A1(n20392), .A2(P1_REIP_REG_3__SCAN_IN), .A3(n14776), .ZN(
        n14774) );
  AOI211_X1 U18299 ( .C1(n20411), .C2(P1_EBX_REG_3__SCAN_IN), .A(n14775), .B(
        n14774), .ZN(n14782) );
  INV_X1 U18300 ( .A(n14776), .ZN(n14777) );
  OAI21_X1 U18301 ( .B1(n20392), .B2(n14777), .A(n20428), .ZN(n14780) );
  NAND2_X1 U18302 ( .A1(n14779), .A2(n14778), .ZN(n20413) );
  INV_X1 U18303 ( .A(n20413), .ZN(n20431) );
  AOI22_X1 U18304 ( .A1(n14780), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20431), 
        .B2(n20893), .ZN(n14781) );
  OAI211_X1 U18305 ( .C1(n14783), .C2(n20402), .A(n14782), .B(n14781), .ZN(
        n14784) );
  AOI21_X1 U18306 ( .B1(n14785), .B2(n20419), .A(n14784), .ZN(n14786) );
  INV_X1 U18307 ( .A(n14786), .ZN(P1_U2837) );
  INV_X1 U18308 ( .A(n20419), .ZN(n20436) );
  AOI22_X1 U18309 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20411), .B1(n20399), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14788) );
  NAND2_X1 U18310 ( .A1(n20430), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14787) );
  OAI211_X1 U18311 ( .C1(n20413), .C2(n14172), .A(n14788), .B(n14787), .ZN(
        n14791) );
  NAND2_X1 U18312 ( .A1(n20425), .A2(n13768), .ZN(n14789) );
  OR2_X1 U18313 ( .A1(n20392), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20429) );
  NAND2_X1 U18314 ( .A1(n14789), .A2(n20429), .ZN(n14790) );
  AOI211_X1 U18315 ( .C1(n20426), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14793) );
  OAI21_X1 U18316 ( .B1(n20436), .B2(n14794), .A(n14793), .ZN(P1_U2839) );
  NAND2_X1 U18317 ( .A1(n20402), .A2(n20394), .ZN(n14800) );
  AOI22_X1 U18318 ( .A1(n20431), .A2(n10782), .B1(n20411), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n14797) );
  INV_X1 U18319 ( .A(n20577), .ZN(n14795) );
  NAND2_X1 U18320 ( .A1(n20425), .A2(n14795), .ZN(n14796) );
  OAI211_X1 U18321 ( .C1(n14798), .C2(n14073), .A(n14797), .B(n14796), .ZN(
        n14799) );
  AOI21_X1 U18322 ( .B1(n14800), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n14799), .ZN(n14801) );
  OAI21_X1 U18323 ( .B1(n20436), .B2(n14802), .A(n14801), .ZN(P1_U2840) );
  INV_X1 U18324 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14804) );
  OAI222_X1 U18325 ( .A1(n14838), .A2(n14805), .B1(n14804), .B2(n20452), .C1(
        n14803), .C2(n14835), .ZN(P1_U2844) );
  INV_X1 U18326 ( .A(n20452), .ZN(n14833) );
  AOI22_X1 U18327 ( .A1(n15175), .A2(n20448), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14833), .ZN(n14806) );
  OAI21_X1 U18328 ( .B1(n14852), .B2(n14838), .A(n14806), .ZN(P1_U2845) );
  INV_X1 U18329 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14808) );
  OAI222_X1 U18330 ( .A1(n14809), .A2(n14838), .B1(n14808), .B2(n20452), .C1(
        n14807), .C2(n14835), .ZN(P1_U2846) );
  OAI222_X1 U18331 ( .A1(n14835), .A2(n14811), .B1(n14810), .B2(n20452), .C1(
        n14865), .C2(n14838), .ZN(P1_U2847) );
  INV_X1 U18332 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14812) );
  OAI222_X1 U18333 ( .A1(n14838), .A2(n14991), .B1(n14812), .B2(n20452), .C1(
        n15209), .C2(n14835), .ZN(P1_U2848) );
  INV_X1 U18334 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14813) );
  OAI222_X1 U18335 ( .A1(n14814), .A2(n14838), .B1(n14813), .B2(n20452), .C1(
        n15214), .C2(n14835), .ZN(P1_U2849) );
  AOI22_X1 U18336 ( .A1(n15231), .A2(n20448), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14833), .ZN(n14815) );
  OAI21_X1 U18337 ( .B1(n14816), .B2(n14838), .A(n14815), .ZN(P1_U2850) );
  INV_X1 U18338 ( .A(n15018), .ZN(n14818) );
  INV_X1 U18339 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14817) );
  OAI222_X1 U18340 ( .A1(n14818), .A2(n14838), .B1(n14817), .B2(n20452), .C1(
        n15238), .C2(n14835), .ZN(P1_U2851) );
  OAI222_X1 U18341 ( .A1(n14820), .A2(n14838), .B1(n14819), .B2(n20452), .C1(
        n15252), .C2(n14835), .ZN(P1_U2852) );
  AOI22_X1 U18342 ( .A1(n15261), .A2(n20448), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14833), .ZN(n14821) );
  OAI21_X1 U18343 ( .B1(n14822), .B2(n14838), .A(n14821), .ZN(P1_U2853) );
  OAI222_X1 U18344 ( .A1(n15279), .A2(n14835), .B1(n21444), .B2(n20452), .C1(
        n15044), .C2(n14838), .ZN(P1_U2854) );
  INV_X1 U18345 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14824) );
  OAI222_X1 U18346 ( .A1(n14825), .A2(n14838), .B1(n14824), .B2(n20452), .C1(
        n14823), .C2(n14835), .ZN(P1_U2855) );
  AOI22_X1 U18347 ( .A1(n15292), .A2(n20448), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14833), .ZN(n14826) );
  OAI21_X1 U18348 ( .B1(n14910), .B2(n14838), .A(n14826), .ZN(P1_U2856) );
  INV_X1 U18349 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14828) );
  OAI222_X1 U18350 ( .A1(n14921), .A2(n14838), .B1(n14828), .B2(n20452), .C1(
        n14827), .C2(n14835), .ZN(P1_U2857) );
  OAI222_X1 U18351 ( .A1(n14923), .A2(n14838), .B1(n14830), .B2(n20452), .C1(
        n14829), .C2(n14835), .ZN(P1_U2858) );
  INV_X1 U18352 ( .A(n15109), .ZN(n14926) );
  OAI222_X1 U18353 ( .A1(n14926), .A2(n14838), .B1(n14831), .B2(n20452), .C1(
        n14835), .C2(n15321), .ZN(P1_U2859) );
  OAI222_X1 U18354 ( .A1(n15335), .A2(n14835), .B1(n21357), .B2(n20452), .C1(
        n15121), .C2(n14838), .ZN(P1_U2860) );
  AOI22_X1 U18355 ( .A1(n15345), .A2(n20448), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14833), .ZN(n14832) );
  OAI21_X1 U18356 ( .B1(n14929), .B2(n14838), .A(n14832), .ZN(P1_U2861) );
  AOI22_X1 U18357 ( .A1(n15355), .A2(n20448), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14833), .ZN(n14834) );
  OAI21_X1 U18358 ( .B1(n14934), .B2(n14838), .A(n14834), .ZN(P1_U2862) );
  INV_X1 U18359 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14837) );
  OAI222_X1 U18360 ( .A1(n14939), .A2(n14838), .B1(n20452), .B2(n14837), .C1(
        n14836), .C2(n14835), .ZN(P1_U2863) );
  NAND2_X1 U18361 ( .A1(n14839), .A2(n14917), .ZN(n14845) );
  INV_X1 U18362 ( .A(DATAI_14_), .ZN(n14841) );
  NAND2_X1 U18363 ( .A1(n14866), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14840) );
  OAI21_X1 U18364 ( .B1(n14866), .B2(n14841), .A(n14840), .ZN(n20496) );
  AOI22_X1 U18365 ( .A1(n14911), .A2(n20496), .B1(n14935), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14844) );
  NAND2_X1 U18366 ( .A1(n14912), .A2(DATAI_30_), .ZN(n14843) );
  NAND2_X1 U18367 ( .A1(n14905), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14842) );
  NAND4_X1 U18368 ( .A1(n14845), .A2(n14844), .A3(n14843), .A4(n14842), .ZN(
        P1_U2874) );
  NAND2_X1 U18369 ( .A1(n14950), .A2(n14917), .ZN(n14851) );
  INV_X1 U18370 ( .A(DATAI_12_), .ZN(n14847) );
  NAND2_X1 U18371 ( .A1(n14866), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14846) );
  OAI21_X1 U18372 ( .B1(n14866), .B2(n14847), .A(n14846), .ZN(n20494) );
  AOI22_X1 U18373 ( .A1(n14911), .A2(n20494), .B1(n14935), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14850) );
  NAND2_X1 U18374 ( .A1(n14912), .A2(DATAI_28_), .ZN(n14849) );
  NAND2_X1 U18375 ( .A1(n14905), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14848) );
  NAND4_X1 U18376 ( .A1(n14851), .A2(n14850), .A3(n14849), .A4(n14848), .ZN(
        P1_U2876) );
  INV_X1 U18377 ( .A(n14852), .ZN(n14960) );
  NAND2_X1 U18378 ( .A1(n14960), .A2(n14917), .ZN(n14858) );
  INV_X1 U18379 ( .A(DATAI_11_), .ZN(n14854) );
  NAND2_X1 U18380 ( .A1(n14866), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14853) );
  OAI21_X1 U18381 ( .B1(n14866), .B2(n14854), .A(n14853), .ZN(n20492) );
  AOI22_X1 U18382 ( .A1(n14911), .A2(n20492), .B1(n14935), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14857) );
  NAND2_X1 U18383 ( .A1(n14912), .A2(DATAI_27_), .ZN(n14856) );
  NAND2_X1 U18384 ( .A1(n14905), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14855) );
  NAND4_X1 U18385 ( .A1(n14858), .A2(n14857), .A3(n14856), .A4(n14855), .ZN(
        P1_U2877) );
  NAND2_X1 U18386 ( .A1(n14971), .A2(n14917), .ZN(n14864) );
  INV_X1 U18387 ( .A(DATAI_10_), .ZN(n14860) );
  NAND2_X1 U18388 ( .A1(n14866), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14859) );
  OAI21_X1 U18389 ( .B1(n14866), .B2(n14860), .A(n14859), .ZN(n20490) );
  AOI22_X1 U18390 ( .A1(n14911), .A2(n20490), .B1(n14935), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14863) );
  NAND2_X1 U18391 ( .A1(n14912), .A2(DATAI_26_), .ZN(n14862) );
  NAND2_X1 U18392 ( .A1(n14905), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14861) );
  NAND4_X1 U18393 ( .A1(n14864), .A2(n14863), .A3(n14862), .A4(n14861), .ZN(
        P1_U2878) );
  INV_X1 U18394 ( .A(n14865), .ZN(n14981) );
  NAND2_X1 U18395 ( .A1(n14981), .A2(n14917), .ZN(n14873) );
  INV_X1 U18396 ( .A(DATAI_9_), .ZN(n14868) );
  NAND2_X1 U18397 ( .A1(n14866), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14867) );
  OAI21_X1 U18398 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n20488) );
  AOI22_X1 U18399 ( .A1(n14911), .A2(n20488), .B1(n14935), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14872) );
  NAND2_X1 U18400 ( .A1(n14912), .A2(DATAI_25_), .ZN(n14871) );
  NAND2_X1 U18401 ( .A1(n14905), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14870) );
  NAND4_X1 U18402 ( .A1(n14873), .A2(n14872), .A3(n14871), .A4(n14870), .ZN(
        P1_U2879) );
  INV_X1 U18403 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U18404 ( .A1(n14911), .A2(n20486), .B1(n14935), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14875) );
  NAND2_X1 U18405 ( .A1(n14912), .A2(DATAI_24_), .ZN(n14874) );
  OAI211_X1 U18406 ( .C1(n20588), .C2(n14915), .A(n14875), .B(n14874), .ZN(
        n14876) );
  AOI21_X1 U18407 ( .B1(n14877), .B2(n14917), .A(n14876), .ZN(n14878) );
  INV_X1 U18408 ( .A(n14878), .ZN(P1_U2880) );
  NAND2_X1 U18409 ( .A1(n14999), .A2(n14917), .ZN(n14882) );
  AOI22_X1 U18410 ( .A1(n14911), .A2(n20652), .B1(n14935), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n14881) );
  NAND2_X1 U18411 ( .A1(n14912), .A2(DATAI_23_), .ZN(n14880) );
  NAND2_X1 U18412 ( .A1(n14905), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14879) );
  NAND4_X1 U18413 ( .A1(n14882), .A2(n14881), .A3(n14880), .A4(n14879), .ZN(
        P1_U2881) );
  INV_X1 U18414 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20635) );
  AOI22_X1 U18415 ( .A1(n14911), .A2(n20639), .B1(n14935), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14884) );
  NAND2_X1 U18416 ( .A1(n14912), .A2(DATAI_22_), .ZN(n14883) );
  OAI211_X1 U18417 ( .C1(n14915), .C2(n20635), .A(n14884), .B(n14883), .ZN(
        n14885) );
  AOI21_X1 U18418 ( .B1(n15007), .B2(n14917), .A(n14885), .ZN(n14886) );
  INV_X1 U18419 ( .A(n14886), .ZN(P1_U2882) );
  NAND2_X1 U18420 ( .A1(n15018), .A2(n14917), .ZN(n14890) );
  AOI22_X1 U18421 ( .A1(n14911), .A2(n20631), .B1(n14935), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U18422 ( .A1(n14912), .A2(DATAI_21_), .ZN(n14888) );
  NAND2_X1 U18423 ( .A1(n14905), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14887) );
  NAND4_X1 U18424 ( .A1(n14890), .A2(n14889), .A3(n14888), .A4(n14887), .ZN(
        P1_U2883) );
  NAND2_X1 U18425 ( .A1(n15027), .A2(n14917), .ZN(n14894) );
  AOI22_X1 U18426 ( .A1(n14911), .A2(n20622), .B1(n14935), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n14893) );
  NAND2_X1 U18427 ( .A1(n14912), .A2(DATAI_20_), .ZN(n14892) );
  NAND2_X1 U18428 ( .A1(n14905), .A2(BUF1_REG_20__SCAN_IN), .ZN(n14891) );
  NAND4_X1 U18429 ( .A1(n14894), .A2(n14893), .A3(n14892), .A4(n14891), .ZN(
        P1_U2884) );
  NAND2_X1 U18430 ( .A1(n15035), .A2(n14917), .ZN(n14898) );
  AOI22_X1 U18431 ( .A1(n14911), .A2(n20614), .B1(n14935), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14897) );
  NAND2_X1 U18432 ( .A1(n14912), .A2(DATAI_19_), .ZN(n14896) );
  NAND2_X1 U18433 ( .A1(n14905), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14895) );
  NAND4_X1 U18434 ( .A1(n14898), .A2(n14897), .A3(n14896), .A4(n14895), .ZN(
        P1_U2885) );
  INV_X1 U18435 ( .A(n15044), .ZN(n14899) );
  NAND2_X1 U18436 ( .A1(n14899), .A2(n14917), .ZN(n14904) );
  AOI22_X1 U18437 ( .A1(n14911), .A2(n14900), .B1(n14935), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14903) );
  NAND2_X1 U18438 ( .A1(n14912), .A2(DATAI_18_), .ZN(n14902) );
  NAND2_X1 U18439 ( .A1(n14905), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14901) );
  NAND4_X1 U18440 ( .A1(n14904), .A2(n14903), .A3(n14902), .A4(n14901), .ZN(
        P1_U2886) );
  NAND2_X1 U18441 ( .A1(n15063), .A2(n14917), .ZN(n14909) );
  AOI22_X1 U18442 ( .A1(n14911), .A2(n20600), .B1(n14935), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14908) );
  NAND2_X1 U18443 ( .A1(n14912), .A2(DATAI_17_), .ZN(n14907) );
  NAND2_X1 U18444 ( .A1(n14905), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14906) );
  NAND4_X1 U18445 ( .A1(n14909), .A2(n14908), .A3(n14907), .A4(n14906), .ZN(
        P1_U2887) );
  INV_X1 U18446 ( .A(n14910), .ZN(n15074) );
  INV_X1 U18447 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20593) );
  AOI22_X1 U18448 ( .A1(n14911), .A2(n20591), .B1(n14935), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14914) );
  NAND2_X1 U18449 ( .A1(n14912), .A2(DATAI_16_), .ZN(n14913) );
  OAI211_X1 U18450 ( .C1(n14915), .C2(n20593), .A(n14914), .B(n14913), .ZN(
        n14916) );
  AOI21_X1 U18451 ( .B1(n15074), .B2(n14917), .A(n14916), .ZN(n14918) );
  INV_X1 U18452 ( .A(n14918), .ZN(P1_U2888) );
  OAI222_X1 U18453 ( .A1(n14938), .A2(n14921), .B1(n14931), .B2(n14920), .C1(
        n14919), .C2(n14932), .ZN(P1_U2889) );
  AOI22_X1 U18454 ( .A1(n14936), .A2(n20496), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14935), .ZN(n14922) );
  OAI21_X1 U18455 ( .B1(n14923), .B2(n14938), .A(n14922), .ZN(P1_U2890) );
  AOI22_X1 U18456 ( .A1(n14936), .A2(n14924), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14935), .ZN(n14925) );
  OAI21_X1 U18457 ( .B1(n14926), .B2(n14938), .A(n14925), .ZN(P1_U2891) );
  AOI22_X1 U18458 ( .A1(n14936), .A2(n20494), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14935), .ZN(n14927) );
  OAI21_X1 U18459 ( .B1(n15121), .B2(n14938), .A(n14927), .ZN(P1_U2892) );
  AOI22_X1 U18460 ( .A1(n14936), .A2(n20492), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14935), .ZN(n14928) );
  OAI21_X1 U18461 ( .B1(n14929), .B2(n14938), .A(n14928), .ZN(P1_U2893) );
  INV_X1 U18462 ( .A(n20490), .ZN(n14930) );
  OAI222_X1 U18463 ( .A1(n14934), .A2(n14938), .B1(n14933), .B2(n14932), .C1(
        n14931), .C2(n14930), .ZN(P1_U2894) );
  AOI22_X1 U18464 ( .A1(n14936), .A2(n20488), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14935), .ZN(n14937) );
  OAI21_X1 U18465 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(P1_U2895) );
  NAND2_X1 U18466 ( .A1(n9623), .A2(n15183), .ZN(n14940) );
  NAND2_X1 U18467 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14941) );
  AND3_X1 U18468 ( .A1(n14975), .A2(n15182), .A3(n14956), .ZN(n14942) );
  NAND4_X1 U18469 ( .A1(n14943), .A2(n14942), .A3(n15203), .A4(n15194), .ZN(
        n14944) );
  NOR2_X1 U18470 ( .A1(n20416), .A2(n14946), .ZN(n15166) );
  AOI21_X1 U18471 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15166), .ZN(n14947) );
  OAI21_X1 U18472 ( .B1(n20524), .B2(n14948), .A(n14947), .ZN(n14949) );
  AOI21_X1 U18473 ( .B1(n14950), .B2(n20519), .A(n14949), .ZN(n14951) );
  OAI21_X1 U18474 ( .B1(n15151), .B2(n15170), .A(n14951), .ZN(P1_U2971) );
  INV_X1 U18475 ( .A(n10712), .ZN(n14952) );
  NAND2_X1 U18476 ( .A1(n14953), .A2(n14952), .ZN(n14954) );
  NOR2_X1 U18477 ( .A1(n20416), .A2(n21269), .ZN(n15173) );
  AOI21_X1 U18478 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15173), .ZN(n14957) );
  OAI21_X1 U18479 ( .B1(n20524), .B2(n14958), .A(n14957), .ZN(n14959) );
  AOI21_X1 U18480 ( .B1(n14960), .B2(n20519), .A(n14959), .ZN(n14961) );
  OAI21_X1 U18481 ( .B1(n15151), .B2(n15178), .A(n14961), .ZN(P1_U2972) );
  OAI21_X1 U18482 ( .B1(n14963), .B2(n15183), .A(n9623), .ZN(n14965) );
  NAND2_X1 U18483 ( .A1(n14962), .A2(n14965), .ZN(n14966) );
  XNOR2_X1 U18484 ( .A(n14966), .B(n15182), .ZN(n15190) );
  NOR2_X1 U18485 ( .A1(n20416), .A2(n14967), .ZN(n15185) );
  AOI21_X1 U18486 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15185), .ZN(n14968) );
  OAI21_X1 U18487 ( .B1(n20524), .B2(n14969), .A(n14968), .ZN(n14970) );
  AOI21_X1 U18488 ( .B1(n14971), .B2(n20519), .A(n14970), .ZN(n14972) );
  OAI21_X1 U18489 ( .B1(n15151), .B2(n15190), .A(n14972), .ZN(P1_U2973) );
  NAND2_X1 U18490 ( .A1(n14973), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14987) );
  MUX2_X1 U18491 ( .A(n14975), .B(n14974), .S(n15049), .Z(n14976) );
  AOI21_X1 U18492 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14987), .A(
        n14976), .ZN(n14977) );
  XNOR2_X1 U18493 ( .A(n14977), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15199) );
  NOR2_X1 U18494 ( .A1(n20416), .A2(n21404), .ZN(n15191) );
  AOI21_X1 U18495 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15191), .ZN(n14978) );
  OAI21_X1 U18496 ( .B1(n20524), .B2(n14979), .A(n14978), .ZN(n14980) );
  AOI21_X1 U18497 ( .B1(n14981), .B2(n20519), .A(n14980), .ZN(n14982) );
  OAI21_X1 U18498 ( .B1(n15151), .B2(n15199), .A(n14982), .ZN(P1_U2974) );
  NOR2_X1 U18499 ( .A1(n20416), .A2(n14983), .ZN(n15205) );
  NOR2_X1 U18500 ( .A1(n20524), .A2(n14984), .ZN(n14985) );
  AOI211_X1 U18501 ( .C1(n17105), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15205), .B(n14985), .ZN(n14990) );
  NAND2_X1 U18502 ( .A1(n14963), .A2(n14987), .ZN(n14986) );
  MUX2_X1 U18503 ( .A(n14987), .B(n14986), .S(n15049), .Z(n14988) );
  XNOR2_X1 U18504 ( .A(n14988), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15200) );
  NAND2_X1 U18505 ( .A1(n15200), .A2(n20518), .ZN(n14989) );
  OAI211_X1 U18506 ( .C1(n14991), .C2(n15122), .A(n14990), .B(n14989), .ZN(
        P1_U2975) );
  XNOR2_X1 U18507 ( .A(n9623), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14992) );
  XNOR2_X1 U18508 ( .A(n14993), .B(n14992), .ZN(n15218) );
  INV_X1 U18509 ( .A(n14994), .ZN(n14997) );
  NOR2_X1 U18510 ( .A1(n20416), .A2(n14995), .ZN(n15212) );
  AOI21_X1 U18511 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15212), .ZN(n14996) );
  OAI21_X1 U18512 ( .B1(n20524), .B2(n14997), .A(n14996), .ZN(n14998) );
  AOI21_X1 U18513 ( .B1(n14999), .B2(n20519), .A(n14998), .ZN(n15000) );
  OAI21_X1 U18514 ( .B1(n15218), .B2(n15151), .A(n15000), .ZN(P1_U2976) );
  NAND2_X1 U18515 ( .A1(n15002), .A2(n15001), .ZN(n15003) );
  XOR2_X1 U18516 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15003), .Z(
        n15234) );
  NOR2_X1 U18517 ( .A1(n20416), .A2(n21264), .ZN(n15229) );
  AOI21_X1 U18518 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15229), .ZN(n15004) );
  OAI21_X1 U18519 ( .B1(n20524), .B2(n15005), .A(n15004), .ZN(n15006) );
  AOI21_X1 U18520 ( .B1(n15007), .B2(n20519), .A(n15006), .ZN(n15008) );
  OAI21_X1 U18521 ( .B1(n15151), .B2(n15234), .A(n15008), .ZN(P1_U2977) );
  NOR3_X1 U18522 ( .A1(n15009), .A2(n15049), .A3(n10709), .ZN(n15021) );
  NOR2_X1 U18523 ( .A1(n15010), .A2(n9623), .ZN(n15020) );
  AOI22_X1 U18524 ( .A1(n15021), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15020), .B2(n15246), .ZN(n15012) );
  XNOR2_X1 U18525 ( .A(n15012), .B(n15011), .ZN(n15242) );
  INV_X1 U18526 ( .A(n15013), .ZN(n15016) );
  NOR2_X1 U18527 ( .A1(n20416), .A2(n15014), .ZN(n15236) );
  AOI21_X1 U18528 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15236), .ZN(n15015) );
  OAI21_X1 U18529 ( .B1(n20524), .B2(n15016), .A(n15015), .ZN(n15017) );
  AOI21_X1 U18530 ( .B1(n15018), .B2(n20519), .A(n15017), .ZN(n15019) );
  OAI21_X1 U18531 ( .B1(n15242), .B2(n15151), .A(n15019), .ZN(P1_U2978) );
  NOR2_X1 U18532 ( .A1(n15021), .A2(n15020), .ZN(n15022) );
  XNOR2_X1 U18533 ( .A(n15022), .B(n15246), .ZN(n15255) );
  NOR2_X1 U18534 ( .A1(n20416), .A2(n15023), .ZN(n15243) );
  AOI21_X1 U18535 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15243), .ZN(n15024) );
  OAI21_X1 U18536 ( .B1(n20524), .B2(n15025), .A(n15024), .ZN(n15026) );
  AOI21_X1 U18537 ( .B1(n15027), .B2(n20519), .A(n15026), .ZN(n15028) );
  OAI21_X1 U18538 ( .B1(n15255), .B2(n15151), .A(n15028), .ZN(P1_U2979) );
  NOR2_X1 U18539 ( .A1(n9623), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15029) );
  MUX2_X1 U18540 ( .A(n9623), .B(n15029), .S(n15009), .Z(n15030) );
  XNOR2_X1 U18541 ( .A(n15030), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15264) );
  NOR2_X1 U18542 ( .A1(n20416), .A2(n15031), .ZN(n15259) );
  AOI21_X1 U18543 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15259), .ZN(n15032) );
  OAI21_X1 U18544 ( .B1(n20524), .B2(n15033), .A(n15032), .ZN(n15034) );
  AOI21_X1 U18545 ( .B1(n15035), .B2(n20519), .A(n15034), .ZN(n15036) );
  OAI21_X1 U18546 ( .B1(n15151), .B2(n15264), .A(n15036), .ZN(P1_U2980) );
  NOR2_X1 U18547 ( .A1(n15037), .A2(n15038), .ZN(n15265) );
  NOR2_X1 U18548 ( .A1(n15265), .A2(n15151), .ZN(n15042) );
  NOR2_X1 U18549 ( .A1(n20416), .A2(n21262), .ZN(n15275) );
  AOI21_X1 U18550 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15275), .ZN(n15039) );
  OAI21_X1 U18551 ( .B1(n20524), .B2(n15040), .A(n15039), .ZN(n15041) );
  AOI21_X1 U18552 ( .B1(n15042), .B2(n15009), .A(n15041), .ZN(n15043) );
  OAI21_X1 U18553 ( .B1(n15044), .B2(n15122), .A(n15043), .ZN(P1_U2981) );
  NAND2_X1 U18554 ( .A1(n9623), .A2(n15352), .ZN(n15047) );
  NAND2_X1 U18555 ( .A1(n15049), .A2(n15048), .ZN(n15050) );
  NAND2_X1 U18556 ( .A1(n15131), .A2(n15050), .ZN(n15052) );
  INV_X1 U18557 ( .A(n15054), .ZN(n15055) );
  NAND2_X1 U18558 ( .A1(n15056), .A2(n15055), .ZN(n15080) );
  NOR2_X1 U18559 ( .A1(n9623), .A2(n15289), .ZN(n15077) );
  NOR2_X1 U18560 ( .A1(n20416), .A2(n15059), .ZN(n15285) );
  AOI21_X1 U18561 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15285), .ZN(n15060) );
  OAI21_X1 U18562 ( .B1(n20524), .B2(n15061), .A(n15060), .ZN(n15062) );
  AOI21_X1 U18563 ( .B1(n15063), .B2(n20519), .A(n15062), .ZN(n15064) );
  OAI21_X1 U18564 ( .B1(n15151), .B2(n15288), .A(n15064), .ZN(P1_U2982) );
  NAND2_X1 U18565 ( .A1(n15076), .A2(n15081), .ZN(n15067) );
  INV_X1 U18566 ( .A(n15065), .ZN(n15066) );
  NAND2_X1 U18567 ( .A1(n15067), .A2(n15066), .ZN(n15069) );
  NAND2_X1 U18568 ( .A1(n15069), .A2(n15068), .ZN(n15298) );
  NOR2_X1 U18569 ( .A1(n20416), .A2(n15070), .ZN(n15291) );
  AOI21_X1 U18570 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15291), .ZN(n15071) );
  OAI21_X1 U18571 ( .B1(n20524), .B2(n15072), .A(n15071), .ZN(n15073) );
  AOI21_X1 U18572 ( .B1(n15074), .B2(n20519), .A(n15073), .ZN(n15075) );
  OAI21_X1 U18573 ( .B1(n15151), .B2(n15298), .A(n15075), .ZN(P1_U2983) );
  INV_X1 U18574 ( .A(n15076), .ZN(n15082) );
  INV_X1 U18575 ( .A(n15077), .ZN(n15078) );
  NAND2_X1 U18576 ( .A1(n15078), .A2(n15081), .ZN(n15079) );
  AOI22_X1 U18577 ( .A1(n15082), .A2(n15081), .B1(n15080), .B2(n15079), .ZN(
        n15305) );
  NOR2_X1 U18578 ( .A1(n20416), .A2(n15083), .ZN(n15299) );
  AOI21_X1 U18579 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15299), .ZN(n15084) );
  OAI21_X1 U18580 ( .B1(n20524), .B2(n15085), .A(n15084), .ZN(n15086) );
  AOI21_X1 U18581 ( .B1(n15087), .B2(n20519), .A(n15086), .ZN(n15088) );
  OAI21_X1 U18582 ( .B1(n15305), .B2(n15151), .A(n15088), .ZN(P1_U2984) );
  XNOR2_X1 U18583 ( .A(n9623), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15090) );
  XNOR2_X1 U18584 ( .A(n15091), .B(n15090), .ZN(n15306) );
  NOR2_X1 U18585 ( .A1(n20416), .A2(n15092), .ZN(n15307) );
  AOI21_X1 U18586 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15307), .ZN(n15093) );
  OAI21_X1 U18587 ( .B1(n20524), .B2(n15094), .A(n15093), .ZN(n15095) );
  AOI21_X1 U18588 ( .B1(n15096), .B2(n20519), .A(n15095), .ZN(n15097) );
  OAI21_X1 U18589 ( .B1(n15306), .B2(n15151), .A(n15097), .ZN(P1_U2985) );
  AOI21_X1 U18590 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15049), .ZN(n15100) );
  OAI22_X1 U18591 ( .A1(n15131), .A2(n15100), .B1(n15099), .B2(n9623), .ZN(
        n15115) );
  NAND2_X1 U18592 ( .A1(n9623), .A2(n15338), .ZN(n15101) );
  OAI21_X1 U18593 ( .B1(n9623), .B2(n15338), .A(n15101), .ZN(n15114) );
  NOR2_X1 U18594 ( .A1(n15115), .A2(n15114), .ZN(n15113) );
  INV_X1 U18595 ( .A(n15101), .ZN(n15102) );
  NOR2_X1 U18596 ( .A1(n15113), .A2(n15102), .ZN(n15104) );
  XNOR2_X1 U18597 ( .A(n15104), .B(n15103), .ZN(n15325) );
  NOR2_X1 U18598 ( .A1(n20416), .A2(n15105), .ZN(n15319) );
  AOI21_X1 U18599 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15319), .ZN(n15106) );
  OAI21_X1 U18600 ( .B1(n20524), .B2(n15107), .A(n15106), .ZN(n15108) );
  AOI21_X1 U18601 ( .B1(n15109), .B2(n20519), .A(n15108), .ZN(n15110) );
  OAI21_X1 U18602 ( .B1(n15151), .B2(n15325), .A(n15110), .ZN(P1_U2986) );
  NAND2_X1 U18603 ( .A1(n20580), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15334) );
  OAI21_X1 U18604 ( .B1(n15112), .B2(n15111), .A(n15334), .ZN(n15117) );
  AOI21_X1 U18605 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15341) );
  NOR2_X1 U18606 ( .A1(n15341), .A2(n15151), .ZN(n15116) );
  AOI211_X1 U18607 ( .C1(n15119), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        n15120) );
  OAI21_X1 U18608 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(P1_U2987) );
  NOR3_X1 U18609 ( .A1(n15131), .A2(n15049), .A3(n15132), .ZN(n15123) );
  NOR3_X1 U18610 ( .A1(n15045), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9623), .ZN(n15136) );
  NOR2_X1 U18611 ( .A1(n15123), .A2(n15136), .ZN(n15124) );
  XNOR2_X1 U18612 ( .A(n15124), .B(n15346), .ZN(n15350) );
  NOR2_X1 U18613 ( .A1(n20416), .A2(n15125), .ZN(n15344) );
  AOI21_X1 U18614 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15344), .ZN(n15126) );
  OAI21_X1 U18615 ( .B1(n20524), .B2(n15127), .A(n15126), .ZN(n15128) );
  AOI21_X1 U18616 ( .B1(n15129), .B2(n20519), .A(n15128), .ZN(n15130) );
  OAI21_X1 U18617 ( .B1(n15350), .B2(n15151), .A(n15130), .ZN(P1_U2988) );
  XNOR2_X1 U18618 ( .A(n15131), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15135) );
  INV_X1 U18619 ( .A(n15045), .ZN(n15133) );
  NOR2_X1 U18620 ( .A1(n15133), .A2(n15132), .ZN(n15134) );
  MUX2_X1 U18621 ( .A(n15135), .B(n15134), .S(n15049), .Z(n15137) );
  NOR2_X1 U18622 ( .A1(n15137), .A2(n15136), .ZN(n15360) );
  NOR2_X1 U18623 ( .A1(n20416), .A2(n15138), .ZN(n15354) );
  AOI21_X1 U18624 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15354), .ZN(n15139) );
  OAI21_X1 U18625 ( .B1(n20524), .B2(n15140), .A(n15139), .ZN(n15141) );
  AOI21_X1 U18626 ( .B1(n15142), .B2(n20519), .A(n15141), .ZN(n15143) );
  OAI21_X1 U18627 ( .B1(n15360), .B2(n15151), .A(n15143), .ZN(P1_U2989) );
  INV_X1 U18628 ( .A(n15144), .ZN(n15145) );
  AOI21_X1 U18629 ( .B1(n17105), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15145), .ZN(n15146) );
  OAI21_X1 U18630 ( .B1(n20524), .B2(n15147), .A(n15146), .ZN(n15148) );
  AOI21_X1 U18631 ( .B1(n15149), .B2(n20519), .A(n15148), .ZN(n15150) );
  OAI21_X1 U18632 ( .B1(n15152), .B2(n15151), .A(n15150), .ZN(P1_U2990) );
  INV_X1 U18633 ( .A(n15153), .ZN(n15159) );
  INV_X1 U18634 ( .A(n15171), .ZN(n15164) );
  AOI21_X1 U18635 ( .B1(n15164), .B2(n15154), .A(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15156) );
  OAI21_X1 U18636 ( .B1(n15157), .B2(n15156), .A(n15155), .ZN(n15158) );
  AOI21_X1 U18637 ( .B1(n15159), .B2(n20544), .A(n15158), .ZN(n15160) );
  OAI21_X1 U18638 ( .B1(n15161), .B2(n20576), .A(n15160), .ZN(P1_U3002) );
  AND3_X1 U18639 ( .A1(n15164), .A2(n15163), .A3(n15162), .ZN(n15165) );
  AOI211_X1 U18640 ( .C1(n15174), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15166), .B(n15165), .ZN(n15169) );
  NAND2_X1 U18641 ( .A1(n15167), .A2(n20544), .ZN(n15168) );
  OAI211_X1 U18642 ( .C1(n15170), .C2(n20576), .A(n15169), .B(n15168), .ZN(
        P1_U3003) );
  NOR2_X1 U18643 ( .A1(n15171), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15172) );
  AOI211_X1 U18644 ( .C1(n15174), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15173), .B(n15172), .ZN(n15177) );
  NAND2_X1 U18645 ( .A1(n15175), .A2(n20544), .ZN(n15176) );
  OAI211_X1 U18646 ( .C1(n15178), .C2(n20576), .A(n15177), .B(n15176), .ZN(
        P1_U3004) );
  INV_X1 U18647 ( .A(n15179), .ZN(n15195) );
  INV_X1 U18648 ( .A(n15210), .ZN(n15181) );
  NAND3_X1 U18649 ( .A1(n15181), .A2(n15180), .A3(n15194), .ZN(n15192) );
  AOI21_X1 U18650 ( .B1(n15195), .B2(n15192), .A(n15182), .ZN(n15186) );
  NOR3_X1 U18651 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15183), .ZN(n15184) );
  NOR3_X1 U18652 ( .A1(n15186), .A2(n15185), .A3(n15184), .ZN(n15189) );
  NAND2_X1 U18653 ( .A1(n15187), .A2(n20544), .ZN(n15188) );
  OAI211_X1 U18654 ( .C1(n15190), .C2(n20576), .A(n15189), .B(n15188), .ZN(
        P1_U3005) );
  INV_X1 U18655 ( .A(n15191), .ZN(n15193) );
  OAI211_X1 U18656 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15196) );
  AOI21_X1 U18657 ( .B1(n15197), .B2(n20544), .A(n15196), .ZN(n15198) );
  OAI21_X1 U18658 ( .B1(n15199), .B2(n20576), .A(n15198), .ZN(P1_U3006) );
  NAND2_X1 U18659 ( .A1(n15200), .A2(n20550), .ZN(n15208) );
  OAI21_X1 U18660 ( .B1(n15202), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15201), .ZN(n15206) );
  NOR3_X1 U18661 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15203), .ZN(n15204) );
  AOI211_X1 U18662 ( .C1(n15206), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15205), .B(n15204), .ZN(n15207) );
  OAI211_X1 U18663 ( .C1(n20578), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        P1_U3007) );
  NOR2_X1 U18664 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15211) );
  AOI211_X1 U18665 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15213), .A(
        n15212), .B(n15211), .ZN(n15217) );
  INV_X1 U18666 ( .A(n15214), .ZN(n15215) );
  NAND2_X1 U18667 ( .A1(n15215), .A2(n20544), .ZN(n15216) );
  OAI211_X1 U18668 ( .C1(n15218), .C2(n20576), .A(n15217), .B(n15216), .ZN(
        P1_U3008) );
  NAND2_X1 U18669 ( .A1(n20573), .A2(n15270), .ZN(n15222) );
  NAND2_X1 U18670 ( .A1(n15219), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15220) );
  OR2_X1 U18671 ( .A1(n20572), .A2(n15220), .ZN(n15221) );
  AND2_X1 U18672 ( .A1(n15222), .A2(n15221), .ZN(n15245) );
  OR2_X1 U18673 ( .A1(n20582), .A2(n15223), .ZN(n15224) );
  NAND2_X1 U18674 ( .A1(n15245), .A2(n15224), .ZN(n15317) );
  NAND2_X1 U18675 ( .A1(n15317), .A2(n15225), .ZN(n15256) );
  NOR3_X1 U18676 ( .A1(n15256), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15226), .ZN(n15235) );
  OR2_X1 U18677 ( .A1(n15235), .A2(n15237), .ZN(n15230) );
  NOR3_X1 U18678 ( .A1(n15256), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15227), .ZN(n15228) );
  AOI211_X1 U18679 ( .C1(n15230), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15229), .B(n15228), .ZN(n15233) );
  NAND2_X1 U18680 ( .A1(n15231), .A2(n20544), .ZN(n15232) );
  OAI211_X1 U18681 ( .C1(n15234), .C2(n20576), .A(n15233), .B(n15232), .ZN(
        P1_U3009) );
  AOI211_X1 U18682 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15237), .A(
        n15236), .B(n15235), .ZN(n15241) );
  INV_X1 U18683 ( .A(n15238), .ZN(n15239) );
  NAND2_X1 U18684 ( .A1(n15239), .A2(n20544), .ZN(n15240) );
  OAI211_X1 U18685 ( .C1(n15242), .C2(n20576), .A(n15241), .B(n15240), .ZN(
        P1_U3010) );
  INV_X1 U18686 ( .A(n15243), .ZN(n15251) );
  INV_X1 U18687 ( .A(n15257), .ZN(n15249) );
  AOI21_X1 U18688 ( .B1(n15245), .B2(n20582), .A(n15244), .ZN(n15248) );
  OAI21_X1 U18689 ( .B1(n15256), .B2(n10709), .A(n15246), .ZN(n15247) );
  OAI21_X1 U18690 ( .B1(n15249), .B2(n15248), .A(n15247), .ZN(n15250) );
  OAI211_X1 U18691 ( .C1(n15252), .C2(n20578), .A(n15251), .B(n15250), .ZN(
        n15253) );
  INV_X1 U18692 ( .A(n15253), .ZN(n15254) );
  OAI21_X1 U18693 ( .B1(n15255), .B2(n20576), .A(n15254), .ZN(P1_U3011) );
  INV_X1 U18694 ( .A(n15256), .ZN(n15260) );
  NOR2_X1 U18695 ( .A1(n15257), .A2(n10709), .ZN(n15258) );
  AOI211_X1 U18696 ( .C1(n15260), .C2(n10709), .A(n15259), .B(n15258), .ZN(
        n15263) );
  NAND2_X1 U18697 ( .A1(n15261), .A2(n20544), .ZN(n15262) );
  OAI211_X1 U18698 ( .C1(n15264), .C2(n20576), .A(n15263), .B(n15262), .ZN(
        P1_U3012) );
  INV_X1 U18699 ( .A(n15265), .ZN(n15266) );
  NAND3_X1 U18700 ( .A1(n15266), .A2(n20550), .A3(n15009), .ZN(n15278) );
  INV_X1 U18701 ( .A(n20573), .ZN(n15328) );
  INV_X1 U18702 ( .A(n15267), .ZN(n15268) );
  NAND2_X1 U18703 ( .A1(n20546), .A2(n15268), .ZN(n15269) );
  OAI211_X1 U18704 ( .C1(n15270), .C2(n15328), .A(n20547), .B(n15269), .ZN(
        n15320) );
  AND2_X1 U18705 ( .A1(n20573), .A2(n15316), .ZN(n15271) );
  OR2_X1 U18706 ( .A1(n15320), .A2(n15271), .ZN(n15311) );
  AOI21_X1 U18707 ( .B1(n15293), .B2(n15272), .A(n15311), .ZN(n15281) );
  INV_X1 U18708 ( .A(n15281), .ZN(n15276) );
  INV_X1 U18709 ( .A(n15280), .ZN(n15273) );
  NOR3_X1 U18710 ( .A1(n15273), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15272), .ZN(n15274) );
  AOI211_X1 U18711 ( .C1(n15276), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15275), .B(n15274), .ZN(n15277) );
  OAI211_X1 U18712 ( .C1(n15279), .C2(n20578), .A(n15278), .B(n15277), .ZN(
        P1_U3013) );
  AND2_X1 U18713 ( .A1(n15280), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15302) );
  NAND3_X1 U18714 ( .A1(n15302), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15282) );
  AOI21_X1 U18715 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(n15284) );
  AOI211_X1 U18716 ( .C1(n15286), .C2(n20544), .A(n15285), .B(n15284), .ZN(
        n15287) );
  OAI21_X1 U18717 ( .B1(n15288), .B2(n20576), .A(n15287), .ZN(P1_U3014) );
  INV_X1 U18718 ( .A(n15302), .ZN(n15295) );
  NOR3_X1 U18719 ( .A1(n15295), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15289), .ZN(n15290) );
  AOI211_X1 U18720 ( .C1(n15292), .C2(n20544), .A(n15291), .B(n15290), .ZN(
        n15297) );
  AOI21_X1 U18721 ( .B1(n15309), .B2(n15293), .A(n15311), .ZN(n15294) );
  OAI21_X1 U18722 ( .B1(n15295), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15294), .ZN(n15301) );
  NAND2_X1 U18723 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15296) );
  OAI211_X1 U18724 ( .C1(n15298), .C2(n20576), .A(n15297), .B(n15296), .ZN(
        P1_U3015) );
  AOI21_X1 U18725 ( .B1(n15300), .B2(n20544), .A(n15299), .ZN(n15304) );
  OAI21_X1 U18726 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15302), .A(
        n15301), .ZN(n15303) );
  OAI211_X1 U18727 ( .C1(n15305), .C2(n20576), .A(n15304), .B(n15303), .ZN(
        P1_U3016) );
  OR2_X1 U18728 ( .A1(n15306), .A2(n20576), .ZN(n15315) );
  AOI21_X1 U18729 ( .B1(n15308), .B2(n20544), .A(n15307), .ZN(n15314) );
  NOR2_X1 U18730 ( .A1(n17123), .A2(n15327), .ZN(n15347) );
  NAND4_X1 U18731 ( .A1(n15347), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15310), .A4(n15309), .ZN(n15313) );
  NAND2_X1 U18732 ( .A1(n15311), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15312) );
  NAND4_X1 U18733 ( .A1(n15315), .A2(n15314), .A3(n15313), .A4(n15312), .ZN(
        P1_U3017) );
  AND2_X1 U18734 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  AOI211_X1 U18735 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15320), .A(
        n15319), .B(n15318), .ZN(n15324) );
  INV_X1 U18736 ( .A(n15321), .ZN(n15322) );
  NAND2_X1 U18737 ( .A1(n15322), .A2(n20544), .ZN(n15323) );
  OAI211_X1 U18738 ( .C1(n15325), .C2(n20576), .A(n15324), .B(n15323), .ZN(
        P1_U3018) );
  INV_X1 U18739 ( .A(n20553), .ZN(n15333) );
  INV_X1 U18740 ( .A(n15326), .ZN(n15332) );
  INV_X1 U18741 ( .A(n15327), .ZN(n15329) );
  AOI21_X1 U18742 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15329), .A(
        n15328), .ZN(n15331) );
  AOI211_X1 U18743 ( .C1(n20546), .C2(n15332), .A(n15331), .B(n15330), .ZN(
        n15342) );
  OAI21_X1 U18744 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15333), .A(
        n15342), .ZN(n15337) );
  OAI21_X1 U18745 ( .B1(n15335), .B2(n20578), .A(n15334), .ZN(n15336) );
  AOI21_X1 U18746 ( .B1(n15337), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15336), .ZN(n15340) );
  NAND3_X1 U18747 ( .A1(n15347), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15338), .ZN(n15339) );
  OAI211_X1 U18748 ( .C1(n15341), .C2(n20576), .A(n15340), .B(n15339), .ZN(
        P1_U3019) );
  NOR2_X1 U18749 ( .A1(n15342), .A2(n15346), .ZN(n15343) );
  AOI211_X1 U18750 ( .C1(n20544), .C2(n15345), .A(n15344), .B(n15343), .ZN(
        n15349) );
  NAND2_X1 U18751 ( .A1(n15347), .A2(n15346), .ZN(n15348) );
  OAI211_X1 U18752 ( .C1(n15350), .C2(n20576), .A(n15349), .B(n15348), .ZN(
        P1_U3020) );
  NOR4_X1 U18753 ( .A1(n17123), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15352), .A4(n15351), .ZN(n15353) );
  AOI211_X1 U18754 ( .C1(n20544), .C2(n15355), .A(n15354), .B(n15353), .ZN(
        n15359) );
  OAI21_X1 U18755 ( .B1(n15357), .B2(n15356), .A(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15358) );
  OAI211_X1 U18756 ( .C1(n15360), .C2(n20576), .A(n15359), .B(n15358), .ZN(
        P1_U3021) );
  NAND2_X1 U18757 ( .A1(n20893), .A2(n15386), .ZN(n15377) );
  NOR2_X1 U18758 ( .A1(n14273), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15362) );
  NOR2_X1 U18759 ( .A1(n15362), .A2(n15361), .ZN(n15364) );
  AND2_X1 U18760 ( .A1(n15364), .A2(n15363), .ZN(n21277) );
  NAND2_X1 U18761 ( .A1(n15378), .A2(n21277), .ZN(n15374) );
  MUX2_X1 U18762 ( .A(n15361), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14273), .Z(n15366) );
  NOR2_X1 U18763 ( .A1(n15366), .A2(n15365), .ZN(n15372) );
  INV_X1 U18764 ( .A(n15367), .ZN(n15369) );
  NAND2_X1 U18765 ( .A1(n15369), .A2(n15368), .ZN(n15382) );
  XNOR2_X1 U18766 ( .A(n15370), .B(n10317), .ZN(n15371) );
  AOI22_X1 U18767 ( .A1(n15372), .A2(n15382), .B1(n17060), .B2(n15371), .ZN(
        n15373) );
  OAI21_X1 U18768 ( .B1(n15386), .B2(n15374), .A(n15373), .ZN(n15375) );
  INV_X1 U18769 ( .A(n15375), .ZN(n15376) );
  NAND2_X1 U18770 ( .A1(n15377), .A2(n15376), .ZN(n21279) );
  MUX2_X1 U18771 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21279), .S(
        n17063), .Z(n17072) );
  NOR2_X1 U18772 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15388), .ZN(n15395) );
  AOI22_X1 U18773 ( .A1(n17072), .A2(n15388), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15395), .ZN(n15390) );
  XNOR2_X1 U18774 ( .A(n14273), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15381) );
  INV_X1 U18775 ( .A(n15381), .ZN(n15420) );
  NAND2_X1 U18776 ( .A1(n15378), .A2(n15420), .ZN(n15384) );
  XNOR2_X1 U18777 ( .A(n15379), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15380) );
  AOI22_X1 U18778 ( .A1(n15382), .A2(n15381), .B1(n17060), .B2(n15380), .ZN(
        n15383) );
  OAI21_X1 U18779 ( .B1(n15386), .B2(n15384), .A(n15383), .ZN(n15385) );
  AOI21_X1 U18780 ( .B1(n21031), .B2(n15386), .A(n15385), .ZN(n15423) );
  NOR2_X1 U18781 ( .A1(n17063), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15387) );
  AOI21_X1 U18782 ( .B1(n15423), .B2(n17063), .A(n15387), .ZN(n17070) );
  AOI22_X1 U18783 ( .A1(n15395), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17070), .B2(n15388), .ZN(n15389) );
  NOR2_X1 U18784 ( .A1(n15390), .A2(n15389), .ZN(n17082) );
  INV_X1 U18785 ( .A(n14272), .ZN(n15391) );
  NAND2_X1 U18786 ( .A1(n17082), .A2(n15391), .ZN(n15399) );
  INV_X1 U18787 ( .A(n17063), .ZN(n15393) );
  AOI21_X1 U18788 ( .B1(n15393), .B2(n15392), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15397) );
  OAI21_X1 U18789 ( .B1(n20412), .B2(n15394), .A(n17063), .ZN(n15396) );
  AOI22_X1 U18790 ( .A1(n15397), .A2(n15396), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15395), .ZN(n17080) );
  NAND3_X1 U18791 ( .A1(n15399), .A2(n17080), .A3(n17131), .ZN(n17086) );
  NAND2_X1 U18792 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21041), .ZN(n15402) );
  NAND2_X1 U18793 ( .A1(n10782), .A2(n15402), .ZN(n15398) );
  OAI211_X1 U18794 ( .C1(n21184), .C2(n21093), .A(n17086), .B(n15398), .ZN(
        n15401) );
  AND3_X1 U18795 ( .A1(n15399), .A2(n17080), .A3(n20354), .ZN(n15400) );
  OAI21_X1 U18796 ( .B1(n17132), .B2(n15400), .A(n20763), .ZN(n20585) );
  MUX2_X1 U18797 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15401), .S(
        n20585), .Z(P1_U3478) );
  INV_X1 U18798 ( .A(n15402), .ZN(n15411) );
  INV_X1 U18799 ( .A(n9622), .ZN(n15409) );
  NOR2_X1 U18800 ( .A1(n21179), .A2(n21184), .ZN(n20719) );
  OAI21_X1 U18801 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9622), .A(n20719), 
        .ZN(n15403) );
  OAI21_X1 U18802 ( .B1(n15411), .B2(n14172), .A(n15403), .ZN(n15404) );
  MUX2_X1 U18803 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15404), .S(
        n20585), .Z(P1_U3477) );
  INV_X1 U18804 ( .A(n21031), .ZN(n20894) );
  NAND2_X1 U18805 ( .A1(n21179), .A2(n21186), .ZN(n21003) );
  NAND2_X1 U18806 ( .A1(n21003), .A2(n14162), .ZN(n20932) );
  OAI21_X1 U18807 ( .B1(n20719), .B2(n14162), .A(n20932), .ZN(n15405) );
  OAI21_X1 U18808 ( .B1(n15411), .B2(n20894), .A(n15405), .ZN(n15406) );
  MUX2_X1 U18809 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15406), .S(
        n20585), .Z(P1_U3476) );
  INV_X1 U18810 ( .A(n21091), .ZN(n15410) );
  OAI21_X1 U18811 ( .B1(n20994), .B2(n21089), .A(n15410), .ZN(n20933) );
  NOR2_X1 U18812 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21184), .ZN(n20961) );
  INV_X1 U18813 ( .A(n20961), .ZN(n20819) );
  INV_X1 U18814 ( .A(n20893), .ZN(n15412) );
  OAI22_X1 U18815 ( .A1(n15413), .A2(n20819), .B1(n15412), .B2(n15411), .ZN(
        n15414) );
  INV_X1 U18816 ( .A(n15414), .ZN(n15415) );
  OAI211_X1 U18817 ( .C1(n21003), .C2(n20866), .A(n20933), .B(n15415), .ZN(
        n15416) );
  MUX2_X1 U18818 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15416), .S(
        n20585), .Z(P1_U3475) );
  INV_X1 U18819 ( .A(n15417), .ZN(n15418) );
  AOI22_X1 U18820 ( .A1(n21276), .A2(n15420), .B1(n15419), .B2(n15418), .ZN(
        n15421) );
  OAI21_X1 U18821 ( .B1(n15423), .B2(n15422), .A(n15421), .ZN(n15424) );
  MUX2_X1 U18822 ( .A(n15424), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n21281), .Z(P1_U3472) );
  INV_X1 U18823 ( .A(n20217), .ZN(n15426) );
  AOI22_X1 U18824 ( .A1(n15426), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n15425), 
        .B2(n16495), .ZN(n15431) );
  NOR2_X1 U18825 ( .A1(n20224), .A2(n20145), .ZN(n15429) );
  NAND2_X1 U18826 ( .A1(n17153), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15427) );
  NAND2_X1 U18827 ( .A1(n15428), .A2(n15427), .ZN(n17156) );
  OAI22_X1 U18828 ( .A1(n15431), .A2(n15430), .B1(n15429), .B2(n17156), .ZN(
        n15437) );
  NAND2_X1 U18829 ( .A1(n15432), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16623) );
  NAND2_X1 U18830 ( .A1(n16623), .A2(n20318), .ZN(n15433) );
  OAI211_X1 U18831 ( .C1(n15435), .C2(n20224), .A(n15434), .B(n15433), .ZN(
        n15436) );
  MUX2_X1 U18832 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n15437), .S(n15436), 
        .Z(P2_U3610) );
  INV_X1 U18833 ( .A(n15791), .ZN(n15438) );
  NAND2_X1 U18834 ( .A1(n15438), .A2(n12854), .ZN(n15451) );
  NAND2_X1 U18835 ( .A1(n15442), .A2(n19532), .ZN(n15447) );
  AOI22_X1 U18836 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19554), .ZN(n15443) );
  OAI21_X1 U18837 ( .B1(n15444), .B2(n19529), .A(n15443), .ZN(n15445) );
  INV_X1 U18838 ( .A(n15445), .ZN(n15446) );
  OAI211_X1 U18839 ( .C1(n19551), .C2(n15903), .A(n15451), .B(n15450), .ZN(
        P2_U2826) );
  NOR2_X1 U18840 ( .A1(n15453), .A2(n15452), .ZN(n15454) );
  AOI21_X1 U18841 ( .B1(n15457), .B2(n9662), .A(n15456), .ZN(n16277) );
  NAND2_X1 U18842 ( .A1(n16277), .A2(n12854), .ZN(n15466) );
  AOI22_X1 U18843 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19554), .ZN(n15458) );
  OAI21_X1 U18844 ( .B1(n15459), .B2(n19529), .A(n15458), .ZN(n15464) );
  INV_X1 U18845 ( .A(n15460), .ZN(n15472) );
  AOI21_X1 U18846 ( .B1(n15772), .B2(n15462), .A(n15461), .ZN(n15463) );
  OAI211_X1 U18847 ( .C1(n19551), .C2(n16275), .A(n15466), .B(n15465), .ZN(
        P2_U2827) );
  INV_X1 U18848 ( .A(n15801), .ZN(n15477) );
  INV_X1 U18849 ( .A(n15467), .ZN(n15916) );
  AOI22_X1 U18850 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19554), .ZN(n15469) );
  NAND2_X1 U18851 ( .A1(n19547), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15468) );
  OAI211_X1 U18852 ( .C1(n15470), .C2(n19549), .A(n15469), .B(n15468), .ZN(
        n15475) );
  OAI21_X1 U18853 ( .B1(n9671), .B2(n15471), .A(n19563), .ZN(n15473) );
  AOI21_X1 U18854 ( .B1(n15772), .B2(n15473), .A(n15472), .ZN(n15474) );
  AOI211_X1 U18855 ( .C1(n15916), .C2(n19542), .A(n15475), .B(n15474), .ZN(
        n15476) );
  OAI21_X1 U18856 ( .B1(n15477), .B2(n19555), .A(n15476), .ZN(P2_U2828) );
  INV_X1 U18857 ( .A(n15812), .ZN(n15489) );
  INV_X1 U18858 ( .A(n15478), .ZN(n15499) );
  OAI21_X1 U18859 ( .B1(n15499), .B2(n15479), .A(n19563), .ZN(n15480) );
  AOI21_X1 U18860 ( .B1(n15772), .B2(n15480), .A(n9671), .ZN(n15487) );
  OAI211_X1 U18861 ( .C1(n15482), .C2(n15485), .A(n15481), .B(n19532), .ZN(
        n15484) );
  AOI22_X1 U18862 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19554), .ZN(n15483) );
  OAI211_X1 U18863 ( .C1(n19529), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15486) );
  AOI211_X1 U18864 ( .C1(n15924), .C2(n19542), .A(n15487), .B(n15486), .ZN(
        n15488) );
  OAI21_X1 U18865 ( .B1(n15489), .B2(n19555), .A(n15488), .ZN(P2_U2829) );
  NAND2_X1 U18866 ( .A1(n15490), .A2(n15491), .ZN(n15492) );
  NAND2_X1 U18867 ( .A1(n15493), .A2(n15492), .ZN(n16290) );
  NAND2_X1 U18868 ( .A1(n12744), .A2(n15494), .ZN(n15510) );
  AOI21_X1 U18869 ( .B1(n15496), .B2(n15510), .A(n15495), .ZN(n16282) );
  NAND2_X1 U18870 ( .A1(n16282), .A2(n12854), .ZN(n15505) );
  AOI22_X1 U18871 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19554), .ZN(n15497) );
  OAI21_X1 U18872 ( .B1(n15818), .B2(n19529), .A(n15497), .ZN(n15502) );
  INV_X1 U18873 ( .A(n15498), .ZN(n15515) );
  OAI21_X1 U18874 ( .B1(n15515), .B2(n16035), .A(n19563), .ZN(n15500) );
  AOI21_X1 U18875 ( .B1(n15772), .B2(n15500), .A(n15499), .ZN(n15501) );
  AOI211_X1 U18876 ( .C1(n19532), .C2(n15503), .A(n15502), .B(n15501), .ZN(
        n15504) );
  OAI211_X1 U18877 ( .C1(n19551), .C2(n16290), .A(n15505), .B(n15504), .ZN(
        P2_U2830) );
  OR2_X1 U18878 ( .A1(n15506), .A2(n15507), .ZN(n15508) );
  NAND2_X1 U18879 ( .A1(n15490), .A2(n15508), .ZN(n16300) );
  NAND2_X1 U18880 ( .A1(n12744), .A2(n15509), .ZN(n15525) );
  INV_X1 U18881 ( .A(n15510), .ZN(n15511) );
  AOI21_X1 U18882 ( .B1(n15512), .B2(n15525), .A(n15511), .ZN(n16303) );
  NAND2_X1 U18883 ( .A1(n16303), .A2(n12854), .ZN(n15521) );
  AOI22_X1 U18884 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19554), .ZN(n15513) );
  OAI21_X1 U18885 ( .B1(n15828), .B2(n19529), .A(n15513), .ZN(n15518) );
  INV_X1 U18886 ( .A(n15514), .ZN(n15532) );
  OAI21_X1 U18887 ( .B1(n15532), .B2(n16043), .A(n19563), .ZN(n15516) );
  AOI21_X1 U18888 ( .B1(n15772), .B2(n15516), .A(n15515), .ZN(n15517) );
  AOI211_X1 U18889 ( .C1(n19532), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n15520) );
  OAI211_X1 U18890 ( .C1(n19551), .C2(n16300), .A(n15521), .B(n15520), .ZN(
        P2_U2831) );
  AOI21_X1 U18891 ( .B1(n15522), .B2(n15545), .A(n15506), .ZN(n15523) );
  INV_X1 U18892 ( .A(n15523), .ZN(n16311) );
  NAND2_X1 U18893 ( .A1(n12744), .A2(n15524), .ZN(n15539) );
  INV_X1 U18894 ( .A(n15525), .ZN(n15526) );
  AOI21_X1 U18895 ( .B1(n15527), .B2(n15539), .A(n15526), .ZN(n16313) );
  NAND2_X1 U18896 ( .A1(n16313), .A2(n12854), .ZN(n15538) );
  AOI22_X1 U18897 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19554), .ZN(n15528) );
  OAI21_X1 U18898 ( .B1(n15529), .B2(n19529), .A(n15528), .ZN(n15535) );
  INV_X1 U18899 ( .A(n15530), .ZN(n15531) );
  OAI21_X1 U18900 ( .B1(n15531), .B2(n16047), .A(n19563), .ZN(n15533) );
  AOI21_X1 U18901 ( .B1(n15772), .B2(n15533), .A(n15532), .ZN(n15534) );
  AOI211_X1 U18902 ( .C1(n19532), .C2(n15536), .A(n15535), .B(n15534), .ZN(
        n15537) );
  OAI211_X1 U18903 ( .C1(n16311), .C2(n19551), .A(n15538), .B(n15537), .ZN(
        P2_U2832) );
  OAI21_X1 U18904 ( .B1(n15541), .B2(n15540), .A(n15539), .ZN(n16062) );
  NAND2_X1 U18905 ( .A1(n15543), .A2(n15542), .ZN(n15544) );
  NAND2_X1 U18906 ( .A1(n15545), .A2(n15544), .ZN(n16327) );
  INV_X1 U18907 ( .A(n16327), .ZN(n15555) );
  NOR2_X1 U18908 ( .A1(n15546), .A2(n19549), .ZN(n15554) );
  INV_X1 U18909 ( .A(n16064), .ZN(n15548) );
  AOI21_X1 U18910 ( .B1(n15547), .B2(n15548), .A(n19537), .ZN(n15549) );
  OAI21_X1 U18911 ( .B1(n15549), .B2(n15773), .A(n15530), .ZN(n15551) );
  AOI22_X1 U18912 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19554), .ZN(n15550) );
  OAI211_X1 U18913 ( .C1(n19529), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        n15553) );
  AOI211_X1 U18914 ( .C1(n15555), .C2(n19542), .A(n15554), .B(n15553), .ZN(
        n15556) );
  OAI21_X1 U18915 ( .B1(n16062), .B2(n19555), .A(n15556), .ZN(P2_U2833) );
  INV_X1 U18916 ( .A(n15845), .ZN(n15566) );
  INV_X1 U18917 ( .A(n15557), .ZN(n15957) );
  OAI211_X1 U18918 ( .C1(n15558), .C2(n15559), .A(n15547), .B(n19563), .ZN(
        n15562) );
  OAI22_X1 U18919 ( .A1(n21452), .A2(n19513), .B1(n19546), .B2(n20264), .ZN(
        n15560) );
  AOI21_X1 U18920 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n19547), .A(n15560), .ZN(
        n15561) );
  OAI211_X1 U18921 ( .C1(n19549), .C2(n15563), .A(n15562), .B(n15561), .ZN(
        n15564) );
  AOI21_X1 U18922 ( .B1(n15957), .B2(n19542), .A(n15564), .ZN(n15565) );
  OAI21_X1 U18923 ( .B1(n15566), .B2(n19555), .A(n15565), .ZN(P2_U2834) );
  NAND2_X1 U18924 ( .A1(n15851), .A2(n12854), .ZN(n15576) );
  OAI21_X1 U18925 ( .B1(n15567), .B2(n15571), .A(n19563), .ZN(n15570) );
  AOI22_X1 U18926 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19554), .ZN(n15569) );
  NAND2_X1 U18927 ( .A1(n19547), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15568) );
  OAI211_X1 U18928 ( .C1(n15558), .C2(n15570), .A(n15569), .B(n15568), .ZN(
        n15573) );
  NOR2_X1 U18929 ( .A1(n15772), .A2(n15571), .ZN(n15572) );
  AOI211_X1 U18930 ( .C1(n19532), .C2(n15574), .A(n15573), .B(n15572), .ZN(
        n15575) );
  OAI211_X1 U18931 ( .C1(n19551), .C2(n15962), .A(n15576), .B(n15575), .ZN(
        P2_U2835) );
  INV_X1 U18932 ( .A(n15578), .ZN(n15577) );
  NOR2_X1 U18933 ( .A1(n15784), .A2(n15577), .ZN(n15581) );
  OAI21_X1 U18934 ( .B1(n19537), .B2(n15578), .A(n15772), .ZN(n15580) );
  MUX2_X1 U18935 ( .A(n15581), .B(n15580), .S(n15579), .Z(n15588) );
  NAND2_X1 U18936 ( .A1(n15582), .A2(n19532), .ZN(n15585) );
  OAI21_X1 U18937 ( .B1(n19546), .B2(n20260), .A(n16032), .ZN(n15583) );
  AOI21_X1 U18938 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19548), .A(
        n15583), .ZN(n15584) );
  OAI211_X1 U18939 ( .C1(n19529), .C2(n15586), .A(n15585), .B(n15584), .ZN(
        n15587) );
  AOI211_X1 U18940 ( .C1(n15972), .C2(n19542), .A(n15588), .B(n15587), .ZN(
        n15589) );
  OAI21_X1 U18941 ( .B1(n15858), .B2(n19555), .A(n15589), .ZN(P2_U2836) );
  NOR2_X1 U18942 ( .A1(n15591), .A2(n15590), .ZN(n15592) );
  OR2_X1 U18943 ( .A1(n15593), .A2(n15592), .ZN(n16339) );
  OAI21_X1 U18944 ( .B1(n19546), .B2(n16074), .A(n16032), .ZN(n15594) );
  AOI21_X1 U18945 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19548), .A(
        n15594), .ZN(n15595) );
  OAI21_X1 U18946 ( .B1(n15596), .B2(n19529), .A(n15595), .ZN(n15602) );
  INV_X1 U18947 ( .A(n15598), .ZN(n15597) );
  NOR2_X1 U18948 ( .A1(n15784), .A2(n15597), .ZN(n15600) );
  OAI21_X1 U18949 ( .B1(n19537), .B2(n15598), .A(n15772), .ZN(n15599) );
  MUX2_X1 U18950 ( .A(n15600), .B(n15599), .S(n16077), .Z(n15601) );
  AOI211_X1 U18951 ( .C1(n19532), .C2(n15603), .A(n15602), .B(n15601), .ZN(
        n15608) );
  NOR2_X1 U18952 ( .A1(n14253), .A2(n15604), .ZN(n15605) );
  OR2_X1 U18953 ( .A1(n9640), .A2(n15605), .ZN(n16333) );
  INV_X1 U18954 ( .A(n16333), .ZN(n15606) );
  NAND2_X1 U18955 ( .A1(n15606), .A2(n12854), .ZN(n15607) );
  OAI211_X1 U18956 ( .C1(n19551), .C2(n16339), .A(n15608), .B(n15607), .ZN(
        P2_U2837) );
  NAND2_X1 U18957 ( .A1(n16087), .A2(n12854), .ZN(n15619) );
  NOR2_X1 U18958 ( .A1(n15683), .A2(n15609), .ZN(n15610) );
  XNOR2_X1 U18959 ( .A(n15610), .B(n16084), .ZN(n15617) );
  NOR2_X1 U18960 ( .A1(n15611), .A2(n19549), .ZN(n15616) );
  INV_X1 U18961 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15614) );
  AOI21_X1 U18962 ( .B1(n19554), .B2(P2_REIP_REG_17__SCAN_IN), .A(n19527), 
        .ZN(n15613) );
  NAND2_X1 U18963 ( .A1(n19547), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15612) );
  OAI211_X1 U18964 ( .C1(n19513), .C2(n15614), .A(n15613), .B(n15612), .ZN(
        n15615) );
  AOI211_X1 U18965 ( .C1(n15617), .C2(n19563), .A(n15616), .B(n15615), .ZN(
        n15618) );
  OAI211_X1 U18966 ( .C1(n19551), .C2(n15620), .A(n15619), .B(n15618), .ZN(
        P2_U2838) );
  NAND2_X1 U18967 ( .A1(n15621), .A2(n15622), .ZN(n15623) );
  NAND2_X1 U18968 ( .A1(n9628), .A2(n15623), .ZN(n16349) );
  INV_X1 U18969 ( .A(n15624), .ZN(n15634) );
  INV_X1 U18970 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15627) );
  AOI21_X1 U18971 ( .B1(n19554), .B2(P2_REIP_REG_16__SCAN_IN), .A(n19553), 
        .ZN(n15626) );
  NAND2_X1 U18972 ( .A1(n19547), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15625) );
  OAI211_X1 U18973 ( .C1(n19513), .C2(n15627), .A(n15626), .B(n15625), .ZN(
        n15633) );
  OAI21_X1 U18974 ( .B1(n19537), .B2(n15628), .A(n15772), .ZN(n15631) );
  INV_X1 U18975 ( .A(n15628), .ZN(n15629) );
  NOR2_X1 U18976 ( .A1(n15784), .A2(n15629), .ZN(n15630) );
  MUX2_X1 U18977 ( .A(n15631), .B(n15630), .S(n16093), .Z(n15632) );
  AOI211_X1 U18978 ( .C1(n19532), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        n15639) );
  INV_X1 U18979 ( .A(n15635), .ZN(n15636) );
  AOI21_X1 U18980 ( .B1(n15637), .B2(n14145), .A(n15636), .ZN(n16347) );
  NAND2_X1 U18981 ( .A1(n16347), .A2(n19542), .ZN(n15638) );
  OAI211_X1 U18982 ( .C1(n19555), .C2(n16349), .A(n15639), .B(n15638), .ZN(
        P2_U2839) );
  OR2_X1 U18983 ( .A1(n15640), .A2(n15641), .ZN(n15642) );
  NAND2_X1 U18984 ( .A1(n15621), .A2(n15642), .ZN(n16357) );
  NAND2_X1 U18985 ( .A1(n15733), .A2(n15643), .ZN(n15646) );
  INV_X1 U18986 ( .A(n15643), .ZN(n15644) );
  AOI21_X1 U18987 ( .B1(n19563), .B2(n15644), .A(n15773), .ZN(n15645) );
  MUX2_X1 U18988 ( .A(n15646), .B(n15645), .S(n16109), .Z(n15650) );
  AOI21_X1 U18989 ( .B1(n19554), .B2(P2_REIP_REG_15__SCAN_IN), .A(n19553), 
        .ZN(n15647) );
  OAI21_X1 U18990 ( .B1(n19513), .B2(n16107), .A(n15647), .ZN(n15648) );
  AOI21_X1 U18991 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n19547), .A(n15648), .ZN(
        n15649) );
  OAI211_X1 U18992 ( .C1(n19549), .C2(n15651), .A(n15650), .B(n15649), .ZN(
        n15652) );
  AOI21_X1 U18993 ( .B1(n16358), .B2(n19542), .A(n15652), .ZN(n15653) );
  OAI21_X1 U18994 ( .B1(n16357), .B2(n19555), .A(n15653), .ZN(P2_U2840) );
  NOR2_X1 U18995 ( .A1(n15655), .A2(n15654), .ZN(n15656) );
  OR2_X1 U18996 ( .A1(n15640), .A2(n15656), .ZN(n16374) );
  AOI21_X1 U18997 ( .B1(n19563), .B2(n15657), .A(n15773), .ZN(n15659) );
  MUX2_X1 U18998 ( .A(n15659), .B(n15658), .S(n16120), .Z(n15667) );
  NAND2_X1 U18999 ( .A1(n15660), .A2(n19532), .ZN(n15663) );
  OAI21_X1 U19000 ( .B1(n19546), .B2(n16119), .A(n16032), .ZN(n15661) );
  AOI21_X1 U19001 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19548), .A(
        n15661), .ZN(n15662) );
  OAI211_X1 U19002 ( .C1(n19529), .C2(n15664), .A(n15663), .B(n15662), .ZN(
        n15665) );
  AOI21_X1 U19003 ( .B1(n16372), .B2(n19542), .A(n15665), .ZN(n15666) );
  OAI211_X1 U19004 ( .C1(n19555), .C2(n16374), .A(n15667), .B(n15666), .ZN(
        P2_U2841) );
  NAND2_X1 U19005 ( .A1(n15669), .A2(n19563), .ZN(n15668) );
  NAND2_X1 U19006 ( .A1(n15772), .A2(n15668), .ZN(n15671) );
  NOR2_X1 U19007 ( .A1(n15784), .A2(n15669), .ZN(n15670) );
  MUX2_X1 U19008 ( .A(n15671), .B(n15670), .S(n16169), .Z(n15681) );
  INV_X1 U19009 ( .A(n15672), .ZN(n15677) );
  AOI21_X1 U19010 ( .B1(n19554), .B2(P2_REIP_REG_10__SCAN_IN), .A(n19553), 
        .ZN(n15674) );
  NAND2_X1 U19011 ( .A1(n19547), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15673) );
  OAI211_X1 U19012 ( .C1(n19513), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        n15676) );
  AOI21_X1 U19013 ( .B1(n15677), .B2(n19532), .A(n15676), .ZN(n15679) );
  NAND2_X1 U19014 ( .A1(n16426), .A2(n19542), .ZN(n15678) );
  OAI211_X1 U19015 ( .C1(n16427), .C2(n19555), .A(n15679), .B(n15678), .ZN(
        n15680) );
  NOR2_X1 U19016 ( .A1(n15683), .A2(n15682), .ZN(n15684) );
  XOR2_X1 U19017 ( .A(n16182), .B(n15684), .Z(n15692) );
  NAND2_X1 U19018 ( .A1(n16440), .A2(n19542), .ZN(n15688) );
  NAND2_X1 U19019 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15685) );
  OAI211_X1 U19020 ( .C1(n20245), .C2(n19546), .A(n15685), .B(n16032), .ZN(
        n15686) );
  AOI21_X1 U19021 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n19547), .A(n15686), .ZN(
        n15687) );
  OAI211_X1 U19022 ( .C1(n19549), .C2(n15689), .A(n15688), .B(n15687), .ZN(
        n15690) );
  AOI21_X1 U19023 ( .B1(n16441), .B2(n12854), .A(n15690), .ZN(n15691) );
  OAI21_X1 U19024 ( .B1(n15692), .B2(n19537), .A(n15691), .ZN(P2_U2846) );
  INV_X1 U19025 ( .A(n15694), .ZN(n15693) );
  NOR2_X1 U19026 ( .A1(n15784), .A2(n15693), .ZN(n15697) );
  OAI21_X1 U19027 ( .B1(n19537), .B2(n15694), .A(n15772), .ZN(n15696) );
  MUX2_X1 U19028 ( .A(n15697), .B(n15696), .S(n15695), .Z(n15710) );
  NAND2_X1 U19029 ( .A1(n13879), .A2(n15698), .ZN(n15699) );
  AND2_X1 U19030 ( .A1(n15700), .A2(n15699), .ZN(n16455) );
  NAND2_X1 U19031 ( .A1(n16455), .A2(n12854), .ZN(n15708) );
  INV_X1 U19032 ( .A(n15701), .ZN(n15706) );
  INV_X1 U19033 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15704) );
  AOI21_X1 U19034 ( .B1(n19554), .B2(P2_REIP_REG_8__SCAN_IN), .A(n19553), .ZN(
        n15703) );
  NAND2_X1 U19035 ( .A1(n19547), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15702) );
  OAI211_X1 U19036 ( .C1(n19513), .C2(n15704), .A(n15703), .B(n15702), .ZN(
        n15705) );
  AOI21_X1 U19037 ( .B1(n15706), .B2(n19532), .A(n15705), .ZN(n15707) );
  OAI211_X1 U19038 ( .C1(n16453), .C2(n19551), .A(n15708), .B(n15707), .ZN(
        n15709) );
  INV_X1 U19039 ( .A(n15711), .ZN(n19538) );
  NOR2_X1 U19040 ( .A1(n15784), .A2(n19538), .ZN(n15713) );
  OAI21_X1 U19041 ( .B1(n19537), .B2(n15711), .A(n15772), .ZN(n15712) );
  MUX2_X1 U19042 ( .A(n15713), .B(n15712), .S(n16199), .Z(n15720) );
  NAND2_X1 U19043 ( .A1(n16209), .A2(n12854), .ZN(n15718) );
  AOI22_X1 U19044 ( .A1(n19547), .A2(P2_EBX_REG_7__SCAN_IN), .B1(n19532), .B2(
        n15714), .ZN(n15715) );
  OAI211_X1 U19045 ( .C1(n20241), .C2(n19546), .A(n15715), .B(n16032), .ZN(
        n15716) );
  AOI21_X1 U19046 ( .B1(n19548), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n15716), .ZN(n15717) );
  OAI211_X1 U19047 ( .C1(n17138), .C2(n19551), .A(n15718), .B(n15717), .ZN(
        n15719) );
  NAND2_X1 U19048 ( .A1(n19559), .A2(n19562), .ZN(n15721) );
  XOR2_X1 U19049 ( .A(n15721), .B(n16219), .Z(n15730) );
  NOR2_X1 U19050 ( .A1(n19529), .A2(n12350), .ZN(n15723) );
  OAI21_X1 U19051 ( .B1(n19546), .B2(n11827), .A(n16032), .ZN(n15722) );
  AOI211_X1 U19052 ( .C1(n19548), .C2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n15723), .B(n15722), .ZN(n15724) );
  OAI21_X1 U19053 ( .B1(n15725), .B2(n19549), .A(n15724), .ZN(n15727) );
  NOR2_X1 U19054 ( .A1(n16223), .A2(n19555), .ZN(n15726) );
  AOI211_X1 U19055 ( .C1(n19542), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        n15729) );
  OAI21_X1 U19056 ( .B1(n15730), .B2(n19537), .A(n15729), .ZN(P2_U2850) );
  AOI21_X1 U19057 ( .B1(n19563), .B2(n15731), .A(n15773), .ZN(n15735) );
  INV_X1 U19058 ( .A(n15731), .ZN(n15732) );
  NAND2_X1 U19059 ( .A1(n15733), .A2(n15732), .ZN(n15734) );
  MUX2_X1 U19060 ( .A(n15735), .B(n15734), .S(n16248), .Z(n15746) );
  AOI22_X1 U19061 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19554), .B2(P2_REIP_REG_3__SCAN_IN), .ZN(n15737) );
  OR2_X1 U19062 ( .A1(n19529), .A2(n12347), .ZN(n15736) );
  OAI211_X1 U19063 ( .C1(n19549), .C2(n15738), .A(n15737), .B(n15736), .ZN(
        n15744) );
  NAND2_X1 U19064 ( .A1(n15741), .A2(n15740), .ZN(n15742) );
  NAND2_X1 U19065 ( .A1(n15739), .A2(n15742), .ZN(n20310) );
  NOR2_X1 U19066 ( .A1(n20310), .A2(n19551), .ZN(n15743) );
  AOI211_X1 U19067 ( .C1(n16257), .C2(n12854), .A(n15744), .B(n15743), .ZN(
        n15745) );
  OAI211_X1 U19068 ( .C1(n19692), .C2(n19556), .A(n15746), .B(n15745), .ZN(
        P2_U2852) );
  NAND2_X1 U19069 ( .A1(n15767), .A2(n19563), .ZN(n15747) );
  NAND2_X1 U19070 ( .A1(n15772), .A2(n15747), .ZN(n15750) );
  NOR2_X1 U19071 ( .A1(n15784), .A2(n15767), .ZN(n15749) );
  MUX2_X1 U19072 ( .A(n15750), .B(n15749), .S(n15748), .Z(n15751) );
  INV_X1 U19073 ( .A(n15751), .ZN(n15758) );
  AOI22_X1 U19074 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19554), .ZN(n15753) );
  NAND2_X1 U19075 ( .A1(n19547), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n15752) );
  OAI211_X1 U19076 ( .C1(n19549), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        n15756) );
  NOR2_X1 U19077 ( .A1(n16572), .A2(n19555), .ZN(n15755) );
  AOI211_X1 U19078 ( .C1(n19542), .C2(n19664), .A(n15756), .B(n15755), .ZN(
        n15757) );
  OAI211_X1 U19079 ( .C1(n19556), .C2(n20299), .A(n15758), .B(n15757), .ZN(
        P2_U2853) );
  AOI22_X1 U19080 ( .A1(n19532), .A2(n16260), .B1(n19554), .B2(
        P2_REIP_REG_1__SCAN_IN), .ZN(n15760) );
  NAND2_X1 U19081 ( .A1(n19547), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n15759) );
  OAI211_X1 U19082 ( .C1(n15761), .C2(n19513), .A(n15760), .B(n15759), .ZN(
        n15762) );
  AOI21_X1 U19083 ( .B1(n19542), .B2(n15763), .A(n15762), .ZN(n15764) );
  OAI21_X1 U19084 ( .B1(n16486), .B2(n19555), .A(n15764), .ZN(n15770) );
  AND2_X1 U19085 ( .A1(n15765), .A2(n16504), .ZN(n15766) );
  NOR2_X1 U19086 ( .A1(n15767), .A2(n15766), .ZN(n15768) );
  NAND2_X1 U19087 ( .A1(n19559), .A2(n15768), .ZN(n16513) );
  NOR2_X1 U19088 ( .A1(n16513), .A2(n19537), .ZN(n15769) );
  AOI211_X1 U19089 ( .C1(n15781), .C2(n20308), .A(n15770), .B(n15769), .ZN(
        n15771) );
  OAI21_X1 U19090 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n15772), .A(
        n15771), .ZN(P2_U2854) );
  INV_X1 U19091 ( .A(n16504), .ZN(n15785) );
  OAI21_X1 U19092 ( .B1(n15773), .B2(n19548), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15783) );
  INV_X1 U19093 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19506) );
  OAI22_X1 U19094 ( .A1(n19546), .A2(n19506), .B1(n19551), .B2(n15774), .ZN(
        n15775) );
  AOI21_X1 U19095 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19547), .A(n15775), .ZN(
        n15778) );
  NAND2_X1 U19096 ( .A1(n19532), .A2(n15776), .ZN(n15777) );
  OAI211_X1 U19097 ( .C1(n15779), .C2(n19555), .A(n15778), .B(n15777), .ZN(
        n15780) );
  AOI21_X1 U19098 ( .B1(n19691), .B2(n15781), .A(n15780), .ZN(n15782) );
  OAI211_X1 U19099 ( .C1(n15785), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        P2_U2855) );
  OR2_X1 U19100 ( .A1(n15787), .A2(n15786), .ZN(n15896) );
  NAND3_X1 U19101 ( .A1(n15896), .A2(n15788), .A3(n15883), .ZN(n15790) );
  NAND2_X1 U19102 ( .A1(n19570), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15789) );
  OAI211_X1 U19103 ( .C1(n15791), .C2(n19570), .A(n15790), .B(n15789), .ZN(
        P2_U2858) );
  NOR2_X1 U19104 ( .A1(n15793), .A2(n15792), .ZN(n15795) );
  XNOR2_X1 U19105 ( .A(n15795), .B(n15794), .ZN(n15910) );
  NAND2_X1 U19106 ( .A1(n16277), .A2(n19575), .ZN(n15797) );
  NAND2_X1 U19107 ( .A1(n19570), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15796) );
  OAI211_X1 U19108 ( .C1(n15910), .C2(n19571), .A(n15797), .B(n15796), .ZN(
        P2_U2859) );
  OAI21_X1 U19109 ( .B1(n15798), .B2(n15800), .A(n15799), .ZN(n15918) );
  NAND2_X1 U19110 ( .A1(n15801), .A2(n19575), .ZN(n15803) );
  NAND2_X1 U19111 ( .A1(n19570), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15802) );
  OAI211_X1 U19112 ( .C1(n15918), .C2(n19571), .A(n15803), .B(n15802), .ZN(
        P2_U2860) );
  AND2_X1 U19113 ( .A1(n15804), .A2(n15817), .ZN(n15815) );
  NOR2_X1 U19114 ( .A1(n15815), .A2(n15805), .ZN(n15811) );
  NOR2_X1 U19115 ( .A1(n15807), .A2(n15806), .ZN(n15808) );
  XNOR2_X1 U19116 ( .A(n15809), .B(n15808), .ZN(n15810) );
  XNOR2_X1 U19117 ( .A(n15811), .B(n15810), .ZN(n15926) );
  NAND2_X1 U19118 ( .A1(n15812), .A2(n19575), .ZN(n15814) );
  NAND2_X1 U19119 ( .A1(n19570), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15813) );
  OAI211_X1 U19120 ( .C1(n15926), .C2(n19571), .A(n15814), .B(n15813), .ZN(
        P2_U2861) );
  INV_X1 U19121 ( .A(n15815), .ZN(n15816) );
  OAI21_X1 U19122 ( .B1(n15817), .B2(n15804), .A(n15816), .ZN(n15933) );
  NOR2_X1 U19123 ( .A1(n19575), .A2(n15818), .ZN(n15819) );
  AOI21_X1 U19124 ( .B1(n16282), .B2(n19575), .A(n15819), .ZN(n15820) );
  OAI21_X1 U19125 ( .B1(n19571), .B2(n15933), .A(n15820), .ZN(P2_U2862) );
  INV_X1 U19126 ( .A(n15821), .ZN(n15839) );
  XOR2_X1 U19127 ( .A(n15823), .B(n15821), .Z(n15833) );
  NAND2_X1 U19128 ( .A1(n12004), .A2(n15822), .ZN(n15832) );
  NOR2_X1 U19129 ( .A1(n15833), .A2(n15832), .ZN(n15831) );
  AOI21_X1 U19130 ( .B1(n15839), .B2(n15823), .A(n15831), .ZN(n15827) );
  XNOR2_X1 U19131 ( .A(n15825), .B(n15824), .ZN(n15826) );
  XNOR2_X1 U19132 ( .A(n15827), .B(n15826), .ZN(n15940) );
  NOR2_X1 U19133 ( .A1(n19575), .A2(n15828), .ZN(n15829) );
  AOI21_X1 U19134 ( .B1(n16303), .B2(n19575), .A(n15829), .ZN(n15830) );
  OAI21_X1 U19135 ( .B1(n15940), .B2(n19571), .A(n15830), .ZN(P2_U2863) );
  INV_X1 U19136 ( .A(n16313), .ZN(n15836) );
  AOI21_X1 U19137 ( .B1(n15833), .B2(n15832), .A(n15831), .ZN(n15944) );
  NAND2_X1 U19138 ( .A1(n15944), .A2(n15883), .ZN(n15835) );
  NAND2_X1 U19139 ( .A1(n19570), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15834) );
  OAI211_X1 U19140 ( .C1(n15836), .C2(n19570), .A(n15835), .B(n15834), .ZN(
        P2_U2864) );
  AOI21_X1 U19141 ( .B1(n15840), .B2(n15838), .A(n15839), .ZN(n15950) );
  NAND2_X1 U19142 ( .A1(n15950), .A2(n15883), .ZN(n15842) );
  NAND2_X1 U19143 ( .A1(n19570), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15841) );
  OAI211_X1 U19144 ( .C1(n16062), .C2(n19570), .A(n15842), .B(n15841), .ZN(
        P2_U2865) );
  OAI21_X1 U19145 ( .B1(n15843), .B2(n15844), .A(n15838), .ZN(n15959) );
  NAND2_X1 U19146 ( .A1(n15845), .A2(n19575), .ZN(n15847) );
  NAND2_X1 U19147 ( .A1(n19570), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15846) );
  OAI211_X1 U19148 ( .C1(n15959), .C2(n19571), .A(n15847), .B(n15846), .ZN(
        P2_U2866) );
  NOR2_X1 U19149 ( .A1(n15848), .A2(n15849), .ZN(n15850) );
  OR2_X1 U19150 ( .A1(n15843), .A2(n15850), .ZN(n15966) );
  NAND2_X1 U19151 ( .A1(n15851), .A2(n19575), .ZN(n15853) );
  NAND2_X1 U19152 ( .A1(n19570), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15852) );
  OAI211_X1 U19153 ( .C1(n15966), .C2(n19571), .A(n15853), .B(n15852), .ZN(
        P2_U2867) );
  AND2_X1 U19154 ( .A1(n15859), .A2(n15854), .ZN(n15855) );
  NOR2_X1 U19155 ( .A1(n15848), .A2(n15855), .ZN(n15967) );
  NAND2_X1 U19156 ( .A1(n15967), .A2(n15883), .ZN(n15857) );
  NAND2_X1 U19157 ( .A1(n19570), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15856) );
  OAI211_X1 U19158 ( .C1(n15858), .C2(n19570), .A(n15857), .B(n15856), .ZN(
        P2_U2868) );
  INV_X1 U19159 ( .A(n15859), .ZN(n15860) );
  AOI21_X1 U19160 ( .B1(n15862), .B2(n15861), .A(n15860), .ZN(n15978) );
  NAND2_X1 U19161 ( .A1(n15978), .A2(n15883), .ZN(n15864) );
  NAND2_X1 U19162 ( .A1(n19570), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15863) );
  OAI211_X1 U19163 ( .C1(n16333), .C2(n19570), .A(n15864), .B(n15863), .ZN(
        P2_U2869) );
  NAND2_X1 U19164 ( .A1(n16087), .A2(n19575), .ZN(n15866) );
  NAND2_X1 U19165 ( .A1(n19570), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15865) );
  OAI211_X1 U19166 ( .C1(n15867), .C2(n19571), .A(n15866), .B(n15865), .ZN(
        P2_U2870) );
  NAND2_X1 U19167 ( .A1(n15886), .A2(n15885), .ZN(n15884) );
  INV_X1 U19168 ( .A(n15879), .ZN(n15868) );
  NOR2_X1 U19169 ( .A1(n15884), .A2(n15868), .ZN(n15877) );
  AOI21_X1 U19170 ( .B1(n15877), .B2(n15874), .A(n15869), .ZN(n15871) );
  NOR2_X1 U19171 ( .A1(n15871), .A2(n15870), .ZN(n15982) );
  NAND2_X1 U19172 ( .A1(n15982), .A2(n15883), .ZN(n15873) );
  NAND2_X1 U19173 ( .A1(n19570), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15872) );
  OAI211_X1 U19174 ( .C1(n16349), .C2(n19570), .A(n15873), .B(n15872), .ZN(
        P2_U2871) );
  XNOR2_X1 U19175 ( .A(n15877), .B(n15874), .ZN(n15876) );
  MUX2_X1 U19176 ( .A(n16357), .B(n12528), .S(n19570), .Z(n15875) );
  OAI21_X1 U19177 ( .B1(n15876), .B2(n19571), .A(n15875), .ZN(P2_U2872) );
  INV_X1 U19178 ( .A(n15884), .ZN(n15880) );
  INV_X1 U19179 ( .A(n15877), .ZN(n15878) );
  OAI211_X1 U19180 ( .C1(n15880), .C2(n15879), .A(n15878), .B(n15883), .ZN(
        n15882) );
  NAND2_X1 U19181 ( .A1(n19570), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15881) );
  OAI211_X1 U19182 ( .C1(n16374), .C2(n19570), .A(n15882), .B(n15881), .ZN(
        P2_U2873) );
  NAND2_X1 U19183 ( .A1(n16130), .A2(n19575), .ZN(n15888) );
  OAI211_X1 U19184 ( .C1(n15886), .C2(n15885), .A(n15884), .B(n15883), .ZN(
        n15887) );
  OAI211_X1 U19185 ( .C1(n19575), .C2(n12360), .A(n15888), .B(n15887), .ZN(
        P2_U2874) );
  INV_X1 U19186 ( .A(n16455), .ZN(n15889) );
  NOR2_X1 U19187 ( .A1(n15889), .A2(n19570), .ZN(n15894) );
  AOI211_X1 U19188 ( .C1(n15892), .C2(n15891), .A(n19571), .B(n15890), .ZN(
        n15893) );
  AOI211_X1 U19189 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19570), .A(n15894), .B(
        n15893), .ZN(n15895) );
  INV_X1 U19190 ( .A(n15895), .ZN(P2_U2879) );
  NAND3_X1 U19191 ( .A1(n15896), .A2(n15788), .A3(n19582), .ZN(n15902) );
  NAND2_X1 U19192 ( .A1(n15984), .A2(BUF2_REG_29__SCAN_IN), .ZN(n15900) );
  NAND2_X1 U19193 ( .A1(n15983), .A2(BUF1_REG_29__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U19194 ( .A1(n15985), .A2(n15897), .B1(n16010), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15898) );
  AND3_X1 U19195 ( .A1(n15900), .A2(n15899), .A3(n15898), .ZN(n15901) );
  OAI211_X1 U19196 ( .C1(n15903), .C2(n15981), .A(n15902), .B(n15901), .ZN(
        P2_U2890) );
  NAND2_X1 U19197 ( .A1(n15983), .A2(BUF1_REG_28__SCAN_IN), .ZN(n15906) );
  AOI22_X1 U19198 ( .A1(n15985), .A2(n15904), .B1(n16010), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15905) );
  NAND2_X1 U19199 ( .A1(n15906), .A2(n15905), .ZN(n15908) );
  NOR2_X1 U19200 ( .A1(n16275), .A2(n15981), .ZN(n15907) );
  OAI21_X1 U19201 ( .B1(n15910), .B2(n16013), .A(n15909), .ZN(P2_U2891) );
  NAND2_X1 U19202 ( .A1(n15984), .A2(BUF2_REG_27__SCAN_IN), .ZN(n15914) );
  NAND2_X1 U19203 ( .A1(n15983), .A2(BUF1_REG_27__SCAN_IN), .ZN(n15913) );
  AOI22_X1 U19204 ( .A1(n15985), .A2(n15911), .B1(n16010), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15912) );
  NAND3_X1 U19205 ( .A1(n15914), .A2(n15913), .A3(n15912), .ZN(n15915) );
  AOI21_X1 U19206 ( .B1(n15916), .B2(n19578), .A(n15915), .ZN(n15917) );
  OAI21_X1 U19207 ( .B1(n16013), .B2(n15918), .A(n15917), .ZN(P2_U2892) );
  NAND2_X1 U19208 ( .A1(n15984), .A2(BUF2_REG_26__SCAN_IN), .ZN(n15922) );
  NAND2_X1 U19209 ( .A1(n15983), .A2(BUF1_REG_26__SCAN_IN), .ZN(n15921) );
  AOI22_X1 U19210 ( .A1(n15985), .A2(n15919), .B1(n16010), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15920) );
  NAND3_X1 U19211 ( .A1(n15922), .A2(n15921), .A3(n15920), .ZN(n15923) );
  AOI21_X1 U19212 ( .B1(n15924), .B2(n19578), .A(n15923), .ZN(n15925) );
  OAI21_X1 U19213 ( .B1(n15926), .B2(n16013), .A(n15925), .ZN(P2_U2893) );
  NAND2_X1 U19214 ( .A1(n15983), .A2(BUF1_REG_25__SCAN_IN), .ZN(n15929) );
  AOI22_X1 U19215 ( .A1(n15985), .A2(n15927), .B1(n16010), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15928) );
  NAND2_X1 U19216 ( .A1(n15929), .A2(n15928), .ZN(n15931) );
  NOR2_X1 U19217 ( .A1(n16290), .A2(n15981), .ZN(n15930) );
  AOI211_X1 U19218 ( .C1(n15984), .C2(BUF2_REG_25__SCAN_IN), .A(n15931), .B(
        n15930), .ZN(n15932) );
  OAI21_X1 U19219 ( .B1(n16013), .B2(n15933), .A(n15932), .ZN(P2_U2894) );
  NAND2_X1 U19220 ( .A1(n15983), .A2(BUF1_REG_24__SCAN_IN), .ZN(n15936) );
  AOI22_X1 U19221 ( .A1(n15985), .A2(n15934), .B1(n16010), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15935) );
  NAND2_X1 U19222 ( .A1(n15936), .A2(n15935), .ZN(n15938) );
  NOR2_X1 U19223 ( .A1(n16300), .A2(n15981), .ZN(n15937) );
  AOI211_X1 U19224 ( .C1(n15984), .C2(BUF2_REG_24__SCAN_IN), .A(n15938), .B(
        n15937), .ZN(n15939) );
  OAI21_X1 U19225 ( .B1(n15940), .B2(n16013), .A(n15939), .ZN(P2_U2895) );
  NAND2_X1 U19226 ( .A1(n15983), .A2(BUF1_REG_23__SCAN_IN), .ZN(n15943) );
  NAND2_X1 U19227 ( .A1(n15984), .A2(BUF2_REG_23__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U19228 ( .A1(n15985), .A2(n16561), .B1(n16010), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15941) );
  AND3_X1 U19229 ( .A1(n15943), .A2(n15942), .A3(n15941), .ZN(n15946) );
  NAND2_X1 U19230 ( .A1(n15944), .A2(n19582), .ZN(n15945) );
  OAI211_X1 U19231 ( .C1(n16311), .C2(n15981), .A(n15946), .B(n15945), .ZN(
        P2_U2896) );
  NAND2_X1 U19232 ( .A1(n15983), .A2(BUF1_REG_22__SCAN_IN), .ZN(n15949) );
  NAND2_X1 U19233 ( .A1(n15984), .A2(BUF2_REG_22__SCAN_IN), .ZN(n15948) );
  AOI22_X1 U19234 ( .A1(n15985), .A2(n16557), .B1(n16010), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15947) );
  AND3_X1 U19235 ( .A1(n15949), .A2(n15948), .A3(n15947), .ZN(n15952) );
  NAND2_X1 U19236 ( .A1(n15950), .A2(n19582), .ZN(n15951) );
  OAI211_X1 U19237 ( .C1(n16327), .C2(n15981), .A(n15952), .B(n15951), .ZN(
        P2_U2897) );
  NAND2_X1 U19238 ( .A1(n15983), .A2(BUF1_REG_21__SCAN_IN), .ZN(n15955) );
  NAND2_X1 U19239 ( .A1(n15984), .A2(BUF2_REG_21__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19240 ( .A1(n15985), .A2(n16552), .B1(n16010), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15953) );
  NAND3_X1 U19241 ( .A1(n15955), .A2(n15954), .A3(n15953), .ZN(n15956) );
  AOI21_X1 U19242 ( .B1(n15957), .B2(n19578), .A(n15956), .ZN(n15958) );
  OAI21_X1 U19243 ( .B1(n16013), .B2(n15959), .A(n15958), .ZN(P2_U2898) );
  NAND2_X1 U19244 ( .A1(n15984), .A2(BUF2_REG_20__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19245 ( .A1(n15985), .A2(n19576), .B1(n16010), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15960) );
  NAND2_X1 U19246 ( .A1(n15961), .A2(n15960), .ZN(n15964) );
  NOR2_X1 U19247 ( .A1(n15962), .A2(n15981), .ZN(n15963) );
  AOI211_X1 U19248 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n15983), .A(n15964), .B(
        n15963), .ZN(n15965) );
  OAI21_X1 U19249 ( .B1(n16013), .B2(n15966), .A(n15965), .ZN(P2_U2899) );
  INV_X1 U19250 ( .A(n15967), .ZN(n15974) );
  NAND2_X1 U19251 ( .A1(n15983), .A2(BUF1_REG_19__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U19252 ( .A1(n15984), .A2(BUF2_REG_19__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19253 ( .A1(n15985), .A2(n16545), .B1(n16010), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15968) );
  NAND3_X1 U19254 ( .A1(n15970), .A2(n15969), .A3(n15968), .ZN(n15971) );
  AOI21_X1 U19255 ( .B1(n15972), .B2(n19578), .A(n15971), .ZN(n15973) );
  OAI21_X1 U19256 ( .B1(n16013), .B2(n15974), .A(n15973), .ZN(P2_U2900) );
  NAND2_X1 U19257 ( .A1(n15983), .A2(BUF1_REG_18__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U19258 ( .A1(n15984), .A2(BUF2_REG_18__SCAN_IN), .ZN(n15976) );
  AOI22_X1 U19259 ( .A1(n15985), .A2(n16541), .B1(n16010), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15975) );
  AND3_X1 U19260 ( .A1(n15977), .A2(n15976), .A3(n15975), .ZN(n15980) );
  NAND2_X1 U19261 ( .A1(n15978), .A2(n19582), .ZN(n15979) );
  OAI211_X1 U19262 ( .C1(n16339), .C2(n15981), .A(n15980), .B(n15979), .ZN(
        P2_U2901) );
  INV_X1 U19263 ( .A(n15982), .ZN(n15991) );
  NAND2_X1 U19264 ( .A1(n15983), .A2(BUF1_REG_16__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U19265 ( .A1(n15984), .A2(BUF2_REG_16__SCAN_IN), .ZN(n15987) );
  AOI22_X1 U19266 ( .A1(n15985), .A2(n16525), .B1(n16010), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n15986) );
  NAND3_X1 U19267 ( .A1(n15988), .A2(n15987), .A3(n15986), .ZN(n15989) );
  AOI21_X1 U19268 ( .B1(n16347), .B2(n19578), .A(n15989), .ZN(n15990) );
  OAI21_X1 U19269 ( .B1(n16013), .B2(n15991), .A(n15990), .ZN(P2_U2903) );
  INV_X1 U19270 ( .A(n15992), .ZN(n15993) );
  NOR2_X1 U19271 ( .A1(n15994), .A2(n15993), .ZN(n16008) );
  XNOR2_X1 U19272 ( .A(n19692), .B(n20310), .ZN(n16009) );
  NOR2_X1 U19273 ( .A1(n16008), .A2(n16009), .ZN(n16007) );
  INV_X1 U19274 ( .A(n20310), .ZN(n16478) );
  NOR2_X1 U19275 ( .A1(n20309), .A2(n16478), .ZN(n15998) );
  NAND2_X1 U19276 ( .A1(n15739), .A2(n15995), .ZN(n15996) );
  NAND2_X1 U19277 ( .A1(n15997), .A2(n15996), .ZN(n19649) );
  OAI21_X1 U19278 ( .B1(n16007), .B2(n15998), .A(n19649), .ZN(n19581) );
  OR2_X1 U19279 ( .A1(n13845), .A2(n15999), .ZN(n16000) );
  NAND2_X1 U19280 ( .A1(n16001), .A2(n16000), .ZN(n19580) );
  INV_X1 U19281 ( .A(n19580), .ZN(n16002) );
  NAND3_X1 U19282 ( .A1(n19581), .A2(n19582), .A3(n16002), .ZN(n16004) );
  AOI22_X1 U19283 ( .A1(n19577), .A2(n16552), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n16010), .ZN(n16003) );
  OAI211_X1 U19284 ( .C1(n16006), .C2(n16005), .A(n16004), .B(n16003), .ZN(
        P2_U2914) );
  AOI21_X1 U19285 ( .B1(n16009), .B2(n16008), .A(n16007), .ZN(n16014) );
  AOI22_X1 U19286 ( .A1(n16478), .A2(n19578), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n16010), .ZN(n16012) );
  NAND2_X1 U19287 ( .A1(n19577), .A2(n16545), .ZN(n16011) );
  OAI211_X1 U19288 ( .C1(n16014), .C2(n16013), .A(n16012), .B(n16011), .ZN(
        P2_U2916) );
  XNOR2_X1 U19289 ( .A(n16015), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16281) );
  XNOR2_X1 U19290 ( .A(n16021), .B(n21443), .ZN(n16022) );
  NAND2_X1 U19291 ( .A1(n16277), .A2(n19642), .ZN(n16024) );
  INV_X1 U19292 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20277) );
  NOR2_X1 U19293 ( .A1(n16032), .A2(n20277), .ZN(n16269) );
  AOI21_X1 U19294 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16269), .ZN(n16023) );
  OAI211_X1 U19295 ( .C1(n16264), .C2(n16025), .A(n16024), .B(n16023), .ZN(
        n16026) );
  NAND2_X1 U19296 ( .A1(n16028), .A2(n16027), .ZN(n16029) );
  XNOR2_X1 U19297 ( .A(n16030), .B(n16029), .ZN(n16294) );
  AOI21_X1 U19298 ( .B1(n16286), .B2(n16044), .A(n16031), .ZN(n16292) );
  NAND2_X1 U19299 ( .A1(n16282), .A2(n19642), .ZN(n16034) );
  INV_X1 U19300 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20272) );
  NOR2_X1 U19301 ( .A1(n16032), .A2(n20272), .ZN(n16284) );
  AOI21_X1 U19302 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16284), .ZN(n16033) );
  OAI211_X1 U19303 ( .C1(n16264), .C2(n16035), .A(n16034), .B(n16033), .ZN(
        n16036) );
  AOI21_X1 U19304 ( .B1(n19636), .B2(n16292), .A(n16036), .ZN(n16037) );
  OAI21_X1 U19305 ( .B1(n19640), .B2(n16294), .A(n16037), .ZN(P2_U2989) );
  NAND2_X1 U19306 ( .A1(n16039), .A2(n16038), .ZN(n16041) );
  INV_X1 U19307 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20270) );
  NOR2_X1 U19308 ( .A1(n16032), .A2(n20270), .ZN(n16295) );
  AOI21_X1 U19309 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16295), .ZN(n16042) );
  OAI21_X1 U19310 ( .B1(n16043), .B2(n16264), .A(n16042), .ZN(n16045) );
  NOR2_X1 U19311 ( .A1(n16061), .A2(n16324), .ZN(n16060) );
  OAI21_X1 U19312 ( .B1(n16060), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9853), .ZN(n16318) );
  INV_X1 U19313 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20268) );
  NOR2_X1 U19314 ( .A1(n16032), .A2(n20268), .ZN(n16304) );
  AOI21_X1 U19315 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16304), .ZN(n16046) );
  OAI21_X1 U19316 ( .B1(n16047), .B2(n16264), .A(n16046), .ZN(n16048) );
  AOI21_X1 U19317 ( .B1(n16313), .B2(n19642), .A(n16048), .ZN(n16053) );
  AND2_X1 U19318 ( .A1(n16049), .A2(n16054), .ZN(n16051) );
  OR2_X1 U19319 ( .A1(n16051), .A2(n16050), .ZN(n16315) );
  NAND3_X1 U19320 ( .A1(n16315), .A2(n16314), .A3(n16263), .ZN(n16052) );
  OAI211_X1 U19321 ( .C1(n16318), .C2(n16253), .A(n16053), .B(n16052), .ZN(
        P2_U2991) );
  NAND2_X1 U19322 ( .A1(n16055), .A2(n16054), .ZN(n16059) );
  NAND2_X1 U19323 ( .A1(n16057), .A2(n16056), .ZN(n16058) );
  XOR2_X1 U19324 ( .A(n16059), .B(n16058), .Z(n16332) );
  AOI21_X1 U19325 ( .B1(n16061), .B2(n16324), .A(n16060), .ZN(n16319) );
  NAND2_X1 U19326 ( .A1(n16319), .A2(n19636), .ZN(n16067) );
  INV_X1 U19327 ( .A(n16062), .ZN(n16329) );
  NAND2_X1 U19328 ( .A1(n19553), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16321) );
  NAND2_X1 U19329 ( .A1(n19634), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16063) );
  OAI211_X1 U19330 ( .C1(n16064), .C2(n16264), .A(n16321), .B(n16063), .ZN(
        n16065) );
  AOI21_X1 U19331 ( .B1(n16329), .B2(n19642), .A(n16065), .ZN(n16066) );
  OAI211_X1 U19332 ( .C1(n16332), .C2(n19640), .A(n16067), .B(n16066), .ZN(
        P2_U2992) );
  OAI21_X1 U19333 ( .B1(n14260), .B2(n16081), .A(n16068), .ZN(n16069) );
  NAND2_X1 U19334 ( .A1(n9698), .A2(n16069), .ZN(n16344) );
  NAND2_X1 U19335 ( .A1(n16071), .A2(n16070), .ZN(n16072) );
  XNOR2_X1 U19336 ( .A(n16073), .B(n16072), .ZN(n16342) );
  NOR2_X1 U19337 ( .A1(n16032), .A2(n16074), .ZN(n16336) );
  NOR2_X1 U19338 ( .A1(n16237), .A2(n16075), .ZN(n16076) );
  AOI211_X1 U19339 ( .C1(n16077), .C2(n16234), .A(n16336), .B(n16076), .ZN(
        n16078) );
  OAI21_X1 U19340 ( .B1(n16333), .B2(n16222), .A(n16078), .ZN(n16079) );
  AOI21_X1 U19341 ( .B1(n16342), .B2(n16263), .A(n16079), .ZN(n16080) );
  OAI21_X1 U19342 ( .B1(n16344), .B2(n16253), .A(n16080), .ZN(P2_U2996) );
  XNOR2_X1 U19343 ( .A(n14260), .B(n16081), .ZN(n16088) );
  NAND2_X1 U19344 ( .A1(n19634), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16082) );
  OAI211_X1 U19345 ( .C1(n16084), .C2(n16264), .A(n16083), .B(n16082), .ZN(
        n16086) );
  XOR2_X1 U19346 ( .A(n16090), .B(n16089), .Z(n16353) );
  INV_X1 U19347 ( .A(n16353), .ZN(n16099) );
  INV_X1 U19348 ( .A(n16349), .ZN(n16095) );
  NOR2_X1 U19349 ( .A1(n16032), .A2(n16091), .ZN(n16346) );
  AOI21_X1 U19350 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16346), .ZN(n16092) );
  OAI21_X1 U19351 ( .B1(n16093), .B2(n16264), .A(n16092), .ZN(n16094) );
  AOI21_X1 U19352 ( .B1(n16095), .B2(n19642), .A(n16094), .ZN(n16098) );
  INV_X1 U19353 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16355) );
  OAI21_X1 U19354 ( .B1(n16114), .B2(n16364), .A(n16355), .ZN(n16096) );
  NAND3_X1 U19355 ( .A1(n16096), .A2(n19636), .A3(n14260), .ZN(n16097) );
  OAI211_X1 U19356 ( .C1(n16099), .C2(n19640), .A(n16098), .B(n16097), .ZN(
        P2_U2998) );
  XNOR2_X1 U19357 ( .A(n16114), .B(n16364), .ZN(n16369) );
  NAND3_X1 U19358 ( .A1(n16100), .A2(n16128), .A3(n16101), .ZN(n16127) );
  OAI21_X1 U19359 ( .B1(n16126), .B2(n16102), .A(n16116), .ZN(n16106) );
  NAND2_X1 U19360 ( .A1(n16104), .A2(n16103), .ZN(n16105) );
  XNOR2_X1 U19361 ( .A(n16106), .B(n16105), .ZN(n16366) );
  NAND2_X1 U19362 ( .A1(n19553), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16360) );
  OAI21_X1 U19363 ( .B1(n16237), .B2(n16107), .A(n16360), .ZN(n16108) );
  AOI21_X1 U19364 ( .B1(n16234), .B2(n16109), .A(n16108), .ZN(n16110) );
  OAI21_X1 U19365 ( .B1(n16357), .B2(n16222), .A(n16110), .ZN(n16111) );
  AOI21_X1 U19366 ( .B1(n16366), .B2(n16263), .A(n16111), .ZN(n16112) );
  OAI21_X1 U19367 ( .B1(n16369), .B2(n16253), .A(n16112), .ZN(P2_U2999) );
  INV_X1 U19368 ( .A(n16113), .ZN(n16397) );
  NAND2_X1 U19369 ( .A1(n16113), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16125) );
  INV_X1 U19370 ( .A(n16125), .ZN(n16115) );
  OAI21_X1 U19371 ( .B1(n16115), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16114), .ZN(n16382) );
  NAND2_X1 U19372 ( .A1(n16117), .A2(n16116), .ZN(n16118) );
  XOR2_X1 U19373 ( .A(n16118), .B(n16126), .Z(n16379) );
  NOR2_X1 U19374 ( .A1(n16032), .A2(n16119), .ZN(n16371) );
  NOR2_X1 U19375 ( .A1(n16264), .A2(n16120), .ZN(n16121) );
  AOI211_X1 U19376 ( .C1(n19634), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16371), .B(n16121), .ZN(n16122) );
  OAI21_X1 U19377 ( .B1(n16374), .B2(n16222), .A(n16122), .ZN(n16123) );
  AOI21_X1 U19378 ( .B1(n16379), .B2(n16263), .A(n16123), .ZN(n16124) );
  OAI21_X1 U19379 ( .B1(n16382), .B2(n16253), .A(n16124), .ZN(P2_U3000) );
  OAI21_X1 U19380 ( .B1(n16113), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16125), .ZN(n16395) );
  INV_X1 U19381 ( .A(n16126), .ZN(n16129) );
  AOI22_X1 U19382 ( .A1(n16129), .A2(n16128), .B1(n16100), .B2(n16127), .ZN(
        n16393) );
  NAND2_X1 U19383 ( .A1(n16130), .A2(n19642), .ZN(n16133) );
  NOR2_X1 U19384 ( .A1(n16032), .A2(n16131), .ZN(n16387) );
  AOI21_X1 U19385 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16387), .ZN(n16132) );
  OAI211_X1 U19386 ( .C1(n16264), .C2(n16134), .A(n16133), .B(n16132), .ZN(
        n16135) );
  AOI21_X1 U19387 ( .B1(n16393), .B2(n16263), .A(n16135), .ZN(n16136) );
  OAI21_X1 U19388 ( .B1(n16253), .B2(n16395), .A(n16136), .ZN(P2_U3001) );
  OAI21_X1 U19389 ( .B1(n16137), .B2(n16139), .A(n16138), .ZN(n16140) );
  INV_X1 U19390 ( .A(n16140), .ZN(n16406) );
  NAND2_X1 U19391 ( .A1(n16147), .A2(n16384), .ZN(n16396) );
  NAND3_X1 U19392 ( .A1(n16397), .A2(n19636), .A3(n16396), .ZN(n16146) );
  NAND2_X1 U19393 ( .A1(n19553), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n16399) );
  OAI21_X1 U19394 ( .B1(n16237), .B2(n16142), .A(n16399), .ZN(n16144) );
  NOR2_X1 U19395 ( .A1(n19521), .A2(n16222), .ZN(n16143) );
  AOI211_X1 U19396 ( .C1(n16234), .C2(n19518), .A(n16144), .B(n16143), .ZN(
        n16145) );
  OAI211_X1 U19397 ( .C1(n16406), .C2(n19640), .A(n16146), .B(n16145), .ZN(
        P2_U3002) );
  NOR2_X1 U19398 ( .A1(n16174), .A2(n16431), .ZN(n16168) );
  OAI21_X1 U19399 ( .B1(n16168), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16147), .ZN(n16423) );
  NAND2_X1 U19400 ( .A1(n16150), .A2(n16149), .ZN(n16151) );
  XNOR2_X1 U19401 ( .A(n16148), .B(n16151), .ZN(n16421) );
  NAND2_X1 U19402 ( .A1(n19553), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16413) );
  OAI21_X1 U19403 ( .B1(n16237), .B2(n16152), .A(n16413), .ZN(n16153) );
  AOI21_X1 U19404 ( .B1(n16234), .B2(n16154), .A(n16153), .ZN(n16155) );
  OAI21_X1 U19405 ( .B1(n16418), .B2(n16222), .A(n16155), .ZN(n16156) );
  AOI21_X1 U19406 ( .B1(n16421), .B2(n16263), .A(n16156), .ZN(n16157) );
  OAI21_X1 U19407 ( .B1(n16423), .B2(n16253), .A(n16157), .ZN(P2_U3003) );
  NAND2_X1 U19408 ( .A1(n16158), .A2(n16159), .ZN(n16204) );
  INV_X1 U19409 ( .A(n16202), .ZN(n16160) );
  INV_X1 U19410 ( .A(n16161), .ZN(n16162) );
  AOI21_X1 U19411 ( .B1(n16206), .B2(n16189), .A(n16162), .ZN(n16179) );
  AOI21_X1 U19412 ( .B1(n16179), .B2(n16176), .A(n16175), .ZN(n16167) );
  INV_X1 U19413 ( .A(n16163), .ZN(n16165) );
  NAND2_X1 U19414 ( .A1(n16165), .A2(n16164), .ZN(n16166) );
  XNOR2_X1 U19415 ( .A(n16167), .B(n16166), .ZN(n16437) );
  AOI21_X1 U19416 ( .B1(n16431), .B2(n16174), .A(n16168), .ZN(n16435) );
  NOR2_X1 U19417 ( .A1(n16032), .A2(n20247), .ZN(n16425) );
  NOR2_X1 U19418 ( .A1(n16264), .A2(n16169), .ZN(n16170) );
  AOI211_X1 U19419 ( .C1(n19634), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16425), .B(n16170), .ZN(n16171) );
  OAI21_X1 U19420 ( .B1(n16427), .B2(n16222), .A(n16171), .ZN(n16172) );
  AOI21_X1 U19421 ( .B1(n16435), .B2(n19636), .A(n16172), .ZN(n16173) );
  OAI21_X1 U19422 ( .B1(n16437), .B2(n19640), .A(n16173), .ZN(P2_U3004) );
  INV_X1 U19423 ( .A(n16175), .ZN(n16177) );
  NAND2_X1 U19424 ( .A1(n16177), .A2(n16176), .ZN(n16178) );
  XNOR2_X1 U19425 ( .A(n16179), .B(n16178), .ZN(n16447) );
  NAND2_X1 U19426 ( .A1(n16441), .A2(n19642), .ZN(n16181) );
  NOR2_X1 U19427 ( .A1(n16032), .A2(n20245), .ZN(n16439) );
  AOI21_X1 U19428 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16439), .ZN(n16180) );
  OAI211_X1 U19429 ( .C1(n16182), .C2(n16264), .A(n16181), .B(n16180), .ZN(
        n16183) );
  AOI21_X1 U19430 ( .B1(n16447), .B2(n16263), .A(n16183), .ZN(n16184) );
  OAI21_X1 U19431 ( .B1(n16253), .B2(n16449), .A(n16184), .ZN(P2_U3005) );
  XNOR2_X1 U19432 ( .A(n16185), .B(n16186), .ZN(n16462) );
  INV_X1 U19433 ( .A(n16205), .ZN(n16187) );
  NOR2_X1 U19434 ( .A1(n16206), .A2(n16187), .ZN(n16191) );
  NAND2_X1 U19435 ( .A1(n16189), .A2(n16188), .ZN(n16190) );
  XNOR2_X1 U19436 ( .A(n16191), .B(n16190), .ZN(n16460) );
  NAND2_X1 U19437 ( .A1(n16460), .A2(n16263), .ZN(n16196) );
  NAND2_X1 U19438 ( .A1(n19553), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16452) );
  NAND2_X1 U19439 ( .A1(n19634), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16192) );
  OAI211_X1 U19440 ( .C1(n16264), .C2(n16193), .A(n16452), .B(n16192), .ZN(
        n16194) );
  AOI21_X1 U19441 ( .B1(n16455), .B2(n19642), .A(n16194), .ZN(n16195) );
  OAI211_X1 U19442 ( .C1(n16462), .C2(n16253), .A(n16196), .B(n16195), .ZN(
        P2_U3006) );
  XNOR2_X1 U19443 ( .A(n16197), .B(n16451), .ZN(n16198) );
  NAND2_X1 U19444 ( .A1(n16234), .A2(n16199), .ZN(n16200) );
  NAND2_X1 U19445 ( .A1(n19553), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n17137) );
  OAI211_X1 U19446 ( .C1(n16237), .C2(n16201), .A(n16200), .B(n17137), .ZN(
        n16208) );
  NAND2_X1 U19447 ( .A1(n16205), .A2(n16202), .ZN(n16203) );
  AOI22_X1 U19448 ( .A1(n16206), .A2(n16205), .B1(n16204), .B2(n16203), .ZN(
        n17139) );
  NOR2_X1 U19449 ( .A1(n17139), .A2(n19640), .ZN(n16207) );
  AOI211_X1 U19450 ( .C1(n19642), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        n16210) );
  OAI21_X1 U19451 ( .B1(n16253), .B2(n17145), .A(n16210), .ZN(P2_U3007) );
  XNOR2_X1 U19452 ( .A(n16212), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16474) );
  XOR2_X1 U19453 ( .A(n16213), .B(n16214), .Z(n16472) );
  NOR2_X1 U19454 ( .A1(n16032), .A2(n20239), .ZN(n16466) );
  NOR2_X1 U19455 ( .A1(n16264), .A2(n19536), .ZN(n16215) );
  AOI211_X1 U19456 ( .C1(n19634), .C2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16466), .B(n16215), .ZN(n16216) );
  OAI21_X1 U19457 ( .B1(n19533), .B2(n16222), .A(n16216), .ZN(n16217) );
  AOI21_X1 U19458 ( .B1(n16472), .B2(n16263), .A(n16217), .ZN(n16218) );
  OAI21_X1 U19459 ( .B1(n16474), .B2(n16253), .A(n16218), .ZN(P2_U3008) );
  AOI22_X1 U19460 ( .A1(n19634), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19553), .ZN(n16221) );
  NAND2_X1 U19461 ( .A1(n16234), .A2(n16219), .ZN(n16220) );
  OAI211_X1 U19462 ( .C1(n16223), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        n16224) );
  AOI21_X1 U19463 ( .B1(n16225), .B2(n19636), .A(n16224), .ZN(n16226) );
  OAI21_X1 U19464 ( .B1(n16227), .B2(n19640), .A(n16226), .ZN(P2_U3009) );
  XNOR2_X1 U19465 ( .A(n16228), .B(n16229), .ZN(n19654) );
  NAND2_X1 U19466 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  AND2_X1 U19467 ( .A1(n16233), .A2(n16232), .ZN(n19651) );
  NAND2_X1 U19468 ( .A1(n16234), .A2(n19561), .ZN(n16235) );
  NAND2_X1 U19469 ( .A1(n19553), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n19647) );
  OAI211_X1 U19470 ( .C1(n16237), .C2(n16236), .A(n16235), .B(n19647), .ZN(
        n16238) );
  AOI21_X1 U19471 ( .B1(n19651), .B2(n19642), .A(n16238), .ZN(n16243) );
  XNOR2_X1 U19472 ( .A(n16239), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16240) );
  XNOR2_X1 U19473 ( .A(n16241), .B(n16240), .ZN(n19656) );
  NAND2_X1 U19474 ( .A1(n19656), .A2(n19636), .ZN(n16242) );
  OAI211_X1 U19475 ( .C1(n19654), .C2(n19640), .A(n16243), .B(n16242), .ZN(
        P2_U3010) );
  XNOR2_X1 U19476 ( .A(n16245), .B(n16476), .ZN(n16246) );
  XNOR2_X1 U19477 ( .A(n16244), .B(n16246), .ZN(n16485) );
  AOI22_X1 U19478 ( .A1(n19634), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19553), .ZN(n16247) );
  OAI21_X1 U19479 ( .B1(n16264), .B2(n16248), .A(n16247), .ZN(n16256) );
  CLKBUF_X1 U19480 ( .A(n16249), .Z(n16251) );
  NOR2_X1 U19481 ( .A1(n16251), .A2(n16250), .ZN(n16475) );
  INV_X1 U19482 ( .A(n16252), .ZN(n16254) );
  NOR3_X1 U19483 ( .A1(n16475), .A2(n16254), .A3(n16253), .ZN(n16255) );
  AOI211_X1 U19484 ( .C1(n19642), .C2(n16257), .A(n16256), .B(n16255), .ZN(
        n16258) );
  OAI21_X1 U19485 ( .B1(n19640), .B2(n16485), .A(n16258), .ZN(P2_U3011) );
  NAND2_X1 U19486 ( .A1(n16516), .A2(n19642), .ZN(n16268) );
  NOR2_X1 U19487 ( .A1(n16032), .A2(n20232), .ZN(n16488) );
  AOI21_X1 U19488 ( .B1(n19634), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16488), .ZN(n16267) );
  XNOR2_X1 U19489 ( .A(n16259), .B(n16514), .ZN(n16491) );
  XNOR2_X1 U19490 ( .A(n16260), .B(n16514), .ZN(n16261) );
  XNOR2_X1 U19491 ( .A(n16262), .B(n16261), .ZN(n16490) );
  AOI22_X1 U19492 ( .A1(n19636), .A2(n16491), .B1(n16263), .B2(n16490), .ZN(
        n16266) );
  OR2_X1 U19493 ( .A1(n16264), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16265) );
  NAND4_X1 U19494 ( .A1(n16268), .A2(n16267), .A3(n16266), .A4(n16265), .ZN(
        P2_U3013) );
  AOI21_X1 U19495 ( .B1(n16270), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16269), .ZN(n16274) );
  XNOR2_X1 U19496 ( .A(n21443), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16271) );
  NAND2_X1 U19497 ( .A1(n16272), .A2(n16271), .ZN(n16273) );
  OAI211_X1 U19498 ( .C1(n16275), .C2(n19648), .A(n16274), .B(n16273), .ZN(
        n16276) );
  AOI21_X1 U19499 ( .B1(n16277), .B2(n19669), .A(n16276), .ZN(n16280) );
  NAND2_X1 U19500 ( .A1(n16278), .A2(n19672), .ZN(n16279) );
  NAND2_X1 U19501 ( .A1(n16282), .A2(n19669), .ZN(n16289) );
  NOR2_X1 U19502 ( .A1(n16283), .A2(n16286), .ZN(n16285) );
  AOI211_X1 U19503 ( .C1(n16287), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        n16288) );
  OAI211_X1 U19504 ( .C1(n19648), .C2(n16290), .A(n16289), .B(n16288), .ZN(
        n16291) );
  AOI21_X1 U19505 ( .B1(n19657), .B2(n16292), .A(n16291), .ZN(n16293) );
  OAI21_X1 U19506 ( .B1(n19653), .B2(n16294), .A(n16293), .ZN(P2_U3021) );
  INV_X1 U19507 ( .A(n16295), .ZN(n16299) );
  OAI21_X1 U19508 ( .B1(n16297), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16296), .ZN(n16298) );
  OAI211_X1 U19509 ( .C1(n16300), .C2(n19648), .A(n16299), .B(n16298), .ZN(
        n16302) );
  AOI21_X1 U19510 ( .B1(n16320), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16304), .ZN(n16310) );
  NOR3_X1 U19511 ( .A1(n16307), .A2(n16306), .A3(n16305), .ZN(n16325) );
  OAI211_X1 U19512 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16325), .B(n16308), .ZN(
        n16309) );
  OAI211_X1 U19513 ( .C1(n16311), .C2(n19648), .A(n16310), .B(n16309), .ZN(
        n16312) );
  AOI21_X1 U19514 ( .B1(n16313), .B2(n19669), .A(n16312), .ZN(n16317) );
  NAND3_X1 U19515 ( .A1(n16315), .A2(n16314), .A3(n19672), .ZN(n16316) );
  OAI211_X1 U19516 ( .C1(n16318), .C2(n19668), .A(n16317), .B(n16316), .ZN(
        P2_U3023) );
  NAND2_X1 U19517 ( .A1(n16319), .A2(n19657), .ZN(n16331) );
  INV_X1 U19518 ( .A(n16320), .ZN(n16322) );
  OAI21_X1 U19519 ( .B1(n16322), .B2(n16324), .A(n16321), .ZN(n16323) );
  AOI21_X1 U19520 ( .B1(n16325), .B2(n16324), .A(n16323), .ZN(n16326) );
  OAI21_X1 U19521 ( .B1(n16327), .B2(n19648), .A(n16326), .ZN(n16328) );
  AOI21_X1 U19522 ( .B1(n16329), .B2(n19669), .A(n16328), .ZN(n16330) );
  OAI211_X1 U19523 ( .C1(n16332), .C2(n19653), .A(n16331), .B(n16330), .ZN(
        P2_U3024) );
  NOR2_X1 U19524 ( .A1(n16333), .A2(n17133), .ZN(n16341) );
  NOR3_X1 U19525 ( .A1(n16438), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16334), .ZN(n16335) );
  AOI211_X1 U19526 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16337), .A(
        n16336), .B(n16335), .ZN(n16338) );
  OAI21_X1 U19527 ( .B1(n19648), .B2(n16339), .A(n16338), .ZN(n16340) );
  OAI21_X1 U19528 ( .B1(n16344), .B2(n19668), .A(n16343), .ZN(P2_U3028) );
  INV_X1 U19529 ( .A(n16345), .ZN(n16356) );
  AOI21_X1 U19530 ( .B1(n16347), .B2(n19665), .A(n16346), .ZN(n16348) );
  OAI21_X1 U19531 ( .B1(n17133), .B2(n16349), .A(n16348), .ZN(n16352) );
  NOR3_X1 U19532 ( .A1(n16350), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16364), .ZN(n16351) );
  AOI211_X1 U19533 ( .C1(n19672), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        n16354) );
  OAI21_X1 U19534 ( .B1(n16356), .B2(n16355), .A(n16354), .ZN(P2_U3030) );
  NOR2_X1 U19535 ( .A1(n16357), .A2(n17133), .ZN(n16363) );
  NAND2_X1 U19536 ( .A1(n16358), .A2(n19665), .ZN(n16359) );
  OAI211_X1 U19537 ( .C1(n16361), .C2(n16364), .A(n16360), .B(n16359), .ZN(
        n16362) );
  AOI211_X1 U19538 ( .C1(n16365), .C2(n16364), .A(n16363), .B(n16362), .ZN(
        n16368) );
  NAND2_X1 U19539 ( .A1(n16366), .A2(n19672), .ZN(n16367) );
  OAI211_X1 U19540 ( .C1(n16369), .C2(n19668), .A(n16368), .B(n16367), .ZN(
        P2_U3031) );
  INV_X1 U19541 ( .A(n16403), .ZN(n16370) );
  OAI21_X1 U19542 ( .B1(n16400), .B2(n16375), .A(n16370), .ZN(n16386) );
  AOI21_X1 U19543 ( .B1(n16372), .B2(n19665), .A(n16371), .ZN(n16373) );
  OAI21_X1 U19544 ( .B1(n16374), .B2(n17133), .A(n16373), .ZN(n16378) );
  INV_X1 U19545 ( .A(n16375), .ZN(n16376) );
  NOR3_X1 U19546 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16376), .ZN(n16377) );
  AOI211_X1 U19547 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16386), .A(
        n16378), .B(n16377), .ZN(n16381) );
  NAND2_X1 U19548 ( .A1(n16379), .A2(n19672), .ZN(n16380) );
  OAI211_X1 U19549 ( .C1(n16382), .C2(n19668), .A(n16381), .B(n16380), .ZN(
        P2_U3032) );
  OAI21_X1 U19550 ( .B1(n16400), .B2(n16384), .A(n16383), .ZN(n16385) );
  NAND2_X1 U19551 ( .A1(n16386), .A2(n16385), .ZN(n16390) );
  AOI21_X1 U19552 ( .B1(n16388), .B2(n19665), .A(n16387), .ZN(n16389) );
  OAI211_X1 U19553 ( .C1(n16391), .C2(n17133), .A(n16390), .B(n16389), .ZN(
        n16392) );
  AOI21_X1 U19554 ( .B1(n16393), .B2(n19672), .A(n16392), .ZN(n16394) );
  OAI21_X1 U19555 ( .B1(n19668), .B2(n16395), .A(n16394), .ZN(P2_U3033) );
  NAND3_X1 U19556 ( .A1(n16397), .A2(n19657), .A3(n16396), .ZN(n16405) );
  NAND2_X1 U19557 ( .A1(n19520), .A2(n19665), .ZN(n16398) );
  OAI211_X1 U19558 ( .C1(n19521), .C2(n17133), .A(n16399), .B(n16398), .ZN(
        n16402) );
  NOR2_X1 U19559 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16401) );
  AOI211_X1 U19560 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16403), .A(
        n16402), .B(n16401), .ZN(n16404) );
  OAI211_X1 U19561 ( .C1(n16406), .C2(n19653), .A(n16405), .B(n16404), .ZN(
        P2_U3034) );
  NOR2_X1 U19562 ( .A1(n16444), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16407) );
  NAND2_X1 U19563 ( .A1(n16411), .A2(n16407), .ZN(n16424) );
  OR2_X1 U19564 ( .A1(n16408), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16409) );
  AND2_X1 U19565 ( .A1(n9631), .A2(n16409), .ZN(n16432) );
  AOI21_X1 U19566 ( .B1(n16424), .B2(n16432), .A(n16410), .ZN(n16420) );
  NAND4_X1 U19567 ( .A1(n16411), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A4(n16410), .ZN(n16417) );
  INV_X1 U19568 ( .A(n16412), .ZN(n16415) );
  INV_X1 U19569 ( .A(n16413), .ZN(n16414) );
  AOI21_X1 U19570 ( .B1(n16415), .B2(n19665), .A(n16414), .ZN(n16416) );
  OAI211_X1 U19571 ( .C1(n16418), .C2(n17133), .A(n16417), .B(n16416), .ZN(
        n16419) );
  AOI211_X1 U19572 ( .C1(n16421), .C2(n19672), .A(n16420), .B(n16419), .ZN(
        n16422) );
  OAI21_X1 U19573 ( .B1(n16423), .B2(n19668), .A(n16422), .ZN(P2_U3035) );
  INV_X1 U19574 ( .A(n16424), .ZN(n16434) );
  AOI21_X1 U19575 ( .B1(n16426), .B2(n19665), .A(n16425), .ZN(n16430) );
  INV_X1 U19576 ( .A(n16427), .ZN(n16428) );
  NAND2_X1 U19577 ( .A1(n16428), .A2(n19669), .ZN(n16429) );
  OAI211_X1 U19578 ( .C1(n16432), .C2(n16431), .A(n16430), .B(n16429), .ZN(
        n16433) );
  AOI211_X1 U19579 ( .C1(n16435), .C2(n19657), .A(n16434), .B(n16433), .ZN(
        n16436) );
  NOR2_X1 U19580 ( .A1(n16438), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16446) );
  AOI21_X1 U19581 ( .B1(n16440), .B2(n19665), .A(n16439), .ZN(n16443) );
  NAND2_X1 U19582 ( .A1(n16441), .A2(n19669), .ZN(n16442) );
  OAI211_X1 U19583 ( .C1(n9631), .C2(n16444), .A(n16443), .B(n16442), .ZN(
        n16445) );
  AOI211_X1 U19584 ( .C1(n16447), .C2(n19672), .A(n16446), .B(n16445), .ZN(
        n16448) );
  OAI21_X1 U19585 ( .B1(n19668), .B2(n16449), .A(n16448), .ZN(P2_U3037) );
  AOI211_X1 U19586 ( .C1(n16451), .C2(n16457), .A(n16450), .B(n17135), .ZN(
        n16459) );
  OAI21_X1 U19587 ( .B1(n16453), .B2(n19648), .A(n16452), .ZN(n16454) );
  AOI21_X1 U19588 ( .B1(n16455), .B2(n19669), .A(n16454), .ZN(n16456) );
  OAI21_X1 U19589 ( .B1(n10023), .B2(n16457), .A(n16456), .ZN(n16458) );
  AOI211_X1 U19590 ( .C1(n16460), .C2(n19672), .A(n16459), .B(n16458), .ZN(
        n16461) );
  OAI21_X1 U19591 ( .B1(n16462), .B2(n19668), .A(n16461), .ZN(P2_U3038) );
  INV_X1 U19592 ( .A(n16463), .ZN(n16470) );
  NAND2_X1 U19593 ( .A1(n16464), .A2(n16469), .ZN(n16468) );
  NOR2_X1 U19594 ( .A1(n19533), .A2(n17133), .ZN(n16465) );
  AOI211_X1 U19595 ( .C1(n19665), .C2(n19543), .A(n16466), .B(n16465), .ZN(
        n16467) );
  OAI211_X1 U19596 ( .C1(n16470), .C2(n16469), .A(n16468), .B(n16467), .ZN(
        n16471) );
  AOI21_X1 U19597 ( .B1(n16472), .B2(n19672), .A(n16471), .ZN(n16473) );
  OAI21_X1 U19598 ( .B1(n16474), .B2(n19668), .A(n16473), .ZN(P2_U3040) );
  NOR2_X1 U19599 ( .A1(n16475), .A2(n19668), .ZN(n16483) );
  AOI22_X1 U19600 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16477), .B1(
        n9687), .B2(n16476), .ZN(n16480) );
  AOI22_X1 U19601 ( .A1(n19665), .A2(n16478), .B1(n19553), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n16479) );
  OAI211_X1 U19602 ( .C1(n16481), .C2(n17133), .A(n16480), .B(n16479), .ZN(
        n16482) );
  AOI21_X1 U19603 ( .B1(n16483), .B2(n16252), .A(n16482), .ZN(n16484) );
  OAI21_X1 U19604 ( .B1(n19653), .B2(n16485), .A(n16484), .ZN(P2_U3043) );
  OAI22_X1 U19605 ( .A1(n17133), .A2(n16486), .B1(n16498), .B2(n19648), .ZN(
        n16487) );
  AOI211_X1 U19606 ( .C1(n16489), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n16488), .B(n16487), .ZN(n16494) );
  AOI22_X1 U19607 ( .A1(n19657), .A2(n16491), .B1(n19672), .B2(n16490), .ZN(
        n16493) );
  OAI211_X1 U19608 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n9986), .B(n19675), .ZN(n16492)
         );
  NAND3_X1 U19609 ( .A1(n16494), .A2(n16493), .A3(n16492), .ZN(P2_U3045) );
  OAI21_X1 U19610 ( .B1(n16495), .B2(n16621), .A(n20306), .ZN(n16496) );
  MUX2_X1 U19611 ( .A(n20303), .B(n16496), .S(n20308), .Z(n16497) );
  OAI21_X1 U19612 ( .B1(n16498), .B2(n20318), .A(n16497), .ZN(n16503) );
  NAND2_X1 U19613 ( .A1(n17156), .A2(n20327), .ZN(n16499) );
  NAND2_X1 U19614 ( .A1(n20338), .A2(n16600), .ZN(n16501) );
  NAND2_X1 U19615 ( .A1(n16501), .A2(n17151), .ZN(n16502) );
  NAND2_X1 U19616 ( .A1(n20101), .A2(n16502), .ZN(n20334) );
  INV_X1 U19617 ( .A(n20334), .ZN(n20333) );
  MUX2_X1 U19618 ( .A(n16503), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n20333), .Z(P2_U3604) );
  MUX2_X1 U19619 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16504), .S(
        n19559), .Z(n16505) );
  NAND2_X1 U19620 ( .A1(n16505), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20296) );
  NAND2_X1 U19621 ( .A1(n16507), .A2(n16506), .ZN(n16520) );
  MUX2_X1 U19622 ( .A(n16520), .B(n12038), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n16508) );
  AOI21_X1 U19623 ( .B1(n19643), .B2(n16515), .A(n16508), .ZN(n16606) );
  OAI21_X1 U19624 ( .B1(n16606), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16621), 
        .ZN(n16510) );
  AOI22_X1 U19625 ( .A1(n20296), .A2(n16510), .B1(n16509), .B2(n17152), .ZN(
        n16512) );
  NAND2_X1 U19626 ( .A1(n20301), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16511) );
  OAI21_X1 U19627 ( .B1(n16512), .B2(n20301), .A(n16511), .ZN(P2_U3601) );
  OAI21_X1 U19628 ( .B1(n19559), .B2(n16514), .A(n16513), .ZN(n20294) );
  NAND2_X1 U19629 ( .A1(n16516), .A2(n16515), .ZN(n16607) );
  NOR2_X1 U19630 ( .A1(n16517), .A2(n16518), .ZN(n16521) );
  AOI22_X1 U19631 ( .A1(n16521), .A2(n16520), .B1(n12038), .B2(n16519), .ZN(
        n16608) );
  AOI21_X1 U19632 ( .B1(n16607), .B2(n16608), .A(n20297), .ZN(n16522) );
  AOI21_X1 U19633 ( .B1(n20308), .B2(n17152), .A(n16522), .ZN(n16523) );
  OAI21_X1 U19634 ( .B1(n20296), .B2(n20294), .A(n16523), .ZN(n16524) );
  MUX2_X1 U19635 ( .A(n16524), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20301), .Z(P2_U3600) );
  INV_X1 U19636 ( .A(n20150), .ZN(n19945) );
  OR2_X1 U19637 ( .A1(n20313), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20095) );
  INV_X1 U19638 ( .A(n16527), .ZN(n16528) );
  NAND2_X1 U19639 ( .A1(n16528), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20144) );
  NOR2_X1 U19640 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19745) );
  INV_X1 U19641 ( .A(n19745), .ZN(n19746) );
  NOR2_X1 U19642 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19746), .ZN(
        n19687) );
  AND2_X1 U19643 ( .A1(n19687), .A2(n20335), .ZN(n16567) );
  OAI21_X1 U19644 ( .B1(n16529), .B2(n20145), .A(n20318), .ZN(n16530) );
  AOI21_X1 U19645 ( .B1(n16531), .B2(n20144), .A(n16530), .ZN(n16532) );
  INV_X1 U19646 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U19647 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16562), .B1(
        n20204), .B2(n20102), .ZN(n16537) );
  INV_X1 U19648 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18870) );
  OAI22_X2 U19649 ( .A1(n20593), .A2(n16564), .B1(n18870), .B2(n16563), .ZN(
        n20159) );
  NOR2_X2 U19650 ( .A1(n16535), .A2(n16553), .ZN(n20149) );
  AOI22_X1 U19651 ( .A1(n20159), .A2(n19711), .B1(n16567), .B2(n20149), .ZN(
        n16536) );
  OAI211_X1 U19652 ( .C1(n19945), .C2(n16570), .A(n16537), .B(n16536), .ZN(
        P2_U3048) );
  NAND2_X1 U19653 ( .A1(n16538), .A2(n20152), .ZN(n19948) );
  INV_X1 U19654 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20601) );
  INV_X1 U19655 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18877) );
  OAI22_X2 U19656 ( .A1(n20601), .A2(n16564), .B1(n18877), .B2(n16563), .ZN(
        n20165) );
  AOI22_X1 U19657 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16562), .B1(
        n19711), .B2(n20165), .ZN(n16540) );
  INV_X1 U19658 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18876) );
  INV_X1 U19659 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20598) );
  OAI22_X1 U19660 ( .A1(n18876), .A2(n16563), .B1(n20598), .B2(n16564), .ZN(
        n20111) );
  AOI22_X1 U19661 ( .A1(n20111), .A2(n20204), .B1(n16567), .B2(n20163), .ZN(
        n16539) );
  OAI211_X1 U19662 ( .C1(n19948), .C2(n16570), .A(n16540), .B(n16539), .ZN(
        P2_U3049) );
  INV_X1 U19663 ( .A(n20170), .ZN(n19951) );
  INV_X1 U19664 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18015) );
  OAI22_X1 U19665 ( .A1(n18015), .A2(n16563), .B1(n21377), .B2(n16564), .ZN(
        n20115) );
  AOI22_X1 U19666 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n16562), .B1(
        n20204), .B2(n20115), .ZN(n16544) );
  INV_X1 U19667 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18882) );
  OAI22_X2 U19668 ( .A1(n17178), .A2(n16564), .B1(n18882), .B2(n16563), .ZN(
        n20171) );
  NOR2_X2 U19669 ( .A1(n16542), .A2(n16553), .ZN(n20169) );
  AOI22_X1 U19670 ( .A1(n20171), .A2(n19711), .B1(n16567), .B2(n20169), .ZN(
        n16543) );
  OAI211_X1 U19671 ( .C1(n16570), .C2(n19951), .A(n16544), .B(n16543), .ZN(
        P2_U3050) );
  NAND2_X1 U19672 ( .A1(n16545), .A2(n20152), .ZN(n19954) );
  INV_X1 U19673 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21324) );
  INV_X1 U19674 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20610) );
  OAI22_X1 U19675 ( .A1(n21324), .A2(n16563), .B1(n20610), .B2(n16564), .ZN(
        n20119) );
  AOI22_X1 U19676 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n16562), .B1(
        n20204), .B2(n20119), .ZN(n16548) );
  INV_X1 U19677 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20608) );
  INV_X1 U19678 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18886) );
  OAI22_X2 U19679 ( .A1(n20608), .A2(n16564), .B1(n18886), .B2(n16563), .ZN(
        n20177) );
  AOI22_X1 U19680 ( .A1(n20177), .A2(n19711), .B1(n16567), .B2(n20175), .ZN(
        n16547) );
  OAI211_X1 U19681 ( .C1(n19954), .C2(n16570), .A(n16548), .B(n16547), .ZN(
        P2_U3051) );
  INV_X1 U19682 ( .A(n20182), .ZN(n19957) );
  INV_X1 U19683 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20620) );
  INV_X1 U19684 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18890) );
  AOI22_X1 U19685 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n16562), .B1(
        n20204), .B2(n20123), .ZN(n16551) );
  INV_X1 U19686 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20618) );
  INV_X1 U19687 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18892) );
  OAI22_X2 U19688 ( .A1(n20618), .A2(n16564), .B1(n18892), .B2(n16563), .ZN(
        n20183) );
  NOR2_X2 U19689 ( .A1(n16549), .A2(n16553), .ZN(n20181) );
  AOI22_X1 U19690 ( .A1(n20183), .A2(n19711), .B1(n16567), .B2(n20181), .ZN(
        n16550) );
  OAI211_X1 U19691 ( .C1(n16570), .C2(n19957), .A(n16551), .B(n16550), .ZN(
        P2_U3052) );
  NAND2_X1 U19692 ( .A1(n16552), .A2(n20152), .ZN(n19960) );
  INV_X1 U19693 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20625) );
  INV_X1 U19694 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18895) );
  OAI22_X2 U19695 ( .A1(n20625), .A2(n16564), .B1(n18895), .B2(n16563), .ZN(
        n20189) );
  AOI22_X1 U19696 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n16562), .B1(
        n19711), .B2(n20189), .ZN(n16556) );
  INV_X1 U19697 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17237) );
  NOR2_X2 U19698 ( .A1(n16554), .A2(n16553), .ZN(n20187) );
  AOI22_X1 U19699 ( .A1(n20127), .A2(n20204), .B1(n16567), .B2(n20187), .ZN(
        n16555) );
  OAI211_X1 U19700 ( .C1(n19960), .C2(n16570), .A(n16556), .B(n16555), .ZN(
        P2_U3053) );
  INV_X1 U19701 ( .A(n20194), .ZN(n19963) );
  INV_X1 U19702 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18903) );
  OAI22_X2 U19703 ( .A1(n20635), .A2(n16564), .B1(n18903), .B2(n16563), .ZN(
        n20195) );
  AOI22_X1 U19704 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16562), .B1(
        n19711), .B2(n20195), .ZN(n16560) );
  INV_X1 U19705 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20637) );
  INV_X1 U19706 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18901) );
  OAI22_X1 U19707 ( .A1(n20637), .A2(n16564), .B1(n18901), .B2(n16563), .ZN(
        n20131) );
  AND2_X1 U19708 ( .A1(n16558), .A2(n16565), .ZN(n20193) );
  AOI22_X1 U19709 ( .A1(n20131), .A2(n20204), .B1(n16567), .B2(n20193), .ZN(
        n16559) );
  OAI211_X1 U19710 ( .C1(n16570), .C2(n19963), .A(n16560), .B(n16559), .ZN(
        P2_U3054) );
  INV_X1 U19711 ( .A(n20201), .ZN(n19969) );
  INV_X1 U19712 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U19713 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n16562), .B1(
        n20204), .B2(n20136), .ZN(n16569) );
  INV_X1 U19714 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20642) );
  INV_X1 U19715 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18907) );
  OAI22_X2 U19716 ( .A1(n20642), .A2(n16564), .B1(n18907), .B2(n16563), .ZN(
        n20203) );
  AOI22_X1 U19717 ( .A1(n20203), .A2(n19711), .B1(n16567), .B2(n20199), .ZN(
        n16568) );
  OAI211_X1 U19718 ( .C1(n16570), .C2(n19969), .A(n16569), .B(n16568), .ZN(
        P2_U3055) );
  OR2_X1 U19719 ( .A1(n16572), .A2(n16571), .ZN(n16584) );
  NAND2_X1 U19720 ( .A1(n9609), .A2(n16573), .ZN(n16575) );
  INV_X1 U19721 ( .A(n16575), .ZN(n16581) );
  NAND2_X1 U19722 ( .A1(n16576), .A2(n16575), .ZN(n16577) );
  OAI21_X1 U19723 ( .B1(n16579), .B2(n16578), .A(n16577), .ZN(n16580) );
  AOI21_X1 U19724 ( .B1(n16582), .B2(n16581), .A(n16580), .ZN(n16583) );
  AND2_X1 U19725 ( .A1(n16584), .A2(n16583), .ZN(n20298) );
  NOR2_X1 U19726 ( .A1(n16610), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16585) );
  AOI21_X1 U19727 ( .B1(n20298), .B2(n16610), .A(n16585), .ZN(n16620) );
  NAND2_X1 U19728 ( .A1(n16586), .A2(n16610), .ZN(n16590) );
  NAND2_X1 U19729 ( .A1(n16610), .A2(n16587), .ZN(n16588) );
  NAND2_X1 U19730 ( .A1(n16588), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16589) );
  NAND2_X1 U19731 ( .A1(n16590), .A2(n16589), .ZN(n16619) );
  INV_X1 U19732 ( .A(n16591), .ZN(n16596) );
  MUX2_X1 U19733 ( .A(n16594), .B(n16593), .S(n16592), .Z(n16595) );
  AOI21_X1 U19734 ( .B1(n16597), .B2(n16596), .A(n16595), .ZN(n20344) );
  INV_X1 U19735 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n16599) );
  AOI21_X1 U19736 ( .B1(n16600), .B2(n16599), .A(n16598), .ZN(n16601) );
  AOI211_X1 U19737 ( .C1(n16603), .C2(n11752), .A(n16602), .B(n16601), .ZN(
        n16604) );
  OAI211_X1 U19738 ( .C1(n16605), .C2(n16610), .A(n20344), .B(n16604), .ZN(
        n16618) );
  AOI22_X1 U19739 ( .A1(n16619), .A2(n20317), .B1(n16620), .B2(n19745), .ZN(
        n16616) );
  INV_X1 U19740 ( .A(n16606), .ZN(n16612) );
  OAI21_X1 U19741 ( .B1(n16612), .B2(n20335), .A(n20034), .ZN(n16609) );
  NAND3_X1 U19742 ( .A1(n16609), .A2(n16608), .A3(n16607), .ZN(n16611) );
  OAI211_X1 U19743 ( .C1(n19747), .C2(n16612), .A(n16611), .B(n16610), .ZN(
        n16613) );
  AOI21_X1 U19744 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20298), .A(
        n16613), .ZN(n16614) );
  OAI21_X1 U19745 ( .B1(n16619), .B2(n20317), .A(n16614), .ZN(n16615) );
  AOI21_X1 U19746 ( .B1(n16616), .B2(n16615), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16617) );
  AOI211_X1 U19747 ( .C1(n16620), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        n17161) );
  AOI21_X1 U19748 ( .B1(n17161), .B2(n16621), .A(n17153), .ZN(n16625) );
  NOR3_X1 U19749 ( .A1(n16622), .A2(n12831), .A3(n15806), .ZN(n16624) );
  NOR3_X1 U19750 ( .A1(n20224), .A2(n17153), .A3(n20297), .ZN(n16627) );
  NOR2_X1 U19751 ( .A1(n16627), .A2(n16626), .ZN(n16630) );
  INV_X1 U19752 ( .A(n17146), .ZN(n16628) );
  OAI211_X1 U19753 ( .C1(n17154), .C2(n16628), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20224), .ZN(n16629) );
  OAI211_X1 U19754 ( .C1(n17154), .C2(n16630), .A(n16629), .B(n19537), .ZN(
        P2_U3177) );
  OAI21_X1 U19755 ( .B1(n17154), .B2(n17153), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n16632) );
  INV_X1 U19756 ( .A(n17151), .ZN(n16631) );
  NAND2_X1 U19757 ( .A1(n16632), .A2(n16631), .ZN(P2_U3593) );
  NOR3_X1 U19758 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17599), .A3(n16639), .ZN(
        n16644) );
  AOI211_X1 U19759 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16656), .A(n17562), .B(
        n17605), .ZN(n16643) );
  AOI22_X1 U19760 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17525), .B1(
        n17518), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16633) );
  INV_X1 U19761 ( .A(n16633), .ZN(n16642) );
  INV_X1 U19762 ( .A(n16634), .ZN(n16635) );
  NOR2_X1 U19763 ( .A1(n16635), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18512) );
  NOR2_X1 U19764 ( .A1(n18561), .A2(n16636), .ZN(n16637) );
  INV_X1 U19765 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17597) );
  AOI21_X1 U19766 ( .B1(n16637), .B2(n17597), .A(n17519), .ZN(n17560) );
  NAND2_X1 U19767 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16634), .ZN(
        n16649) );
  INV_X1 U19768 ( .A(n16649), .ZN(n16638) );
  INV_X1 U19769 ( .A(n16637), .ZN(n17557) );
  OAI21_X1 U19770 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16638), .A(
        n17557), .ZN(n18522) );
  AOI22_X1 U19771 ( .A1(n17579), .A2(n18512), .B1(n17560), .B2(n18522), .ZN(
        n16640) );
  AOI21_X1 U19772 ( .B1(n17581), .B2(n16639), .A(n17593), .ZN(n16651) );
  OAI22_X1 U19773 ( .A1(n16640), .A2(n19355), .B1(n19382), .B2(n16651), .ZN(
        n16641) );
  NOR4_X1 U19774 ( .A1(n16644), .A2(n16643), .A3(n16642), .A4(n16641), .ZN(
        n16647) );
  OAI21_X1 U19775 ( .B1(n17858), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19489), .ZN(n16646) );
  NAND2_X1 U19776 ( .A1(n17558), .A2(n17519), .ZN(n17572) );
  OR2_X1 U19777 ( .A1(n18522), .A2(n17572), .ZN(n16645) );
  NAND4_X1 U19778 ( .A1(n16647), .A2(n18748), .A3(n16646), .A4(n16645), .ZN(
        P3_U2667) );
  INV_X1 U19779 ( .A(n16930), .ZN(n16648) );
  AOI21_X1 U19780 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16648), .A(
        n17872), .ZN(n16661) );
  NAND2_X1 U19781 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17571) );
  INV_X1 U19782 ( .A(n17571), .ZN(n17577) );
  AOI21_X1 U19783 ( .B1(n17577), .B2(n17597), .A(n17519), .ZN(n16650) );
  OAI21_X1 U19784 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17577), .A(
        n16649), .ZN(n18535) );
  XNOR2_X1 U19785 ( .A(n16650), .B(n18535), .ZN(n16655) );
  INV_X1 U19786 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19380) );
  NAND2_X1 U19787 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17580) );
  AOI221_X1 U19788 ( .B1(n17599), .B2(n19380), .C1(n17580), .C2(n19380), .A(
        n16651), .ZN(n16654) );
  OAI22_X1 U19789 ( .A1(n16652), .A2(n17595), .B1(n17598), .B2(n16657), .ZN(
        n16653) );
  AOI211_X1 U19790 ( .C1(n16655), .C2(n17558), .A(n16654), .B(n16653), .ZN(
        n16659) );
  OAI211_X1 U19791 ( .C1(n17582), .C2(n16657), .A(n17584), .B(n16656), .ZN(
        n16658) );
  OAI211_X1 U19792 ( .C1(n16661), .C2(n16660), .A(n16659), .B(n16658), .ZN(
        P3_U2668) );
  AOI21_X1 U19793 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n16662), .A(
        P3_EAX_REG_2__SCAN_IN), .ZN(n16665) );
  NAND3_X1 U19794 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n18125) );
  AOI21_X1 U19795 ( .B1(n18910), .B2(n18125), .A(n13921), .ZN(n18130) );
  AOI22_X1 U19796 ( .A1(n18128), .A2(BUF2_REG_2__SCAN_IN), .B1(n18127), .B2(
        n16663), .ZN(n16664) );
  OAI21_X1 U19797 ( .B1(n16665), .B2(n18130), .A(n16664), .ZN(P3_U2733) );
  INV_X1 U19798 ( .A(n13921), .ZN(n16666) );
  NAND2_X1 U19799 ( .A1(n18910), .A2(n16666), .ZN(n18124) );
  NAND2_X1 U19800 ( .A1(n18128), .A2(BUF2_REG_0__SCAN_IN), .ZN(n16669) );
  AOI22_X1 U19801 ( .A1(n13921), .A2(P3_EAX_REG_0__SCAN_IN), .B1(n18127), .B2(
        n16667), .ZN(n16668) );
  OAI211_X1 U19802 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(n18124), .A(n16669), .B(
        n16668), .ZN(P3_U2735) );
  NAND2_X1 U19803 ( .A1(n18369), .A2(n16808), .ZN(n16670) );
  INV_X1 U19804 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U19805 ( .A1(n16694), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16693) );
  XNOR2_X1 U19806 ( .A(n18369), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16674) );
  NAND2_X1 U19807 ( .A1(n16671), .A2(n18369), .ZN(n16672) );
  NAND3_X1 U19808 ( .A1(n16693), .A2(n16674), .A3(n16672), .ZN(n16678) );
  INV_X1 U19809 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16895) );
  NAND2_X1 U19810 ( .A1(n16895), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16780) );
  NAND3_X1 U19811 ( .A1(n16673), .A2(n16672), .A3(n16780), .ZN(n16676) );
  INV_X1 U19812 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16799) );
  NAND2_X1 U19813 ( .A1(n16799), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16778) );
  INV_X1 U19814 ( .A(n16674), .ZN(n16675) );
  NAND3_X1 U19815 ( .A1(n16676), .A2(n16778), .A3(n16675), .ZN(n16677) );
  NAND2_X1 U19816 ( .A1(n16678), .A2(n16677), .ZN(n16792) );
  AND2_X1 U19817 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16814) );
  NAND2_X1 U19818 ( .A1(n16814), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16783) );
  NOR2_X1 U19819 ( .A1(n16679), .A2(n16783), .ZN(n16695) );
  NAND2_X1 U19820 ( .A1(n16695), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16680) );
  XNOR2_X1 U19821 ( .A(n16680), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16790) );
  XOR2_X1 U19822 ( .A(n10147), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16690) );
  NAND2_X1 U19823 ( .A1(n18398), .A2(n16681), .ZN(n16702) );
  INV_X1 U19824 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19433) );
  NOR2_X1 U19825 ( .A1(n18748), .A2(n19433), .ZN(n16785) );
  NOR2_X1 U19826 ( .A1(n18277), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16714) );
  INV_X1 U19827 ( .A(n16682), .ZN(n16684) );
  OR2_X1 U19828 ( .A1(n18906), .A2(n16681), .ZN(n16710) );
  INV_X1 U19829 ( .A(n16710), .ZN(n16683) );
  AOI21_X1 U19830 ( .B1(n18396), .B2(n16684), .A(n16683), .ZN(n16685) );
  NAND2_X1 U19831 ( .A1(n18547), .A2(n16685), .ZN(n16712) );
  NOR2_X1 U19832 ( .A1(n16714), .A2(n16712), .ZN(n16697) );
  NOR2_X1 U19833 ( .A1(n16697), .A2(n10147), .ZN(n16686) );
  AOI211_X1 U19834 ( .C1(n18417), .C2(n17508), .A(n16785), .B(n16686), .ZN(
        n16689) );
  INV_X1 U19835 ( .A(n16796), .ZN(n16845) );
  INV_X1 U19836 ( .A(n16783), .ZN(n16775) );
  NAND2_X1 U19837 ( .A1(n16845), .A2(n16775), .ZN(n16797) );
  NAND2_X1 U19838 ( .A1(n16797), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16687) );
  OAI211_X1 U19839 ( .C1(n16797), .C2(n16780), .A(n16778), .B(n16687), .ZN(
        n16777) );
  NAND2_X1 U19840 ( .A1(n16777), .A2(n18557), .ZN(n16688) );
  OAI211_X1 U19841 ( .C1(n16690), .C2(n16702), .A(n16689), .B(n16688), .ZN(
        n16691) );
  AOI21_X1 U19842 ( .B1(n16790), .B2(n18426), .A(n16691), .ZN(n16692) );
  OAI21_X1 U19843 ( .B1(n16792), .B2(n18464), .A(n16692), .ZN(P3_U2799) );
  OAI21_X1 U19844 ( .B1(n16694), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16693), .ZN(n16805) );
  INV_X1 U19845 ( .A(n16695), .ZN(n16798) );
  NAND2_X1 U19846 ( .A1(n16798), .A2(n18426), .ZN(n16719) );
  NAND2_X1 U19847 ( .A1(n16797), .A2(n18557), .ZN(n16717) );
  AOI21_X1 U19848 ( .B1(n16719), .B2(n16717), .A(n16799), .ZN(n16704) );
  NOR2_X1 U19849 ( .A1(n18748), .A2(n19436), .ZN(n16802) );
  NOR2_X1 U19850 ( .A1(n16697), .A2(n16696), .ZN(n16698) );
  AOI211_X1 U19851 ( .C1(n18417), .C2(n12923), .A(n16802), .B(n16698), .ZN(
        n16701) );
  NOR2_X1 U19852 ( .A1(n16783), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16803) );
  INV_X1 U19853 ( .A(n16853), .ZN(n16699) );
  NAND3_X1 U19854 ( .A1(n18268), .A2(n16803), .A3(n16699), .ZN(n16700) );
  OAI211_X1 U19855 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n16702), .A(
        n16701), .B(n16700), .ZN(n16703) );
  NOR2_X1 U19856 ( .A1(n16704), .A2(n16703), .ZN(n16705) );
  OAI21_X1 U19857 ( .B1(n18464), .B2(n16805), .A(n16705), .ZN(P3_U2800) );
  NOR2_X1 U19858 ( .A1(n16707), .A2(n16706), .ZN(n16708) );
  XNOR2_X1 U19859 ( .A(n16708), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16812) );
  INV_X1 U19860 ( .A(n16814), .ZN(n16709) );
  NOR2_X1 U19861 ( .A1(n16796), .A2(n16709), .ZN(n16822) );
  NOR2_X1 U19862 ( .A1(n16822), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16718) );
  NAND2_X1 U19863 ( .A1(n18846), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16817) );
  OAI21_X1 U19864 ( .B1(n12899), .B2(n16710), .A(n16817), .ZN(n16711) );
  AOI21_X1 U19865 ( .B1(n16712), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16711), .ZN(n16716) );
  INV_X1 U19866 ( .A(n17290), .ZN(n16713) );
  OAI21_X1 U19867 ( .B1(n16714), .B2(n18417), .A(n16713), .ZN(n16715) );
  OAI211_X1 U19868 ( .C1(n16718), .C2(n16717), .A(n16716), .B(n16715), .ZN(
        n16721) );
  NAND2_X1 U19869 ( .A1(n16846), .A2(n16814), .ZN(n16824) );
  AOI21_X1 U19870 ( .B1(n16813), .B2(n16824), .A(n16719), .ZN(n16720) );
  AOI211_X1 U19871 ( .C1(n18436), .C2(n16812), .A(n16721), .B(n16720), .ZN(
        n16722) );
  INV_X1 U19872 ( .A(n16722), .ZN(P3_U2801) );
  NOR2_X1 U19873 ( .A1(n16724), .A2(n16723), .ZN(n16725) );
  XNOR2_X1 U19874 ( .A(n16725), .B(n18369), .ZN(n16860) );
  OAI21_X1 U19875 ( .B1(n16758), .B2(n16853), .A(n16854), .ZN(n16731) );
  NAND2_X1 U19876 ( .A1(n16726), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16728) );
  INV_X1 U19877 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19427) );
  NOR2_X1 U19878 ( .A1(n18748), .A2(n19427), .ZN(n16856) );
  INV_X1 U19879 ( .A(n16856), .ZN(n16727) );
  OAI211_X1 U19880 ( .C1(n18402), .C2(n17312), .A(n16728), .B(n16727), .ZN(
        n16729) );
  AOI211_X1 U19881 ( .C1(n16732), .C2(n16731), .A(n16730), .B(n16729), .ZN(
        n16733) );
  OAI21_X1 U19882 ( .B1(n16860), .B2(n18464), .A(n16733), .ZN(P3_U2803) );
  XOR2_X1 U19883 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n16734), .Z(
        n16866) );
  INV_X1 U19884 ( .A(n16735), .ZN(n16745) );
  NOR2_X1 U19885 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18241), .ZN(
        n16862) );
  INV_X1 U19886 ( .A(n16862), .ZN(n16743) );
  AOI21_X1 U19887 ( .B1(n19188), .B2(n11623), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16736) );
  OAI22_X1 U19888 ( .A1(n16737), .A2(n16736), .B1(n18748), .B2(n19426), .ZN(
        n16738) );
  INV_X1 U19889 ( .A(n16738), .ZN(n16742) );
  INV_X1 U19890 ( .A(n18277), .ZN(n16740) );
  INV_X1 U19891 ( .A(n17321), .ZN(n16739) );
  OAI21_X1 U19892 ( .B1(n18417), .B2(n16740), .A(n16739), .ZN(n16741) );
  OAI211_X1 U19893 ( .C1(n18360), .C2(n16743), .A(n16742), .B(n16741), .ZN(
        n16744) );
  AOI21_X1 U19894 ( .B1(n16745), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16744), .ZN(n16746) );
  OAI21_X1 U19895 ( .B1(n18464), .B2(n16866), .A(n16746), .ZN(P3_U2804) );
  OAI21_X1 U19896 ( .B1(n16749), .B2(n16748), .A(n16747), .ZN(n16876) );
  INV_X1 U19897 ( .A(n16876), .ZN(n16761) );
  INV_X1 U19898 ( .A(n18426), .ZN(n18256) );
  INV_X1 U19899 ( .A(n18671), .ZN(n18372) );
  NAND2_X1 U19900 ( .A1(n16750), .A2(n18372), .ZN(n18250) );
  INV_X1 U19901 ( .A(n18250), .ZN(n16751) );
  OAI22_X1 U19902 ( .A1(n16869), .A2(n18256), .B1(n16751), .B2(n18484), .ZN(
        n18266) );
  OR2_X1 U19903 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18267), .ZN(
        n16872) );
  INV_X1 U19904 ( .A(n18398), .ZN(n18316) );
  NOR2_X1 U19905 ( .A1(n18316), .A2(n16752), .ZN(n16756) );
  NOR2_X1 U19906 ( .A1(n18748), .A2(n19423), .ZN(n16875) );
  INV_X1 U19907 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U19908 ( .A1(n19188), .A2(n16752), .B1(n18396), .B2(n16753), .ZN(
        n16754) );
  NAND2_X1 U19909 ( .A1(n16754), .A2(n18547), .ZN(n18260) );
  AOI21_X1 U19910 ( .B1(n16740), .B2(n17346), .A(n18260), .ZN(n18246) );
  OAI22_X1 U19911 ( .A1(n18246), .A2(n18243), .B1(n18402), .B2(n17342), .ZN(
        n16755) );
  AOI211_X1 U19912 ( .C1(n16756), .C2(n18243), .A(n16875), .B(n16755), .ZN(
        n16757) );
  OAI21_X1 U19913 ( .B1(n16758), .B2(n16872), .A(n16757), .ZN(n16759) );
  AOI21_X1 U19914 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18266), .A(
        n16759), .ZN(n16760) );
  OAI21_X1 U19915 ( .B1(n16761), .B2(n18464), .A(n16760), .ZN(P3_U2806) );
  NAND2_X1 U19916 ( .A1(n18368), .A2(n11633), .ZN(n18755) );
  INV_X1 U19917 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16765) );
  INV_X1 U19918 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18465) );
  NOR2_X1 U19919 ( .A1(n16762), .A2(n18465), .ZN(n16763) );
  NAND2_X1 U19920 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16763), .ZN(
        n17529) );
  NOR2_X1 U19921 ( .A1(n16765), .A2(n17529), .ZN(n17503) );
  AOI21_X1 U19922 ( .B1(n16765), .B2(n17529), .A(n17503), .ZN(n17521) );
  NOR2_X1 U19923 ( .A1(n16740), .A2(n18417), .ZN(n18264) );
  INV_X1 U19924 ( .A(n18547), .ZN(n18530) );
  AOI21_X1 U19925 ( .B1(n18859), .B2(n16762), .A(n18530), .ZN(n18467) );
  NAND2_X1 U19926 ( .A1(n18846), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18780) );
  OAI211_X1 U19927 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n16763), .A(
        n19188), .B(n18440), .ZN(n16764) );
  OAI211_X1 U19928 ( .C1(n18467), .C2(n16765), .A(n18780), .B(n16764), .ZN(
        n16769) );
  XNOR2_X1 U19929 ( .A(n18755), .B(n18367), .ZN(n18758) );
  OAI21_X1 U19930 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16767), .A(
        n16766), .ZN(n18763) );
  OAI22_X1 U19931 ( .A1(n18758), .A2(n18464), .B1(n18484), .B2(n18763), .ZN(
        n16768) );
  AOI211_X1 U19932 ( .C1(n17521), .C2(n18558), .A(n16769), .B(n16768), .ZN(
        n16770) );
  OAI21_X1 U19933 ( .B1(n18256), .B2(n18755), .A(n16770), .ZN(P3_U2822) );
  NOR2_X1 U19934 ( .A1(n16772), .A2(n18104), .ZN(n18757) );
  NAND2_X1 U19935 ( .A1(n16903), .A2(n16842), .ZN(n18769) );
  INV_X1 U19936 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18776) );
  INV_X1 U19937 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18840) );
  INV_X1 U19938 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18849) );
  NOR2_X1 U19939 ( .A1(n18840), .A2(n18849), .ZN(n18768) );
  NAND3_X1 U19940 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18789) );
  NOR3_X1 U19941 ( .A1(n11379), .A2(n18765), .A3(n18789), .ZN(n18777) );
  NAND2_X1 U19942 ( .A1(n18768), .A2(n18777), .ZN(n18743) );
  OR2_X1 U19943 ( .A1(n18776), .A2(n18743), .ZN(n18695) );
  NOR2_X1 U19944 ( .A1(n16850), .A2(n18695), .ZN(n18626) );
  NAND2_X1 U19945 ( .A1(n16852), .A2(n18626), .ZN(n16843) );
  OAI21_X1 U19946 ( .B1(n16843), .B2(n16836), .A(n16903), .ZN(n16774) );
  OAI21_X1 U19947 ( .B1(n16843), .B2(n16853), .A(n18851), .ZN(n16773) );
  OAI21_X1 U19948 ( .B1(n18849), .B2(n16842), .A(n18840), .ZN(n18775) );
  NAND3_X1 U19949 ( .A1(n18775), .A2(n18777), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18678) );
  INV_X1 U19950 ( .A(n18678), .ZN(n18650) );
  NAND2_X1 U19951 ( .A1(n16835), .A2(n18650), .ZN(n18628) );
  OR2_X1 U19952 ( .A1(n16873), .A2(n18628), .ZN(n18565) );
  OAI21_X1 U19953 ( .B1(n18565), .B2(n16853), .A(n19300), .ZN(n16841) );
  NAND4_X1 U19954 ( .A1(n18769), .A2(n16774), .A3(n16773), .A4(n16841), .ZN(
        n16807) );
  OR2_X1 U19955 ( .A1(n18773), .A2(n18834), .ZN(n18806) );
  NOR2_X1 U19956 ( .A1(n18806), .A2(n16775), .ZN(n16776) );
  AOI211_X1 U19957 ( .C1(n18813), .C2(n16807), .A(n18848), .B(n16776), .ZN(
        n16800) );
  NAND2_X1 U19958 ( .A1(n16777), .A2(n18845), .ZN(n16788) );
  INV_X1 U19959 ( .A(n16778), .ZN(n16786) );
  INV_X1 U19960 ( .A(n18806), .ZN(n18850) );
  INV_X1 U19961 ( .A(n19300), .ZN(n18766) );
  AOI21_X1 U19962 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16903), .A(
        n18851), .ZN(n18823) );
  OAI22_X1 U19963 ( .A1(n18766), .A2(n18565), .B1(n18823), .B2(n16843), .ZN(
        n16779) );
  NAND2_X1 U19964 ( .A1(n18563), .A2(n16779), .ZN(n18568) );
  INV_X1 U19965 ( .A(n16780), .ZN(n16781) );
  NAND2_X1 U19966 ( .A1(n16781), .A2(n16844), .ZN(n16782) );
  NOR4_X1 U19967 ( .A1(n18568), .A2(n18834), .A3(n16783), .A4(n16782), .ZN(
        n16784) );
  AOI211_X1 U19968 ( .C1(n16786), .C2(n18850), .A(n16785), .B(n16784), .ZN(
        n16787) );
  OAI211_X1 U19969 ( .C1(n16800), .C2(n16895), .A(n16788), .B(n16787), .ZN(
        n16789) );
  AOI21_X1 U19970 ( .B1(n16790), .B2(n18757), .A(n16789), .ZN(n16791) );
  OAI21_X1 U19971 ( .B1(n16792), .B2(n18753), .A(n16791), .ZN(P3_U2831) );
  NAND2_X1 U19972 ( .A1(n16846), .A2(n18757), .ZN(n16795) );
  INV_X1 U19973 ( .A(n18568), .ZN(n16793) );
  NAND3_X1 U19974 ( .A1(n16793), .A2(n18813), .A3(n16844), .ZN(n16794) );
  OAI211_X1 U19975 ( .C1(n16796), .C2(n18833), .A(n16795), .B(n16794), .ZN(
        n16815) );
  AOI22_X1 U19976 ( .A1(n16798), .A2(n18757), .B1(n18845), .B2(n16797), .ZN(
        n16806) );
  AOI21_X1 U19977 ( .B1(n16806), .B2(n16800), .A(n16799), .ZN(n16801) );
  AOI211_X1 U19978 ( .C1(n16803), .C2(n16815), .A(n16802), .B(n16801), .ZN(
        n16804) );
  OAI21_X1 U19979 ( .B1(n18753), .B2(n16805), .A(n16804), .ZN(P3_U2832) );
  INV_X1 U19980 ( .A(n16806), .ZN(n16811) );
  INV_X1 U19981 ( .A(n18736), .ZN(n18652) );
  AOI21_X1 U19982 ( .B1(n16854), .B2(n18652), .A(n16807), .ZN(n16821) );
  INV_X1 U19983 ( .A(n18773), .ZN(n18771) );
  NAND3_X1 U19984 ( .A1(n18771), .A2(n16808), .A3(n18748), .ZN(n16809) );
  OAI211_X1 U19985 ( .C1(n16821), .C2(n18846), .A(n16809), .B(n18839), .ZN(
        n16810) );
  OAI21_X1 U19986 ( .B1(n16811), .B2(n16810), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16819) );
  NAND2_X1 U19987 ( .A1(n16812), .A2(n18760), .ZN(n16818) );
  NAND3_X1 U19988 ( .A1(n16815), .A2(n16814), .A3(n16813), .ZN(n16816) );
  NAND4_X1 U19989 ( .A1(n16819), .A2(n16818), .A3(n16817), .A4(n16816), .ZN(
        P3_U2833) );
  INV_X1 U19990 ( .A(n19295), .ZN(n18829) );
  OAI211_X1 U19991 ( .C1(n16820), .C2(n16830), .A(n18829), .B(n18104), .ZN(
        n16826) );
  INV_X1 U19992 ( .A(n19298), .ZN(n18700) );
  OAI211_X1 U19993 ( .C1(n16822), .C2(n18700), .A(n16821), .B(n18839), .ZN(
        n16823) );
  AOI21_X1 U19994 ( .B1(n18661), .B2(n16824), .A(n16823), .ZN(n16825) );
  OAI21_X1 U19995 ( .B1(n16828), .B2(n16826), .A(n16825), .ZN(n16827) );
  NAND3_X1 U19996 ( .A1(n16827), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18748), .ZN(n16840) );
  INV_X1 U19997 ( .A(n16828), .ZN(n16832) );
  OAI21_X1 U19998 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16830), .A(
        n16829), .ZN(n16831) );
  NAND3_X1 U19999 ( .A1(n16832), .A2(n18760), .A3(n16831), .ZN(n16839) );
  INV_X1 U20000 ( .A(n18373), .ZN(n18721) );
  INV_X1 U20001 ( .A(n18768), .ZN(n16833) );
  OAI21_X1 U20002 ( .B1(n18823), .B2(n16833), .A(n18766), .ZN(n18774) );
  NAND2_X1 U20003 ( .A1(n18650), .A2(n18774), .ZN(n18684) );
  OAI21_X1 U20004 ( .B1(n18721), .B2(n18700), .A(n18684), .ZN(n16834) );
  OR4_X1 U20005 ( .A1(n18659), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16873), .A4(n16836), .ZN(n16838) );
  NAND4_X1 U20006 ( .A1(n16840), .A2(n16839), .A3(n16838), .A4(n16837), .ZN(
        P3_U2834) );
  INV_X1 U20007 ( .A(n16841), .ZN(n16849) );
  NOR2_X1 U20008 ( .A1(n18851), .A2(n16903), .ZN(n18767) );
  INV_X1 U20009 ( .A(n18767), .ZN(n18634) );
  NOR2_X1 U20010 ( .A1(n16842), .A2(n18695), .ZN(n18747) );
  INV_X1 U20011 ( .A(n18747), .ZN(n18676) );
  NOR2_X1 U20012 ( .A1(n16850), .A2(n18676), .ZN(n18649) );
  AOI21_X1 U20013 ( .B1(n18273), .B2(n18649), .A(n18746), .ZN(n18596) );
  AOI21_X1 U20014 ( .B1(n18634), .B2(n16843), .A(n18596), .ZN(n16868) );
  OAI21_X1 U20015 ( .B1(n18563), .B2(n18767), .A(n16868), .ZN(n18564) );
  OAI22_X1 U20016 ( .A1(n18585), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18746), .B2(n16844), .ZN(n16848) );
  OAI22_X1 U20017 ( .A1(n16846), .A2(n18723), .B1(n16845), .B2(n18700), .ZN(
        n16847) );
  NOR4_X1 U20018 ( .A1(n16849), .A2(n18564), .A3(n16848), .A4(n16847), .ZN(
        n16861) );
  OAI211_X1 U20019 ( .C1(n18585), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n16861), .ZN(n16858) );
  NOR2_X1 U20020 ( .A1(n16851), .A2(n16850), .ZN(n18590) );
  NAND2_X1 U20021 ( .A1(n16852), .A2(n18590), .ZN(n18578) );
  AOI221_X1 U20022 ( .B1(n16853), .B2(n16854), .C1(n18578), .C2(n16854), .A(
        n18834), .ZN(n16857) );
  NOR2_X1 U20023 ( .A1(n18839), .A2(n16854), .ZN(n16855) );
  AOI211_X1 U20024 ( .C1(n16858), .C2(n16857), .A(n16856), .B(n16855), .ZN(
        n16859) );
  OAI21_X1 U20025 ( .B1(n16860), .B2(n18753), .A(n16859), .ZN(P3_U2835) );
  INV_X1 U20026 ( .A(n16861), .ZN(n16863) );
  INV_X1 U20027 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16864) );
  OAI22_X1 U20028 ( .A1(n18839), .A2(n16864), .B1(n18748), .B2(n19426), .ZN(
        n16865) );
  AOI21_X1 U20029 ( .B1(n19298), .B2(n18250), .A(n18848), .ZN(n16867) );
  OAI211_X1 U20030 ( .C1(n16869), .C2(n18723), .A(n16868), .B(n16867), .ZN(
        n16871) );
  AOI211_X1 U20031 ( .C1(n19300), .C2(n18565), .A(n18267), .B(n16871), .ZN(
        n16870) );
  NOR2_X1 U20032 ( .A1(n18846), .A2(n16870), .ZN(n18579) );
  OAI211_X1 U20033 ( .C1(n16871), .C2(n18771), .A(n18579), .B(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16878) );
  NOR3_X1 U20034 ( .A1(n18659), .A2(n16873), .A3(n16872), .ZN(n16874) );
  AOI211_X1 U20035 ( .C1(n16876), .C2(n18760), .A(n16875), .B(n16874), .ZN(
        n16877) );
  NAND2_X1 U20036 ( .A1(n16878), .A2(n16877), .ZN(P3_U2838) );
  NOR3_X1 U20037 ( .A1(n19472), .A2(n19475), .A3(n16879), .ZN(n19448) );
  NOR2_X1 U20038 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19452), .ZN(n19449) );
  NOR2_X1 U20039 ( .A1(n19471), .A2(n18189), .ZN(n19339) );
  OAI21_X1 U20040 ( .B1(n9892), .B2(n19339), .A(n19470), .ZN(n18132) );
  OAI21_X1 U20041 ( .B1(n16881), .B2(n18132), .A(n16880), .ZN(n16882) );
  NOR3_X1 U20042 ( .A1(n16884), .A2(n16883), .A3(n16882), .ZN(n19319) );
  INV_X1 U20043 ( .A(n19469), .ZN(n19337) );
  NOR2_X1 U20044 ( .A1(n19319), .A2(n19337), .ZN(n16885) );
  AOI211_X2 U20045 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n19448), .A(n19449), .B(
        n16885), .ZN(n16935) );
  NAND2_X1 U20046 ( .A1(n19342), .A2(n16909), .ZN(n16890) );
  INV_X1 U20047 ( .A(n16935), .ZN(n17055) );
  NAND2_X1 U20048 ( .A1(n18746), .A2(n16886), .ZN(n16891) );
  MUX2_X1 U20049 ( .A(n18851), .B(n16891), .S(n16909), .Z(n19316) );
  AOI21_X1 U20050 ( .B1(n19316), .B2(n19452), .A(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n16887) );
  NAND2_X1 U20051 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16920) );
  INV_X1 U20052 ( .A(n16920), .ZN(n16896) );
  OAI21_X1 U20053 ( .B1(n16887), .B2(n16896), .A(n17055), .ZN(n16888) );
  OAI21_X1 U20054 ( .B1(n17055), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n16888), .ZN(n16889) );
  OAI21_X1 U20055 ( .B1(n16935), .B2(n16890), .A(n16889), .ZN(P3_U3290) );
  XNOR2_X1 U20056 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17591) );
  INV_X1 U20057 ( .A(n16891), .ZN(n16894) );
  NOR2_X1 U20058 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18851), .ZN(
        n16923) );
  INV_X1 U20059 ( .A(n16923), .ZN(n16892) );
  NAND2_X1 U20060 ( .A1(n16900), .A2(n16892), .ZN(n16893) );
  OAI21_X1 U20061 ( .B1(n17591), .B2(n16894), .A(n16893), .ZN(n19312) );
  INV_X1 U20062 ( .A(n19342), .ZN(n16929) );
  AOI22_X1 U20063 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18849), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16895), .ZN(n16919) );
  NAND2_X1 U20064 ( .A1(n16896), .A2(n16919), .ZN(n16897) );
  OAI211_X1 U20065 ( .C1(n16929), .C2(n17591), .A(n17055), .B(n16897), .ZN(
        n16898) );
  AOI21_X1 U20066 ( .B1(n17052), .B2(n19312), .A(n16898), .ZN(n16899) );
  AOI21_X1 U20067 ( .B1(n16935), .B2(n16900), .A(n16899), .ZN(P3_U3289) );
  NOR2_X1 U20068 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16901) );
  OR2_X1 U20069 ( .A1(n16902), .A2(n16901), .ZN(n16927) );
  NOR2_X1 U20070 ( .A1(n16927), .A2(n16930), .ZN(n17576) );
  NAND2_X1 U20071 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n16903), .ZN(
        n16905) );
  INV_X1 U20072 ( .A(n16904), .ZN(n16912) );
  AOI21_X1 U20073 ( .B1(n16905), .B2(n16914), .A(n16912), .ZN(n16918) );
  AOI21_X1 U20074 ( .B1(n16908), .B2(n16907), .A(n16906), .ZN(n16925) );
  AOI21_X1 U20075 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n16909), .A(
        n16911), .ZN(n16910) );
  NOR2_X1 U20076 ( .A1(n16925), .A2(n16910), .ZN(n16917) );
  INV_X1 U20077 ( .A(n16911), .ZN(n16913) );
  AOI21_X1 U20078 ( .B1(n16913), .B2(n16912), .A(n17051), .ZN(n16916) );
  OAI22_X1 U20079 ( .A1(n16914), .A2(n16913), .B1(n18766), .B2(n17576), .ZN(
        n16915) );
  NOR4_X1 U20080 ( .A1(n16918), .A2(n16917), .A3(n16916), .A4(n16915), .ZN(
        n19320) );
  OAI22_X1 U20081 ( .A1(n19320), .A2(n16931), .B1(n16920), .B2(n16919), .ZN(
        n16921) );
  AOI211_X1 U20082 ( .C1(n19342), .C2(n17576), .A(n16921), .B(n16935), .ZN(
        n16922) );
  AOI21_X1 U20083 ( .B1(n16935), .B2(n9896), .A(n16922), .ZN(P3_U3288) );
  INV_X1 U20084 ( .A(n17046), .ZN(n16928) );
  OAI22_X1 U20085 ( .A1(n16923), .A2(n16928), .B1(n18766), .B2(n16927), .ZN(
        n19303) );
  NOR2_X1 U20086 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n16931), .ZN(
        n16924) );
  AOI22_X1 U20087 ( .A1(n19303), .A2(n16924), .B1(n17872), .B2(n19342), .ZN(
        n16934) );
  NOR2_X1 U20088 ( .A1(n16925), .A2(n16930), .ZN(n16926) );
  AOI211_X1 U20089 ( .C1(n18851), .C2(n16928), .A(n16927), .B(n16926), .ZN(
        n19304) );
  OAI22_X1 U20090 ( .A1(n19304), .A2(n16931), .B1(n16930), .B2(n16929), .ZN(
        n16932) );
  OAI21_X1 U20091 ( .B1(n16935), .B2(n16932), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16933) );
  OAI21_X1 U20092 ( .B1(n16935), .B2(n16934), .A(n16933), .ZN(P3_U3285) );
  INV_X1 U20093 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17608) );
  INV_X1 U20094 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17606) );
  INV_X1 U20095 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17375) );
  NAND2_X1 U20096 ( .A1(n19471), .A2(n19469), .ZN(n16936) );
  NOR3_X4 U20097 ( .A1(n18873), .A2(n16937), .A3(n16936), .ZN(n17981) );
  NAND3_X1 U20098 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .ZN(n17773) );
  INV_X1 U20099 ( .A(n17773), .ZN(n16940) );
  INV_X1 U20100 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17585) );
  NAND2_X1 U20101 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17976) );
  NOR2_X1 U20102 ( .A1(n17585), .A2(n17976), .ZN(n17969) );
  NAND3_X1 U20103 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17969), .ZN(n17968) );
  NAND2_X1 U20104 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17958) );
  NAND4_X1 U20105 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n16938) );
  NOR4_X1 U20106 ( .A1(n17457), .A2(n17968), .A3(n17958), .A4(n16938), .ZN(
        n16939) );
  NAND4_X1 U20107 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(n16940), .A4(n16939), .ZN(n17788) );
  NOR3_X1 U20108 ( .A1(n17415), .A2(n17984), .A3(n17788), .ZN(n17757) );
  NAND2_X1 U20109 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17757), .ZN(n17737) );
  NAND2_X1 U20110 ( .A1(n18910), .A2(n17756), .ZN(n17733) );
  NOR2_X1 U20111 ( .A1(n17375), .A2(n17733), .ZN(n17718) );
  NAND2_X1 U20112 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17718), .ZN(n17695) );
  NAND2_X1 U20113 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17673), .ZN(n17667) );
  NAND2_X1 U20114 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17666), .ZN(n17657) );
  NAND2_X1 U20115 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17662), .ZN(n17031) );
  NOR2_X2 U20116 ( .A1(n18910), .A2(n17984), .ZN(n17985) );
  NOR2_X1 U20117 ( .A1(n17985), .A2(n17651), .ZN(n17652) );
  AOI22_X1 U20118 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16941) );
  OAI21_X1 U20119 ( .B1(n16942), .B2(n17708), .A(n16941), .ZN(n16943) );
  AOI21_X1 U20120 ( .B1(n17872), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n16943), .ZN(n16946) );
  AOI22_X1 U20121 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20122 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16944) );
  NAND3_X1 U20123 ( .A1(n16946), .A2(n16945), .A3(n16944), .ZN(n16955) );
  AOI22_X1 U20124 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16948) );
  NAND2_X1 U20125 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n16947) );
  OAI211_X1 U20126 ( .C1(n16949), .C2(n17950), .A(n16948), .B(n16947), .ZN(
        n16953) );
  INV_X1 U20127 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16950) );
  OAI22_X1 U20128 ( .A1(n9754), .A2(n16950), .B1(n17818), .B2(n17711), .ZN(
        n16952) );
  INV_X1 U20129 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17698) );
  INV_X1 U20130 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17707) );
  OAI22_X1 U20131 ( .A1(n9668), .A2(n17698), .B1(n17918), .B2(n17707), .ZN(
        n16951) );
  OR3_X1 U20132 ( .A1(n16953), .A2(n16952), .A3(n16951), .ZN(n16954) );
  NOR2_X1 U20133 ( .A1(n16955), .A2(n16954), .ZN(n17029) );
  AOI22_X1 U20134 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16959) );
  AOI22_X1 U20135 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20136 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20137 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16956) );
  NAND4_X1 U20138 ( .A1(n16959), .A2(n16958), .A3(n16957), .A4(n16956), .ZN(
        n16968) );
  INV_X1 U20139 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16966) );
  INV_X1 U20140 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17746) );
  OAI22_X1 U20141 ( .A1(n17709), .A2(n16960), .B1(n17799), .B2(n17746), .ZN(
        n16963) );
  INV_X1 U20142 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17745) );
  OAI22_X1 U20143 ( .A1(n9754), .A2(n16961), .B1(n17943), .B2(n17745), .ZN(
        n16962) );
  AOI211_X1 U20144 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n16963), .B(n16962), .ZN(n16965) );
  AOI22_X1 U20145 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16964) );
  OAI211_X1 U20146 ( .C1(n17950), .C2(n16966), .A(n16965), .B(n16964), .ZN(
        n16967) );
  NOR2_X1 U20147 ( .A1(n16968), .A2(n16967), .ZN(n17659) );
  INV_X1 U20148 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16973) );
  INV_X1 U20149 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17908) );
  INV_X1 U20150 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17907) );
  OAI22_X1 U20151 ( .A1(n11436), .A2(n17908), .B1(n9668), .B2(n17907), .ZN(
        n16970) );
  INV_X1 U20152 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17781) );
  OAI22_X1 U20153 ( .A1(n9666), .A2(n17909), .B1(n9754), .B2(n17781), .ZN(
        n16969) );
  AOI211_X1 U20154 ( .C1(n17872), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n16970), .B(n16969), .ZN(n16972) );
  AOI22_X1 U20155 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16971) );
  OAI211_X1 U20156 ( .C1(n17950), .C2(n16973), .A(n16972), .B(n16971), .ZN(
        n16979) );
  AOI22_X1 U20157 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20158 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20159 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20160 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16974) );
  NAND4_X1 U20161 ( .A1(n16977), .A2(n16976), .A3(n16975), .A4(n16974), .ZN(
        n16978) );
  NOR2_X1 U20162 ( .A1(n16979), .A2(n16978), .ZN(n17669) );
  INV_X1 U20163 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17801) );
  OAI22_X1 U20164 ( .A1(n17941), .A2(n17801), .B1(n17939), .B2(n16980), .ZN(
        n16982) );
  INV_X1 U20165 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17944) );
  OAI22_X1 U20166 ( .A1(n17747), .A2(n17944), .B1(n17799), .B2(n17800), .ZN(
        n16981) );
  AOI211_X1 U20167 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n16982), .B(n16981), .ZN(n16990) );
  AOI22_X1 U20168 ( .A1(n11447), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20169 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20170 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20171 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16983) );
  AND4_X1 U20172 ( .A1(n16986), .A2(n16985), .A3(n16984), .A4(n16983), .ZN(
        n16989) );
  AOI22_X1 U20173 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16988) );
  NAND2_X1 U20174 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n16987) );
  NAND4_X1 U20175 ( .A1(n16990), .A2(n16989), .A3(n16988), .A4(n16987), .ZN(
        n17675) );
  INV_X1 U20176 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17629) );
  INV_X1 U20177 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16991) );
  OAI22_X1 U20178 ( .A1(n17629), .A2(n17941), .B1(n17939), .B2(n16991), .ZN(
        n16995) );
  INV_X1 U20179 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16993) );
  INV_X1 U20180 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16992) );
  OAI22_X1 U20181 ( .A1(n16993), .A2(n17747), .B1(n17799), .B2(n16992), .ZN(
        n16994) );
  AOI211_X1 U20182 ( .C1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .C2(n17872), .A(
        n16995), .B(n16994), .ZN(n17004) );
  AOI22_X1 U20183 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20184 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17878), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20185 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n17921), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20186 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16997) );
  AND4_X1 U20187 ( .A1(n17000), .A2(n16999), .A3(n16998), .A4(n16997), .ZN(
        n17003) );
  AOI22_X1 U20188 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17002) );
  NAND2_X1 U20189 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n17001) );
  NAND4_X1 U20190 ( .A1(n17004), .A2(n17003), .A3(n17002), .A4(n17001), .ZN(
        n17676) );
  NAND2_X1 U20191 ( .A1(n17675), .A2(n17676), .ZN(n17674) );
  NOR2_X1 U20192 ( .A1(n17669), .A2(n17674), .ZN(n17668) );
  INV_X1 U20193 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17766) );
  INV_X1 U20194 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17890) );
  OAI22_X1 U20195 ( .A1(n17941), .A2(n17766), .B1(n17939), .B2(n17890), .ZN(
        n17007) );
  INV_X1 U20196 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17759) );
  INV_X1 U20197 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17005) );
  OAI22_X1 U20198 ( .A1(n17747), .A2(n17759), .B1(n17799), .B2(n17005), .ZN(
        n17006) );
  AOI211_X1 U20199 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17007), .B(n17006), .ZN(n17015) );
  AOI22_X1 U20200 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20201 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20202 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20203 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17008) );
  AND4_X1 U20204 ( .A1(n17011), .A2(n17010), .A3(n17009), .A4(n17008), .ZN(
        n17014) );
  AOI22_X1 U20205 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17013) );
  NAND2_X1 U20206 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n17012) );
  NAND4_X1 U20207 ( .A1(n17015), .A2(n17014), .A3(n17013), .A4(n17012), .ZN(
        n17664) );
  NAND2_X1 U20208 ( .A1(n17668), .A2(n17664), .ZN(n17663) );
  NOR2_X1 U20209 ( .A1(n17659), .A2(n17663), .ZN(n17658) );
  INV_X1 U20210 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17016) );
  OAI22_X1 U20211 ( .A1(n17941), .A2(n17017), .B1(n17939), .B2(n17016), .ZN(
        n17019) );
  INV_X1 U20212 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21429) );
  INV_X1 U20213 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17856) );
  OAI22_X1 U20214 ( .A1(n21429), .A2(n17747), .B1(n17799), .B2(n17856), .ZN(
        n17018) );
  AOI211_X1 U20215 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17019), .B(n17018), .ZN(n17028) );
  AOI22_X1 U20216 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20217 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20218 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20219 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17021) );
  AND4_X1 U20220 ( .A1(n17024), .A2(n17023), .A3(n17022), .A4(n17021), .ZN(
        n17027) );
  AOI22_X1 U20221 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17026) );
  NAND2_X1 U20222 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n17025) );
  NAND4_X1 U20223 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17655) );
  NAND2_X1 U20224 ( .A1(n17658), .A2(n17655), .ZN(n17654) );
  NOR2_X1 U20225 ( .A1(n17029), .A2(n17654), .ZN(n17649) );
  AOI21_X1 U20226 ( .B1(n17029), .B2(n17654), .A(n17649), .ZN(n18002) );
  AOI22_X1 U20227 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17652), .B1(n18002), 
        .B2(n17985), .ZN(n17030) );
  OAI21_X1 U20228 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17031), .A(n17030), .ZN(
        P3_U2675) );
  INV_X1 U20229 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17953) );
  NAND2_X1 U20230 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17967), .ZN(n17957) );
  NAND3_X1 U20231 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(n17906), .ZN(n17032) );
  AOI21_X1 U20232 ( .B1(n17457), .B2(n17032), .A(n17844), .ZN(n17045) );
  INV_X1 U20233 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17696) );
  OAI22_X1 U20234 ( .A1(n17941), .A2(n17696), .B1(n17939), .B2(n17707), .ZN(
        n17035) );
  INV_X1 U20235 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17697) );
  INV_X1 U20236 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17033) );
  OAI22_X1 U20237 ( .A1(n17747), .A2(n17697), .B1(n17799), .B2(n17033), .ZN(
        n17034) );
  AOI211_X1 U20238 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n17035), .B(n17034), .ZN(n17044) );
  AOI22_X1 U20239 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20240 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17878), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20241 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20242 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17037) );
  AND4_X1 U20243 ( .A1(n17040), .A2(n17039), .A3(n17038), .A4(n17037), .ZN(
        n17043) );
  AOI22_X1 U20244 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17867), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17042) );
  NAND2_X1 U20245 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n17041) );
  NAND4_X1 U20246 ( .A1(n17044), .A2(n17043), .A3(n17042), .A4(n17041), .ZN(
        n18080) );
  MUX2_X1 U20247 ( .A(n17045), .B(n18080), .S(n17985), .Z(P3_U2690) );
  NOR2_X1 U20248 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19452), .ZN(
        n18915) );
  AOI21_X1 U20249 ( .B1(n17046), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17050) );
  NAND2_X1 U20250 ( .A1(n9668), .A2(n17050), .ZN(n18857) );
  INV_X1 U20251 ( .A(n18857), .ZN(n17047) );
  INV_X1 U20252 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17258) );
  NAND2_X1 U20253 ( .A1(n17047), .A2(n17258), .ZN(n17048) );
  AOI21_X1 U20254 ( .B1(n19448), .B2(n17048), .A(n19216), .ZN(n18869) );
  NOR2_X1 U20255 ( .A1(n18915), .A2(n18869), .ZN(n18860) );
  INV_X1 U20256 ( .A(n19159), .ZN(n19214) );
  INV_X1 U20257 ( .A(n18869), .ZN(n18863) );
  OAI22_X1 U20258 ( .A1(n19468), .A2(n18859), .B1(n11545), .B2(n19452), .ZN(
        n18864) );
  NAND3_X1 U20259 ( .A1(n19311), .A2(n18863), .A3(n18864), .ZN(n17049) );
  OAI221_X1 U20260 ( .B1(n19311), .B2(n18860), .C1(n19311), .C2(n19214), .A(
        n17049), .ZN(P3_U2864) );
  NOR2_X1 U20261 ( .A1(n17051), .A2(n17050), .ZN(n19302) );
  NAND3_X1 U20262 ( .A1(n17055), .A2(n17052), .A3(n19302), .ZN(n17053) );
  OAI21_X1 U20263 ( .B1(n17055), .B2(n17054), .A(n17053), .ZN(P3_U3284) );
  NOR2_X1 U20264 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17056), .ZN(n17091) );
  NOR3_X1 U20265 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21246), .A3(n21293), 
        .ZN(n17059) );
  OAI22_X1 U20266 ( .A1(n17084), .A2(n17059), .B1(n17058), .B2(n17057), .ZN(
        n17130) );
  OAI21_X1 U20267 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21293), .A(n17127), 
        .ZN(n17089) );
  INV_X1 U20268 ( .A(n17060), .ZN(n17062) );
  OAI211_X1 U20269 ( .C1(n10429), .C2(n17062), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17061), .ZN(n17065) );
  OAI211_X1 U20270 ( .C1(n21033), .C2(n17065), .A(n17064), .B(n17063), .ZN(
        n17067) );
  NAND2_X1 U20271 ( .A1(n21033), .A2(n17065), .ZN(n17066) );
  NAND2_X1 U20272 ( .A1(n17067), .A2(n17066), .ZN(n17068) );
  AND2_X1 U20273 ( .A1(n10743), .A2(n17068), .ZN(n17069) );
  OAI22_X1 U20274 ( .A1(n17070), .A2(n17069), .B1(n10743), .B2(n17068), .ZN(
        n17075) );
  NOR2_X1 U20275 ( .A1(n17072), .A2(n17071), .ZN(n17074) );
  INV_X1 U20276 ( .A(n17072), .ZN(n17073) );
  OAI22_X1 U20277 ( .A1(n17075), .A2(n17074), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17073), .ZN(n17083) );
  OAI21_X1 U20278 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17076), .ZN(n17077) );
  NAND4_X1 U20279 ( .A1(n17080), .A2(n17079), .A3(n17078), .A4(n17077), .ZN(
        n17081) );
  AOI211_X1 U20280 ( .C1(n17083), .C2(n20586), .A(n17082), .B(n17081), .ZN(
        n17087) );
  INV_X1 U20281 ( .A(n17084), .ZN(n21244) );
  INV_X1 U20282 ( .A(n17130), .ZN(n17085) );
  AOI21_X1 U20283 ( .B1(n17085), .B2(n17087), .A(n20351), .ZN(n21247) );
  OAI211_X1 U20284 ( .C1(n17087), .C2(n21244), .A(n21247), .B(n17086), .ZN(
        n17088) );
  OAI22_X1 U20285 ( .A1(n17125), .A2(n17130), .B1(n17089), .B2(n17088), .ZN(
        n17090) );
  AOI21_X1 U20286 ( .B1(n21296), .B2(n17091), .A(n17090), .ZN(P1_U3161) );
  AND2_X1 U20287 ( .A1(n20471), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U20288 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17092) );
  NOR2_X1 U20289 ( .A1(n17092), .A2(n20334), .ZN(P2_U3047) );
  AOI22_X1 U20290 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20580), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17098) );
  NAND2_X1 U20291 ( .A1(n17095), .A2(n17094), .ZN(n17096) );
  XNOR2_X1 U20292 ( .A(n17093), .B(n17096), .ZN(n17110) );
  AOI22_X1 U20293 ( .A1(n17110), .A2(n20518), .B1(n20376), .B2(n20519), .ZN(
        n17097) );
  OAI211_X1 U20294 ( .C1(n20524), .C2(n20374), .A(n17098), .B(n17097), .ZN(
        P1_U2992) );
  AOI22_X1 U20295 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20580), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17104) );
  XNOR2_X1 U20296 ( .A(n17101), .B(n17100), .ZN(n17102) );
  XNOR2_X1 U20297 ( .A(n17099), .B(n17102), .ZN(n17120) );
  AOI22_X1 U20298 ( .A1(n20445), .A2(n20519), .B1(n20518), .B2(n17120), .ZN(
        n17103) );
  OAI211_X1 U20299 ( .C1(n20524), .C2(n20391), .A(n17104), .B(n17103), .ZN(
        P1_U2993) );
  AOI22_X1 U20300 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20580), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17109) );
  INV_X1 U20301 ( .A(n17106), .ZN(n20404) );
  AOI22_X1 U20302 ( .A1(n17107), .A2(n20518), .B1(n20519), .B2(n20404), .ZN(
        n17108) );
  OAI211_X1 U20303 ( .C1(n20524), .C2(n20401), .A(n17109), .B(n17108), .ZN(
        P1_U2994) );
  INV_X1 U20304 ( .A(n20373), .ZN(n17111) );
  AOI222_X1 U20305 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20580), .B1(n20544), 
        .B2(n17111), .C1(n17110), .C2(n20550), .ZN(n17112) );
  OAI221_X1 U20306 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17115), .C1(
        n17114), .C2(n17113), .A(n17112), .ZN(P1_U3024) );
  AOI21_X1 U20307 ( .B1(n17117), .B2(n17116), .A(n9722), .ZN(n20444) );
  AOI22_X1 U20308 ( .A1(n20444), .A2(n20544), .B1(n20580), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n17122) );
  INV_X1 U20309 ( .A(n17118), .ZN(n17119) );
  AOI22_X1 U20310 ( .A1(n17120), .A2(n20550), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17119), .ZN(n17121) );
  OAI211_X1 U20311 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17123), .A(
        n17122), .B(n17121), .ZN(P1_U3025) );
  NAND4_X1 U20312 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21246), .A4(n21293), .ZN(n17124) );
  OAI21_X1 U20313 ( .B1(n17125), .B2(n20900), .A(n17124), .ZN(n21243) );
  NAND2_X1 U20314 ( .A1(n17126), .A2(n21246), .ZN(n17128) );
  OAI221_X1 U20315 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n21247), .C1(
        P1_STATE2_REG_1__SCAN_IN), .C2(n17128), .A(n17127), .ZN(n17129) );
  AOI221_X1 U20316 ( .B1(n17131), .B2(n17130), .C1(n21243), .C2(n17130), .A(
        n17129), .ZN(P1_U3162) );
  OAI21_X1 U20317 ( .B1(n21247), .B2(n21041), .A(n17132), .ZN(P1_U3466) );
  OAI22_X1 U20318 ( .A1(n17135), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n17134), .B2(n17133), .ZN(n17136) );
  INV_X1 U20319 ( .A(n17136), .ZN(n17144) );
  OAI21_X1 U20320 ( .B1(n17138), .B2(n19648), .A(n17137), .ZN(n17141) );
  NOR2_X1 U20321 ( .A1(n17139), .A2(n19653), .ZN(n17140) );
  AOI211_X1 U20322 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17142), .A(
        n17141), .B(n17140), .ZN(n17143) );
  OAI211_X1 U20323 ( .C1(n19668), .C2(n17145), .A(n17144), .B(n17143), .ZN(
        P2_U3039) );
  NOR2_X1 U20324 ( .A1(n17147), .A2(n17146), .ZN(n17150) );
  INV_X1 U20325 ( .A(n17148), .ZN(n17149) );
  AOI211_X1 U20326 ( .C1(n20338), .C2(n17151), .A(n17150), .B(n17149), .ZN(
        n17159) );
  INV_X1 U20327 ( .A(n17152), .ZN(n20300) );
  MUX2_X1 U20328 ( .A(n20300), .B(n17154), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n17157) );
  NAND3_X1 U20329 ( .A1(n17154), .A2(n17153), .A3(n20224), .ZN(n17155) );
  OAI21_X1 U20330 ( .B1(n17157), .B2(n17156), .A(n17155), .ZN(n17158) );
  OAI211_X1 U20331 ( .C1(n17161), .C2(n17160), .A(n17159), .B(n17158), .ZN(
        P2_U3176) );
  NOR3_X1 U20332 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n17163) );
  NOR4_X1 U20333 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17162) );
  INV_X2 U20334 ( .A(n17241), .ZN(U215) );
  NAND4_X1 U20335 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17163), .A3(n17162), .A4(
        U215), .ZN(U213) );
  INV_X1 U20336 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19587) );
  INV_X2 U20337 ( .A(U214), .ZN(n17204) );
  INV_X1 U20338 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17243) );
  OAI222_X1 U20339 ( .A1(U212), .A2(n19587), .B1(n17206), .B2(n20645), .C1(
        U214), .C2(n17243), .ZN(U216) );
  AOI222_X1 U20340 ( .A1(n17203), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17201), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17204), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17165) );
  INV_X1 U20341 ( .A(n17165), .ZN(U217) );
  AOI22_X1 U20342 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17203), .ZN(n17166) );
  OAI21_X1 U20343 ( .B1(n20628), .B2(n17206), .A(n17166), .ZN(U218) );
  AOI22_X1 U20344 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17203), .ZN(n17167) );
  OAI21_X1 U20345 ( .B1(n20620), .B2(n17206), .A(n17167), .ZN(U219) );
  AOI22_X1 U20346 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17203), .ZN(n17168) );
  OAI21_X1 U20347 ( .B1(n20610), .B2(n17206), .A(n17168), .ZN(U220) );
  AOI22_X1 U20348 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17203), .ZN(n17169) );
  OAI21_X1 U20349 ( .B1(n21377), .B2(n17206), .A(n17169), .ZN(U221) );
  INV_X1 U20350 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n21332) );
  INV_X1 U20351 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n17170) );
  OAI222_X1 U20352 ( .A1(U212), .A2(n21332), .B1(n17206), .B2(n20598), .C1(
        U214), .C2(n17170), .ZN(U222) );
  AOI22_X1 U20353 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17203), .ZN(n17171) );
  OAI21_X1 U20354 ( .B1(n20588), .B2(n17206), .A(n17171), .ZN(U223) );
  AOI22_X1 U20355 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17203), .ZN(n17172) );
  OAI21_X1 U20356 ( .B1(n20642), .B2(n17206), .A(n17172), .ZN(U224) );
  AOI22_X1 U20357 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17203), .ZN(n17173) );
  OAI21_X1 U20358 ( .B1(n20635), .B2(n17206), .A(n17173), .ZN(U225) );
  AOI22_X1 U20359 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17203), .ZN(n17174) );
  OAI21_X1 U20360 ( .B1(n20625), .B2(n17206), .A(n17174), .ZN(U226) );
  AOI22_X1 U20361 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17203), .ZN(n17175) );
  OAI21_X1 U20362 ( .B1(n20618), .B2(n17206), .A(n17175), .ZN(U227) );
  AOI22_X1 U20363 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17203), .ZN(n17176) );
  OAI21_X1 U20364 ( .B1(n20608), .B2(n17206), .A(n17176), .ZN(U228) );
  AOI22_X1 U20365 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17203), .ZN(n17177) );
  OAI21_X1 U20366 ( .B1(n17178), .B2(n17206), .A(n17177), .ZN(U229) );
  AOI22_X1 U20367 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17203), .ZN(n17179) );
  OAI21_X1 U20368 ( .B1(n20601), .B2(n17206), .A(n17179), .ZN(U230) );
  AOI22_X1 U20369 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17203), .ZN(n17180) );
  OAI21_X1 U20370 ( .B1(n20593), .B2(n17206), .A(n17180), .ZN(U231) );
  AOI22_X1 U20371 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17203), .ZN(n17181) );
  OAI21_X1 U20372 ( .B1(n13978), .B2(n17206), .A(n17181), .ZN(U232) );
  INV_X1 U20373 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20374 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17203), .ZN(n17182) );
  OAI21_X1 U20375 ( .B1(n17183), .B2(n17206), .A(n17182), .ZN(U233) );
  INV_X1 U20376 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n21321) );
  AOI22_X1 U20377 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17201), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17203), .ZN(n17184) );
  OAI21_X1 U20378 ( .B1(n21321), .B2(U214), .A(n17184), .ZN(U234) );
  INV_X1 U20379 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17219) );
  INV_X1 U20380 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17185) );
  INV_X1 U20381 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n21323) );
  OAI222_X1 U20382 ( .A1(U212), .A2(n17219), .B1(n17206), .B2(n17185), .C1(
        U214), .C2(n21323), .ZN(U235) );
  INV_X1 U20383 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20384 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17201), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17204), .ZN(n17186) );
  OAI21_X1 U20385 ( .B1(n17218), .B2(U212), .A(n17186), .ZN(U236) );
  INV_X1 U20386 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20387 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17203), .ZN(n17187) );
  OAI21_X1 U20388 ( .B1(n17188), .B2(n17206), .A(n17187), .ZN(U237) );
  INV_X1 U20389 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20390 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17201), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17204), .ZN(n17189) );
  OAI21_X1 U20391 ( .B1(n17216), .B2(U212), .A(n17189), .ZN(U238) );
  INV_X1 U20392 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n21405) );
  INV_X1 U20393 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17191) );
  INV_X1 U20394 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n17190) );
  OAI222_X1 U20395 ( .A1(U212), .A2(n21405), .B1(n17206), .B2(n17191), .C1(
        U214), .C2(n17190), .ZN(U239) );
  INV_X1 U20396 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20397 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17201), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17204), .ZN(n17192) );
  OAI21_X1 U20398 ( .B1(n17215), .B2(U212), .A(n17192), .ZN(U240) );
  INV_X1 U20399 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20400 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17203), .ZN(n17193) );
  OAI21_X1 U20401 ( .B1(n17194), .B2(n17206), .A(n17193), .ZN(U241) );
  INV_X1 U20402 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20403 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17201), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17204), .ZN(n17195) );
  OAI21_X1 U20404 ( .B1(n17213), .B2(U212), .A(n17195), .ZN(U242) );
  INV_X1 U20405 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20406 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17203), .ZN(n17196) );
  OAI21_X1 U20407 ( .B1(n17197), .B2(n17206), .A(n17196), .ZN(U243) );
  INV_X1 U20408 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20409 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17201), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17204), .ZN(n17198) );
  OAI21_X1 U20410 ( .B1(n17211), .B2(U212), .A(n17198), .ZN(U244) );
  INV_X1 U20411 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20412 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17203), .ZN(n17199) );
  OAI21_X1 U20413 ( .B1(n17200), .B2(n17206), .A(n17199), .ZN(U245) );
  INV_X1 U20414 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20415 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17201), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17204), .ZN(n17202) );
  OAI21_X1 U20416 ( .B1(n17209), .B2(U212), .A(n17202), .ZN(U246) );
  INV_X1 U20417 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20418 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17204), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17203), .ZN(n17205) );
  OAI21_X1 U20419 ( .B1(n17207), .B2(n17206), .A(n17205), .ZN(U247) );
  INV_X1 U20420 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20421 ( .A1(n17241), .A2(n17208), .B1(n18871), .B2(U215), .ZN(U251) );
  AOI22_X1 U20422 ( .A1(n17227), .A2(n17209), .B1(n13926), .B2(U215), .ZN(U252) );
  INV_X1 U20423 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20424 ( .A1(n17241), .A2(n17210), .B1(n18881), .B2(U215), .ZN(U253) );
  AOI22_X1 U20425 ( .A1(n17241), .A2(n17211), .B1(n13585), .B2(U215), .ZN(U254) );
  INV_X1 U20426 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20427 ( .A1(n17241), .A2(n17212), .B1(n18891), .B2(U215), .ZN(U255) );
  AOI22_X1 U20428 ( .A1(n17227), .A2(n17213), .B1(n13582), .B2(U215), .ZN(U256) );
  INV_X1 U20429 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20430 ( .A1(n17241), .A2(n17214), .B1(n18902), .B2(U215), .ZN(U257) );
  AOI22_X1 U20431 ( .A1(n17227), .A2(n17215), .B1(n13588), .B2(U215), .ZN(U258) );
  AOI22_X1 U20432 ( .A1(n17227), .A2(n21405), .B1(n18222), .B2(U215), .ZN(U259) );
  AOI22_X1 U20433 ( .A1(n17227), .A2(n17216), .B1(n13579), .B2(U215), .ZN(U260) );
  INV_X1 U20434 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20435 ( .A1(n17227), .A2(n17217), .B1(n18225), .B2(U215), .ZN(U261) );
  AOI22_X1 U20436 ( .A1(n17227), .A2(n17218), .B1(n13620), .B2(U215), .ZN(U262) );
  AOI22_X1 U20437 ( .A1(n17227), .A2(n17219), .B1(n18231), .B2(U215), .ZN(U263) );
  OAI22_X1 U20438 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17241), .ZN(n17220) );
  INV_X1 U20439 ( .A(n17220), .ZN(U264) );
  OAI22_X1 U20440 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17241), .ZN(n17221) );
  INV_X1 U20441 ( .A(n17221), .ZN(U265) );
  OAI22_X1 U20442 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17241), .ZN(n17222) );
  INV_X1 U20443 ( .A(n17222), .ZN(U266) );
  INV_X1 U20444 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20445 ( .A1(n17241), .A2(n17223), .B1(n18870), .B2(U215), .ZN(U267) );
  INV_X1 U20446 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20447 ( .A1(n17227), .A2(n17224), .B1(n18877), .B2(U215), .ZN(U268) );
  INV_X1 U20448 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20449 ( .A1(n17241), .A2(n17225), .B1(n18882), .B2(U215), .ZN(U269) );
  INV_X1 U20450 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20451 ( .A1(n17227), .A2(n17226), .B1(n18886), .B2(U215), .ZN(U270) );
  INV_X1 U20452 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20453 ( .A1(n17241), .A2(n17228), .B1(n18892), .B2(U215), .ZN(U271) );
  INV_X1 U20454 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20455 ( .A1(n17241), .A2(n17229), .B1(n18895), .B2(U215), .ZN(U272) );
  INV_X1 U20456 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20457 ( .A1(n17241), .A2(n17230), .B1(n18903), .B2(U215), .ZN(U273) );
  INV_X1 U20458 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20459 ( .A1(n17241), .A2(n17231), .B1(n18907), .B2(U215), .ZN(U274) );
  INV_X1 U20460 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20461 ( .A1(n17241), .A2(n17233), .B1(n17232), .B2(U215), .ZN(U275) );
  AOI22_X1 U20462 ( .A1(n17241), .A2(n21332), .B1(n18876), .B2(U215), .ZN(U276) );
  INV_X1 U20463 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20464 ( .A1(n17241), .A2(n17234), .B1(n18015), .B2(U215), .ZN(U277) );
  INV_X1 U20465 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20466 ( .A1(n17241), .A2(n17235), .B1(n21324), .B2(U215), .ZN(U278) );
  INV_X1 U20467 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20468 ( .A1(n17241), .A2(n17236), .B1(n18890), .B2(U215), .ZN(U279) );
  INV_X1 U20469 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20470 ( .A1(n17241), .A2(n17238), .B1(n17237), .B2(U215), .ZN(U280) );
  INV_X1 U20471 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19591) );
  AOI22_X1 U20472 ( .A1(n17241), .A2(n19591), .B1(n18901), .B2(U215), .ZN(U281) );
  AOI22_X1 U20473 ( .A1(n17241), .A2(n19587), .B1(n17240), .B2(U215), .ZN(U282) );
  INV_X1 U20474 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17242) );
  AOI222_X1 U20475 ( .A1(n17243), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17242), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17244) );
  INV_X2 U20476 ( .A(n17246), .ZN(n17245) );
  INV_X1 U20477 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19395) );
  INV_X1 U20478 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20248) );
  AOI22_X1 U20479 ( .A1(n17245), .A2(n19395), .B1(n20248), .B2(n17246), .ZN(
        U347) );
  INV_X1 U20480 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19393) );
  INV_X1 U20481 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20246) );
  AOI22_X1 U20482 ( .A1(n17245), .A2(n19393), .B1(n20246), .B2(n17246), .ZN(
        U348) );
  INV_X1 U20483 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19390) );
  INV_X1 U20484 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20244) );
  AOI22_X1 U20485 ( .A1(n17245), .A2(n19390), .B1(n20244), .B2(n17246), .ZN(
        U349) );
  INV_X1 U20486 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19389) );
  INV_X1 U20487 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20242) );
  AOI22_X1 U20488 ( .A1(n17245), .A2(n19389), .B1(n20242), .B2(n17246), .ZN(
        U350) );
  INV_X1 U20489 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19387) );
  INV_X1 U20490 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20240) );
  AOI22_X1 U20491 ( .A1(n17245), .A2(n19387), .B1(n20240), .B2(n17246), .ZN(
        U351) );
  INV_X1 U20492 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19384) );
  INV_X1 U20493 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20238) );
  AOI22_X1 U20494 ( .A1(n17245), .A2(n19384), .B1(n20238), .B2(n17246), .ZN(
        U352) );
  INV_X1 U20495 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19383) );
  AOI22_X1 U20496 ( .A1(n17245), .A2(n19383), .B1(n20237), .B2(n17246), .ZN(
        U353) );
  INV_X1 U20497 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19381) );
  INV_X1 U20498 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20236) );
  AOI22_X1 U20499 ( .A1(n17245), .A2(n19381), .B1(n20236), .B2(n17246), .ZN(
        U354) );
  INV_X1 U20500 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19435) );
  INV_X1 U20501 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20283) );
  AOI22_X1 U20502 ( .A1(n17245), .A2(n19435), .B1(n20283), .B2(n17246), .ZN(
        U355) );
  INV_X1 U20503 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19432) );
  INV_X1 U20504 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20280) );
  AOI22_X1 U20505 ( .A1(n17245), .A2(n19432), .B1(n20280), .B2(n17246), .ZN(
        U356) );
  INV_X1 U20506 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19429) );
  INV_X1 U20507 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20278) );
  AOI22_X1 U20508 ( .A1(n17245), .A2(n19429), .B1(n20278), .B2(n17246), .ZN(
        U357) );
  INV_X1 U20509 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19428) );
  INV_X1 U20510 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21349) );
  AOI22_X1 U20511 ( .A1(n17245), .A2(n19428), .B1(n21349), .B2(n17246), .ZN(
        U358) );
  INV_X1 U20512 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19425) );
  INV_X1 U20513 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20275) );
  AOI22_X1 U20514 ( .A1(n17245), .A2(n19425), .B1(n20275), .B2(n17246), .ZN(
        U359) );
  INV_X1 U20515 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19424) );
  INV_X1 U20516 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20273) );
  AOI22_X1 U20517 ( .A1(n17245), .A2(n19424), .B1(n20273), .B2(n17246), .ZN(
        U360) );
  INV_X1 U20518 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19422) );
  INV_X1 U20519 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20271) );
  AOI22_X1 U20520 ( .A1(n17245), .A2(n19422), .B1(n20271), .B2(n17246), .ZN(
        U361) );
  INV_X1 U20521 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19420) );
  INV_X1 U20522 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20269) );
  AOI22_X1 U20523 ( .A1(n17245), .A2(n19420), .B1(n20269), .B2(n17246), .ZN(
        U362) );
  INV_X1 U20524 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19418) );
  INV_X1 U20525 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20267) );
  AOI22_X1 U20526 ( .A1(n17245), .A2(n19418), .B1(n20267), .B2(n17246), .ZN(
        U363) );
  INV_X1 U20527 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19416) );
  INV_X1 U20528 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20265) );
  AOI22_X1 U20529 ( .A1(n17245), .A2(n19416), .B1(n20265), .B2(n17246), .ZN(
        U364) );
  INV_X1 U20530 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19378) );
  INV_X1 U20531 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n21345) );
  AOI22_X1 U20532 ( .A1(n17245), .A2(n19378), .B1(n21345), .B2(n17246), .ZN(
        U365) );
  INV_X1 U20533 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19414) );
  INV_X1 U20534 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20263) );
  AOI22_X1 U20535 ( .A1(n17245), .A2(n19414), .B1(n20263), .B2(n17246), .ZN(
        U366) );
  INV_X1 U20536 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19413) );
  INV_X1 U20537 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20261) );
  AOI22_X1 U20538 ( .A1(n17245), .A2(n19413), .B1(n20261), .B2(n17246), .ZN(
        U367) );
  INV_X1 U20539 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19411) );
  INV_X1 U20540 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20259) );
  AOI22_X1 U20541 ( .A1(n17245), .A2(n19411), .B1(n20259), .B2(n17246), .ZN(
        U368) );
  INV_X1 U20542 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19409) );
  INV_X1 U20543 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20258) );
  AOI22_X1 U20544 ( .A1(n17245), .A2(n19409), .B1(n20258), .B2(n17246), .ZN(
        U369) );
  INV_X1 U20545 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19407) );
  INV_X1 U20546 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20256) );
  AOI22_X1 U20547 ( .A1(n17245), .A2(n19407), .B1(n20256), .B2(n17246), .ZN(
        U370) );
  INV_X1 U20548 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19405) );
  INV_X1 U20549 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U20550 ( .A1(n17245), .A2(n19405), .B1(n20255), .B2(n17246), .ZN(
        U371) );
  INV_X1 U20551 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19403) );
  INV_X1 U20552 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20253) );
  AOI22_X1 U20553 ( .A1(n17245), .A2(n19403), .B1(n20253), .B2(n17246), .ZN(
        U372) );
  INV_X1 U20554 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19401) );
  INV_X1 U20555 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20252) );
  AOI22_X1 U20556 ( .A1(n17245), .A2(n19401), .B1(n20252), .B2(n17246), .ZN(
        U373) );
  INV_X1 U20557 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19399) );
  INV_X1 U20558 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20251) );
  AOI22_X1 U20559 ( .A1(n17245), .A2(n19399), .B1(n20251), .B2(n17246), .ZN(
        U374) );
  INV_X1 U20560 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19397) );
  INV_X1 U20561 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20249) );
  AOI22_X1 U20562 ( .A1(n17245), .A2(n19397), .B1(n20249), .B2(n17246), .ZN(
        U375) );
  INV_X1 U20563 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19376) );
  INV_X1 U20564 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20233) );
  AOI22_X1 U20565 ( .A1(n17245), .A2(n19376), .B1(n20233), .B2(n17246), .ZN(
        U376) );
  INV_X1 U20566 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17247) );
  INV_X1 U20567 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19375) );
  NAND2_X1 U20568 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19375), .ZN(n19364) );
  AOI22_X1 U20569 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19364), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19373), .ZN(n19446) );
  OAI21_X1 U20570 ( .B1(n19373), .B2(n17247), .A(n19443), .ZN(P3_U2633) );
  AOI21_X1 U20571 ( .B1(n17249), .B2(n18189), .A(n17248), .ZN(n17256) );
  INV_X1 U20572 ( .A(n17256), .ZN(n17250) );
  OAI21_X1 U20573 ( .B1(n19337), .B2(n17250), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17251) );
  OAI21_X1 U20574 ( .B1(n17252), .B2(n19349), .A(n17251), .ZN(P3_U2634) );
  AOI21_X1 U20575 ( .B1(n19373), .B2(n19375), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17253) );
  AOI22_X1 U20576 ( .A1(n19434), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17253), 
        .B2(n19482), .ZN(P3_U2635) );
  OAI21_X1 U20577 ( .B1(n19361), .B2(BS16), .A(n19446), .ZN(n19444) );
  OAI21_X1 U20578 ( .B1(n19446), .B2(n17254), .A(n19444), .ZN(P3_U2636) );
  AND2_X1 U20579 ( .A1(n17256), .A2(n17255), .ZN(n19333) );
  NOR2_X1 U20580 ( .A1(n19333), .A2(n19337), .ZN(n19462) );
  OAI21_X1 U20581 ( .B1(n19462), .B2(n17258), .A(n17257), .ZN(P3_U2637) );
  NOR4_X1 U20582 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17262) );
  NOR4_X1 U20583 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17261) );
  NOR4_X1 U20584 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17260) );
  NOR4_X1 U20585 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17259) );
  NAND4_X1 U20586 ( .A1(n17262), .A2(n17261), .A3(n17260), .A4(n17259), .ZN(
        n17268) );
  NOR4_X1 U20587 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17266) );
  AOI211_X1 U20588 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_24__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17265) );
  NOR4_X1 U20589 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17264) );
  NOR4_X1 U20590 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17263) );
  NAND4_X1 U20591 ( .A1(n17266), .A2(n17265), .A3(n17264), .A4(n17263), .ZN(
        n17267) );
  NOR2_X1 U20592 ( .A1(n17268), .A2(n17267), .ZN(n19454) );
  INV_X1 U20593 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19439) );
  NOR3_X1 U20594 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17270) );
  OAI21_X1 U20595 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17270), .A(n19454), .ZN(
        n17269) );
  OAI21_X1 U20596 ( .B1(n19454), .B2(n19439), .A(n17269), .ZN(P3_U2638) );
  NAND2_X1 U20597 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n19454), .ZN(n19456) );
  NOR2_X1 U20598 ( .A1(n17270), .A2(n19456), .ZN(n17272) );
  NOR2_X1 U20599 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n19454), .ZN(n17271)
         );
  AOI211_X1 U20600 ( .C1(n19454), .C2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n17272), 
        .B(n17271), .ZN(P3_U2639) );
  INV_X1 U20601 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17617) );
  NOR3_X1 U20602 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19436), .A3(n17273), 
        .ZN(n17276) );
  INV_X1 U20603 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n17274) );
  OAI22_X1 U20604 ( .A1(n10147), .A2(n17595), .B1(n17274), .B2(n17598), .ZN(
        n17275) );
  AOI211_X1 U20605 ( .C1(n17277), .C2(n17617), .A(n17276), .B(n17275), .ZN(
        n17284) );
  INV_X1 U20606 ( .A(n17278), .ZN(n17287) );
  OAI21_X1 U20607 ( .B1(n17279), .B2(n17287), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n17283) );
  NOR2_X1 U20608 ( .A1(n17519), .A2(n19355), .ZN(n17594) );
  NAND3_X1 U20609 ( .A1(n17594), .A2(n17281), .A3(n17280), .ZN(n17282) );
  NAND3_X1 U20610 ( .A1(n17284), .A2(n17283), .A3(n17282), .ZN(P3_U2640) );
  NOR2_X1 U20611 ( .A1(n17296), .A2(n17650), .ZN(n17295) );
  OAI22_X1 U20612 ( .A1(n17285), .A2(n17595), .B1(n17598), .B2(n17650), .ZN(
        n17286) );
  AOI221_X1 U20613 ( .B1(n17288), .B2(n19431), .C1(n17287), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n17286), .ZN(n17293) );
  OAI211_X1 U20614 ( .C1(n17291), .C2(n17290), .A(n17558), .B(n17289), .ZN(
        n17292) );
  OAI211_X1 U20615 ( .C1(n17295), .C2(n17294), .A(n17293), .B(n17292), .ZN(
        P3_U2642) );
  AOI22_X1 U20616 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17525), .B1(
        n17518), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17305) );
  NOR2_X1 U20617 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17301), .ZN(n17307) );
  AOI211_X1 U20618 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17308), .A(n17296), .B(
        n17605), .ZN(n17297) );
  AOI221_X1 U20619 ( .B1(n17318), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n17307), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n17297), .ZN(n17304) );
  OAI211_X1 U20620 ( .C1(n17300), .C2(n17298), .A(n17558), .B(n17299), .ZN(
        n17303) );
  OR3_X1 U20621 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17301), .A3(n19427), .ZN(
        n17302) );
  NAND4_X1 U20622 ( .A1(n17305), .A2(n17304), .A3(n17303), .A4(n17302), .ZN(
        P3_U2643) );
  OAI22_X1 U20623 ( .A1(n11625), .A2(n17595), .B1(n17598), .B2(n17309), .ZN(
        n17306) );
  AOI211_X1 U20624 ( .C1(n17318), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17307), 
        .B(n17306), .ZN(n17315) );
  OAI211_X1 U20625 ( .C1(n17316), .C2(n17309), .A(n17584), .B(n17308), .ZN(
        n17314) );
  OAI211_X1 U20626 ( .C1(n17312), .C2(n17310), .A(n17558), .B(n17311), .ZN(
        n17313) );
  NAND3_X1 U20627 ( .A1(n17315), .A2(n17314), .A3(n17313), .ZN(P3_U2644) );
  AOI22_X1 U20628 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17525), .B1(
        n17518), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17325) );
  AOI211_X1 U20629 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17329), .A(n17316), .B(
        n17605), .ZN(n17317) );
  AOI21_X1 U20630 ( .B1(n17318), .B2(P3_REIP_REG_26__SCAN_IN), .A(n17317), 
        .ZN(n17324) );
  OAI211_X1 U20631 ( .C1(n17321), .C2(n17320), .A(n17558), .B(n17319), .ZN(
        n17323) );
  NAND3_X1 U20632 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17328), .A3(n19426), 
        .ZN(n17322) );
  NAND4_X1 U20633 ( .A1(n17325), .A2(n17324), .A3(n17323), .A4(n17322), .ZN(
        P3_U2645) );
  OAI21_X1 U20634 ( .B1(n17593), .B2(n17337), .A(n17450), .ZN(n17345) );
  OAI21_X1 U20635 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17599), .A(n17345), 
        .ZN(n17327) );
  INV_X1 U20636 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18245) );
  OAI22_X1 U20637 ( .A1(n18245), .A2(n17595), .B1(n17598), .B2(n17610), .ZN(
        n17326) );
  AOI221_X1 U20638 ( .B1(n17328), .B2(n21348), .C1(n17327), .C2(
        P3_REIP_REG_25__SCAN_IN), .A(n17326), .ZN(n17334) );
  OAI211_X1 U20639 ( .C1(n17335), .C2(n17610), .A(n17584), .B(n17329), .ZN(
        n17333) );
  OAI211_X1 U20640 ( .C1(n18244), .C2(n17330), .A(n17558), .B(n17331), .ZN(
        n17332) );
  NAND3_X1 U20641 ( .A1(n17334), .A2(n17333), .A3(n17332), .ZN(P3_U2646) );
  AOI211_X1 U20642 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17350), .A(n17335), .B(
        n17605), .ZN(n17339) );
  NAND2_X1 U20643 ( .A1(n17581), .A2(n19423), .ZN(n17336) );
  OAI22_X1 U20644 ( .A1(n18243), .A2(n17595), .B1(n17337), .B2(n17336), .ZN(
        n17338) );
  AOI211_X1 U20645 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17518), .A(n17339), .B(
        n17338), .ZN(n17344) );
  OAI211_X1 U20646 ( .C1(n17342), .C2(n17340), .A(n17558), .B(n17341), .ZN(
        n17343) );
  OAI211_X1 U20647 ( .C1(n17345), .C2(n19423), .A(n17344), .B(n17343), .ZN(
        P3_U2647) );
  INV_X1 U20648 ( .A(n17345), .ZN(n17349) );
  NOR3_X1 U20649 ( .A1(n17599), .A2(n17360), .A3(n17361), .ZN(n17348) );
  OAI22_X1 U20650 ( .A1(n17346), .A2(n17595), .B1(n17598), .B2(n17607), .ZN(
        n17347) );
  AOI221_X1 U20651 ( .B1(n17349), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n17348), 
        .C2(n19419), .A(n17347), .ZN(n17354) );
  OAI211_X1 U20652 ( .C1(n17356), .C2(n17607), .A(n17584), .B(n17350), .ZN(
        n17353) );
  NAND3_X1 U20653 ( .A1(n17354), .A2(n17353), .A3(n17352), .ZN(P3_U2648) );
  AOI22_X1 U20654 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17525), .B1(
        n17518), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n17365) );
  AOI21_X1 U20655 ( .B1(n17360), .B2(n17581), .A(n17593), .ZN(n17355) );
  INV_X1 U20656 ( .A(n17355), .ZN(n17378) );
  AOI211_X1 U20657 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17368), .A(n17356), .B(
        n17605), .ZN(n17357) );
  AOI21_X1 U20658 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n17378), .A(n17357), 
        .ZN(n17364) );
  OAI211_X1 U20659 ( .C1(n18281), .C2(n17358), .A(n17558), .B(n17359), .ZN(
        n17363) );
  NOR2_X1 U20660 ( .A1(n17599), .A2(n17360), .ZN(n17367) );
  OAI211_X1 U20661 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(P3_REIP_REG_22__SCAN_IN), .A(n17367), .B(n17361), .ZN(n17362) );
  NAND4_X1 U20662 ( .A1(n17365), .A2(n17364), .A3(n17363), .A4(n17362), .ZN(
        P3_U2649) );
  INV_X1 U20663 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21391) );
  OAI22_X1 U20664 ( .A1(n18292), .A2(n17595), .B1(n17598), .B2(n17717), .ZN(
        n17366) );
  AOI221_X1 U20665 ( .B1(n17378), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17367), 
        .C2(n21391), .A(n17366), .ZN(n17373) );
  OAI211_X1 U20666 ( .C1(n17374), .C2(n17717), .A(n17584), .B(n17368), .ZN(
        n17372) );
  OAI211_X1 U20667 ( .C1(n18289), .C2(n17369), .A(n17558), .B(n17370), .ZN(
        n17371) );
  NAND3_X1 U20668 ( .A1(n17373), .A2(n17372), .A3(n17371), .ZN(P3_U2650) );
  NAND4_X1 U20669 ( .A1(n17581), .A2(P3_REIP_REG_19__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .A4(n17406), .ZN(n17383) );
  AOI211_X1 U20670 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17387), .A(n17374), .B(
        n17605), .ZN(n17377) );
  INV_X1 U20671 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18303) );
  OAI22_X1 U20672 ( .A1(n18303), .A2(n17595), .B1(n17598), .B2(n17375), .ZN(
        n17376) );
  AOI211_X1 U20673 ( .C1(n17378), .C2(P3_REIP_REG_20__SCAN_IN), .A(n17377), 
        .B(n17376), .ZN(n17382) );
  OAI211_X1 U20674 ( .C1(n18305), .C2(n17380), .A(n17558), .B(n17379), .ZN(
        n17381) );
  OAI211_X1 U20675 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n17383), .A(n17382), 
        .B(n17381), .ZN(P3_U2651) );
  NOR2_X1 U20676 ( .A1(n17397), .A2(n17384), .ZN(n17385) );
  OAI22_X1 U20677 ( .A1(n17605), .A2(n17385), .B1(n17598), .B2(n17384), .ZN(
        n17386) );
  AOI22_X1 U20678 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17525), .B1(
        n17387), .B2(n17386), .ZN(n17395) );
  INV_X1 U20680 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19410) );
  NAND2_X1 U20681 ( .A1(n17581), .A2(n17406), .ZN(n17388) );
  NOR2_X1 U20682 ( .A1(n19410), .A2(n17388), .ZN(n17389) );
  INV_X1 U20683 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19412) );
  NOR2_X1 U20684 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17388), .ZN(n17398) );
  OAI21_X1 U20685 ( .B1(n17406), .B2(n17599), .A(n17573), .ZN(n17396) );
  OAI33_X1 U20686 ( .A1(1'b0), .A2(n17389), .A3(P3_REIP_REG_19__SCAN_IN), .B1(
        n19412), .B2(n17398), .B3(n17396), .ZN(n17394) );
  OAI211_X1 U20687 ( .C1(n18320), .C2(n17391), .A(n17558), .B(n17392), .ZN(
        n17393) );
  NAND4_X1 U20688 ( .A1(n17395), .A2(n17394), .A3(n18748), .A4(n17393), .ZN(
        P3_U2652) );
  INV_X1 U20689 ( .A(n17396), .ZN(n17419) );
  AOI211_X1 U20690 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17412), .A(n17397), .B(
        n17605), .ZN(n17401) );
  INV_X1 U20691 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17774) );
  INV_X1 U20692 ( .A(n17398), .ZN(n17399) );
  OAI211_X1 U20693 ( .C1(n17598), .C2(n17774), .A(n18748), .B(n17399), .ZN(
        n17400) );
  AOI211_X1 U20694 ( .C1(n17525), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17401), .B(n17400), .ZN(n17405) );
  OAI211_X1 U20695 ( .C1(n18325), .C2(n17402), .A(n17558), .B(n17403), .ZN(
        n17404) );
  OAI211_X1 U20696 ( .C1(n17419), .C2(n19410), .A(n17405), .B(n17404), .ZN(
        P3_U2653) );
  OR2_X1 U20697 ( .A1(n17599), .A2(n17406), .ZN(n17407) );
  OAI22_X1 U20698 ( .A1(n18339), .A2(n17595), .B1(n17408), .B2(n17407), .ZN(
        n17417) );
  OAI211_X1 U20699 ( .C1(n17411), .C2(n17410), .A(n17558), .B(n17409), .ZN(
        n17414) );
  OAI211_X1 U20700 ( .C1(n17420), .C2(n17415), .A(n17584), .B(n17412), .ZN(
        n17413) );
  OAI211_X1 U20701 ( .C1(n17415), .C2(n17598), .A(n17414), .B(n17413), .ZN(
        n17416) );
  NOR3_X1 U20702 ( .A1(n18846), .A2(n17417), .A3(n17416), .ZN(n17418) );
  OAI21_X1 U20703 ( .B1(n17419), .B2(n19408), .A(n17418), .ZN(P3_U2654) );
  INV_X1 U20704 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19404) );
  NAND2_X1 U20705 ( .A1(n17428), .A2(n17573), .ZN(n17449) );
  OAI21_X1 U20706 ( .B1(n19404), .B2(n17449), .A(n17450), .ZN(n17434) );
  INV_X1 U20707 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19406) );
  AOI211_X1 U20708 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17436), .A(n17420), .B(
        n17605), .ZN(n17423) );
  INV_X1 U20709 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18355) );
  NAND4_X1 U20710 ( .A1(n17581), .A2(P3_REIP_REG_15__SCAN_IN), .A3(n17428), 
        .A4(n19406), .ZN(n17421) );
  OAI211_X1 U20711 ( .C1(n18355), .C2(n17595), .A(n18748), .B(n17421), .ZN(
        n17422) );
  AOI211_X1 U20712 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17518), .A(n17423), .B(
        n17422), .ZN(n17427) );
  OAI211_X1 U20713 ( .C1(n18353), .C2(n17424), .A(n17558), .B(n17425), .ZN(
        n17426) );
  OAI211_X1 U20714 ( .C1(n17434), .C2(n19406), .A(n17427), .B(n17426), .ZN(
        P3_U2655) );
  AOI21_X1 U20715 ( .B1(n17581), .B2(n17428), .A(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17433) );
  AOI21_X1 U20716 ( .B1(n18363), .B2(n18354), .A(n17429), .ZN(n18366) );
  NAND2_X1 U20717 ( .A1(n17508), .A2(n17430), .ZN(n17431) );
  XOR2_X1 U20718 ( .A(n18366), .B(n17431), .Z(n17432) );
  OAI22_X1 U20719 ( .A1(n17434), .A2(n17433), .B1(n19355), .B2(n17432), .ZN(
        n17435) );
  AOI211_X1 U20720 ( .C1(n17518), .C2(P3_EBX_REG_15__SCAN_IN), .A(n18846), .B(
        n17435), .ZN(n17439) );
  OAI211_X1 U20721 ( .C1(n17446), .C2(n17437), .A(n17584), .B(n17436), .ZN(
        n17438) );
  OAI211_X1 U20722 ( .C1(n17595), .C2(n18363), .A(n17439), .B(n17438), .ZN(
        P3_U2656) );
  OR2_X1 U20723 ( .A1(n17599), .A2(n17440), .ZN(n17465) );
  NOR2_X1 U20724 ( .A1(n19400), .A2(n17465), .ZN(n17441) );
  AOI22_X1 U20725 ( .A1(n17518), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n17441), 
        .B2(n17449), .ZN(n17453) );
  AOI21_X1 U20726 ( .B1(n18379), .B2(n17454), .A(n17442), .ZN(n18381) );
  INV_X1 U20727 ( .A(n18380), .ZN(n17443) );
  AOI21_X1 U20728 ( .B1(n17443), .B2(n17579), .A(n17519), .ZN(n17462) );
  INV_X1 U20729 ( .A(n18381), .ZN(n17445) );
  INV_X1 U20730 ( .A(n17462), .ZN(n17444) );
  AOI221_X1 U20731 ( .B1(n18381), .B2(n17462), .C1(n17445), .C2(n17444), .A(
        n19355), .ZN(n17448) );
  AOI211_X1 U20732 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17456), .A(n17446), .B(
        n17605), .ZN(n17447) );
  AOI211_X1 U20733 ( .C1(n17525), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17448), .B(n17447), .ZN(n17452) );
  NAND3_X1 U20734 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17450), .A3(n17449), 
        .ZN(n17451) );
  NAND4_X1 U20735 ( .A1(n17453), .A2(n17452), .A3(n18748), .A4(n17451), .ZN(
        P3_U2657) );
  OAI21_X1 U20736 ( .B1(n17469), .B2(n17599), .A(n17573), .ZN(n17487) );
  NOR2_X1 U20737 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17599), .ZN(n17468) );
  AOI22_X1 U20738 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17525), .B1(
        n17518), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20739 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17470), .A(
        n17454), .ZN(n18401) );
  INV_X1 U20740 ( .A(n18401), .ZN(n17455) );
  AOI21_X1 U20741 ( .B1(n17508), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19355), .ZN(n17601) );
  OAI211_X1 U20742 ( .C1(n17470), .C2(n17519), .A(n17455), .B(n17601), .ZN(
        n17459) );
  OAI211_X1 U20743 ( .C1(n17466), .C2(n17457), .A(n17584), .B(n17456), .ZN(
        n17458) );
  NAND4_X1 U20744 ( .A1(n17460), .A2(n18748), .A3(n17459), .A4(n17458), .ZN(
        n17461) );
  AOI221_X1 U20745 ( .B1(n17487), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17468), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17461), .ZN(n17464) );
  NAND3_X1 U20746 ( .A1(n17558), .A2(n17462), .A3(n18401), .ZN(n17463) );
  OAI211_X1 U20747 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17465), .A(n17464), 
        .B(n17463), .ZN(P3_U2658) );
  AOI211_X1 U20748 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17481), .A(n17466), .B(
        n17605), .ZN(n17467) );
  AOI21_X1 U20749 ( .B1(n17525), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17467), .ZN(n17476) );
  AOI22_X1 U20750 ( .A1(n17518), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n17469), 
        .B2(n17468), .ZN(n17475) );
  AOI21_X1 U20751 ( .B1(n18400), .B2(n18395), .A(n17470), .ZN(n18416) );
  AOI21_X1 U20752 ( .B1(n17471), .B2(n17579), .A(n17519), .ZN(n17472) );
  XOR2_X1 U20753 ( .A(n18416), .B(n17472), .Z(n17473) );
  AOI22_X1 U20754 ( .A1(n17558), .A2(n17473), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n17487), .ZN(n17474) );
  NAND4_X1 U20755 ( .A1(n17476), .A2(n17475), .A3(n17474), .A4(n18748), .ZN(
        P3_U2659) );
  NOR2_X1 U20756 ( .A1(n17599), .A2(n17492), .ZN(n17537) );
  INV_X1 U20757 ( .A(n17537), .ZN(n17545) );
  OAI21_X1 U20758 ( .B1(n17477), .B2(n17545), .A(n19396), .ZN(n17486) );
  NAND2_X1 U20759 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17503), .ZN(
        n17502) );
  NOR2_X1 U20760 ( .A1(n17478), .A2(n17502), .ZN(n17494) );
  OAI21_X1 U20761 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17494), .A(
        n18395), .ZN(n18431) );
  NAND2_X1 U20762 ( .A1(n17597), .A2(n17543), .ZN(n17544) );
  OAI21_X1 U20763 ( .B1(n18429), .B2(n17544), .A(n17508), .ZN(n17480) );
  AOI21_X1 U20764 ( .B1(n18431), .B2(n17480), .A(n19355), .ZN(n17479) );
  OAI21_X1 U20765 ( .B1(n18431), .B2(n17480), .A(n17479), .ZN(n17483) );
  OAI211_X1 U20766 ( .C1(n17490), .C2(n17489), .A(n17584), .B(n17481), .ZN(
        n17482) );
  OAI211_X1 U20767 ( .C1(n17595), .C2(n17484), .A(n17483), .B(n17482), .ZN(
        n17485) );
  AOI21_X1 U20768 ( .B1(n17487), .B2(n17486), .A(n17485), .ZN(n17488) );
  OAI211_X1 U20769 ( .C1(n17598), .C2(n17489), .A(n17488), .B(n18748), .ZN(
        P3_U2660) );
  AOI211_X1 U20770 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17509), .A(n17490), .B(
        n17605), .ZN(n17491) );
  AOI211_X1 U20771 ( .C1(n17518), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18846), .B(
        n17491), .ZN(n17500) );
  AOI21_X1 U20772 ( .B1(n17581), .B2(n17492), .A(n17593), .ZN(n17555) );
  OAI21_X1 U20773 ( .B1(n17496), .B2(n17493), .A(n17555), .ZN(n17501) );
  AOI21_X1 U20774 ( .B1(n17478), .B2(n17502), .A(n17494), .ZN(n18447) );
  AND2_X1 U20775 ( .A1(n17597), .A2(n17503), .ZN(n17505) );
  AOI21_X1 U20776 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17505), .A(
        n17519), .ZN(n17506) );
  OAI21_X1 U20777 ( .B1(n18447), .B2(n17506), .A(n17558), .ZN(n17495) );
  AOI21_X1 U20778 ( .B1(n18447), .B2(n17506), .A(n17495), .ZN(n17498) );
  INV_X1 U20779 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19394) );
  INV_X1 U20780 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19392) );
  NAND2_X1 U20781 ( .A1(n17496), .A2(n17537), .ZN(n17512) );
  AOI221_X1 U20782 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n19394), .C2(n19392), .A(n17512), .ZN(n17497) );
  AOI211_X1 U20783 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n17501), .A(n17498), 
        .B(n17497), .ZN(n17499) );
  OAI211_X1 U20784 ( .C1(n17478), .C2(n17595), .A(n17500), .B(n17499), .ZN(
        P3_U2661) );
  INV_X1 U20785 ( .A(n17501), .ZN(n17528) );
  OAI21_X1 U20786 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17503), .A(
        n17502), .ZN(n18459) );
  AOI22_X1 U20787 ( .A1(n17506), .A2(n18459), .B1(n17505), .B2(n17504), .ZN(
        n17507) );
  OAI21_X1 U20788 ( .B1(n17508), .B2(n18459), .A(n17507), .ZN(n17514) );
  AOI22_X1 U20789 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17525), .B1(
        n17518), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n17511) );
  OAI211_X1 U20790 ( .C1(n17522), .C2(n17928), .A(n17584), .B(n17509), .ZN(
        n17510) );
  OAI211_X1 U20791 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n17512), .A(n17511), .B(
        n17510), .ZN(n17513) );
  AOI211_X1 U20792 ( .C1(n17558), .C2(n17514), .A(n18846), .B(n17513), .ZN(
        n17515) );
  OAI21_X1 U20793 ( .B1(n17528), .B2(n19392), .A(n17515), .ZN(P3_U2662) );
  NOR3_X1 U20794 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17516), .A3(n17545), .ZN(
        n17517) );
  AOI211_X1 U20795 ( .C1(n17518), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18846), .B(
        n17517), .ZN(n17527) );
  INV_X1 U20796 ( .A(n17544), .ZN(n17531) );
  AOI21_X1 U20797 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17531), .A(
        n17519), .ZN(n17530) );
  OAI21_X1 U20798 ( .B1(n17521), .B2(n17530), .A(n17558), .ZN(n17520) );
  AOI21_X1 U20799 ( .B1(n17521), .B2(n17530), .A(n17520), .ZN(n17524) );
  AOI211_X1 U20800 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17538), .A(n17522), .B(
        n17605), .ZN(n17523) );
  AOI211_X1 U20801 ( .C1(n17525), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17524), .B(n17523), .ZN(n17526) );
  OAI211_X1 U20802 ( .C1(n17528), .C2(n19391), .A(n17527), .B(n17526), .ZN(
        P3_U2663) );
  OAI21_X1 U20803 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17545), .A(n17555), .ZN(
        n17536) );
  OAI21_X1 U20804 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17543), .A(
        n17529), .ZN(n18477) );
  INV_X1 U20805 ( .A(n17530), .ZN(n17533) );
  OAI21_X1 U20806 ( .B1(n17531), .B2(n18477), .A(n17558), .ZN(n17532) );
  AOI22_X1 U20807 ( .A1(n18477), .A2(n17533), .B1(n17572), .B2(n17532), .ZN(
        n17535) );
  OAI22_X1 U20808 ( .A1(n18465), .A2(n17595), .B1(n17598), .B2(n17962), .ZN(
        n17534) );
  AOI211_X1 U20809 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n17536), .A(n17535), .B(
        n17534), .ZN(n17541) );
  INV_X1 U20810 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19388) );
  NAND3_X1 U20811 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17537), .A3(n19388), 
        .ZN(n17540) );
  OAI211_X1 U20812 ( .C1(n17542), .C2(n17962), .A(n17584), .B(n17538), .ZN(
        n17539) );
  NAND4_X1 U20813 ( .A1(n17541), .A2(n18748), .A3(n17540), .A4(n17539), .ZN(
        P3_U2664) );
  INV_X1 U20814 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19386) );
  AOI211_X1 U20815 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17561), .A(n17542), .B(
        n17605), .ZN(n17550) );
  AOI21_X1 U20816 ( .B1(n18494), .B2(n17551), .A(n17543), .ZN(n18491) );
  NAND2_X1 U20817 ( .A1(n17594), .A2(n17544), .ZN(n17546) );
  OAI22_X1 U20818 ( .A1(n18491), .A2(n17546), .B1(P3_REIP_REG_6__SCAN_IN), 
        .B2(n17545), .ZN(n17549) );
  INV_X1 U20819 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17547) );
  OAI22_X1 U20820 ( .A1(n18494), .A2(n17595), .B1(n17598), .B2(n17547), .ZN(
        n17548) );
  NOR4_X1 U20821 ( .A1(n18846), .A2(n17550), .A3(n17549), .A4(n17548), .ZN(
        n17554) );
  INV_X1 U20822 ( .A(n17551), .ZN(n17556) );
  INV_X1 U20823 ( .A(n17572), .ZN(n17552) );
  OAI211_X1 U20824 ( .C1(n17556), .C2(n17552), .A(n18491), .B(n17601), .ZN(
        n17553) );
  OAI211_X1 U20825 ( .C1(n17555), .C2(n19386), .A(n17554), .B(n17553), .ZN(
        P3_U2665) );
  INV_X1 U20826 ( .A(n17555), .ZN(n17567) );
  AOI21_X1 U20827 ( .B1(n18495), .B2(n17557), .A(n17556), .ZN(n18503) );
  OAI21_X1 U20828 ( .B1(n18503), .B2(n17560), .A(n17558), .ZN(n17559) );
  AOI21_X1 U20829 ( .B1(n18503), .B2(n17560), .A(n17559), .ZN(n17566) );
  OAI211_X1 U20830 ( .C1(n17562), .C2(n17564), .A(n17584), .B(n17561), .ZN(
        n17563) );
  OAI211_X1 U20831 ( .C1(n17598), .C2(n17564), .A(n18748), .B(n17563), .ZN(
        n17565) );
  AOI211_X1 U20832 ( .C1(n17567), .C2(P3_REIP_REG_5__SCAN_IN), .A(n17566), .B(
        n17565), .ZN(n17570) );
  INV_X1 U20833 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19385) );
  NAND3_X1 U20834 ( .A1(n17581), .A2(n17568), .A3(n19385), .ZN(n17569) );
  OAI211_X1 U20835 ( .C1(n17595), .C2(n18495), .A(n17570), .B(n17569), .ZN(
        P3_U2666) );
  OAI22_X1 U20836 ( .A1(n18548), .A2(n17595), .B1(n17598), .B2(n17585), .ZN(
        n17575) );
  INV_X1 U20837 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19377) );
  OAI21_X1 U20838 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17571), .ZN(n18543) );
  OAI22_X1 U20839 ( .A1(n19377), .A2(n17573), .B1(n18543), .B2(n17572), .ZN(
        n17574) );
  AOI211_X1 U20840 ( .C1(n17576), .C2(n19489), .A(n17575), .B(n17574), .ZN(
        n17590) );
  NAND2_X1 U20841 ( .A1(n17577), .A2(n17597), .ZN(n17578) );
  OAI211_X1 U20842 ( .C1(n17579), .C2(n18543), .A(n17594), .B(n17578), .ZN(
        n17589) );
  OAI211_X1 U20843 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17581), .B(n17580), .ZN(n17588) );
  NOR2_X1 U20844 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17586) );
  INV_X1 U20845 ( .A(n17582), .ZN(n17583) );
  OAI211_X1 U20846 ( .C1(n17586), .C2(n17585), .A(n17584), .B(n17583), .ZN(
        n17587) );
  NAND4_X1 U20847 ( .A1(n17590), .A2(n17589), .A3(n17588), .A4(n17587), .ZN(
        P3_U2669) );
  OAI21_X1 U20848 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17976), .ZN(n17983) );
  INV_X1 U20849 ( .A(n17591), .ZN(n17592) );
  AOI22_X1 U20850 ( .A1(n17593), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n19489), 
        .B2(n17592), .ZN(n17604) );
  INV_X1 U20851 ( .A(n17594), .ZN(n17596) );
  OAI21_X1 U20852 ( .B1(n17597), .B2(n17596), .A(n17595), .ZN(n17602) );
  INV_X1 U20853 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17982) );
  OAI22_X1 U20854 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17599), .B1(n17598), 
        .B2(n17982), .ZN(n17600) );
  AOI221_X1 U20855 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17602), .C1(
        n18561), .C2(n17601), .A(n17600), .ZN(n17603) );
  OAI211_X1 U20856 ( .C1(n17605), .C2(n17983), .A(n17604), .B(n17603), .ZN(
        P3_U2670) );
  NOR4_X1 U20857 ( .A1(n17608), .A2(n17607), .A3(n17606), .A4(n17717), .ZN(
        n17613) );
  INV_X1 U20858 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17611) );
  NAND2_X1 U20859 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17609) );
  NOR4_X1 U20860 ( .A1(n17650), .A2(n17611), .A3(n17610), .A4(n17609), .ZN(
        n17612) );
  NAND4_X1 U20861 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17756), .A3(n17613), 
        .A4(n17612), .ZN(n17616) );
  NOR2_X1 U20862 ( .A1(n17617), .A2(n17616), .ZN(n17646) );
  NAND2_X1 U20863 ( .A1(n17980), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17615) );
  NAND2_X1 U20864 ( .A1(n17646), .A2(n18910), .ZN(n17614) );
  OAI22_X1 U20865 ( .A1(n17646), .A2(n17615), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17614), .ZN(P3_U2672) );
  NAND2_X1 U20866 ( .A1(n17617), .A2(n17616), .ZN(n17618) );
  NAND2_X1 U20867 ( .A1(n17618), .A2(n17980), .ZN(n17645) );
  AOI22_X1 U20868 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U20869 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U20870 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n9608), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U20871 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17619) );
  NAND4_X1 U20872 ( .A1(n17622), .A2(n17621), .A3(n17620), .A4(n17619), .ZN(
        n17631) );
  OAI22_X1 U20873 ( .A1(n17891), .A2(n17816), .B1(n17939), .B2(n17623), .ZN(
        n17626) );
  INV_X1 U20874 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17624) );
  OAI22_X1 U20875 ( .A1(n11436), .A2(n17624), .B1(n17918), .B2(n17815), .ZN(
        n17625) );
  AOI211_X1 U20876 ( .C1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .C2(n17872), .A(
        n17626), .B(n17625), .ZN(n17628) );
  AOI22_X1 U20877 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n17933), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17627) );
  OAI211_X1 U20878 ( .C1(n17950), .C2(n17629), .A(n17628), .B(n17627), .ZN(
        n17630) );
  NOR2_X1 U20879 ( .A1(n17631), .A2(n17630), .ZN(n17644) );
  INV_X1 U20880 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17633) );
  INV_X1 U20881 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17632) );
  OAI22_X1 U20882 ( .A1(n17941), .A2(n17633), .B1(n17939), .B2(n17632), .ZN(
        n17635) );
  INV_X1 U20883 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17685) );
  INV_X1 U20884 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17830) );
  OAI22_X1 U20885 ( .A1(n17747), .A2(n17685), .B1(n17799), .B2(n17830), .ZN(
        n17634) );
  AOI211_X1 U20886 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17635), .B(n17634), .ZN(n17643) );
  AOI22_X1 U20887 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17639) );
  AOI22_X1 U20888 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U20889 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17637) );
  AOI22_X1 U20890 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17636) );
  AND4_X1 U20891 ( .A1(n17639), .A2(n17638), .A3(n17637), .A4(n17636), .ZN(
        n17642) );
  AOI22_X1 U20892 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17641) );
  NAND2_X1 U20893 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n17640) );
  NAND4_X1 U20894 ( .A1(n17643), .A2(n17642), .A3(n17641), .A4(n17640), .ZN(
        n17648) );
  NAND2_X1 U20895 ( .A1(n17649), .A2(n17648), .ZN(n17647) );
  XNOR2_X1 U20896 ( .A(n17644), .B(n17647), .ZN(n17997) );
  OAI22_X1 U20897 ( .A1(n17646), .A2(n17645), .B1(n17997), .B2(n17980), .ZN(
        P3_U2673) );
  OAI21_X1 U20898 ( .B1(n17649), .B2(n17648), .A(n17647), .ZN(n18001) );
  AOI22_X1 U20899 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17652), .B1(n17651), 
        .B2(n17650), .ZN(n17653) );
  OAI21_X1 U20900 ( .B1(n18001), .B2(n17980), .A(n17653), .ZN(P3_U2674) );
  OAI21_X1 U20901 ( .B1(n17658), .B2(n17655), .A(n17654), .ZN(n18009) );
  NAND3_X1 U20902 ( .A1(n17657), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17980), 
        .ZN(n17656) );
  OAI221_X1 U20903 ( .B1(n17657), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17980), 
        .C2(n18009), .A(n17656), .ZN(P3_U2676) );
  AOI21_X1 U20904 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17980), .A(n17666), .ZN(
        n17661) );
  AOI21_X1 U20905 ( .B1(n17659), .B2(n17663), .A(n17658), .ZN(n18010) );
  INV_X1 U20906 ( .A(n18010), .ZN(n17660) );
  OAI22_X1 U20907 ( .A1(n17662), .A2(n17661), .B1(n17660), .B2(n17980), .ZN(
        P3_U2677) );
  AOI21_X1 U20908 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17980), .A(n17672), .ZN(
        n17665) );
  OAI21_X1 U20909 ( .B1(n17668), .B2(n17664), .A(n17663), .ZN(n18020) );
  OAI22_X1 U20910 ( .A1(n17666), .A2(n17665), .B1(n18020), .B2(n17980), .ZN(
        P3_U2678) );
  INV_X1 U20911 ( .A(n17667), .ZN(n17678) );
  AOI21_X1 U20912 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17980), .A(n17678), .ZN(
        n17671) );
  AOI21_X1 U20913 ( .B1(n17669), .B2(n17674), .A(n17668), .ZN(n18021) );
  INV_X1 U20914 ( .A(n18021), .ZN(n17670) );
  OAI22_X1 U20915 ( .A1(n17672), .A2(n17671), .B1(n17980), .B2(n17670), .ZN(
        P3_U2679) );
  AOI21_X1 U20916 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17980), .A(n17673), .ZN(
        n17677) );
  OAI21_X1 U20917 ( .B1(n17676), .B2(n17675), .A(n17674), .ZN(n18030) );
  OAI22_X1 U20918 ( .A1(n17678), .A2(n17677), .B1(n17980), .B2(n18030), .ZN(
        P3_U2680) );
  AOI22_X1 U20919 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U20920 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17912), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17681) );
  AOI22_X1 U20921 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U20922 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17793), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17679) );
  NAND4_X1 U20923 ( .A1(n17682), .A2(n17681), .A3(n17680), .A4(n17679), .ZN(
        n17693) );
  INV_X1 U20924 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17691) );
  INV_X1 U20925 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17684) );
  INV_X1 U20926 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17683) );
  OAI22_X1 U20927 ( .A1(n17818), .A2(n17684), .B1(n17939), .B2(n17683), .ZN(
        n17688) );
  INV_X1 U20928 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17686) );
  OAI22_X1 U20929 ( .A1(n17891), .A2(n17686), .B1(n17918), .B2(n17685), .ZN(
        n17687) );
  AOI211_X1 U20930 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17688), .B(n17687), .ZN(n17690) );
  AOI22_X1 U20931 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17689) );
  OAI211_X1 U20932 ( .C1(n17950), .C2(n17691), .A(n17690), .B(n17689), .ZN(
        n17692) );
  NOR2_X1 U20933 ( .A1(n17693), .A2(n17692), .ZN(n18033) );
  NAND3_X1 U20934 ( .A1(n17695), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17980), 
        .ZN(n17694) );
  OAI221_X1 U20935 ( .B1(n17695), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17980), 
        .C2(n18033), .A(n17694), .ZN(P3_U2681) );
  NOR2_X1 U20936 ( .A1(n17950), .A2(n17696), .ZN(n17700) );
  OAI22_X1 U20937 ( .A1(n11436), .A2(n17698), .B1(n17799), .B2(n17697), .ZN(
        n17699) );
  AOI211_X1 U20938 ( .C1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .C2(n17933), .A(
        n17700), .B(n17699), .ZN(n17703) );
  AOI22_X1 U20939 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17793), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17702) );
  AOI22_X1 U20940 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17701) );
  NAND3_X1 U20941 ( .A1(n17703), .A2(n17702), .A3(n17701), .ZN(n17716) );
  AOI22_X1 U20942 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17705) );
  NAND2_X1 U20943 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n17704) );
  OAI211_X1 U20944 ( .C1(n11488), .C2(n17706), .A(n17705), .B(n17704), .ZN(
        n17714) );
  OAI22_X1 U20945 ( .A1(n17709), .A2(n17708), .B1(n9754), .B2(n17707), .ZN(
        n17713) );
  INV_X1 U20946 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17710) );
  OAI22_X1 U20947 ( .A1(n9666), .A2(n17711), .B1(n17918), .B2(n17710), .ZN(
        n17712) );
  OR3_X1 U20948 ( .A1(n17714), .A2(n17713), .A3(n17712), .ZN(n17715) );
  NOR2_X1 U20949 ( .A1(n17716), .A2(n17715), .ZN(n18039) );
  AOI21_X1 U20950 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17756), .A(n17985), .ZN(
        n17734) );
  AOI22_X1 U20951 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17734), .B1(n17718), 
        .B2(n17717), .ZN(n17719) );
  OAI21_X1 U20952 ( .B1(n18039), .B2(n17980), .A(n17719), .ZN(P3_U2682) );
  INV_X1 U20953 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17726) );
  INV_X1 U20954 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17850) );
  INV_X1 U20955 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17720) );
  OAI22_X1 U20956 ( .A1(n17941), .A2(n17850), .B1(n17939), .B2(n17720), .ZN(
        n17723) );
  INV_X1 U20957 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17721) );
  OAI22_X1 U20958 ( .A1(n17891), .A2(n17721), .B1(n17747), .B2(n17856), .ZN(
        n17722) );
  AOI211_X1 U20959 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17723), .B(n17722), .ZN(n17725) );
  AOI22_X1 U20960 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17724) );
  OAI211_X1 U20961 ( .C1(n17950), .C2(n17726), .A(n17725), .B(n17724), .ZN(
        n17732) );
  AOI22_X1 U20962 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17730) );
  AOI22_X1 U20963 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17729) );
  AOI22_X1 U20964 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17728) );
  AOI22_X1 U20965 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17727) );
  NAND4_X1 U20966 ( .A1(n17730), .A2(n17729), .A3(n17728), .A4(n17727), .ZN(
        n17731) );
  NOR2_X1 U20967 ( .A1(n17732), .A2(n17731), .ZN(n18044) );
  INV_X1 U20968 ( .A(n17733), .ZN(n17735) );
  OAI21_X1 U20969 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17735), .A(n17734), .ZN(
        n17736) );
  OAI21_X1 U20970 ( .B1(n18044), .B2(n17980), .A(n17736), .ZN(P3_U2683) );
  INV_X1 U20971 ( .A(n17737), .ZN(n17738) );
  OAI21_X1 U20972 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17738), .A(n17980), .ZN(
        n17755) );
  AOI22_X1 U20973 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17739) );
  OAI21_X1 U20974 ( .B1(n9668), .B2(n17740), .A(n17739), .ZN(n17741) );
  AOI21_X1 U20975 ( .B1(n17858), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n17741), .ZN(n17744) );
  AOI22_X1 U20976 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17743) );
  AOI22_X1 U20977 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17742) );
  NAND3_X1 U20978 ( .A1(n17744), .A2(n17743), .A3(n17742), .ZN(n17754) );
  OAI22_X1 U20979 ( .A1(n17747), .A2(n17746), .B1(n17799), .B2(n17745), .ZN(
        n17748) );
  AOI21_X1 U20980 ( .B1(n17932), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17748), .ZN(n17752) );
  AOI22_X1 U20981 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U20982 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17750) );
  NAND2_X1 U20983 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n17749) );
  NAND4_X1 U20984 ( .A1(n17752), .A2(n17751), .A3(n17750), .A4(n17749), .ZN(
        n17753) );
  NOR2_X1 U20985 ( .A1(n17754), .A2(n17753), .ZN(n18052) );
  OAI22_X1 U20986 ( .A1(n17756), .A2(n17755), .B1(n18052), .B2(n17980), .ZN(
        P3_U2684) );
  OR2_X1 U20987 ( .A1(n17774), .A2(n17757), .ZN(n17776) );
  AOI22_X1 U20988 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17758) );
  OAI21_X1 U20989 ( .B1(n17918), .B2(n17759), .A(n17758), .ZN(n17760) );
  AOI21_X1 U20990 ( .B1(n17858), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17760), .ZN(n17763) );
  AOI22_X1 U20991 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17762) );
  AOI22_X1 U20992 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17761) );
  NAND3_X1 U20993 ( .A1(n17763), .A2(n17762), .A3(n17761), .ZN(n17772) );
  AOI22_X1 U20994 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17765) );
  NAND2_X1 U20995 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n17764) );
  OAI211_X1 U20996 ( .C1(n17766), .C2(n17943), .A(n17765), .B(n17764), .ZN(
        n17767) );
  INV_X1 U20997 ( .A(n17767), .ZN(n17770) );
  AOI22_X1 U20998 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U20999 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17768) );
  NAND3_X1 U21000 ( .A1(n17770), .A2(n17769), .A3(n17768), .ZN(n17771) );
  NOR2_X1 U21001 ( .A1(n17772), .A2(n17771), .ZN(n18057) );
  NAND2_X1 U21002 ( .A1(n18910), .A2(n17844), .ZN(n17843) );
  NOR2_X1 U21003 ( .A1(n17773), .A2(n17843), .ZN(n17791) );
  NAND3_X1 U21004 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17791), .A3(n17774), 
        .ZN(n17775) );
  OAI221_X1 U21005 ( .B1(n17985), .B2(n17776), .C1(n17980), .C2(n18057), .A(
        n17775), .ZN(P3_U2685) );
  AOI22_X1 U21006 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U21007 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U21008 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U21009 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17793), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17777) );
  NAND4_X1 U21010 ( .A1(n17780), .A2(n17779), .A3(n17778), .A4(n17777), .ZN(
        n17787) );
  OAI22_X1 U21011 ( .A1(n9668), .A2(n17909), .B1(n17939), .B2(n17781), .ZN(
        n17783) );
  INV_X1 U21012 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21446) );
  INV_X1 U21013 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17919) );
  OAI22_X1 U21014 ( .A1(n17943), .A2(n21446), .B1(n17747), .B2(n17919), .ZN(
        n17782) );
  AOI211_X1 U21015 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17783), .B(n17782), .ZN(n17785) );
  AOI22_X1 U21016 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17784) );
  OAI211_X1 U21017 ( .C1(n17950), .C2(n17908), .A(n17785), .B(n17784), .ZN(
        n17786) );
  NOR2_X1 U21018 ( .A1(n17787), .A2(n17786), .ZN(n18062) );
  NAND2_X1 U21019 ( .A1(n18910), .A2(n17788), .ZN(n17809) );
  INV_X1 U21020 ( .A(n17809), .ZN(n17790) );
  NAND2_X1 U21021 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17981), .ZN(n17789) );
  OAI22_X1 U21022 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17791), .B1(n17790), 
        .B2(n17789), .ZN(n17792) );
  OAI21_X1 U21023 ( .B1(n18062), .B2(n17980), .A(n17792), .ZN(P3_U2686) );
  NAND3_X1 U21024 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17844), .ZN(n17810) );
  AOI22_X1 U21025 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17912), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17797) );
  AOI22_X1 U21026 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17796) );
  AOI22_X1 U21027 ( .A1(n17793), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17795) );
  AOI22_X1 U21028 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17794) );
  NAND4_X1 U21029 ( .A1(n17797), .A2(n17796), .A3(n17795), .A4(n17794), .ZN(
        n17807) );
  INV_X1 U21030 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17938) );
  INV_X1 U21031 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17798) );
  OAI22_X1 U21032 ( .A1(n9754), .A2(n17938), .B1(n17799), .B2(n17798), .ZN(
        n17803) );
  OAI22_X1 U21033 ( .A1(n17943), .A2(n17801), .B1(n17747), .B2(n17800), .ZN(
        n17802) );
  AOI211_X1 U21034 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17803), .B(n17802), .ZN(n17805) );
  AOI22_X1 U21035 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17804) );
  OAI211_X1 U21036 ( .C1(n17950), .C2(n17940), .A(n17805), .B(n17804), .ZN(
        n17806) );
  NOR2_X1 U21037 ( .A1(n17807), .A2(n17806), .ZN(n18069) );
  INV_X1 U21038 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17808) );
  NAND2_X1 U21039 ( .A1(n17980), .A2(n17810), .ZN(n17827) );
  OAI222_X1 U21040 ( .A1(n17810), .A2(n17809), .B1(n17980), .B2(n18069), .C1(
        n17808), .C2(n17827), .ZN(P3_U2687) );
  AOI22_X1 U21041 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11322), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17814) );
  AOI22_X1 U21042 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U21043 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17812) );
  AOI22_X1 U21044 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17811) );
  NAND4_X1 U21045 ( .A1(n17814), .A2(n17813), .A3(n17812), .A4(n17811), .ZN(
        n17826) );
  INV_X1 U21046 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17824) );
  OAI22_X1 U21047 ( .A1(n17709), .A2(n17816), .B1(n17939), .B2(n17815), .ZN(
        n17821) );
  INV_X1 U21048 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17819) );
  INV_X1 U21049 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17817) );
  OAI22_X1 U21050 ( .A1(n9754), .A2(n17819), .B1(n17818), .B2(n17817), .ZN(
        n17820) );
  AOI211_X1 U21051 ( .C1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .C2(n17872), .A(
        n17821), .B(n17820), .ZN(n17823) );
  AOI22_X1 U21052 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17822) );
  OAI211_X1 U21053 ( .C1(n17950), .C2(n17824), .A(n17823), .B(n17822), .ZN(
        n17825) );
  NOR2_X1 U21054 ( .A1(n17826), .A2(n17825), .ZN(n18074) );
  AOI21_X1 U21055 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17844), .A(
        P3_EBX_REG_15__SCAN_IN), .ZN(n17828) );
  OAI22_X1 U21056 ( .A1(n18074), .A2(n17980), .B1(n17828), .B2(n17827), .ZN(
        P3_U2688) );
  AOI22_X1 U21057 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17829) );
  OAI21_X1 U21058 ( .B1(n17918), .B2(n17830), .A(n17829), .ZN(n17831) );
  AOI21_X1 U21059 ( .B1(n17858), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17831), .ZN(n17834) );
  AOI22_X1 U21060 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11322), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U21061 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17832) );
  NAND3_X1 U21062 ( .A1(n17834), .A2(n17833), .A3(n17832), .ZN(n17842) );
  AOI22_X1 U21063 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17835) );
  OAI21_X1 U21064 ( .B1(n9668), .B2(n17836), .A(n17835), .ZN(n17837) );
  AOI21_X1 U21065 ( .B1(n17894), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17837), .ZN(n17840) );
  AOI22_X1 U21066 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U21067 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17921), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17838) );
  NAND3_X1 U21068 ( .A1(n17840), .A2(n17839), .A3(n17838), .ZN(n17841) );
  NOR2_X1 U21069 ( .A1(n17842), .A2(n17841), .ZN(n18079) );
  INV_X1 U21070 ( .A(n17843), .ZN(n17846) );
  NAND2_X1 U21071 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17844), .ZN(n17845) );
  OAI21_X1 U21072 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17846), .A(n17845), .ZN(
        n17847) );
  AOI22_X1 U21073 ( .A1(n17985), .A2(n18079), .B1(n17847), .B2(n17980), .ZN(
        P3_U2689) );
  AOI22_X1 U21074 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U21075 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n17848) );
  OAI211_X1 U21076 ( .C1(n17850), .C2(n17943), .A(n17849), .B(n17848), .ZN(
        n17851) );
  INV_X1 U21077 ( .A(n17851), .ZN(n17854) );
  AOI22_X1 U21078 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U21079 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17852) );
  NAND3_X1 U21080 ( .A1(n17854), .A2(n17853), .A3(n17852), .ZN(n17863) );
  AOI22_X1 U21081 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17855) );
  OAI21_X1 U21082 ( .B1(n17918), .B2(n17856), .A(n17855), .ZN(n17857) );
  AOI21_X1 U21083 ( .B1(n17858), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17857), .ZN(n17861) );
  AOI22_X1 U21084 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17860) );
  AOI22_X1 U21085 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17859) );
  NAND3_X1 U21086 ( .A1(n17861), .A2(n17860), .A3(n17859), .ZN(n17862) );
  NOR2_X1 U21087 ( .A1(n17863), .A2(n17862), .ZN(n18085) );
  AOI21_X1 U21088 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17906), .A(n17985), .ZN(
        n17885) );
  NAND2_X1 U21089 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17885), .ZN(n17866) );
  INV_X1 U21090 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17864) );
  NAND4_X1 U21091 ( .A1(n18910), .A2(P3_EBX_REG_11__SCAN_IN), .A3(n17906), 
        .A4(n17864), .ZN(n17865) );
  OAI211_X1 U21092 ( .C1(n18085), .C2(n17980), .A(n17866), .B(n17865), .ZN(
        P3_U2691) );
  NAND2_X1 U21093 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n17869) );
  NAND2_X1 U21094 ( .A1(n17867), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n17868) );
  OAI211_X1 U21095 ( .C1(n17950), .C2(n17870), .A(n17869), .B(n17868), .ZN(
        n17871) );
  INV_X1 U21096 ( .A(n17871), .ZN(n17876) );
  AOI22_X1 U21097 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17875) );
  AOI22_X1 U21098 ( .A1(n17898), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17874) );
  NAND2_X1 U21099 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n17873) );
  NAND4_X1 U21100 ( .A1(n17876), .A2(n17875), .A3(n17874), .A4(n17873), .ZN(
        n17884) );
  AOI22_X1 U21101 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17882) );
  AOI22_X1 U21102 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9625), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17881) );
  INV_X1 U21103 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n21397) );
  AOI22_X1 U21104 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17933), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17880) );
  AOI22_X1 U21105 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17879) );
  NAND4_X1 U21106 ( .A1(n17882), .A2(n17881), .A3(n17880), .A4(n17879), .ZN(
        n17883) );
  OR2_X1 U21107 ( .A1(n17884), .A2(n17883), .ZN(n18088) );
  INV_X1 U21108 ( .A(n18088), .ZN(n17887) );
  OAI21_X1 U21109 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17906), .A(n17885), .ZN(
        n17886) );
  OAI21_X1 U21110 ( .B1(n17887), .B2(n17980), .A(n17886), .ZN(P3_U2692) );
  OAI21_X1 U21111 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17927), .A(n17980), .ZN(
        n17905) );
  INV_X1 U21112 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17897) );
  INV_X1 U21113 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17889) );
  INV_X1 U21114 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17888) );
  OAI22_X1 U21115 ( .A1(n9666), .A2(n17889), .B1(n17943), .B2(n17888), .ZN(
        n17893) );
  OAI22_X1 U21116 ( .A1(n11436), .A2(n21374), .B1(n17891), .B2(n17890), .ZN(
        n17892) );
  AOI211_X1 U21117 ( .C1(n17894), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17893), .B(n17892), .ZN(n17896) );
  AOI22_X1 U21118 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17895) );
  OAI211_X1 U21119 ( .C1(n17950), .C2(n17897), .A(n17896), .B(n17895), .ZN(
        n17904) );
  AOI22_X1 U21120 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11322), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17902) );
  AOI22_X1 U21121 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17901) );
  AOI22_X1 U21122 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17898), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17900) );
  AOI22_X1 U21123 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17899) );
  NAND4_X1 U21124 ( .A1(n17902), .A2(n17901), .A3(n17900), .A4(n17899), .ZN(
        n17903) );
  NOR2_X1 U21125 ( .A1(n17904), .A2(n17903), .ZN(n18091) );
  OAI22_X1 U21126 ( .A1(n17906), .A2(n17905), .B1(n18091), .B2(n17980), .ZN(
        P3_U2693) );
  NOR2_X1 U21127 ( .A1(n17950), .A2(n17907), .ZN(n17911) );
  OAI22_X1 U21128 ( .A1(n11436), .A2(n17909), .B1(n17941), .B2(n17908), .ZN(
        n17910) );
  AOI211_X1 U21129 ( .C1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .C2(n17933), .A(
        n17911), .B(n17910), .ZN(n17915) );
  AOI22_X1 U21130 ( .A1(n17912), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17914) );
  AOI22_X1 U21131 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17913) );
  NAND3_X1 U21132 ( .A1(n17915), .A2(n17914), .A3(n17913), .ZN(n17926) );
  AOI22_X1 U21133 ( .A1(n17931), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11411), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17917) );
  NAND2_X1 U21134 ( .A1(n17872), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n17916) );
  OAI211_X1 U21135 ( .C1(n17919), .C2(n17918), .A(n17917), .B(n17916), .ZN(
        n17920) );
  INV_X1 U21136 ( .A(n17920), .ZN(n17924) );
  AOI22_X1 U21137 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11322), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U21138 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17922) );
  NAND3_X1 U21139 ( .A1(n17924), .A2(n17923), .A3(n17922), .ZN(n17925) );
  NOR2_X1 U21140 ( .A1(n17926), .A2(n17925), .ZN(n18096) );
  AOI221_X1 U21141 ( .B1(n17928), .B2(n17953), .C1(n17928), .C2(n17954), .A(
        n17927), .ZN(n17929) );
  INV_X1 U21142 ( .A(n17929), .ZN(n17930) );
  AOI22_X1 U21143 ( .A1(n17985), .A2(n18096), .B1(n17930), .B2(n17980), .ZN(
        P3_U2694) );
  AOI22_X1 U21144 ( .A1(n11322), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17931), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U21145 ( .A1(n17877), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17912), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17936) );
  AOI22_X1 U21146 ( .A1(n17921), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17935) );
  AOI22_X1 U21147 ( .A1(n17933), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17934) );
  NAND4_X1 U21148 ( .A1(n17937), .A2(n17936), .A3(n17935), .A4(n17934), .ZN(
        n17952) );
  INV_X1 U21149 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17949) );
  OAI22_X1 U21150 ( .A1(n17941), .A2(n17940), .B1(n17939), .B2(n17938), .ZN(
        n17946) );
  OAI22_X1 U21151 ( .A1(n9754), .A2(n17944), .B1(n17943), .B2(n17942), .ZN(
        n17945) );
  AOI211_X1 U21152 ( .C1(n17872), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n17946), .B(n17945), .ZN(n17948) );
  AOI22_X1 U21153 ( .A1(n9625), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17947) );
  OAI211_X1 U21154 ( .C1(n17950), .C2(n17949), .A(n17948), .B(n17947), .ZN(
        n17951) );
  NOR2_X1 U21155 ( .A1(n17952), .A2(n17951), .ZN(n18103) );
  OAI33_X1 U21156 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18031), .A3(n17954), .B1(
        n17953), .B2(n17985), .B3(n17959), .ZN(n17955) );
  INV_X1 U21157 ( .A(n17955), .ZN(n17956) );
  OAI21_X1 U21158 ( .B1(n18103), .B2(n17980), .A(n17956), .ZN(P3_U2695) );
  NAND2_X1 U21159 ( .A1(n17980), .A2(n17957), .ZN(n17963) );
  NAND2_X1 U21160 ( .A1(n18910), .A2(n17981), .ZN(n17987) );
  NOR4_X1 U21161 ( .A1(n17959), .A2(n17958), .A3(n17968), .A4(n17987), .ZN(
        n17960) );
  AOI21_X1 U21162 ( .B1(n17985), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n17960), .ZN(n17961) );
  OAI21_X1 U21163 ( .B1(n17962), .B2(n17963), .A(n17961), .ZN(P3_U2696) );
  NOR2_X1 U21164 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17967), .ZN(n17964) );
  OAI22_X1 U21165 ( .A1(n17964), .A2(n17963), .B1(n11320), .B2(n17980), .ZN(
        P3_U2697) );
  NOR2_X1 U21166 ( .A1(n17984), .A2(n17968), .ZN(n17965) );
  OAI21_X1 U21167 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17965), .A(n17980), .ZN(
        n17966) );
  OAI22_X1 U21168 ( .A1(n17967), .A2(n17966), .B1(n11466), .B2(n17980), .ZN(
        P3_U2698) );
  NOR2_X1 U21169 ( .A1(n17968), .A2(n17987), .ZN(n17973) );
  INV_X1 U21170 ( .A(n17969), .ZN(n17970) );
  NOR2_X1 U21171 ( .A1(n17970), .A2(n17987), .ZN(n17978) );
  AND2_X1 U21172 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17978), .ZN(n17975) );
  AOI21_X1 U21173 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17980), .A(n17975), .ZN(
        n17972) );
  INV_X1 U21174 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17971) );
  OAI22_X1 U21175 ( .A1(n17973), .A2(n17972), .B1(n17971), .B2(n17980), .ZN(
        P3_U2699) );
  AOI21_X1 U21176 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17980), .A(n17978), .ZN(
        n17974) );
  OAI22_X1 U21177 ( .A1(n17975), .A2(n17974), .B1(n17740), .B2(n17980), .ZN(
        P3_U2700) );
  INV_X1 U21178 ( .A(n17976), .ZN(n17977) );
  AOI221_X1 U21179 ( .B1(n17977), .B2(n17981), .C1(n18031), .C2(n17981), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17979) );
  AOI211_X1 U21180 ( .C1(n17985), .C2(n21374), .A(n17979), .B(n17978), .ZN(
        P3_U2701) );
  OAI222_X1 U21181 ( .A1(n17987), .A2(n17983), .B1(n17982), .B2(n17981), .C1(
        n17909), .C2(n17980), .ZN(P3_U2702) );
  AOI22_X1 U21182 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17985), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17984), .ZN(n17986) );
  OAI21_X1 U21183 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17987), .A(n17986), .ZN(
        P3_U2703) );
  INV_X1 U21184 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18137) );
  INV_X1 U21185 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18140) );
  INV_X1 U21186 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18240) );
  INV_X1 U21187 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18170) );
  INV_X1 U21188 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18215) );
  NOR2_X1 U21189 ( .A1(n18215), .A2(n18125), .ZN(n17988) );
  NAND4_X1 U21190 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n17988), .ZN(n18109) );
  INV_X1 U21191 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18235) );
  INV_X1 U21192 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18227) );
  INV_X1 U21193 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18166) );
  INV_X1 U21194 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18168) );
  NOR3_X1 U21195 ( .A1(n18227), .A2(n18166), .A3(n18168), .ZN(n18084) );
  NAND3_X1 U21196 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(n18084), .ZN(n18076) );
  NOR2_X1 U21197 ( .A1(n18235), .A2(n18076), .ZN(n18071) );
  NOR2_X2 U21198 ( .A1(n18240), .A2(n18070), .ZN(n18066) );
  NAND2_X1 U21199 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18066), .ZN(n18065) );
  NAND3_X1 U21200 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .ZN(n18032) );
  NAND3_X1 U21201 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n17989) );
  NOR3_X2 U21202 ( .A1(n18065), .A2(n18032), .A3(n17989), .ZN(n18027) );
  NAND2_X1 U21203 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18027), .ZN(n18026) );
  NAND2_X1 U21204 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17994), .ZN(n17993) );
  NAND2_X1 U21205 ( .A1(n17993), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17992) );
  NAND2_X1 U21206 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18063), .ZN(n17991) );
  OAI221_X1 U21207 ( .B1(n17993), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17992), 
        .C2(n18100), .A(n17991), .ZN(P3_U2704) );
  NAND2_X1 U21208 ( .A1(n18896), .A2(n18100), .ZN(n18038) );
  AOI22_X1 U21209 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18063), .ZN(n17996) );
  OAI211_X1 U21210 ( .C1(n17994), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18118), .B(
        n17993), .ZN(n17995) );
  OAI211_X1 U21211 ( .C1(n17997), .C2(n18120), .A(n17996), .B(n17995), .ZN(
        P3_U2705) );
  AOI22_X1 U21212 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18063), .ZN(n18000) );
  OAI211_X1 U21213 ( .C1(n9674), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18118), .B(
        n17998), .ZN(n17999) );
  OAI211_X1 U21214 ( .C1(n18001), .C2(n18120), .A(n18000), .B(n17999), .ZN(
        P3_U2706) );
  INV_X1 U21215 ( .A(n18063), .ZN(n18043) );
  AOI22_X1 U21216 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18064), .B1(n18127), .B2(
        n18002), .ZN(n18005) );
  AOI211_X1 U21217 ( .C1(n18137), .C2(n18006), .A(n9674), .B(n18100), .ZN(
        n18003) );
  INV_X1 U21218 ( .A(n18003), .ZN(n18004) );
  OAI211_X1 U21219 ( .C1(n18043), .C2(n18890), .A(n18005), .B(n18004), .ZN(
        P3_U2707) );
  AOI22_X1 U21220 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18063), .ZN(n18008) );
  OAI211_X1 U21221 ( .C1(n18011), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18118), .B(
        n18006), .ZN(n18007) );
  OAI211_X1 U21222 ( .C1(n18009), .C2(n18120), .A(n18008), .B(n18007), .ZN(
        P3_U2708) );
  AOI22_X1 U21223 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18064), .B1(n18127), .B2(
        n18010), .ZN(n18014) );
  AOI211_X1 U21224 ( .C1(n18140), .C2(n18016), .A(n18011), .B(n18100), .ZN(
        n18012) );
  INV_X1 U21225 ( .A(n18012), .ZN(n18013) );
  OAI211_X1 U21226 ( .C1(n18043), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        P3_U2709) );
  AOI22_X1 U21227 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18063), .ZN(n18019) );
  OAI211_X1 U21228 ( .C1(n18017), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18118), .B(
        n18016), .ZN(n18018) );
  OAI211_X1 U21229 ( .C1(n18020), .C2(n18120), .A(n18019), .B(n18018), .ZN(
        P3_U2710) );
  AOI22_X1 U21230 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18063), .B1(n18127), .B2(
        n18021), .ZN(n18025) );
  OAI211_X1 U21231 ( .C1(n18023), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18118), .B(
        n18022), .ZN(n18024) );
  OAI211_X1 U21232 ( .C1(n18038), .C2(n18222), .A(n18025), .B(n18024), .ZN(
        P3_U2711) );
  AOI22_X1 U21233 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18063), .ZN(n18029) );
  OAI211_X1 U21234 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18027), .A(n18118), .B(
        n18026), .ZN(n18028) );
  OAI211_X1 U21235 ( .C1(n18030), .C2(n18120), .A(n18029), .B(n18028), .ZN(
        P3_U2712) );
  INV_X1 U21236 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18154) );
  NAND2_X1 U21237 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18059), .ZN(n18058) );
  NAND3_X1 U21238 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n18049), .ZN(n18042) );
  NAND2_X1 U21239 ( .A1(n18118), .A2(n18042), .ZN(n18047) );
  OAI21_X1 U21240 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18124), .A(n18047), .ZN(
        n18036) );
  INV_X1 U21241 ( .A(n18049), .ZN(n18053) );
  NOR3_X1 U21242 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18032), .A3(n18053), .ZN(
        n18035) );
  OAI22_X1 U21243 ( .A1(n18033), .A2(n18120), .B1(n18903), .B2(n18043), .ZN(
        n18034) );
  AOI211_X1 U21244 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n18036), .A(n18035), .B(
        n18034), .ZN(n18037) );
  OAI21_X1 U21245 ( .B1(n18902), .B2(n18038), .A(n18037), .ZN(P3_U2713) );
  INV_X1 U21246 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18149) );
  OAI22_X1 U21247 ( .A1(n18039), .A2(n18120), .B1(n18895), .B2(n18043), .ZN(
        n18040) );
  AOI21_X1 U21248 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18064), .A(n18040), .ZN(
        n18041) );
  OAI221_X1 U21249 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18042), .C1(n18149), 
        .C2(n18047), .A(n18041), .ZN(P3_U2714) );
  NAND2_X1 U21250 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18049), .ZN(n18048) );
  INV_X1 U21251 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18151) );
  OAI22_X1 U21252 ( .A1(n18044), .A2(n18120), .B1(n18892), .B2(n18043), .ZN(
        n18045) );
  AOI21_X1 U21253 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n18064), .A(n18045), .ZN(
        n18046) );
  OAI221_X1 U21254 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n18048), .C1(n18151), 
        .C2(n18047), .A(n18046), .ZN(P3_U2715) );
  AOI22_X1 U21255 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18063), .ZN(n18051) );
  OAI211_X1 U21256 ( .C1(n18049), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18118), .B(
        n18048), .ZN(n18050) );
  OAI211_X1 U21257 ( .C1(n18052), .C2(n18120), .A(n18051), .B(n18050), .ZN(
        P3_U2716) );
  AOI22_X1 U21258 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18063), .ZN(n18056) );
  INV_X1 U21259 ( .A(n18058), .ZN(n18054) );
  OAI211_X1 U21260 ( .C1(n18054), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18118), .B(
        n18053), .ZN(n18055) );
  OAI211_X1 U21261 ( .C1(n18057), .C2(n18120), .A(n18056), .B(n18055), .ZN(
        P3_U2717) );
  AOI22_X1 U21262 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18063), .ZN(n18061) );
  OAI211_X1 U21263 ( .C1(n18059), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18118), .B(
        n18058), .ZN(n18060) );
  OAI211_X1 U21264 ( .C1(n18062), .C2(n18120), .A(n18061), .B(n18060), .ZN(
        P3_U2718) );
  AOI22_X1 U21265 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18064), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18063), .ZN(n18068) );
  OAI211_X1 U21266 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18066), .A(n18118), .B(
        n18065), .ZN(n18067) );
  OAI211_X1 U21267 ( .C1(n18069), .C2(n18120), .A(n18068), .B(n18067), .ZN(
        P3_U2719) );
  AND2_X1 U21268 ( .A1(n18118), .A2(n18070), .ZN(n18075) );
  AOI22_X1 U21269 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n18075), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18128), .ZN(n18073) );
  NAND2_X1 U21270 ( .A1(n18910), .A2(n18099), .ZN(n18094) );
  NAND3_X1 U21271 ( .A1(n18071), .A2(n18095), .A3(n18240), .ZN(n18072) );
  OAI211_X1 U21272 ( .C1(n18074), .C2(n18120), .A(n18073), .B(n18072), .ZN(
        P3_U2720) );
  AOI22_X1 U21273 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18128), .B1(
        P3_EAX_REG_14__SCAN_IN), .B2(n18075), .ZN(n18078) );
  OR3_X1 U21274 ( .A1(n18076), .A2(n18094), .A3(P3_EAX_REG_14__SCAN_IN), .ZN(
        n18077) );
  OAI211_X1 U21275 ( .C1(n18079), .C2(n18120), .A(n18078), .B(n18077), .ZN(
        P3_U2721) );
  NAND3_X1 U21276 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18084), .A3(n18095), 
        .ZN(n18083) );
  NAND2_X1 U21277 ( .A1(n18083), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n18082) );
  AOI22_X1 U21278 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18128), .B1(n18127), .B2(
        n18080), .ZN(n18081) );
  OAI221_X1 U21279 ( .B1(n18083), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n18082), 
        .C2(n18100), .A(n18081), .ZN(P3_U2722) );
  INV_X1 U21280 ( .A(n18083), .ZN(n18087) );
  AOI22_X1 U21281 ( .A1(n18095), .A2(n18084), .B1(P3_EAX_REG_12__SCAN_IN), 
        .B2(n18118), .ZN(n18086) );
  OAI222_X1 U21282 ( .A1(n18123), .A2(n18231), .B1(n18087), .B2(n18086), .C1(
        n18120), .C2(n18085), .ZN(P3_U2723) );
  NAND3_X1 U21283 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n18095), .ZN(n18090) );
  NAND2_X1 U21284 ( .A1(n18118), .A2(n18090), .ZN(n18093) );
  AOI22_X1 U21285 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18128), .B1(n18127), .B2(
        n18088), .ZN(n18089) );
  OAI221_X1 U21286 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18090), .C1(n18227), 
        .C2(n18093), .A(n18089), .ZN(P3_U2724) );
  AOI21_X1 U21287 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18095), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n18092) );
  OAI222_X1 U21288 ( .A1(n18123), .A2(n18225), .B1(n18093), .B2(n18092), .C1(
        n18120), .C2(n18091), .ZN(P3_U2725) );
  NOR2_X1 U21289 ( .A1(n18168), .A2(n18094), .ZN(n18098) );
  AOI21_X1 U21290 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18118), .A(n18095), .ZN(
        n18097) );
  OAI222_X1 U21291 ( .A1(n18123), .A2(n13579), .B1(n18098), .B2(n18097), .C1(
        n18120), .C2(n18096), .ZN(P3_U2726) );
  AOI211_X1 U21292 ( .C1(n18170), .C2(n18105), .A(n18100), .B(n18099), .ZN(
        n18101) );
  AOI21_X1 U21293 ( .B1(n18128), .B2(BUF2_REG_8__SCAN_IN), .A(n18101), .ZN(
        n18102) );
  OAI21_X1 U21294 ( .B1(n18103), .B2(n18120), .A(n18102), .ZN(P3_U2727) );
  AOI22_X1 U21295 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18128), .B1(n18127), .B2(
        n18104), .ZN(n18108) );
  OAI211_X1 U21296 ( .C1(P3_EAX_REG_7__SCAN_IN), .C2(n18106), .A(n18118), .B(
        n18105), .ZN(n18107) );
  NAND2_X1 U21297 ( .A1(n18108), .A2(n18107), .ZN(P3_U2728) );
  NOR2_X1 U21298 ( .A1(n18109), .A2(n18124), .ZN(n18112) );
  INV_X1 U21299 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18177) );
  NOR3_X1 U21300 ( .A1(n18215), .A2(n18125), .A3(n18124), .ZN(n18117) );
  NAND2_X1 U21301 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18117), .ZN(n18113) );
  NOR2_X1 U21302 ( .A1(n18177), .A2(n18113), .ZN(n18115) );
  AOI21_X1 U21303 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18118), .A(n18115), .ZN(
        n18111) );
  OAI222_X1 U21304 ( .A1(n18123), .A2(n18902), .B1(n18112), .B2(n18111), .C1(
        n18120), .C2(n18110), .ZN(P3_U2729) );
  INV_X1 U21305 ( .A(n18113), .ZN(n18122) );
  AOI21_X1 U21306 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18118), .A(n18122), .ZN(
        n18116) );
  OAI222_X1 U21307 ( .A1(n18123), .A2(n13582), .B1(n18116), .B2(n18115), .C1(
        n18120), .C2(n18114), .ZN(P3_U2730) );
  AOI21_X1 U21308 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18118), .A(n18117), .ZN(
        n18121) );
  OAI222_X1 U21309 ( .A1(n18891), .A2(n18123), .B1(n18122), .B2(n18121), .C1(
        n18120), .C2(n18119), .ZN(P3_U2731) );
  OR2_X1 U21310 ( .A1(n18125), .A2(n18124), .ZN(n18131) );
  AOI22_X1 U21311 ( .A1(n18128), .A2(BUF2_REG_3__SCAN_IN), .B1(n18127), .B2(
        n18126), .ZN(n18129) );
  OAI221_X1 U21312 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18131), .C1(n18215), 
        .C2(n18130), .A(n18129), .ZN(P3_U2732) );
  NAND2_X1 U21313 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18396), .ZN(n19341) );
  INV_X2 U21314 ( .A(n19341), .ZN(n18184) );
  AND2_X1 U21315 ( .A1(n18175), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21316 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18210) );
  NAND2_X1 U21317 ( .A1(n18171), .A2(n18133), .ZN(n18157) );
  AOI22_X1 U21318 ( .A1(n18184), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18134) );
  OAI21_X1 U21319 ( .B1(n18210), .B2(n18157), .A(n18134), .ZN(P3_U2737) );
  INV_X1 U21320 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18208) );
  AOI22_X1 U21321 ( .A1(n18184), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18135) );
  OAI21_X1 U21322 ( .B1(n18208), .B2(n18157), .A(n18135), .ZN(P3_U2738) );
  AOI22_X1 U21323 ( .A1(n18184), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18136) );
  OAI21_X1 U21324 ( .B1(n18137), .B2(n18157), .A(n18136), .ZN(P3_U2739) );
  INV_X1 U21325 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U21326 ( .A1(n18184), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18138) );
  OAI21_X1 U21327 ( .B1(n18205), .B2(n18157), .A(n18138), .ZN(P3_U2740) );
  AOI22_X1 U21328 ( .A1(n18184), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18139) );
  OAI21_X1 U21329 ( .B1(n18140), .B2(n18157), .A(n18139), .ZN(P3_U2741) );
  INV_X1 U21330 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U21331 ( .A1(n18184), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18141) );
  OAI21_X1 U21332 ( .B1(n18142), .B2(n18157), .A(n18141), .ZN(P3_U2742) );
  INV_X1 U21333 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18144) );
  AOI22_X1 U21334 ( .A1(n18184), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18143) );
  OAI21_X1 U21335 ( .B1(n18144), .B2(n18157), .A(n18143), .ZN(P3_U2743) );
  INV_X1 U21336 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U21337 ( .A1(n18184), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18145) );
  OAI21_X1 U21338 ( .B1(n18200), .B2(n18157), .A(n18145), .ZN(P3_U2744) );
  INV_X1 U21339 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18147) );
  AOI22_X1 U21340 ( .A1(n18184), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18146) );
  OAI21_X1 U21341 ( .B1(n18147), .B2(n18157), .A(n18146), .ZN(P3_U2745) );
  AOI22_X1 U21342 ( .A1(n18184), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18148) );
  OAI21_X1 U21343 ( .B1(n18149), .B2(n18157), .A(n18148), .ZN(P3_U2746) );
  AOI22_X1 U21344 ( .A1(n18184), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18150) );
  OAI21_X1 U21345 ( .B1(n18151), .B2(n18157), .A(n18150), .ZN(P3_U2747) );
  INV_X1 U21346 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18195) );
  AOI22_X1 U21347 ( .A1(n18184), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18152) );
  OAI21_X1 U21348 ( .B1(n18195), .B2(n18157), .A(n18152), .ZN(P3_U2748) );
  AOI22_X1 U21349 ( .A1(n18184), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18153) );
  OAI21_X1 U21350 ( .B1(n18154), .B2(n18157), .A(n18153), .ZN(P3_U2749) );
  INV_X1 U21351 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18192) );
  AOI22_X1 U21352 ( .A1(n18184), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18155) );
  OAI21_X1 U21353 ( .B1(n18192), .B2(n18157), .A(n18155), .ZN(P3_U2750) );
  INV_X1 U21354 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18158) );
  AOI22_X1 U21355 ( .A1(n18184), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18156) );
  OAI21_X1 U21356 ( .B1(n18158), .B2(n18157), .A(n18156), .ZN(P3_U2751) );
  AOI22_X1 U21357 ( .A1(n18184), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18159) );
  OAI21_X1 U21358 ( .B1(n18240), .B2(n18186), .A(n18159), .ZN(P3_U2752) );
  AOI22_X1 U21359 ( .A1(n18184), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18160) );
  OAI21_X1 U21360 ( .B1(n18235), .B2(n18186), .A(n18160), .ZN(P3_U2753) );
  INV_X1 U21361 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U21362 ( .A1(n18184), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18161) );
  OAI21_X1 U21363 ( .B1(n18233), .B2(n18186), .A(n18161), .ZN(P3_U2754) );
  INV_X1 U21364 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18163) );
  AOI22_X1 U21365 ( .A1(n18184), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18162) );
  OAI21_X1 U21366 ( .B1(n18163), .B2(n18186), .A(n18162), .ZN(P3_U2755) );
  AOI22_X1 U21367 ( .A1(n18184), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18164) );
  OAI21_X1 U21368 ( .B1(n18227), .B2(n18186), .A(n18164), .ZN(P3_U2756) );
  AOI22_X1 U21369 ( .A1(n18184), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18165) );
  OAI21_X1 U21370 ( .B1(n18166), .B2(n18186), .A(n18165), .ZN(P3_U2757) );
  AOI22_X1 U21371 ( .A1(n18184), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18167) );
  OAI21_X1 U21372 ( .B1(n18168), .B2(n18186), .A(n18167), .ZN(P3_U2758) );
  AOI22_X1 U21373 ( .A1(n18184), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18169) );
  OAI21_X1 U21374 ( .B1(n18170), .B2(n18186), .A(n18169), .ZN(P3_U2759) );
  INV_X1 U21375 ( .A(P3_LWORD_REG_7__SCAN_IN), .ZN(n21354) );
  AOI22_X1 U21376 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18171), .B1(n18183), .B2(
        P3_DATAO_REG_7__SCAN_IN), .ZN(n18172) );
  OAI21_X1 U21377 ( .B1(n19341), .B2(n21354), .A(n18172), .ZN(P3_U2760) );
  INV_X1 U21378 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U21379 ( .A1(n18184), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18173) );
  OAI21_X1 U21380 ( .B1(n18174), .B2(n18186), .A(n18173), .ZN(P3_U2761) );
  AOI22_X1 U21381 ( .A1(n18184), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18175), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18176) );
  OAI21_X1 U21382 ( .B1(n18177), .B2(n18186), .A(n18176), .ZN(P3_U2762) );
  INV_X1 U21383 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21428) );
  AOI22_X1 U21384 ( .A1(n18184), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18178) );
  OAI21_X1 U21385 ( .B1(n21428), .B2(n18186), .A(n18178), .ZN(P3_U2763) );
  AOI22_X1 U21386 ( .A1(n18184), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18179) );
  OAI21_X1 U21387 ( .B1(n18215), .B2(n18186), .A(n18179), .ZN(P3_U2764) );
  INV_X1 U21388 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18181) );
  AOI22_X1 U21389 ( .A1(n18184), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18180) );
  OAI21_X1 U21390 ( .B1(n18181), .B2(n18186), .A(n18180), .ZN(P3_U2765) );
  AOI22_X1 U21391 ( .A1(n18184), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18182) );
  OAI21_X1 U21392 ( .B1(n21450), .B2(n18186), .A(n18182), .ZN(P3_U2766) );
  AOI22_X1 U21393 ( .A1(n18184), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18183), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18185) );
  OAI21_X1 U21394 ( .B1(n18187), .B2(n18186), .A(n18185), .ZN(P3_U2767) );
  NOR3_X4 U21395 ( .A1(n19471), .A2(n18189), .A3(n18188), .ZN(n18228) );
  INV_X2 U21396 ( .A(n18220), .ZN(n18236) );
  AOI22_X1 U21397 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18236), .ZN(n18190) );
  OAI21_X1 U21398 ( .B1(n18871), .B2(n18230), .A(n18190), .ZN(P3_U2768) );
  INV_X1 U21399 ( .A(n18228), .ZN(n18239) );
  AOI22_X1 U21400 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18237), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18236), .ZN(n18191) );
  OAI21_X1 U21401 ( .B1(n18192), .B2(n18239), .A(n18191), .ZN(P3_U2769) );
  AOI22_X1 U21402 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18236), .ZN(n18193) );
  OAI21_X1 U21403 ( .B1(n18881), .B2(n18230), .A(n18193), .ZN(P3_U2770) );
  AOI22_X1 U21404 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18237), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18236), .ZN(n18194) );
  OAI21_X1 U21405 ( .B1(n18195), .B2(n18239), .A(n18194), .ZN(P3_U2771) );
  AOI22_X1 U21406 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18236), .ZN(n18196) );
  OAI21_X1 U21407 ( .B1(n18891), .B2(n18230), .A(n18196), .ZN(P3_U2772) );
  AOI22_X1 U21408 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18236), .ZN(n18197) );
  OAI21_X1 U21409 ( .B1(n13582), .B2(n18230), .A(n18197), .ZN(P3_U2773) );
  AOI22_X1 U21410 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18236), .ZN(n18198) );
  OAI21_X1 U21411 ( .B1(n18902), .B2(n18230), .A(n18198), .ZN(P3_U2774) );
  AOI22_X1 U21412 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18237), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18236), .ZN(n18199) );
  OAI21_X1 U21413 ( .B1(n18200), .B2(n18239), .A(n18199), .ZN(P3_U2775) );
  AOI22_X1 U21414 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18236), .ZN(n18201) );
  OAI21_X1 U21415 ( .B1(n18222), .B2(n18230), .A(n18201), .ZN(P3_U2776) );
  AOI22_X1 U21416 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18236), .ZN(n18202) );
  OAI21_X1 U21417 ( .B1(n13579), .B2(n18230), .A(n18202), .ZN(P3_U2777) );
  AOI22_X1 U21418 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18236), .ZN(n18203) );
  OAI21_X1 U21419 ( .B1(n18225), .B2(n18230), .A(n18203), .ZN(P3_U2778) );
  AOI22_X1 U21420 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18237), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18236), .ZN(n18204) );
  OAI21_X1 U21421 ( .B1(n18205), .B2(n18239), .A(n18204), .ZN(P3_U2779) );
  AOI22_X1 U21422 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18228), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18236), .ZN(n18206) );
  OAI21_X1 U21423 ( .B1(n18231), .B2(n18230), .A(n18206), .ZN(P3_U2780) );
  AOI22_X1 U21424 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18237), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18236), .ZN(n18207) );
  OAI21_X1 U21425 ( .B1(n18208), .B2(n18239), .A(n18207), .ZN(P3_U2781) );
  AOI22_X1 U21426 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18237), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18236), .ZN(n18209) );
  OAI21_X1 U21427 ( .B1(n18210), .B2(n18239), .A(n18209), .ZN(P3_U2782) );
  AOI22_X1 U21428 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18236), .ZN(n18211) );
  OAI21_X1 U21429 ( .B1(n18871), .B2(n18230), .A(n18211), .ZN(P3_U2783) );
  AOI22_X1 U21430 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18237), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18236), .ZN(n18212) );
  OAI21_X1 U21431 ( .B1(n21450), .B2(n18239), .A(n18212), .ZN(P3_U2784) );
  AOI22_X1 U21432 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18236), .ZN(n18213) );
  OAI21_X1 U21433 ( .B1(n18881), .B2(n18230), .A(n18213), .ZN(P3_U2785) );
  AOI22_X1 U21434 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18237), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18236), .ZN(n18214) );
  OAI21_X1 U21435 ( .B1(n18215), .B2(n18239), .A(n18214), .ZN(P3_U2786) );
  AOI22_X1 U21436 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18236), .ZN(n18216) );
  OAI21_X1 U21437 ( .B1(n18891), .B2(n18230), .A(n18216), .ZN(P3_U2787) );
  AOI22_X1 U21438 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18236), .ZN(n18217) );
  OAI21_X1 U21439 ( .B1(n13582), .B2(n18230), .A(n18217), .ZN(P3_U2788) );
  AOI22_X1 U21440 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18236), .ZN(n18218) );
  OAI21_X1 U21441 ( .B1(n18902), .B2(n18230), .A(n18218), .ZN(P3_U2789) );
  AOI22_X1 U21442 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18237), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n18228), .ZN(n18219) );
  OAI21_X1 U21443 ( .B1(n18220), .B2(n21354), .A(n18219), .ZN(P3_U2790) );
  AOI22_X1 U21444 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18236), .ZN(n18221) );
  OAI21_X1 U21445 ( .B1(n18222), .B2(n18230), .A(n18221), .ZN(P3_U2791) );
  AOI22_X1 U21446 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18236), .ZN(n18223) );
  OAI21_X1 U21447 ( .B1(n13579), .B2(n18230), .A(n18223), .ZN(P3_U2792) );
  AOI22_X1 U21448 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18236), .ZN(n18224) );
  OAI21_X1 U21449 ( .B1(n18225), .B2(n18230), .A(n18224), .ZN(P3_U2793) );
  AOI22_X1 U21450 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18237), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18236), .ZN(n18226) );
  OAI21_X1 U21451 ( .B1(n18227), .B2(n18239), .A(n18226), .ZN(P3_U2794) );
  AOI22_X1 U21452 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18236), .ZN(n18229) );
  OAI21_X1 U21453 ( .B1(n18231), .B2(n18230), .A(n18229), .ZN(P3_U2795) );
  AOI22_X1 U21454 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18237), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18236), .ZN(n18232) );
  OAI21_X1 U21455 ( .B1(n18233), .B2(n18239), .A(n18232), .ZN(P3_U2796) );
  AOI22_X1 U21456 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18237), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18236), .ZN(n18234) );
  OAI21_X1 U21457 ( .B1(n18235), .B2(n18239), .A(n18234), .ZN(P3_U2797) );
  AOI22_X1 U21458 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18237), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18236), .ZN(n18238) );
  OAI21_X1 U21459 ( .B1(n18240), .B2(n18239), .A(n18238), .ZN(P3_U2798) );
  OAI22_X1 U21460 ( .A1(n18242), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18660), .B2(n18241), .ZN(n18576) );
  AOI211_X1 U21461 ( .C1(n18243), .C2(n18245), .A(n18316), .B(n16752), .ZN(
        n18249) );
  NOR2_X1 U21462 ( .A1(n18748), .A2(n21348), .ZN(n18571) );
  OAI22_X1 U21463 ( .A1(n18246), .A2(n18245), .B1(n18402), .B2(n18244), .ZN(
        n18247) );
  AOI211_X1 U21464 ( .C1(n18249), .C2(n18248), .A(n18571), .B(n18247), .ZN(
        n18255) );
  INV_X1 U21465 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18567) );
  AOI221_X1 U21466 ( .B1(n16748), .B2(n18567), .C1(n18250), .C2(n18567), .A(
        n9686), .ZN(n18573) );
  NAND2_X1 U21467 ( .A1(n18252), .A2(n18251), .ZN(n18253) );
  XNOR2_X1 U21468 ( .A(n18253), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18572) );
  AOI22_X1 U21469 ( .A1(n18557), .A2(n18573), .B1(n18436), .B2(n18572), .ZN(
        n18254) );
  OAI211_X1 U21470 ( .C1(n18256), .C2(n18576), .A(n18255), .B(n18254), .ZN(
        P3_U2805) );
  AND2_X1 U21471 ( .A1(n18285), .A2(n18587), .ZN(n18271) );
  NAND2_X1 U21472 ( .A1(n18369), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18257) );
  OAI211_X1 U21473 ( .C1(n18258), .C2(n18271), .A(n18299), .B(n18257), .ZN(
        n18259) );
  XNOR2_X1 U21474 ( .A(n18259), .B(n18267), .ZN(n18583) );
  OAI221_X1 U21475 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19188), .C1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18261), .A(n18260), .ZN(
        n18262) );
  NAND2_X1 U21476 ( .A1(n18846), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18582) );
  OAI211_X1 U21477 ( .C1(n18264), .C2(n18263), .A(n18262), .B(n18582), .ZN(
        n18265) );
  AOI221_X1 U21478 ( .B1(n18268), .B2(n18267), .C1(n18266), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18265), .ZN(n18269) );
  OAI21_X1 U21479 ( .B1(n18464), .B2(n18583), .A(n18269), .ZN(P3_U2807) );
  INV_X1 U21480 ( .A(n18273), .ZN(n18593) );
  NOR2_X1 U21481 ( .A1(n18660), .A2(n18593), .ZN(n18270) );
  OAI21_X1 U21482 ( .B1(n18271), .B2(n18270), .A(n18299), .ZN(n18272) );
  XNOR2_X1 U21483 ( .A(n18272), .B(n18591), .ZN(n18599) );
  NOR2_X1 U21484 ( .A1(n18593), .A2(n18360), .ZN(n18283) );
  NOR2_X1 U21485 ( .A1(n18426), .A2(n18557), .ZN(n18308) );
  AOI22_X1 U21486 ( .A1(n18426), .A2(n18660), .B1(n18557), .B2(n18671), .ZN(
        n18359) );
  OAI21_X1 U21487 ( .B1(n18273), .B2(n18308), .A(n18359), .ZN(n18295) );
  OAI21_X1 U21488 ( .B1(n18275), .B2(n19360), .A(n18547), .ZN(n18276) );
  AOI21_X1 U21489 ( .B1(n18859), .B2(n18274), .A(n18276), .ZN(n18302) );
  OAI21_X1 U21490 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18277), .A(
        n18302), .ZN(n18291) );
  AOI22_X1 U21491 ( .A1(n18846), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18291), .ZN(n18280) );
  NOR2_X1 U21492 ( .A1(n18316), .A2(n18274), .ZN(n18293) );
  OAI211_X1 U21493 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18293), .B(n18278), .ZN(n18279) );
  OAI211_X1 U21494 ( .C1(n18281), .C2(n18402), .A(n18280), .B(n18279), .ZN(
        n18282) );
  AOI221_X1 U21495 ( .B1(n18283), .B2(n18591), .C1(n18295), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18282), .ZN(n18284) );
  OAI21_X1 U21496 ( .B1(n18464), .B2(n18599), .A(n18284), .ZN(P3_U2808) );
  INV_X1 U21497 ( .A(n18285), .ZN(n18287) );
  INV_X1 U21498 ( .A(n18606), .ZN(n18294) );
  NAND2_X1 U21499 ( .A1(n18367), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18333) );
  OAI22_X1 U21500 ( .A1(n18334), .A2(n18287), .B1(n18294), .B2(n18312), .ZN(
        n18288) );
  XNOR2_X1 U21501 ( .A(n18288), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18610) );
  OAI22_X1 U21502 ( .A1(n18748), .A2(n21391), .B1(n18402), .B2(n18289), .ZN(
        n18290) );
  AOI221_X1 U21503 ( .B1(n18293), .B2(n18292), .C1(n18291), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18290), .ZN(n18297) );
  NOR2_X1 U21504 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18294), .ZN(
        n18601) );
  NOR2_X1 U21505 ( .A1(n18600), .A2(n18360), .ZN(n18323) );
  AOI22_X1 U21506 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18295), .B1(
        n18601), .B2(n18323), .ZN(n18296) );
  OAI211_X1 U21507 ( .C1(n18610), .C2(n18464), .A(n18297), .B(n18296), .ZN(
        P3_U2809) );
  NAND2_X1 U21508 ( .A1(n18312), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18298) );
  OAI211_X1 U21509 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18329), .A(
        n18299), .B(n18298), .ZN(n18300) );
  XOR2_X1 U21510 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18300), .Z(
        n18619) );
  OR2_X1 U21511 ( .A1(n18906), .A2(n18301), .ZN(n18338) );
  AOI221_X1 U21512 ( .B1(n18304), .B2(n18303), .C1(n18338), .C2(n18303), .A(
        n18302), .ZN(n18307) );
  AOI21_X1 U21513 ( .B1(n18402), .B2(n18277), .A(n18305), .ZN(n18306) );
  AOI211_X1 U21514 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n18846), .A(n18307), 
        .B(n18306), .ZN(n18310) );
  NOR2_X1 U21515 ( .A1(n18600), .A2(n18620), .ZN(n18614) );
  OAI21_X1 U21516 ( .B1(n18308), .B2(n18614), .A(n18359), .ZN(n18322) );
  NOR2_X1 U21517 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18620), .ZN(
        n18611) );
  AOI22_X1 U21518 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18322), .B1(
        n18323), .B2(n18611), .ZN(n18309) );
  OAI211_X1 U21519 ( .C1(n18464), .C2(n18619), .A(n18310), .B(n18309), .ZN(
        P3_U2810) );
  INV_X1 U21520 ( .A(n18334), .ZN(n18311) );
  NAND2_X1 U21521 ( .A1(n18311), .A2(n18329), .ZN(n18332) );
  NAND2_X1 U21522 ( .A1(n18332), .A2(n18312), .ZN(n18313) );
  XOR2_X1 U21523 ( .A(n18620), .B(n18313), .Z(n18625) );
  INV_X1 U21524 ( .A(n11620), .ZN(n18315) );
  AOI21_X1 U21525 ( .B1(n18859), .B2(n18315), .A(n18530), .ZN(n18337) );
  OAI21_X1 U21526 ( .B1(n18314), .B2(n19360), .A(n18337), .ZN(n18327) );
  AOI22_X1 U21527 ( .A1(n18846), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18327), .ZN(n18319) );
  NOR2_X1 U21528 ( .A1(n18316), .A2(n18315), .ZN(n18328) );
  NAND2_X1 U21529 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18317) );
  OAI211_X1 U21530 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18328), .B(n18317), .ZN(n18318) );
  OAI211_X1 U21531 ( .C1(n18320), .C2(n18402), .A(n18319), .B(n18318), .ZN(
        n18321) );
  AOI221_X1 U21532 ( .B1(n18323), .B2(n18620), .C1(n18322), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n18321), .ZN(n18324) );
  OAI21_X1 U21533 ( .B1(n18625), .B2(n18464), .A(n18324), .ZN(P3_U2811) );
  NAND2_X1 U21534 ( .A1(n18631), .A2(n18635), .ZN(n18641) );
  NAND2_X1 U21535 ( .A1(n18846), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18639) );
  OAI21_X1 U21536 ( .B1(n18325), .B2(n18402), .A(n18639), .ZN(n18326) );
  AOI221_X1 U21537 ( .B1(n18328), .B2(n21318), .C1(n18327), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18326), .ZN(n18336) );
  OAI21_X1 U21538 ( .B1(n18631), .B2(n18360), .A(n18359), .ZN(n18345) );
  INV_X1 U21539 ( .A(n18329), .ZN(n18330) );
  NAND3_X1 U21540 ( .A1(n18334), .A2(n18330), .A3(n18333), .ZN(n18331) );
  OAI211_X1 U21541 ( .C1(n18334), .C2(n18333), .A(n18332), .B(n18331), .ZN(
        n18636) );
  AOI22_X1 U21542 ( .A1(n18345), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n18436), .B2(n18636), .ZN(n18335) );
  OAI211_X1 U21543 ( .C1(n18360), .C2(n18641), .A(n18336), .B(n18335), .ZN(
        P3_U2812) );
  INV_X1 U21544 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18642) );
  NAND2_X1 U21545 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18642), .ZN(
        n18648) );
  NOR2_X1 U21546 ( .A1(n18748), .A2(n19408), .ZN(n18645) );
  AOI21_X1 U21547 ( .B1(n18339), .B2(n18338), .A(n18337), .ZN(n18340) );
  AOI211_X1 U21548 ( .C1(n18341), .C2(n18558), .A(n18645), .B(n18340), .ZN(
        n18347) );
  AOI22_X1 U21549 ( .A1(n18342), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18631), .B2(n18660), .ZN(n18344) );
  NAND2_X1 U21550 ( .A1(n18344), .A2(n18343), .ZN(n18646) );
  AOI22_X1 U21551 ( .A1(n18345), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18436), .B2(n18646), .ZN(n18346) );
  OAI211_X1 U21552 ( .C1(n18360), .C2(n18648), .A(n18347), .B(n18346), .ZN(
        P3_U2813) );
  INV_X1 U21553 ( .A(n18660), .ZN(n18349) );
  OAI21_X1 U21554 ( .B1(n18349), .B2(n18369), .A(n18348), .ZN(n18350) );
  XNOR2_X1 U21555 ( .A(n18350), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18655) );
  NAND2_X1 U21556 ( .A1(n9734), .A2(n18398), .ZN(n18364) );
  OAI21_X1 U21557 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18351), .ZN(n18352) );
  OAI22_X1 U21558 ( .A1(n18402), .A2(n18353), .B1(n18364), .B2(n18352), .ZN(
        n18357) );
  OAI21_X1 U21559 ( .B1(n9734), .B2(n18519), .A(n18547), .ZN(n18383) );
  AOI21_X1 U21560 ( .B1(n18396), .B2(n18354), .A(n18383), .ZN(n18362) );
  OAI22_X1 U21561 ( .A1(n18362), .A2(n18355), .B1(n18748), .B2(n19406), .ZN(
        n18356) );
  AOI211_X1 U21562 ( .C1(n18436), .C2(n18655), .A(n18357), .B(n18356), .ZN(
        n18358) );
  OAI221_X1 U21563 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18360), 
        .C1(n18658), .C2(n18359), .A(n18358), .ZN(P3_U2814) );
  INV_X1 U21564 ( .A(n18663), .ZN(n18361) );
  NOR2_X1 U21565 ( .A1(n11633), .A2(n18361), .ZN(n18384) );
  NOR2_X1 U21566 ( .A1(n18384), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18667) );
  NAND2_X1 U21567 ( .A1(n18426), .A2(n18660), .ZN(n18378) );
  NAND2_X1 U21568 ( .A1(n18846), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18674) );
  OAI221_X1 U21569 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18364), .C1(
        n18363), .C2(n18362), .A(n18674), .ZN(n18365) );
  AOI21_X1 U21570 ( .B1(n18417), .B2(n18366), .A(n18365), .ZN(n18377) );
  NOR2_X1 U21571 ( .A1(n18368), .A2(n18367), .ZN(n18452) );
  AND2_X1 U21572 ( .A1(n18452), .A2(n18445), .ZN(n18433) );
  NAND2_X1 U21573 ( .A1(n18433), .A2(n11390), .ZN(n18412) );
  NOR2_X1 U21574 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18412), .ZN(
        n18389) );
  NOR2_X1 U21575 ( .A1(n11633), .A2(n18369), .ZN(n18451) );
  INV_X1 U21576 ( .A(n18677), .ZN(n18370) );
  AND2_X1 U21577 ( .A1(n18451), .A2(n18370), .ZN(n18406) );
  NAND2_X1 U21578 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n11388), .ZN(
        n18707) );
  OAI221_X1 U21579 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18389), 
        .C1(n18680), .C2(n18406), .A(n18707), .ZN(n18371) );
  XNOR2_X1 U21580 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18371), .ZN(
        n18668) );
  NOR2_X1 U21581 ( .A1(n18372), .A2(n18484), .ZN(n18375) );
  INV_X1 U21582 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18374) );
  NAND3_X1 U21583 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18386), .A3(
        n18373), .ZN(n18387) );
  NAND2_X1 U21584 ( .A1(n18374), .A2(n18387), .ZN(n18670) );
  AOI22_X1 U21585 ( .A1(n18436), .A2(n18668), .B1(n18375), .B2(n18670), .ZN(
        n18376) );
  OAI211_X1 U21586 ( .C1(n18667), .C2(n18378), .A(n18377), .B(n18376), .ZN(
        P3_U2815) );
  OAI21_X1 U21587 ( .B1(n18906), .B2(n18380), .A(n18379), .ZN(n18382) );
  AOI22_X1 U21588 ( .A1(n18383), .A2(n18382), .B1(n18381), .B2(n18558), .ZN(
        n18393) );
  AOI21_X1 U21589 ( .B1(n18724), .B2(n18386), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18385) );
  NOR2_X1 U21590 ( .A1(n18385), .A2(n18384), .ZN(n18691) );
  INV_X1 U21591 ( .A(n18386), .ZN(n18685) );
  NOR2_X1 U21592 ( .A1(n18721), .A2(n18685), .ZN(n18388) );
  OAI21_X1 U21593 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18388), .A(
        n18387), .ZN(n18689) );
  OAI21_X1 U21594 ( .B1(n18406), .B2(n18389), .A(n18707), .ZN(n18390) );
  XNOR2_X1 U21595 ( .A(n18390), .B(n18680), .ZN(n18688) );
  OAI22_X1 U21596 ( .A1(n18484), .A2(n18689), .B1(n18464), .B2(n18688), .ZN(
        n18391) );
  AOI21_X1 U21597 ( .B1(n18426), .B2(n18691), .A(n18391), .ZN(n18392) );
  OAI211_X1 U21598 ( .C1(n18748), .C2(n19402), .A(n18393), .B(n18392), .ZN(
        P3_U2816) );
  NAND2_X1 U21599 ( .A1(n18462), .A2(n18697), .ZN(n18424) );
  AOI22_X1 U21600 ( .A1(n18396), .A2(n18395), .B1(n18859), .B2(n18394), .ZN(
        n18397) );
  NAND2_X1 U21601 ( .A1(n18467), .A2(n18397), .ZN(n18418) );
  INV_X1 U21602 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18399) );
  NAND2_X1 U21603 ( .A1(n17471), .A2(n18398), .ZN(n18420) );
  AOI221_X1 U21604 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C1(n18400), .C2(n18399), .A(
        n18420), .ZN(n18404) );
  OAI22_X1 U21605 ( .A1(n18748), .A2(n19400), .B1(n18402), .B2(n18401), .ZN(
        n18403) );
  AOI211_X1 U21606 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18418), .A(
        n18404), .B(n18403), .ZN(n18411) );
  OR2_X1 U21607 ( .A1(n11633), .A2(n18677), .ZN(n18698) );
  NOR2_X1 U21608 ( .A1(n18721), .A2(n18677), .ZN(n18701) );
  NOR2_X1 U21609 ( .A1(n18484), .A2(n18701), .ZN(n18405) );
  AOI21_X1 U21610 ( .B1(n18426), .B2(n18698), .A(n18405), .ZN(n18423) );
  INV_X1 U21611 ( .A(n18423), .ZN(n18409) );
  INV_X1 U21612 ( .A(n18406), .ZN(n18407) );
  OAI21_X1 U21613 ( .B1(n18412), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18407), .ZN(n18408) );
  XNOR2_X1 U21614 ( .A(n18408), .B(n11388), .ZN(n18694) );
  AOI22_X1 U21615 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18409), .B1(
        n18436), .B2(n18694), .ZN(n18410) );
  OAI211_X1 U21616 ( .C1(n18707), .C2(n18424), .A(n18411), .B(n18410), .ZN(
        P3_U2817) );
  INV_X1 U21617 ( .A(n18697), .ZN(n18414) );
  INV_X1 U21618 ( .A(n18451), .ZN(n18413) );
  OAI21_X1 U21619 ( .B1(n18414), .B2(n18413), .A(n18412), .ZN(n18415) );
  XNOR2_X1 U21620 ( .A(n18415), .B(n11389), .ZN(n18714) );
  AOI22_X1 U21621 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18418), .B1(
        n18417), .B2(n18416), .ZN(n18419) );
  NAND2_X1 U21622 ( .A1(n18846), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18715) );
  OAI211_X1 U21623 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18420), .A(
        n18419), .B(n18715), .ZN(n18421) );
  AOI21_X1 U21624 ( .B1(n18436), .B2(n18714), .A(n18421), .ZN(n18422) );
  OAI221_X1 U21625 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18424), 
        .C1(n11389), .C2(n18423), .A(n18422), .ZN(P3_U2818) );
  INV_X1 U21626 ( .A(n18462), .ZN(n18425) );
  INV_X1 U21627 ( .A(n18727), .ZN(n18434) );
  NOR2_X1 U21628 ( .A1(n18425), .A2(n18434), .ZN(n18442) );
  NAND2_X1 U21629 ( .A1(n18426), .A2(n11633), .ZN(n18428) );
  NAND2_X1 U21630 ( .A1(n18721), .A2(n18557), .ZN(n18427) );
  NAND2_X1 U21631 ( .A1(n18428), .A2(n18427), .ZN(n18454) );
  NOR2_X1 U21632 ( .A1(n18442), .A2(n18454), .ZN(n18439) );
  NAND3_X1 U21633 ( .A1(n19188), .A2(n12900), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18466) );
  NOR2_X1 U21634 ( .A1(n18429), .A2(n18466), .ZN(n18450) );
  NOR2_X1 U21635 ( .A1(n18562), .A2(n18450), .ZN(n18441) );
  NOR2_X1 U21636 ( .A1(n18748), .A2(n19396), .ZN(n18719) );
  INV_X1 U21637 ( .A(n18450), .ZN(n18430) );
  OAI22_X1 U21638 ( .A1(n18264), .A2(n18431), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18430), .ZN(n18432) );
  AOI211_X1 U21639 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18441), .A(
        n18719), .B(n18432), .ZN(n18438) );
  NOR2_X1 U21640 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18727), .ZN(
        n18717) );
  AOI21_X1 U21641 ( .B1(n18451), .B2(n18434), .A(n18433), .ZN(n18435) );
  XNOR2_X1 U21642 ( .A(n18435), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18718) );
  AOI22_X1 U21643 ( .A1(n18462), .A2(n18717), .B1(n18436), .B2(n18718), .ZN(
        n18437) );
  OAI211_X1 U21644 ( .C1(n18439), .C2(n11390), .A(n18438), .B(n18437), .ZN(
        P3_U2819) );
  NOR2_X1 U21645 ( .A1(n18440), .A2(n18466), .ZN(n18456) );
  NAND2_X1 U21646 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18456), .ZN(
        n18455) );
  AOI22_X1 U21647 ( .A1(n18846), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18441), .ZN(n18449) );
  AOI21_X1 U21648 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18454), .A(
        n18442), .ZN(n18444) );
  INV_X1 U21649 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18741) );
  AOI22_X1 U21650 ( .A1(n18452), .A2(n18741), .B1(n18451), .B2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18443) );
  XOR2_X1 U21651 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18443), .Z(
        n18740) );
  OAI22_X1 U21652 ( .A1(n18445), .A2(n18444), .B1(n18740), .B2(n18464), .ZN(
        n18446) );
  AOI21_X1 U21653 ( .B1(n18447), .B2(n18558), .A(n18446), .ZN(n18448) );
  OAI211_X1 U21654 ( .C1(n18450), .C2(n18455), .A(n18449), .B(n18448), .ZN(
        P3_U2820) );
  NOR2_X1 U21655 ( .A1(n18452), .A2(n18451), .ZN(n18453) );
  XNOR2_X1 U21656 ( .A(n18453), .B(n18741), .ZN(n18754) );
  AND2_X1 U21657 ( .A1(n18454), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18461) );
  OAI211_X1 U21658 ( .C1(n18456), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n18478), .B(n18455), .ZN(n18458) );
  NAND2_X1 U21659 ( .A1(n18846), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18457) );
  OAI211_X1 U21660 ( .C1(n18264), .C2(n18459), .A(n18458), .B(n18457), .ZN(
        n18460) );
  AOI211_X1 U21661 ( .C1(n18741), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        n18463) );
  OAI21_X1 U21662 ( .B1(n18754), .B2(n18464), .A(n18463), .ZN(P3_U2821) );
  AOI22_X1 U21663 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18467), .B1(
        n18466), .B2(n18465), .ZN(n18468) );
  AOI21_X1 U21664 ( .B1(n18846), .B2(P3_REIP_REG_7__SCAN_IN), .A(n18468), .ZN(
        n18476) );
  NOR2_X1 U21665 ( .A1(n18470), .A2(n18469), .ZN(n18471) );
  XNOR2_X1 U21666 ( .A(n18471), .B(n18765), .ZN(n18783) );
  OAI21_X1 U21667 ( .B1(n18473), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18472), .ZN(n18474) );
  INV_X1 U21668 ( .A(n18474), .ZN(n18782) );
  AOI22_X1 U21669 ( .A1(n18557), .A2(n18783), .B1(n18515), .B2(n18782), .ZN(
        n18475) );
  OAI211_X1 U21670 ( .C1(n18264), .C2(n18477), .A(n18476), .B(n18475), .ZN(
        P3_U2823) );
  NAND2_X1 U21671 ( .A1(n19188), .A2(n12900), .ZN(n18485) );
  NAND2_X1 U21672 ( .A1(n18478), .A2(n18485), .ZN(n18506) );
  INV_X1 U21673 ( .A(n18481), .ZN(n18479) );
  AOI22_X1 U21674 ( .A1(n18481), .A2(n18497), .B1(n18480), .B2(n18479), .ZN(
        n18483) );
  XNOR2_X1 U21675 ( .A(n18483), .B(n18482), .ZN(n18795) );
  OAI22_X1 U21676 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18485), .B1(
        n18795), .B2(n18484), .ZN(n18486) );
  AOI21_X1 U21677 ( .B1(n18846), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18486), .ZN(
        n18493) );
  OAI21_X1 U21678 ( .B1(n18489), .B2(n18488), .A(n18487), .ZN(n18490) );
  INV_X1 U21679 ( .A(n18490), .ZN(n18792) );
  AOI22_X1 U21680 ( .A1(n18558), .A2(n18491), .B1(n18515), .B2(n18792), .ZN(
        n18492) );
  OAI211_X1 U21681 ( .C1(n18494), .C2(n18506), .A(n18493), .B(n18492), .ZN(
        P3_U2824) );
  OAI21_X1 U21682 ( .B1(n16636), .B2(n18530), .A(n18495), .ZN(n18496) );
  INV_X1 U21683 ( .A(n18496), .ZN(n18507) );
  AOI21_X1 U21684 ( .B1(n18499), .B2(n18498), .A(n18497), .ZN(n18796) );
  AOI22_X1 U21685 ( .A1(n18557), .A2(n18796), .B1(n18846), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18505) );
  OAI21_X1 U21686 ( .B1(n18501), .B2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n18500), .ZN(n18502) );
  INV_X1 U21687 ( .A(n18502), .ZN(n18797) );
  AOI22_X1 U21688 ( .A1(n18558), .A2(n18503), .B1(n18515), .B2(n18797), .ZN(
        n18504) );
  OAI211_X1 U21689 ( .C1(n18507), .C2(n18506), .A(n18505), .B(n18504), .ZN(
        P3_U2825) );
  OR2_X1 U21690 ( .A1(n18509), .A2(n18508), .ZN(n18510) );
  AND2_X1 U21691 ( .A1(n18511), .A2(n18510), .ZN(n18807) );
  INV_X1 U21692 ( .A(n18512), .ZN(n18513) );
  OAI22_X1 U21693 ( .A1(n18906), .A2(n18513), .B1(n19382), .B2(n18748), .ZN(
        n18514) );
  AOI21_X1 U21694 ( .B1(n18515), .B2(n18807), .A(n18514), .ZN(n18521) );
  AOI21_X1 U21695 ( .B1(n18518), .B2(n18517), .A(n18516), .ZN(n18803) );
  OAI21_X1 U21696 ( .B1(n16634), .B2(n18519), .A(n18547), .ZN(n18532) );
  AOI22_X1 U21697 ( .A1(n18557), .A2(n18803), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18532), .ZN(n18520) );
  OAI211_X1 U21698 ( .C1(n18264), .C2(n18522), .A(n18521), .B(n18520), .ZN(
        P3_U2826) );
  OR2_X1 U21699 ( .A1(n18524), .A2(n18523), .ZN(n18525) );
  NAND2_X1 U21700 ( .A1(n18526), .A2(n18525), .ZN(n18815) );
  OAI22_X1 U21701 ( .A1(n18552), .A2(n18815), .B1(n18748), .B2(n19380), .ZN(
        n18527) );
  INV_X1 U21702 ( .A(n18527), .ZN(n18534) );
  AOI21_X1 U21703 ( .B1(n18529), .B2(n18528), .A(n9757), .ZN(n18817) );
  OAI21_X1 U21704 ( .B1(n18530), .B2(n18548), .A(n16652), .ZN(n18531) );
  AOI22_X1 U21705 ( .A1(n18557), .A2(n18817), .B1(n18532), .B2(n18531), .ZN(
        n18533) );
  OAI211_X1 U21706 ( .C1(n18264), .C2(n18535), .A(n18534), .B(n18533), .ZN(
        P3_U2827) );
  AOI21_X1 U21707 ( .B1(n18538), .B2(n18537), .A(n18536), .ZN(n18831) );
  OAI21_X1 U21708 ( .B1(n18541), .B2(n18540), .A(n18539), .ZN(n18822) );
  NOR2_X1 U21709 ( .A1(n18748), .A2(n19377), .ZN(n18836) );
  INV_X1 U21710 ( .A(n18836), .ZN(n18542) );
  OAI21_X1 U21711 ( .B1(n18552), .B2(n18822), .A(n18542), .ZN(n18545) );
  NOR2_X1 U21712 ( .A1(n18264), .A2(n18543), .ZN(n18544) );
  AOI211_X1 U21713 ( .C1(n18557), .C2(n18831), .A(n18545), .B(n18544), .ZN(
        n18546) );
  OAI221_X1 U21714 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18906), .C1(
        n18548), .C2(n18547), .A(n18546), .ZN(P3_U2828) );
  OAI21_X1 U21715 ( .B1(n18550), .B2(n10308), .A(n18549), .ZN(n18841) );
  INV_X1 U21716 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18551) );
  OAI22_X1 U21717 ( .A1(n18552), .A2(n18841), .B1(n18748), .B2(n18551), .ZN(
        n18553) );
  INV_X1 U21718 ( .A(n18553), .ZN(n18560) );
  OAI21_X1 U21719 ( .B1(n18556), .B2(n18555), .A(n18554), .ZN(n18844) );
  AOI22_X1 U21720 ( .A1(n18558), .A2(n18561), .B1(n18557), .B2(n18844), .ZN(
        n18559) );
  OAI211_X1 U21721 ( .C1(n18562), .C2(n18561), .A(n18560), .B(n18559), .ZN(
        P3_U2829) );
  INV_X1 U21722 ( .A(n18757), .ZN(n18577) );
  INV_X1 U21723 ( .A(n18563), .ZN(n18566) );
  AOI221_X1 U21724 ( .B1(n18566), .B2(n19300), .C1(n18565), .C2(n19300), .A(
        n18564), .ZN(n18569) );
  AOI221_X1 U21725 ( .B1(n18569), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n18568), .C2(n18567), .A(n18834), .ZN(n18570) );
  AOI211_X1 U21726 ( .C1(n18848), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18571), .B(n18570), .ZN(n18575) );
  AOI22_X1 U21727 ( .A1(n18845), .A2(n18573), .B1(n18760), .B2(n18572), .ZN(
        n18574) );
  OAI211_X1 U21728 ( .C1(n18577), .C2(n18576), .A(n18575), .B(n18574), .ZN(
        P3_U2837) );
  NOR2_X1 U21729 ( .A1(n18848), .A2(n18578), .ZN(n18580) );
  OAI21_X1 U21730 ( .B1(n18580), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18579), .ZN(n18581) );
  OAI211_X1 U21731 ( .C1(n18583), .C2(n18753), .A(n18582), .B(n18581), .ZN(
        P3_U2839) );
  AOI22_X1 U21732 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18848), .B1(
        n18846), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n18598) );
  AOI22_X1 U21733 ( .A1(n19298), .A2(n18671), .B1(n18661), .B2(n18660), .ZN(
        n18603) );
  NAND2_X1 U21734 ( .A1(n18700), .A2(n18723), .ZN(n18726) );
  AOI21_X1 U21735 ( .B1(n18626), .B2(n18614), .A(n18585), .ZN(n18584) );
  AOI221_X1 U21736 ( .B1(n18600), .B2(n19300), .C1(n18628), .C2(n19300), .A(
        n18584), .ZN(n18613) );
  OAI21_X1 U21737 ( .B1(n18585), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n18613), .ZN(n18586) );
  AOI21_X1 U21738 ( .B1(n18593), .B2(n18726), .A(n18586), .ZN(n18605) );
  AOI22_X1 U21739 ( .A1(n19300), .A2(n18588), .B1(n18851), .B2(n18587), .ZN(
        n18589) );
  NAND4_X1 U21740 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18603), .A3(
        n18605), .A4(n18589), .ZN(n18595) );
  INV_X1 U21741 ( .A(n18590), .ZN(n18592) );
  OAI21_X1 U21742 ( .B1(n18593), .B2(n18592), .A(n18591), .ZN(n18594) );
  OAI211_X1 U21743 ( .C1(n18596), .C2(n18595), .A(n18813), .B(n18594), .ZN(
        n18597) );
  OAI211_X1 U21744 ( .C1(n18599), .C2(n18753), .A(n18598), .B(n18597), .ZN(
        P3_U2840) );
  NOR2_X1 U21745 ( .A1(n18600), .A2(n18659), .ZN(n18621) );
  AOI22_X1 U21746 ( .A1(n18846), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18601), 
        .B2(n18621), .ZN(n18609) );
  AOI21_X1 U21747 ( .B1(n18602), .B2(n18649), .A(n18746), .ZN(n18604) );
  NAND2_X1 U21748 ( .A1(n18813), .A2(n18603), .ZN(n18654) );
  NOR2_X1 U21749 ( .A1(n18604), .A2(n18654), .ZN(n18612) );
  OAI211_X1 U21750 ( .C1(n18606), .C2(n18681), .A(n18605), .B(n18612), .ZN(
        n18607) );
  NAND3_X1 U21751 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18748), .A3(
        n18607), .ZN(n18608) );
  OAI211_X1 U21752 ( .C1(n18610), .C2(n18753), .A(n18609), .B(n18608), .ZN(
        P3_U2841) );
  AOI22_X1 U21753 ( .A1(n18846), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18621), 
        .B2(n18611), .ZN(n18618) );
  INV_X1 U21754 ( .A(n18726), .ZN(n18630) );
  OAI211_X1 U21755 ( .C1(n18614), .C2(n18630), .A(n18613), .B(n18612), .ZN(
        n18615) );
  NOR3_X1 U21756 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18681), .A3(
        n19472), .ZN(n18616) );
  OAI21_X1 U21757 ( .B1(n18622), .B2(n18616), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18617) );
  OAI211_X1 U21758 ( .C1(n18619), .C2(n18753), .A(n18618), .B(n18617), .ZN(
        P3_U2842) );
  AOI22_X1 U21759 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18622), .B1(
        n18621), .B2(n18620), .ZN(n18624) );
  NAND2_X1 U21760 ( .A1(n18846), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18623) );
  OAI211_X1 U21761 ( .C1(n18625), .C2(n18753), .A(n18624), .B(n18623), .ZN(
        P3_U2843) );
  NAND3_X1 U21762 ( .A1(n18626), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18769), .ZN(n18633) );
  NOR2_X1 U21763 ( .A1(n18628), .A2(n18627), .ZN(n18629) );
  OAI22_X1 U21764 ( .A1(n18631), .A2(n18630), .B1(n18629), .B2(n18766), .ZN(
        n18632) );
  AOI211_X1 U21765 ( .C1(n18634), .C2(n18633), .A(n18632), .B(n18654), .ZN(
        n18643) );
  OAI21_X1 U21766 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18767), .A(
        n18643), .ZN(n18638) );
  NOR2_X1 U21767 ( .A1(n18846), .A2(n18635), .ZN(n18637) );
  AOI22_X1 U21768 ( .A1(n18638), .A2(n18637), .B1(n18760), .B2(n18636), .ZN(
        n18640) );
  OAI211_X1 U21769 ( .C1(n18659), .C2(n18641), .A(n18640), .B(n18639), .ZN(
        P3_U2844) );
  NOR3_X1 U21770 ( .A1(n18643), .A2(n18846), .A3(n18642), .ZN(n18644) );
  AOI211_X1 U21771 ( .C1(n18760), .C2(n18646), .A(n18645), .B(n18644), .ZN(
        n18647) );
  OAI21_X1 U21772 ( .B1(n18659), .B2(n18648), .A(n18647), .ZN(P3_U2845) );
  OAI21_X1 U21773 ( .B1(n18776), .B2(n18743), .A(n18851), .ZN(n18735) );
  NAND2_X1 U21774 ( .A1(n18663), .A2(n18735), .ZN(n18679) );
  AOI21_X1 U21775 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18746), .A(
        n18649), .ZN(n18651) );
  NOR2_X1 U21776 ( .A1(n18650), .A2(n18766), .ZN(n18720) );
  AOI211_X1 U21777 ( .C1(n18652), .C2(n18679), .A(n18651), .B(n18720), .ZN(
        n18665) );
  NOR2_X1 U21778 ( .A1(n18773), .A2(n18665), .ZN(n18653) );
  OAI21_X1 U21779 ( .B1(n18654), .B2(n18653), .A(n18748), .ZN(n18657) );
  AOI22_X1 U21780 ( .A1(n18846), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18760), 
        .B2(n18655), .ZN(n18656) );
  OAI221_X1 U21781 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18659), 
        .C1(n18658), .C2(n18657), .A(n18656), .ZN(P3_U2846) );
  NAND2_X1 U21782 ( .A1(n18661), .A2(n18660), .ZN(n18666) );
  INV_X1 U21783 ( .A(n18684), .ZN(n18662) );
  AOI21_X1 U21784 ( .B1(n18663), .B2(n18662), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18664) );
  OAI22_X1 U21785 ( .A1(n18667), .A2(n18666), .B1(n18665), .B2(n18664), .ZN(
        n18669) );
  AOI22_X1 U21786 ( .A1(n18813), .A2(n18669), .B1(n18760), .B2(n18668), .ZN(
        n18675) );
  NAND3_X1 U21787 ( .A1(n18845), .A2(n18671), .A3(n18670), .ZN(n18673) );
  NAND2_X1 U21788 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18848), .ZN(
        n18672) );
  NAND4_X1 U21789 ( .A1(n18675), .A2(n18674), .A3(n18673), .A4(n18672), .ZN(
        P3_U2847) );
  NOR2_X1 U21790 ( .A1(n18677), .A2(n18676), .ZN(n18710) );
  NOR2_X1 U21791 ( .A1(n18746), .A2(n18710), .ZN(n18704) );
  NOR3_X1 U21792 ( .A1(n18704), .A2(n18678), .A3(n18685), .ZN(n18683) );
  OAI21_X1 U21793 ( .B1(n18680), .B2(n18851), .A(n18679), .ZN(n18682) );
  AOI221_X1 U21794 ( .B1(n18683), .B2(n18682), .C1(n18681), .C2(n18682), .A(
        n18834), .ZN(n18687) );
  NOR2_X1 U21795 ( .A1(n18685), .A2(n18684), .ZN(n18686) );
  AOI222_X1 U21796 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18687), 
        .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18848), .C1(n18687), 
        .C2(n18686), .ZN(n18693) );
  OAI22_X1 U21797 ( .A1(n18833), .A2(n18689), .B1(n18753), .B2(n18688), .ZN(
        n18690) );
  AOI21_X1 U21798 ( .B1(n18757), .B2(n18691), .A(n18690), .ZN(n18692) );
  OAI211_X1 U21799 ( .C1(n18748), .C2(n19402), .A(n18693), .B(n18692), .ZN(
        P3_U2848) );
  NAND2_X1 U21800 ( .A1(n18697), .A2(n18742), .ZN(n18711) );
  AOI22_X1 U21801 ( .A1(n18846), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18760), 
        .B2(n18694), .ZN(n18706) );
  AOI21_X1 U21802 ( .B1(n18851), .B2(n11390), .A(n11389), .ZN(n18709) );
  OAI21_X1 U21803 ( .B1(n18727), .B2(n18695), .A(n18851), .ZN(n18696) );
  OAI21_X1 U21804 ( .B1(n18697), .B2(n18766), .A(n18696), .ZN(n18729) );
  INV_X1 U21805 ( .A(n18698), .ZN(n18699) );
  OAI22_X1 U21806 ( .A1(n18701), .A2(n18700), .B1(n18723), .B2(n18699), .ZN(
        n18702) );
  NOR3_X1 U21807 ( .A1(n18720), .A2(n18729), .A3(n18702), .ZN(n18708) );
  OAI211_X1 U21808 ( .C1(n18736), .C2(n18709), .A(n18813), .B(n18708), .ZN(
        n18703) );
  OAI211_X1 U21809 ( .C1(n18704), .C2(n18703), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18748), .ZN(n18705) );
  OAI211_X1 U21810 ( .C1(n18707), .C2(n18711), .A(n18706), .B(n18705), .ZN(
        P3_U2849) );
  OAI211_X1 U21811 ( .C1(n18710), .C2(n18746), .A(n18709), .B(n18708), .ZN(
        n18713) );
  OAI21_X1 U21812 ( .B1(n18834), .B2(n11389), .A(n18711), .ZN(n18712) );
  AOI22_X1 U21813 ( .A1(n18760), .A2(n18714), .B1(n18713), .B2(n18712), .ZN(
        n18716) );
  OAI211_X1 U21814 ( .C1(n18839), .C2(n11389), .A(n18716), .B(n18715), .ZN(
        P3_U2850) );
  AOI22_X1 U21815 ( .A1(n18760), .A2(n18718), .B1(n18742), .B2(n18717), .ZN(
        n18732) );
  INV_X1 U21816 ( .A(n18719), .ZN(n18731) );
  AOI21_X1 U21817 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18747), .A(
        n18746), .ZN(n18725) );
  AOI211_X1 U21818 ( .C1(n18721), .C2(n19298), .A(n18720), .B(n18834), .ZN(
        n18722) );
  OAI21_X1 U21819 ( .B1(n18724), .B2(n18723), .A(n18722), .ZN(n18750) );
  AOI211_X1 U21820 ( .C1(n18727), .C2(n18726), .A(n18725), .B(n18750), .ZN(
        n18734) );
  OAI21_X1 U21821 ( .B1(n18746), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18734), .ZN(n18728) );
  OAI211_X1 U21822 ( .C1(n18729), .C2(n18728), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18748), .ZN(n18730) );
  NAND3_X1 U21823 ( .A1(n18732), .A2(n18731), .A3(n18730), .ZN(P3_U2851) );
  NOR2_X1 U21824 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18741), .ZN(
        n18733) );
  AOI22_X1 U21825 ( .A1(n18846), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18742), 
        .B2(n18733), .ZN(n18739) );
  OAI211_X1 U21826 ( .C1(n18736), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18735), .B(n18734), .ZN(n18737) );
  NAND3_X1 U21827 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18748), .A3(
        n18737), .ZN(n18738) );
  OAI211_X1 U21828 ( .C1(n18740), .C2(n18753), .A(n18739), .B(n18738), .ZN(
        P3_U2852) );
  AOI22_X1 U21829 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18846), .B1(n18742), 
        .B2(n18741), .ZN(n18752) );
  NAND2_X1 U21830 ( .A1(n18851), .A2(n18776), .ZN(n18745) );
  NAND2_X1 U21831 ( .A1(n18851), .A2(n18743), .ZN(n18744) );
  OAI211_X1 U21832 ( .C1(n18747), .C2(n18746), .A(n18745), .B(n18744), .ZN(
        n18749) );
  OAI211_X1 U21833 ( .C1(n18750), .C2(n18749), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18748), .ZN(n18751) );
  OAI211_X1 U21834 ( .C1(n18754), .C2(n18753), .A(n18752), .B(n18751), .ZN(
        P3_U2853) );
  INV_X1 U21835 ( .A(n18755), .ZN(n18756) );
  NAND2_X1 U21836 ( .A1(n18757), .A2(n18756), .ZN(n18762) );
  INV_X1 U21837 ( .A(n18758), .ZN(n18759) );
  NAND2_X1 U21838 ( .A1(n18760), .A2(n18759), .ZN(n18761) );
  OAI211_X1 U21839 ( .C1(n18763), .C2(n18833), .A(n18762), .B(n18761), .ZN(
        n18764) );
  INV_X1 U21840 ( .A(n18764), .ZN(n18781) );
  NOR2_X1 U21841 ( .A1(n11379), .A2(n18765), .ZN(n18772) );
  OR2_X1 U21842 ( .A1(n18766), .A2(n18775), .ZN(n18824) );
  AOI21_X1 U21843 ( .B1(n18769), .B2(n18768), .A(n18767), .ZN(n18770) );
  INV_X1 U21844 ( .A(n18770), .ZN(n18826) );
  NAND2_X1 U21845 ( .A1(n18824), .A2(n18826), .ZN(n18804) );
  AOI21_X1 U21846 ( .B1(n18771), .B2(n18789), .A(n18804), .ZN(n18791) );
  OAI21_X1 U21847 ( .B1(n18773), .B2(n18772), .A(n18791), .ZN(n18784) );
  OAI221_X1 U21848 ( .B1(n18848), .B2(n18850), .C1(n18848), .C2(n18784), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18779) );
  NAND2_X1 U21849 ( .A1(n18775), .A2(n18774), .ZN(n18812) );
  NOR2_X1 U21850 ( .A1(n18834), .A2(n18812), .ZN(n18802) );
  NAND3_X1 U21851 ( .A1(n18777), .A2(n18802), .A3(n18776), .ZN(n18778) );
  NAND4_X1 U21852 ( .A1(n18781), .A2(n18780), .A3(n18779), .A4(n18778), .ZN(
        P3_U2854) );
  AOI22_X1 U21853 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18848), .B1(
        n18846), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18788) );
  AOI22_X1 U21854 ( .A1(n18845), .A2(n18783), .B1(n18843), .B2(n18782), .ZN(
        n18787) );
  NOR3_X1 U21855 ( .A1(n11379), .A2(n18789), .A3(n18812), .ZN(n18785) );
  OAI211_X1 U21856 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18785), .A(
        n18813), .B(n18784), .ZN(n18786) );
  NAND3_X1 U21857 ( .A1(n18788), .A2(n18787), .A3(n18786), .ZN(P3_U2855) );
  NOR2_X1 U21858 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18789), .ZN(
        n18790) );
  AOI22_X1 U21859 ( .A1(n18846), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18802), 
        .B2(n18790), .ZN(n18794) );
  OAI21_X1 U21860 ( .B1(n18791), .B2(n18846), .A(n18839), .ZN(n18798) );
  AOI22_X1 U21861 ( .A1(n18798), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18843), .B2(n18792), .ZN(n18793) );
  OAI211_X1 U21862 ( .C1(n18795), .C2(n18833), .A(n18794), .B(n18793), .ZN(
        P3_U2856) );
  AOI22_X1 U21863 ( .A1(n18846), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18845), 
        .B2(n18796), .ZN(n18801) );
  AOI22_X1 U21864 ( .A1(n18798), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n18843), .B2(n18797), .ZN(n18800) );
  NAND4_X1 U21865 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18802), .A4(n9918), .ZN(
        n18799) );
  NAND3_X1 U21866 ( .A1(n18801), .A2(n18800), .A3(n18799), .ZN(P3_U2857) );
  NAND2_X1 U21867 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18802), .ZN(
        n18811) );
  AOI22_X1 U21868 ( .A1(n18846), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18845), 
        .B2(n18803), .ZN(n18810) );
  NOR2_X1 U21869 ( .A1(n18805), .A2(n18804), .ZN(n18821) );
  OAI21_X1 U21870 ( .B1(n18821), .B2(n18806), .A(n18839), .ZN(n18808) );
  AOI22_X1 U21871 ( .A1(n18808), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n18843), .B2(n18807), .ZN(n18809) );
  OAI211_X1 U21872 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18811), .A(
        n18810), .B(n18809), .ZN(P3_U2858) );
  INV_X1 U21873 ( .A(n18812), .ZN(n18814) );
  OAI21_X1 U21874 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18814), .A(
        n18813), .ZN(n18820) );
  AOI22_X1 U21875 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18848), .B1(
        n18846), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18819) );
  INV_X1 U21876 ( .A(n18815), .ZN(n18816) );
  AOI22_X1 U21877 ( .A1(n18845), .A2(n18817), .B1(n18843), .B2(n18816), .ZN(
        n18818) );
  OAI211_X1 U21878 ( .C1(n18821), .C2(n18820), .A(n18819), .B(n18818), .ZN(
        P3_U2859) );
  INV_X1 U21879 ( .A(n18822), .ZN(n18830) );
  NOR3_X1 U21880 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18849), .A3(
        n18823), .ZN(n18828) );
  NAND3_X1 U21881 ( .A1(n19300), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18825) );
  OAI221_X1 U21882 ( .B1(n18840), .B2(n18826), .C1(n18840), .C2(n18825), .A(
        n18824), .ZN(n18827) );
  AOI211_X1 U21883 ( .C1(n18830), .C2(n18829), .A(n18828), .B(n18827), .ZN(
        n18835) );
  INV_X1 U21884 ( .A(n18831), .ZN(n18832) );
  OAI22_X1 U21885 ( .A1(n18835), .A2(n18834), .B1(n18833), .B2(n18832), .ZN(
        n18837) );
  NOR2_X1 U21886 ( .A1(n18837), .A2(n18836), .ZN(n18838) );
  OAI21_X1 U21887 ( .B1(n18840), .B2(n18839), .A(n18838), .ZN(P3_U2860) );
  INV_X1 U21888 ( .A(n18841), .ZN(n18842) );
  AOI22_X1 U21889 ( .A1(n18845), .A2(n18844), .B1(n18843), .B2(n18842), .ZN(
        n18855) );
  NAND2_X1 U21890 ( .A1(n18846), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18854) );
  OAI21_X1 U21891 ( .B1(n18848), .B2(n18847), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18853) );
  OAI211_X1 U21892 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18851), .A(
        n18850), .B(n18849), .ZN(n18852) );
  NAND4_X1 U21893 ( .A1(n18855), .A2(n18854), .A3(n18853), .A4(n18852), .ZN(
        P3_U2861) );
  NAND2_X1 U21894 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18856) );
  AOI21_X1 U21895 ( .B1(n18857), .B2(n17258), .A(n18856), .ZN(n19340) );
  OAI21_X1 U21896 ( .B1(n19340), .B2(n18915), .A(n18863), .ZN(n18858) );
  OAI221_X1 U21897 ( .B1(n11545), .B2(n19468), .C1(n11545), .C2(n18863), .A(
        n18858), .ZN(P3_U2863) );
  NAND2_X1 U21898 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19244) );
  NOR2_X1 U21899 ( .A1(n19468), .A2(n18859), .ZN(n18862) );
  INV_X1 U21900 ( .A(n18860), .ZN(n18861) );
  AOI221_X1 U21901 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19244), .C1(n18862), 
        .C2(n19244), .A(n18861), .ZN(n18868) );
  OAI221_X1 U21902 ( .B1(n19159), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19159), .C2(n18864), .A(n18863), .ZN(n18866) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18868), .B1(
        n18866), .B2(n18865), .ZN(P3_U2865) );
  NOR2_X1 U21904 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19326), .ZN(
        n19158) );
  NOR2_X1 U21905 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18865), .ZN(
        n19046) );
  NOR2_X1 U21906 ( .A1(n19158), .A2(n19046), .ZN(n18867) );
  OAI22_X1 U21907 ( .A1(n18868), .A2(n19326), .B1(n18867), .B2(n18866), .ZN(
        P3_U2866) );
  AND2_X1 U21908 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18869), .ZN(
        P3_U2867) );
  NAND2_X1 U21909 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19212) );
  NAND2_X1 U21910 ( .A1(n19311), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19091) );
  NOR2_X2 U21911 ( .A1(n19212), .A2(n19091), .ZN(n21306) );
  INV_X1 U21912 ( .A(n21306), .ZN(n19292) );
  NAND2_X1 U21913 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19188), .ZN(n19221) );
  NOR2_X1 U21914 ( .A1(n18906), .A2(n18870), .ZN(n19213) );
  NAND2_X1 U21915 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n11545), .ZN(
        n19112) );
  NOR2_X2 U21916 ( .A1(n19212), .A2(n19112), .ZN(n19240) );
  NOR2_X2 U21917 ( .A1(n18914), .A2(n18871), .ZN(n19245) );
  NOR2_X1 U21918 ( .A1(n19311), .A2(n11545), .ZN(n19309) );
  INV_X1 U21919 ( .A(n19212), .ZN(n19186) );
  NAND2_X1 U21920 ( .A1(n19309), .A2(n19186), .ZN(n21309) );
  NOR2_X1 U21921 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19156) );
  NOR2_X1 U21922 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18956) );
  NAND2_X1 U21923 ( .A1(n19156), .A2(n18956), .ZN(n18969) );
  INV_X1 U21924 ( .A(n19350), .ZN(n19163) );
  AOI21_X1 U21925 ( .B1(n21309), .B2(n18969), .A(n19163), .ZN(n18908) );
  AOI22_X1 U21926 ( .A1(n19213), .A2(n19240), .B1(n19245), .B2(n18908), .ZN(
        n18875) );
  NOR2_X1 U21927 ( .A1(n18906), .A2(n19212), .ZN(n19247) );
  NAND2_X1 U21928 ( .A1(n19091), .A2(n19112), .ZN(n19157) );
  AOI21_X1 U21929 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18914), .ZN(n18935) );
  INV_X1 U21930 ( .A(n18935), .ZN(n19022) );
  AOI21_X1 U21931 ( .B1(n21309), .B2(n18969), .A(n19022), .ZN(n18936) );
  AOI21_X1 U21932 ( .B1(n19247), .B2(n19157), .A(n18936), .ZN(n18911) );
  INV_X1 U21933 ( .A(n18969), .ZN(n18973) );
  NAND2_X1 U21934 ( .A1(n18872), .A2(n19449), .ZN(n18909) );
  NOR2_X2 U21935 ( .A1(n18873), .A2(n18909), .ZN(n19250) );
  AOI22_X1 U21936 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18911), .B1(
        n18973), .B2(n19250), .ZN(n18874) );
  OAI211_X1 U21937 ( .C1(n19292), .C2(n19221), .A(n18875), .B(n18874), .ZN(
        P3_U2868) );
  INV_X1 U21938 ( .A(n18909), .ZN(n18900) );
  NAND2_X1 U21939 ( .A1(n18900), .A2(n19471), .ZN(n19259) );
  NOR2_X2 U21940 ( .A1(n18876), .A2(n18906), .ZN(n19255) );
  NOR2_X2 U21941 ( .A1(n18914), .A2(n13926), .ZN(n19254) );
  AOI22_X1 U21942 ( .A1(n21306), .A2(n19255), .B1(n18908), .B2(n19254), .ZN(
        n18879) );
  NOR2_X2 U21943 ( .A1(n18906), .A2(n18877), .ZN(n19256) );
  AOI22_X1 U21944 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18911), .B1(
        n19240), .B2(n19256), .ZN(n18878) );
  OAI211_X1 U21945 ( .C1(n18969), .C2(n19259), .A(n18879), .B(n18878), .ZN(
        P3_U2869) );
  NAND2_X1 U21946 ( .A1(n18900), .A2(n18880), .ZN(n21310) );
  NAND2_X1 U21947 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19188), .ZN(n21311) );
  NOR2_X2 U21948 ( .A1(n18914), .A2(n18881), .ZN(n21304) );
  AOI22_X1 U21949 ( .A1(n19224), .A2(n21306), .B1(n21304), .B2(n18908), .ZN(
        n18884) );
  NOR2_X2 U21950 ( .A1(n18906), .A2(n18882), .ZN(n21307) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18911), .B1(
        n21307), .B2(n19240), .ZN(n18883) );
  OAI211_X1 U21952 ( .C1(n21310), .C2(n18969), .A(n18884), .B(n18883), .ZN(
        P3_U2870) );
  NAND2_X1 U21953 ( .A1(n18900), .A2(n18885), .ZN(n19265) );
  NOR2_X2 U21954 ( .A1(n21324), .A2(n18906), .ZN(n19262) );
  NOR2_X2 U21955 ( .A1(n18914), .A2(n13585), .ZN(n19260) );
  AOI22_X1 U21956 ( .A1(n21306), .A2(n19262), .B1(n18908), .B2(n19260), .ZN(
        n18888) );
  NOR2_X2 U21957 ( .A1(n18906), .A2(n18886), .ZN(n19261) );
  AOI22_X1 U21958 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18911), .B1(
        n19240), .B2(n19261), .ZN(n18887) );
  OAI211_X1 U21959 ( .C1(n18969), .C2(n19265), .A(n18888), .B(n18887), .ZN(
        P3_U2871) );
  NAND2_X1 U21960 ( .A1(n18900), .A2(n18889), .ZN(n19271) );
  NOR2_X2 U21961 ( .A1(n18890), .A2(n18906), .ZN(n19267) );
  NOR2_X2 U21962 ( .A1(n18914), .A2(n18891), .ZN(n19266) );
  AOI22_X1 U21963 ( .A1(n21306), .A2(n19267), .B1(n18908), .B2(n19266), .ZN(
        n18894) );
  NOR2_X2 U21964 ( .A1(n18906), .A2(n18892), .ZN(n19268) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18911), .B1(
        n19240), .B2(n19268), .ZN(n18893) );
  OAI211_X1 U21966 ( .C1(n18969), .C2(n19271), .A(n18894), .B(n18893), .ZN(
        P3_U2872) );
  NAND2_X1 U21967 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19188), .ZN(n19277) );
  NOR2_X1 U21968 ( .A1(n18895), .A2(n18906), .ZN(n19273) );
  NOR2_X2 U21969 ( .A1(n13582), .A2(n18914), .ZN(n19272) );
  AOI22_X1 U21970 ( .A1(n19240), .A2(n19273), .B1(n18908), .B2(n19272), .ZN(
        n18898) );
  NOR2_X2 U21971 ( .A1(n18896), .A2(n18909), .ZN(n19274) );
  AOI22_X1 U21972 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18911), .B1(
        n18973), .B2(n19274), .ZN(n18897) );
  OAI211_X1 U21973 ( .C1(n19292), .C2(n19277), .A(n18898), .B(n18897), .ZN(
        P3_U2873) );
  NAND2_X1 U21974 ( .A1(n18900), .A2(n18899), .ZN(n19283) );
  NOR2_X2 U21975 ( .A1(n18901), .A2(n18906), .ZN(n19280) );
  NOR2_X2 U21976 ( .A1(n18902), .A2(n18914), .ZN(n19278) );
  AOI22_X1 U21977 ( .A1(n21306), .A2(n19280), .B1(n18908), .B2(n19278), .ZN(
        n18905) );
  NOR2_X2 U21978 ( .A1(n18903), .A2(n18906), .ZN(n19279) );
  AOI22_X1 U21979 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18911), .B1(
        n19240), .B2(n19279), .ZN(n18904) );
  OAI211_X1 U21980 ( .C1(n18969), .C2(n19283), .A(n18905), .B(n18904), .ZN(
        P3_U2874) );
  NAND2_X1 U21981 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n19188), .ZN(n19210) );
  NOR2_X1 U21982 ( .A1(n18907), .A2(n18906), .ZN(n19205) );
  NOR2_X2 U21983 ( .A1(n13588), .A2(n18914), .ZN(n19284) );
  AOI22_X1 U21984 ( .A1(n19240), .A2(n19205), .B1(n18908), .B2(n19284), .ZN(
        n18913) );
  NOR2_X2 U21985 ( .A1(n18910), .A2(n18909), .ZN(n19287) );
  AOI22_X1 U21986 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18911), .B1(
        n18973), .B2(n19287), .ZN(n18912) );
  OAI211_X1 U21987 ( .C1(n19292), .C2(n19210), .A(n18913), .B(n18912), .ZN(
        P3_U2875) );
  INV_X1 U21988 ( .A(n19213), .ZN(n19253) );
  INV_X1 U21989 ( .A(n19221), .ZN(n19246) );
  INV_X1 U21990 ( .A(n18956), .ZN(n18999) );
  NAND2_X1 U21991 ( .A1(n19311), .A2(n19350), .ZN(n19184) );
  NOR2_X1 U21992 ( .A1(n18999), .A2(n19184), .ZN(n18930) );
  AOI22_X1 U21993 ( .A1(n19246), .A2(n19240), .B1(n19245), .B2(n18930), .ZN(
        n18917) );
  NOR2_X1 U21994 ( .A1(n18915), .A2(n18914), .ZN(n19249) );
  INV_X1 U21995 ( .A(n19249), .ZN(n18955) );
  NOR2_X1 U21996 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18955), .ZN(
        n19185) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19247), .B1(
        n18956), .B2(n19185), .ZN(n18931) );
  NOR2_X2 U21998 ( .A1(n19091), .A2(n18999), .ZN(n18995) );
  AOI22_X1 U21999 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18931), .B1(
        n19250), .B2(n18995), .ZN(n18916) );
  OAI211_X1 U22000 ( .C1(n21309), .C2(n19253), .A(n18917), .B(n18916), .ZN(
        P3_U2876) );
  INV_X1 U22001 ( .A(n18995), .ZN(n18977) );
  INV_X1 U22002 ( .A(n21309), .ZN(n19288) );
  AOI22_X1 U22003 ( .A1(n19288), .A2(n19256), .B1(n19254), .B2(n18930), .ZN(
        n18919) );
  AOI22_X1 U22004 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18931), .B1(
        n19240), .B2(n19255), .ZN(n18918) );
  OAI211_X1 U22005 ( .C1(n19259), .C2(n18977), .A(n18919), .B(n18918), .ZN(
        P3_U2877) );
  AOI22_X1 U22006 ( .A1(n19288), .A2(n21307), .B1(n21304), .B2(n18930), .ZN(
        n18921) );
  AOI22_X1 U22007 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18931), .B1(
        n19224), .B2(n19240), .ZN(n18920) );
  OAI211_X1 U22008 ( .C1(n21310), .C2(n18977), .A(n18921), .B(n18920), .ZN(
        P3_U2878) );
  AOI22_X1 U22009 ( .A1(n19288), .A2(n19261), .B1(n19260), .B2(n18930), .ZN(
        n18923) );
  AOI22_X1 U22010 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18931), .B1(
        n19240), .B2(n19262), .ZN(n18922) );
  OAI211_X1 U22011 ( .C1(n19265), .C2(n18977), .A(n18923), .B(n18922), .ZN(
        P3_U2879) );
  AOI22_X1 U22012 ( .A1(n19240), .A2(n19267), .B1(n19266), .B2(n18930), .ZN(
        n18925) );
  AOI22_X1 U22013 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18931), .B1(
        n19288), .B2(n19268), .ZN(n18924) );
  OAI211_X1 U22014 ( .C1(n19271), .C2(n18977), .A(n18925), .B(n18924), .ZN(
        P3_U2880) );
  INV_X1 U22015 ( .A(n19240), .ZN(n19237) );
  AOI22_X1 U22016 ( .A1(n19288), .A2(n19273), .B1(n19272), .B2(n18930), .ZN(
        n18927) );
  AOI22_X1 U22017 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18931), .B1(
        n19274), .B2(n18995), .ZN(n18926) );
  OAI211_X1 U22018 ( .C1(n19237), .C2(n19277), .A(n18927), .B(n18926), .ZN(
        P3_U2881) );
  AOI22_X1 U22019 ( .A1(n19288), .A2(n19279), .B1(n19278), .B2(n18930), .ZN(
        n18929) );
  AOI22_X1 U22020 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18931), .B1(
        n19240), .B2(n19280), .ZN(n18928) );
  OAI211_X1 U22021 ( .C1(n19283), .C2(n18977), .A(n18929), .B(n18928), .ZN(
        P3_U2882) );
  INV_X1 U22022 ( .A(n19205), .ZN(n19291) );
  INV_X1 U22023 ( .A(n19210), .ZN(n19285) );
  AOI22_X1 U22024 ( .A1(n19240), .A2(n19285), .B1(n19284), .B2(n18930), .ZN(
        n18933) );
  AOI22_X1 U22025 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18931), .B1(
        n19287), .B2(n18995), .ZN(n18932) );
  OAI211_X1 U22026 ( .C1(n21309), .C2(n19291), .A(n18933), .B(n18932), .ZN(
        P3_U2883) );
  NOR2_X2 U22027 ( .A1(n18999), .A2(n19112), .ZN(n19017) );
  NOR2_X1 U22028 ( .A1(n18995), .A2(n19017), .ZN(n18978) );
  NOR2_X1 U22029 ( .A1(n19163), .A2(n18978), .ZN(n18951) );
  AOI22_X1 U22030 ( .A1(n19288), .A2(n19246), .B1(n19245), .B2(n18951), .ZN(
        n18938) );
  INV_X1 U22031 ( .A(n18978), .ZN(n18934) );
  AOI22_X1 U22032 ( .A1(n19159), .A2(n18936), .B1(n18935), .B2(n18934), .ZN(
        n18952) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18952), .B1(
        n19250), .B2(n19017), .ZN(n18937) );
  OAI211_X1 U22034 ( .C1(n18969), .C2(n19253), .A(n18938), .B(n18937), .ZN(
        P3_U2884) );
  INV_X1 U22035 ( .A(n19017), .ZN(n19013) );
  AOI22_X1 U22036 ( .A1(n18973), .A2(n19256), .B1(n19254), .B2(n18951), .ZN(
        n18940) );
  AOI22_X1 U22037 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18952), .B1(
        n19288), .B2(n19255), .ZN(n18939) );
  OAI211_X1 U22038 ( .C1(n19259), .C2(n19013), .A(n18940), .B(n18939), .ZN(
        P3_U2885) );
  AOI22_X1 U22039 ( .A1(n19224), .A2(n19288), .B1(n21304), .B2(n18951), .ZN(
        n18942) );
  AOI22_X1 U22040 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18952), .B1(
        n21307), .B2(n18973), .ZN(n18941) );
  OAI211_X1 U22041 ( .C1(n21310), .C2(n19013), .A(n18942), .B(n18941), .ZN(
        P3_U2886) );
  AOI22_X1 U22042 ( .A1(n19288), .A2(n19262), .B1(n19260), .B2(n18951), .ZN(
        n18944) );
  AOI22_X1 U22043 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18952), .B1(
        n18973), .B2(n19261), .ZN(n18943) );
  OAI211_X1 U22044 ( .C1(n19265), .C2(n19013), .A(n18944), .B(n18943), .ZN(
        P3_U2887) );
  AOI22_X1 U22045 ( .A1(n18973), .A2(n19268), .B1(n19266), .B2(n18951), .ZN(
        n18946) );
  AOI22_X1 U22046 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18952), .B1(
        n19288), .B2(n19267), .ZN(n18945) );
  OAI211_X1 U22047 ( .C1(n19271), .C2(n19013), .A(n18946), .B(n18945), .ZN(
        P3_U2888) );
  INV_X1 U22048 ( .A(n19273), .ZN(n19234) );
  INV_X1 U22049 ( .A(n19277), .ZN(n19231) );
  AOI22_X1 U22050 ( .A1(n19288), .A2(n19231), .B1(n19272), .B2(n18951), .ZN(
        n18948) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18952), .B1(
        n19274), .B2(n19017), .ZN(n18947) );
  OAI211_X1 U22052 ( .C1(n18969), .C2(n19234), .A(n18948), .B(n18947), .ZN(
        P3_U2889) );
  AOI22_X1 U22053 ( .A1(n18973), .A2(n19279), .B1(n19278), .B2(n18951), .ZN(
        n18950) );
  AOI22_X1 U22054 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18952), .B1(
        n19288), .B2(n19280), .ZN(n18949) );
  OAI211_X1 U22055 ( .C1(n19283), .C2(n19013), .A(n18950), .B(n18949), .ZN(
        P3_U2890) );
  AOI22_X1 U22056 ( .A1(n19288), .A2(n19285), .B1(n19284), .B2(n18951), .ZN(
        n18954) );
  AOI22_X1 U22057 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18952), .B1(
        n19287), .B2(n19017), .ZN(n18953) );
  OAI211_X1 U22058 ( .C1(n18969), .C2(n19291), .A(n18954), .B(n18953), .ZN(
        P3_U2891) );
  AOI22_X1 U22059 ( .A1(n18973), .A2(n19246), .B1(n19245), .B2(n18972), .ZN(
        n18958) );
  AOI21_X1 U22060 ( .B1(n19311), .B2(n19214), .A(n18955), .ZN(n19045) );
  NAND2_X1 U22061 ( .A1(n18956), .A2(n19045), .ZN(n18974) );
  NAND2_X1 U22062 ( .A1(n19309), .A2(n18956), .ZN(n19037) );
  AOI22_X1 U22063 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18974), .B1(
        n19250), .B2(n19042), .ZN(n18957) );
  OAI211_X1 U22064 ( .C1(n19253), .C2(n18977), .A(n18958), .B(n18957), .ZN(
        P3_U2892) );
  AOI22_X1 U22065 ( .A1(n19256), .A2(n18995), .B1(n19254), .B2(n18972), .ZN(
        n18960) );
  AOI22_X1 U22066 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18974), .B1(
        n18973), .B2(n19255), .ZN(n18959) );
  OAI211_X1 U22067 ( .C1(n19259), .C2(n19037), .A(n18960), .B(n18959), .ZN(
        P3_U2893) );
  AOI22_X1 U22068 ( .A1(n21307), .A2(n18995), .B1(n21304), .B2(n18972), .ZN(
        n18962) );
  AOI22_X1 U22069 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18974), .B1(
        n19224), .B2(n18973), .ZN(n18961) );
  OAI211_X1 U22070 ( .C1(n21310), .C2(n19037), .A(n18962), .B(n18961), .ZN(
        P3_U2894) );
  AOI22_X1 U22071 ( .A1(n18973), .A2(n19262), .B1(n19260), .B2(n18972), .ZN(
        n18964) );
  AOI22_X1 U22072 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18974), .B1(
        n19261), .B2(n18995), .ZN(n18963) );
  OAI211_X1 U22073 ( .C1(n19265), .C2(n19037), .A(n18964), .B(n18963), .ZN(
        P3_U2895) );
  AOI22_X1 U22074 ( .A1(n18973), .A2(n19267), .B1(n19266), .B2(n18972), .ZN(
        n18966) );
  AOI22_X1 U22075 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18974), .B1(
        n19268), .B2(n18995), .ZN(n18965) );
  OAI211_X1 U22076 ( .C1(n19271), .C2(n19037), .A(n18966), .B(n18965), .ZN(
        P3_U2896) );
  AOI22_X1 U22077 ( .A1(n19273), .A2(n18995), .B1(n19272), .B2(n18972), .ZN(
        n18968) );
  AOI22_X1 U22078 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18974), .B1(
        n19274), .B2(n19042), .ZN(n18967) );
  OAI211_X1 U22079 ( .C1(n18969), .C2(n19277), .A(n18968), .B(n18967), .ZN(
        P3_U2897) );
  AOI22_X1 U22080 ( .A1(n18973), .A2(n19280), .B1(n19278), .B2(n18972), .ZN(
        n18971) );
  AOI22_X1 U22081 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18974), .B1(
        n19279), .B2(n18995), .ZN(n18970) );
  OAI211_X1 U22082 ( .C1(n19283), .C2(n19037), .A(n18971), .B(n18970), .ZN(
        P3_U2898) );
  AOI22_X1 U22083 ( .A1(n18973), .A2(n19285), .B1(n19284), .B2(n18972), .ZN(
        n18976) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18974), .B1(
        n19287), .B2(n19042), .ZN(n18975) );
  OAI211_X1 U22085 ( .C1(n19291), .C2(n18977), .A(n18976), .B(n18975), .ZN(
        P3_U2899) );
  INV_X1 U22086 ( .A(n19156), .ZN(n19317) );
  INV_X1 U22087 ( .A(n19046), .ZN(n19021) );
  NOR2_X2 U22088 ( .A1(n19317), .A2(n19021), .ZN(n19063) );
  NOR2_X1 U22089 ( .A1(n19042), .A2(n19063), .ZN(n19023) );
  NOR2_X1 U22090 ( .A1(n19163), .A2(n19023), .ZN(n18994) );
  AOI22_X1 U22091 ( .A1(n19246), .A2(n18995), .B1(n19245), .B2(n18994), .ZN(
        n18981) );
  OAI21_X1 U22092 ( .B1(n18978), .B2(n19214), .A(n19023), .ZN(n18979) );
  OAI211_X1 U22093 ( .C1(n19063), .C2(n19452), .A(n19216), .B(n18979), .ZN(
        n18996) );
  AOI22_X1 U22094 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18996), .B1(
        n19250), .B2(n19063), .ZN(n18980) );
  OAI211_X1 U22095 ( .C1(n19253), .C2(n19013), .A(n18981), .B(n18980), .ZN(
        P3_U2900) );
  INV_X1 U22096 ( .A(n19063), .ZN(n19059) );
  AOI22_X1 U22097 ( .A1(n19256), .A2(n19017), .B1(n19254), .B2(n18994), .ZN(
        n18983) );
  AOI22_X1 U22098 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18996), .B1(
        n19255), .B2(n18995), .ZN(n18982) );
  OAI211_X1 U22099 ( .C1(n19259), .C2(n19059), .A(n18983), .B(n18982), .ZN(
        P3_U2901) );
  AOI22_X1 U22100 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18996), .B1(
        n21304), .B2(n18994), .ZN(n18985) );
  AOI22_X1 U22101 ( .A1(n19224), .A2(n18995), .B1(n21307), .B2(n19017), .ZN(
        n18984) );
  OAI211_X1 U22102 ( .C1(n21310), .C2(n19059), .A(n18985), .B(n18984), .ZN(
        P3_U2902) );
  AOI22_X1 U22103 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18996), .B1(
        n19260), .B2(n18994), .ZN(n18987) );
  AOI22_X1 U22104 ( .A1(n19261), .A2(n19017), .B1(n19262), .B2(n18995), .ZN(
        n18986) );
  OAI211_X1 U22105 ( .C1(n19265), .C2(n19059), .A(n18987), .B(n18986), .ZN(
        P3_U2903) );
  AOI22_X1 U22106 ( .A1(n19268), .A2(n19017), .B1(n19266), .B2(n18994), .ZN(
        n18989) );
  AOI22_X1 U22107 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18996), .B1(
        n19267), .B2(n18995), .ZN(n18988) );
  OAI211_X1 U22108 ( .C1(n19271), .C2(n19059), .A(n18989), .B(n18988), .ZN(
        P3_U2904) );
  AOI22_X1 U22109 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18996), .B1(
        n19272), .B2(n18994), .ZN(n18991) );
  AOI22_X1 U22110 ( .A1(n19231), .A2(n18995), .B1(n19274), .B2(n19063), .ZN(
        n18990) );
  OAI211_X1 U22111 ( .C1(n19234), .C2(n19013), .A(n18991), .B(n18990), .ZN(
        P3_U2905) );
  AOI22_X1 U22112 ( .A1(n19280), .A2(n18995), .B1(n19278), .B2(n18994), .ZN(
        n18993) );
  AOI22_X1 U22113 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18996), .B1(
        n19279), .B2(n19017), .ZN(n18992) );
  OAI211_X1 U22114 ( .C1(n19283), .C2(n19059), .A(n18993), .B(n18992), .ZN(
        P3_U2906) );
  AOI22_X1 U22115 ( .A1(n19285), .A2(n18995), .B1(n19284), .B2(n18994), .ZN(
        n18998) );
  AOI22_X1 U22116 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18996), .B1(
        n19287), .B2(n19063), .ZN(n18997) );
  OAI211_X1 U22117 ( .C1(n19291), .C2(n19013), .A(n18998), .B(n18997), .ZN(
        P3_U2907) );
  NOR2_X1 U22118 ( .A1(n19021), .A2(n19184), .ZN(n19016) );
  AOI22_X1 U22119 ( .A1(n19213), .A2(n19042), .B1(n19245), .B2(n19016), .ZN(
        n19002) );
  NOR2_X1 U22120 ( .A1(n19311), .A2(n18999), .ZN(n19000) );
  AOI22_X1 U22121 ( .A1(n19188), .A2(n19000), .B1(n19046), .B2(n19185), .ZN(
        n19018) );
  NOR2_X2 U22122 ( .A1(n19091), .A2(n19021), .ZN(n19081) );
  AOI22_X1 U22123 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19018), .B1(
        n19250), .B2(n19081), .ZN(n19001) );
  OAI211_X1 U22124 ( .C1(n19221), .C2(n19013), .A(n19002), .B(n19001), .ZN(
        P3_U2908) );
  INV_X1 U22125 ( .A(n19081), .ZN(n19088) );
  AOI22_X1 U22126 ( .A1(n19255), .A2(n19017), .B1(n19254), .B2(n19016), .ZN(
        n19004) );
  AOI22_X1 U22127 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19018), .B1(
        n19256), .B2(n19042), .ZN(n19003) );
  OAI211_X1 U22128 ( .C1(n19259), .C2(n19088), .A(n19004), .B(n19003), .ZN(
        P3_U2909) );
  AOI22_X1 U22129 ( .A1(n21307), .A2(n19042), .B1(n21304), .B2(n19016), .ZN(
        n19006) );
  AOI22_X1 U22130 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19018), .B1(
        n19224), .B2(n19017), .ZN(n19005) );
  OAI211_X1 U22131 ( .C1(n21310), .C2(n19088), .A(n19006), .B(n19005), .ZN(
        P3_U2910) );
  AOI22_X1 U22132 ( .A1(n19261), .A2(n19042), .B1(n19260), .B2(n19016), .ZN(
        n19008) );
  AOI22_X1 U22133 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19018), .B1(
        n19262), .B2(n19017), .ZN(n19007) );
  OAI211_X1 U22134 ( .C1(n19265), .C2(n19088), .A(n19008), .B(n19007), .ZN(
        P3_U2911) );
  AOI22_X1 U22135 ( .A1(n19268), .A2(n19042), .B1(n19266), .B2(n19016), .ZN(
        n19010) );
  AOI22_X1 U22136 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19018), .B1(
        n19267), .B2(n19017), .ZN(n19009) );
  OAI211_X1 U22137 ( .C1(n19271), .C2(n19088), .A(n19010), .B(n19009), .ZN(
        P3_U2912) );
  AOI22_X1 U22138 ( .A1(n19273), .A2(n19042), .B1(n19272), .B2(n19016), .ZN(
        n19012) );
  AOI22_X1 U22139 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19018), .B1(
        n19274), .B2(n19081), .ZN(n19011) );
  OAI211_X1 U22140 ( .C1(n19277), .C2(n19013), .A(n19012), .B(n19011), .ZN(
        P3_U2913) );
  AOI22_X1 U22141 ( .A1(n19279), .A2(n19042), .B1(n19278), .B2(n19016), .ZN(
        n19015) );
  AOI22_X1 U22142 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19018), .B1(
        n19280), .B2(n19017), .ZN(n19014) );
  OAI211_X1 U22143 ( .C1(n19283), .C2(n19088), .A(n19015), .B(n19014), .ZN(
        P3_U2914) );
  AOI22_X1 U22144 ( .A1(n19285), .A2(n19017), .B1(n19284), .B2(n19016), .ZN(
        n19020) );
  AOI22_X1 U22145 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19018), .B1(
        n19287), .B2(n19081), .ZN(n19019) );
  OAI211_X1 U22146 ( .C1(n19291), .C2(n19037), .A(n19020), .B(n19019), .ZN(
        P3_U2915) );
  NOR2_X2 U22147 ( .A1(n19021), .A2(n19112), .ZN(n19104) );
  NOR2_X1 U22148 ( .A1(n19081), .A2(n19104), .ZN(n19067) );
  NOR2_X1 U22149 ( .A1(n19163), .A2(n19067), .ZN(n19040) );
  AOI22_X1 U22150 ( .A1(n19213), .A2(n19063), .B1(n19245), .B2(n19040), .ZN(
        n19026) );
  AOI221_X1 U22151 ( .B1(n19067), .B2(n19214), .C1(n19067), .C2(n19023), .A(
        n19022), .ZN(n19024) );
  INV_X1 U22152 ( .A(n19024), .ZN(n19041) );
  AOI22_X1 U22153 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19041), .B1(
        n19250), .B2(n19104), .ZN(n19025) );
  OAI211_X1 U22154 ( .C1(n19221), .C2(n19037), .A(n19026), .B(n19025), .ZN(
        P3_U2916) );
  INV_X1 U22155 ( .A(n19104), .ZN(n19111) );
  AOI22_X1 U22156 ( .A1(n19255), .A2(n19042), .B1(n19254), .B2(n19040), .ZN(
        n19028) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19041), .B1(
        n19256), .B2(n19063), .ZN(n19027) );
  OAI211_X1 U22158 ( .C1(n19259), .C2(n19111), .A(n19028), .B(n19027), .ZN(
        P3_U2917) );
  AOI22_X1 U22159 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19041), .B1(
        n21304), .B2(n19040), .ZN(n19030) );
  AOI22_X1 U22160 ( .A1(n19224), .A2(n19042), .B1(n21307), .B2(n19063), .ZN(
        n19029) );
  OAI211_X1 U22161 ( .C1(n21310), .C2(n19111), .A(n19030), .B(n19029), .ZN(
        P3_U2918) );
  AOI22_X1 U22162 ( .A1(n19262), .A2(n19042), .B1(n19260), .B2(n19040), .ZN(
        n19032) );
  AOI22_X1 U22163 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19041), .B1(
        n19261), .B2(n19063), .ZN(n19031) );
  OAI211_X1 U22164 ( .C1(n19265), .C2(n19111), .A(n19032), .B(n19031), .ZN(
        P3_U2919) );
  AOI22_X1 U22165 ( .A1(n19268), .A2(n19063), .B1(n19266), .B2(n19040), .ZN(
        n19034) );
  AOI22_X1 U22166 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19041), .B1(
        n19267), .B2(n19042), .ZN(n19033) );
  OAI211_X1 U22167 ( .C1(n19271), .C2(n19111), .A(n19034), .B(n19033), .ZN(
        P3_U2920) );
  AOI22_X1 U22168 ( .A1(n19273), .A2(n19063), .B1(n19272), .B2(n19040), .ZN(
        n19036) );
  AOI22_X1 U22169 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19041), .B1(
        n19274), .B2(n19104), .ZN(n19035) );
  OAI211_X1 U22170 ( .C1(n19277), .C2(n19037), .A(n19036), .B(n19035), .ZN(
        P3_U2921) );
  AOI22_X1 U22171 ( .A1(n19279), .A2(n19063), .B1(n19278), .B2(n19040), .ZN(
        n19039) );
  AOI22_X1 U22172 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19041), .B1(
        n19280), .B2(n19042), .ZN(n19038) );
  OAI211_X1 U22173 ( .C1(n19283), .C2(n19111), .A(n19039), .B(n19038), .ZN(
        P3_U2922) );
  AOI22_X1 U22174 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19041), .B1(
        n19284), .B2(n19040), .ZN(n19044) );
  AOI22_X1 U22175 ( .A1(n19285), .A2(n19042), .B1(n19287), .B2(n19104), .ZN(
        n19043) );
  OAI211_X1 U22176 ( .C1(n19291), .C2(n19059), .A(n19044), .B(n19043), .ZN(
        P3_U2923) );
  AOI22_X1 U22177 ( .A1(n19213), .A2(n19081), .B1(n19245), .B2(n19062), .ZN(
        n19048) );
  NAND2_X1 U22178 ( .A1(n19046), .A2(n19045), .ZN(n19064) );
  NAND2_X1 U22179 ( .A1(n19309), .A2(n19046), .ZN(n19117) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19064), .B1(
        n19250), .B2(n19131), .ZN(n19047) );
  OAI211_X1 U22181 ( .C1(n19221), .C2(n19059), .A(n19048), .B(n19047), .ZN(
        P3_U2924) );
  AOI22_X1 U22182 ( .A1(n19256), .A2(n19081), .B1(n19254), .B2(n19062), .ZN(
        n19050) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19064), .B1(
        n19255), .B2(n19063), .ZN(n19049) );
  OAI211_X1 U22184 ( .C1(n19259), .C2(n19117), .A(n19050), .B(n19049), .ZN(
        P3_U2925) );
  AOI22_X1 U22185 ( .A1(n21307), .A2(n19081), .B1(n21304), .B2(n19062), .ZN(
        n19052) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19064), .B1(
        n19224), .B2(n19063), .ZN(n19051) );
  OAI211_X1 U22187 ( .C1(n21310), .C2(n19117), .A(n19052), .B(n19051), .ZN(
        P3_U2926) );
  AOI22_X1 U22188 ( .A1(n19262), .A2(n19063), .B1(n19260), .B2(n19062), .ZN(
        n19054) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19064), .B1(
        n19261), .B2(n19081), .ZN(n19053) );
  OAI211_X1 U22190 ( .C1(n19265), .C2(n19117), .A(n19054), .B(n19053), .ZN(
        P3_U2927) );
  AOI22_X1 U22191 ( .A1(n19266), .A2(n19062), .B1(n19267), .B2(n19063), .ZN(
        n19056) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19064), .B1(
        n19268), .B2(n19081), .ZN(n19055) );
  OAI211_X1 U22193 ( .C1(n19271), .C2(n19117), .A(n19056), .B(n19055), .ZN(
        P3_U2928) );
  AOI22_X1 U22194 ( .A1(n19273), .A2(n19081), .B1(n19272), .B2(n19062), .ZN(
        n19058) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19064), .B1(
        n19274), .B2(n19131), .ZN(n19057) );
  OAI211_X1 U22196 ( .C1(n19277), .C2(n19059), .A(n19058), .B(n19057), .ZN(
        P3_U2929) );
  AOI22_X1 U22197 ( .A1(n19279), .A2(n19081), .B1(n19278), .B2(n19062), .ZN(
        n19061) );
  AOI22_X1 U22198 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19064), .B1(
        n19280), .B2(n19063), .ZN(n19060) );
  OAI211_X1 U22199 ( .C1(n19283), .C2(n19117), .A(n19061), .B(n19060), .ZN(
        P3_U2930) );
  AOI22_X1 U22200 ( .A1(n19285), .A2(n19063), .B1(n19284), .B2(n19062), .ZN(
        n19066) );
  AOI22_X1 U22201 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19064), .B1(
        n19287), .B2(n19131), .ZN(n19065) );
  OAI211_X1 U22202 ( .C1(n19291), .C2(n19088), .A(n19066), .B(n19065), .ZN(
        P3_U2931) );
  NOR2_X2 U22203 ( .A1(n19317), .A2(n19135), .ZN(n19148) );
  NOR2_X1 U22204 ( .A1(n19131), .A2(n19148), .ZN(n19113) );
  NOR2_X1 U22205 ( .A1(n19163), .A2(n19113), .ZN(n19084) );
  AOI22_X1 U22206 ( .A1(n19213), .A2(n19104), .B1(n19245), .B2(n19084), .ZN(
        n19070) );
  OAI21_X1 U22207 ( .B1(n19067), .B2(n19214), .A(n19113), .ZN(n19068) );
  OAI211_X1 U22208 ( .C1(n19148), .C2(n19452), .A(n19216), .B(n19068), .ZN(
        n19085) );
  AOI22_X1 U22209 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19085), .B1(
        n19250), .B2(n19148), .ZN(n19069) );
  OAI211_X1 U22210 ( .C1(n19221), .C2(n19088), .A(n19070), .B(n19069), .ZN(
        P3_U2932) );
  INV_X1 U22211 ( .A(n19148), .ZN(n19155) );
  AOI22_X1 U22212 ( .A1(n19256), .A2(n19104), .B1(n19254), .B2(n19084), .ZN(
        n19072) );
  AOI22_X1 U22213 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19085), .B1(
        n19255), .B2(n19081), .ZN(n19071) );
  OAI211_X1 U22214 ( .C1(n19259), .C2(n19155), .A(n19072), .B(n19071), .ZN(
        P3_U2933) );
  AOI22_X1 U22215 ( .A1(n19224), .A2(n19081), .B1(n21304), .B2(n19084), .ZN(
        n19074) );
  AOI22_X1 U22216 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19085), .B1(
        n21307), .B2(n19104), .ZN(n19073) );
  OAI211_X1 U22217 ( .C1(n21310), .C2(n19155), .A(n19074), .B(n19073), .ZN(
        P3_U2934) );
  AOI22_X1 U22218 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19085), .B1(
        n19260), .B2(n19084), .ZN(n19076) );
  AOI22_X1 U22219 ( .A1(n19261), .A2(n19104), .B1(n19262), .B2(n19081), .ZN(
        n19075) );
  OAI211_X1 U22220 ( .C1(n19265), .C2(n19155), .A(n19076), .B(n19075), .ZN(
        P3_U2935) );
  AOI22_X1 U22221 ( .A1(n19266), .A2(n19084), .B1(n19267), .B2(n19081), .ZN(
        n19078) );
  AOI22_X1 U22222 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19085), .B1(
        n19268), .B2(n19104), .ZN(n19077) );
  OAI211_X1 U22223 ( .C1(n19271), .C2(n19155), .A(n19078), .B(n19077), .ZN(
        P3_U2936) );
  AOI22_X1 U22224 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19085), .B1(
        n19272), .B2(n19084), .ZN(n19080) );
  AOI22_X1 U22225 ( .A1(n19274), .A2(n19148), .B1(n19273), .B2(n19104), .ZN(
        n19079) );
  OAI211_X1 U22226 ( .C1(n19277), .C2(n19088), .A(n19080), .B(n19079), .ZN(
        P3_U2937) );
  AOI22_X1 U22227 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19085), .B1(
        n19278), .B2(n19084), .ZN(n19083) );
  AOI22_X1 U22228 ( .A1(n19279), .A2(n19104), .B1(n19280), .B2(n19081), .ZN(
        n19082) );
  OAI211_X1 U22229 ( .C1(n19283), .C2(n19155), .A(n19083), .B(n19082), .ZN(
        P3_U2938) );
  AOI22_X1 U22230 ( .A1(n19205), .A2(n19104), .B1(n19284), .B2(n19084), .ZN(
        n19087) );
  AOI22_X1 U22231 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19085), .B1(
        n19287), .B2(n19148), .ZN(n19086) );
  OAI211_X1 U22232 ( .C1(n19210), .C2(n19088), .A(n19087), .B(n19086), .ZN(
        P3_U2939) );
  NOR2_X1 U22233 ( .A1(n19135), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19089) );
  AND2_X1 U22234 ( .A1(n19350), .A2(n19089), .ZN(n19107) );
  AOI22_X1 U22235 ( .A1(n19213), .A2(n19131), .B1(n19245), .B2(n19107), .ZN(
        n19093) );
  NOR2_X1 U22236 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19244), .ZN(
        n19090) );
  AOI22_X1 U22237 ( .A1(n19188), .A2(n19090), .B1(n19249), .B2(n19089), .ZN(
        n19108) );
  NOR2_X2 U22238 ( .A1(n19091), .A2(n19135), .ZN(n19180) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19108), .B1(
        n19250), .B2(n19180), .ZN(n19092) );
  OAI211_X1 U22240 ( .C1(n19221), .C2(n19111), .A(n19093), .B(n19092), .ZN(
        P3_U2940) );
  INV_X1 U22241 ( .A(n19180), .ZN(n19176) );
  AOI22_X1 U22242 ( .A1(n19256), .A2(n19131), .B1(n19254), .B2(n19107), .ZN(
        n19095) );
  AOI22_X1 U22243 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19108), .B1(
        n19255), .B2(n19104), .ZN(n19094) );
  OAI211_X1 U22244 ( .C1(n19259), .C2(n19176), .A(n19095), .B(n19094), .ZN(
        P3_U2941) );
  AOI22_X1 U22245 ( .A1(n21307), .A2(n19131), .B1(n21304), .B2(n19107), .ZN(
        n19097) );
  AOI22_X1 U22246 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19108), .B1(
        n19224), .B2(n19104), .ZN(n19096) );
  OAI211_X1 U22247 ( .C1(n21310), .C2(n19176), .A(n19097), .B(n19096), .ZN(
        P3_U2942) );
  AOI22_X1 U22248 ( .A1(n19261), .A2(n19131), .B1(n19260), .B2(n19107), .ZN(
        n19099) );
  AOI22_X1 U22249 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19108), .B1(
        n19262), .B2(n19104), .ZN(n19098) );
  OAI211_X1 U22250 ( .C1(n19265), .C2(n19176), .A(n19099), .B(n19098), .ZN(
        P3_U2943) );
  AOI22_X1 U22251 ( .A1(n19266), .A2(n19107), .B1(n19267), .B2(n19104), .ZN(
        n19101) );
  AOI22_X1 U22252 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19108), .B1(
        n19268), .B2(n19131), .ZN(n19100) );
  OAI211_X1 U22253 ( .C1(n19271), .C2(n19176), .A(n19101), .B(n19100), .ZN(
        P3_U2944) );
  AOI22_X1 U22254 ( .A1(n19273), .A2(n19131), .B1(n19272), .B2(n19107), .ZN(
        n19103) );
  AOI22_X1 U22255 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19108), .B1(
        n19274), .B2(n19180), .ZN(n19102) );
  OAI211_X1 U22256 ( .C1(n19277), .C2(n19111), .A(n19103), .B(n19102), .ZN(
        P3_U2945) );
  AOI22_X1 U22257 ( .A1(n19279), .A2(n19131), .B1(n19278), .B2(n19107), .ZN(
        n19106) );
  AOI22_X1 U22258 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19108), .B1(
        n19280), .B2(n19104), .ZN(n19105) );
  OAI211_X1 U22259 ( .C1(n19283), .C2(n19176), .A(n19106), .B(n19105), .ZN(
        P3_U2946) );
  AOI22_X1 U22260 ( .A1(n19205), .A2(n19131), .B1(n19284), .B2(n19107), .ZN(
        n19110) );
  AOI22_X1 U22261 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19108), .B1(
        n19287), .B2(n19180), .ZN(n19109) );
  OAI211_X1 U22262 ( .C1(n19210), .C2(n19111), .A(n19110), .B(n19109), .ZN(
        P3_U2947) );
  NAND2_X1 U22263 ( .A1(n19350), .A2(n19157), .ZN(n19211) );
  NOR2_X1 U22264 ( .A1(n19135), .A2(n19211), .ZN(n19130) );
  AOI22_X1 U22265 ( .A1(n19213), .A2(n19148), .B1(n19245), .B2(n19130), .ZN(
        n19116) );
  NOR2_X2 U22266 ( .A1(n19135), .A2(n19112), .ZN(n19201) );
  AOI221_X1 U22267 ( .B1(n19113), .B2(n19176), .C1(n19214), .C2(n19176), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19114) );
  OAI21_X1 U22268 ( .B1(n19201), .B2(n19114), .A(n19216), .ZN(n19132) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19132), .B1(
        n19250), .B2(n19201), .ZN(n19115) );
  OAI211_X1 U22270 ( .C1(n19221), .C2(n19117), .A(n19116), .B(n19115), .ZN(
        P3_U2948) );
  INV_X1 U22271 ( .A(n19201), .ZN(n19209) );
  AOI22_X1 U22272 ( .A1(n19255), .A2(n19131), .B1(n19254), .B2(n19130), .ZN(
        n19119) );
  AOI22_X1 U22273 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19132), .B1(
        n19256), .B2(n19148), .ZN(n19118) );
  OAI211_X1 U22274 ( .C1(n19259), .C2(n19209), .A(n19119), .B(n19118), .ZN(
        P3_U2949) );
  AOI22_X1 U22275 ( .A1(n21307), .A2(n19148), .B1(n21304), .B2(n19130), .ZN(
        n19121) );
  AOI22_X1 U22276 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19132), .B1(
        n19224), .B2(n19131), .ZN(n19120) );
  OAI211_X1 U22277 ( .C1(n21310), .C2(n19209), .A(n19121), .B(n19120), .ZN(
        P3_U2950) );
  AOI22_X1 U22278 ( .A1(n19261), .A2(n19148), .B1(n19260), .B2(n19130), .ZN(
        n19123) );
  AOI22_X1 U22279 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19132), .B1(
        n19262), .B2(n19131), .ZN(n19122) );
  OAI211_X1 U22280 ( .C1(n19265), .C2(n19209), .A(n19123), .B(n19122), .ZN(
        P3_U2951) );
  AOI22_X1 U22281 ( .A1(n19266), .A2(n19130), .B1(n19267), .B2(n19131), .ZN(
        n19125) );
  AOI22_X1 U22282 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19132), .B1(
        n19268), .B2(n19148), .ZN(n19124) );
  OAI211_X1 U22283 ( .C1(n19271), .C2(n19209), .A(n19125), .B(n19124), .ZN(
        P3_U2952) );
  AOI22_X1 U22284 ( .A1(n19231), .A2(n19131), .B1(n19272), .B2(n19130), .ZN(
        n19127) );
  AOI22_X1 U22285 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19132), .B1(
        n19274), .B2(n19201), .ZN(n19126) );
  OAI211_X1 U22286 ( .C1(n19234), .C2(n19155), .A(n19127), .B(n19126), .ZN(
        P3_U2953) );
  AOI22_X1 U22287 ( .A1(n19280), .A2(n19131), .B1(n19278), .B2(n19130), .ZN(
        n19129) );
  AOI22_X1 U22288 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19132), .B1(
        n19279), .B2(n19148), .ZN(n19128) );
  OAI211_X1 U22289 ( .C1(n19283), .C2(n19209), .A(n19129), .B(n19128), .ZN(
        P3_U2954) );
  AOI22_X1 U22290 ( .A1(n19285), .A2(n19131), .B1(n19284), .B2(n19130), .ZN(
        n19134) );
  AOI22_X1 U22291 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19132), .B1(
        n19287), .B2(n19201), .ZN(n19133) );
  OAI211_X1 U22292 ( .C1(n19291), .C2(n19155), .A(n19134), .B(n19133), .ZN(
        P3_U2955) );
  NOR2_X1 U22293 ( .A1(n19311), .A2(n19135), .ZN(n19187) );
  AND2_X1 U22294 ( .A1(n19350), .A2(n19187), .ZN(n19151) );
  AOI22_X1 U22295 ( .A1(n19246), .A2(n19148), .B1(n19245), .B2(n19151), .ZN(
        n19137) );
  OAI211_X1 U22296 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19188), .A(
        n19249), .B(n19158), .ZN(n19152) );
  NAND2_X1 U22297 ( .A1(n19309), .A2(n19158), .ZN(n19220) );
  INV_X1 U22298 ( .A(n19220), .ZN(n19239) );
  AOI22_X1 U22299 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19152), .B1(
        n19250), .B2(n19239), .ZN(n19136) );
  OAI211_X1 U22300 ( .C1(n19253), .C2(n19176), .A(n19137), .B(n19136), .ZN(
        P3_U2956) );
  AOI22_X1 U22301 ( .A1(n19255), .A2(n19148), .B1(n19254), .B2(n19151), .ZN(
        n19139) );
  AOI22_X1 U22302 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19152), .B1(
        n19256), .B2(n19180), .ZN(n19138) );
  OAI211_X1 U22303 ( .C1(n19259), .C2(n19220), .A(n19139), .B(n19138), .ZN(
        P3_U2957) );
  AOI22_X1 U22304 ( .A1(n21307), .A2(n19180), .B1(n21304), .B2(n19151), .ZN(
        n19141) );
  AOI22_X1 U22305 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19152), .B1(
        n19224), .B2(n19148), .ZN(n19140) );
  OAI211_X1 U22306 ( .C1(n21310), .C2(n19220), .A(n19141), .B(n19140), .ZN(
        P3_U2958) );
  AOI22_X1 U22307 ( .A1(n19261), .A2(n19180), .B1(n19260), .B2(n19151), .ZN(
        n19143) );
  AOI22_X1 U22308 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19152), .B1(
        n19262), .B2(n19148), .ZN(n19142) );
  OAI211_X1 U22309 ( .C1(n19265), .C2(n19220), .A(n19143), .B(n19142), .ZN(
        P3_U2959) );
  AOI22_X1 U22310 ( .A1(n19266), .A2(n19151), .B1(n19267), .B2(n19148), .ZN(
        n19145) );
  AOI22_X1 U22311 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19152), .B1(
        n19268), .B2(n19180), .ZN(n19144) );
  OAI211_X1 U22312 ( .C1(n19271), .C2(n19220), .A(n19145), .B(n19144), .ZN(
        P3_U2960) );
  AOI22_X1 U22313 ( .A1(n19273), .A2(n19180), .B1(n19272), .B2(n19151), .ZN(
        n19147) );
  AOI22_X1 U22314 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19152), .B1(
        n19274), .B2(n19239), .ZN(n19146) );
  OAI211_X1 U22315 ( .C1(n19277), .C2(n19155), .A(n19147), .B(n19146), .ZN(
        P3_U2961) );
  AOI22_X1 U22316 ( .A1(n19279), .A2(n19180), .B1(n19278), .B2(n19151), .ZN(
        n19150) );
  AOI22_X1 U22317 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19152), .B1(
        n19280), .B2(n19148), .ZN(n19149) );
  OAI211_X1 U22318 ( .C1(n19283), .C2(n19220), .A(n19150), .B(n19149), .ZN(
        P3_U2962) );
  AOI22_X1 U22319 ( .A1(n19205), .A2(n19180), .B1(n19284), .B2(n19151), .ZN(
        n19154) );
  AOI22_X1 U22320 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19152), .B1(
        n19287), .B2(n19239), .ZN(n19153) );
  OAI211_X1 U22321 ( .C1(n19210), .C2(n19155), .A(n19154), .B(n19153), .ZN(
        P3_U2963) );
  NAND2_X1 U22322 ( .A1(n19156), .A2(n19186), .ZN(n21312) );
  INV_X1 U22323 ( .A(n21312), .ZN(n19286) );
  INV_X1 U22324 ( .A(n19157), .ZN(n19161) );
  NAND2_X1 U22325 ( .A1(n19159), .A2(n19158), .ZN(n19160) );
  OAI211_X1 U22326 ( .C1(n19161), .C2(n19160), .A(n21312), .B(n19220), .ZN(
        n19162) );
  OAI211_X1 U22327 ( .C1(n19286), .C2(n19452), .A(n19216), .B(n19162), .ZN(
        n19181) );
  AOI21_X1 U22328 ( .B1(n21312), .B2(n19220), .A(n19163), .ZN(n19179) );
  AOI22_X1 U22329 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19181), .B1(
        n19245), .B2(n19179), .ZN(n19165) );
  AOI22_X1 U22330 ( .A1(n19286), .A2(n19250), .B1(n19213), .B2(n19201), .ZN(
        n19164) );
  OAI211_X1 U22331 ( .C1(n19221), .C2(n19176), .A(n19165), .B(n19164), .ZN(
        P3_U2964) );
  AOI22_X1 U22332 ( .A1(n19256), .A2(n19201), .B1(n19254), .B2(n19179), .ZN(
        n19167) );
  AOI22_X1 U22333 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19181), .B1(
        n19255), .B2(n19180), .ZN(n19166) );
  OAI211_X1 U22334 ( .C1(n21312), .C2(n19259), .A(n19167), .B(n19166), .ZN(
        P3_U2965) );
  AOI22_X1 U22335 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19181), .B1(
        n21304), .B2(n19179), .ZN(n19169) );
  AOI22_X1 U22336 ( .A1(n19224), .A2(n19180), .B1(n21307), .B2(n19201), .ZN(
        n19168) );
  OAI211_X1 U22337 ( .C1(n21312), .C2(n21310), .A(n19169), .B(n19168), .ZN(
        P3_U2966) );
  AOI22_X1 U22338 ( .A1(n19261), .A2(n19201), .B1(n19260), .B2(n19179), .ZN(
        n19171) );
  AOI22_X1 U22339 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19181), .B1(
        n19262), .B2(n19180), .ZN(n19170) );
  OAI211_X1 U22340 ( .C1(n21312), .C2(n19265), .A(n19171), .B(n19170), .ZN(
        P3_U2967) );
  AOI22_X1 U22341 ( .A1(n19268), .A2(n19201), .B1(n19266), .B2(n19179), .ZN(
        n19173) );
  AOI22_X1 U22342 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19181), .B1(
        n19267), .B2(n19180), .ZN(n19172) );
  OAI211_X1 U22343 ( .C1(n21312), .C2(n19271), .A(n19173), .B(n19172), .ZN(
        P3_U2968) );
  AOI22_X1 U22344 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19181), .B1(
        n19272), .B2(n19179), .ZN(n19175) );
  AOI22_X1 U22345 ( .A1(n19286), .A2(n19274), .B1(n19273), .B2(n19201), .ZN(
        n19174) );
  OAI211_X1 U22346 ( .C1(n19277), .C2(n19176), .A(n19175), .B(n19174), .ZN(
        P3_U2969) );
  AOI22_X1 U22347 ( .A1(n19280), .A2(n19180), .B1(n19278), .B2(n19179), .ZN(
        n19178) );
  AOI22_X1 U22348 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19181), .B1(
        n19279), .B2(n19201), .ZN(n19177) );
  OAI211_X1 U22349 ( .C1(n21312), .C2(n19283), .A(n19178), .B(n19177), .ZN(
        P3_U2970) );
  AOI22_X1 U22350 ( .A1(n19285), .A2(n19180), .B1(n19284), .B2(n19179), .ZN(
        n19183) );
  AOI22_X1 U22351 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19181), .B1(
        n19286), .B2(n19287), .ZN(n19182) );
  OAI211_X1 U22352 ( .C1(n19291), .C2(n19209), .A(n19183), .B(n19182), .ZN(
        P3_U2971) );
  NOR2_X1 U22353 ( .A1(n19212), .A2(n19184), .ZN(n19204) );
  AOI22_X1 U22354 ( .A1(n19246), .A2(n19201), .B1(n19245), .B2(n19204), .ZN(
        n19190) );
  AOI22_X1 U22355 ( .A1(n19188), .A2(n19187), .B1(n19186), .B2(n19185), .ZN(
        n19206) );
  AOI22_X1 U22356 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19206), .B1(
        n21306), .B2(n19250), .ZN(n19189) );
  OAI211_X1 U22357 ( .C1(n19253), .C2(n19220), .A(n19190), .B(n19189), .ZN(
        P3_U2972) );
  AOI22_X1 U22358 ( .A1(n19256), .A2(n19239), .B1(n19254), .B2(n19204), .ZN(
        n19192) );
  AOI22_X1 U22359 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19206), .B1(
        n19255), .B2(n19201), .ZN(n19191) );
  OAI211_X1 U22360 ( .C1(n19292), .C2(n19259), .A(n19192), .B(n19191), .ZN(
        P3_U2973) );
  AOI22_X1 U22361 ( .A1(n19224), .A2(n19201), .B1(n21304), .B2(n19204), .ZN(
        n19194) );
  AOI22_X1 U22362 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19206), .B1(
        n21307), .B2(n19239), .ZN(n19193) );
  OAI211_X1 U22363 ( .C1(n21310), .C2(n19292), .A(n19194), .B(n19193), .ZN(
        P3_U2974) );
  AOI22_X1 U22364 ( .A1(n19261), .A2(n19239), .B1(n19260), .B2(n19204), .ZN(
        n19196) );
  AOI22_X1 U22365 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19206), .B1(
        n19262), .B2(n19201), .ZN(n19195) );
  OAI211_X1 U22366 ( .C1(n19292), .C2(n19265), .A(n19196), .B(n19195), .ZN(
        P3_U2975) );
  AOI22_X1 U22367 ( .A1(n19266), .A2(n19204), .B1(n19267), .B2(n19201), .ZN(
        n19198) );
  AOI22_X1 U22368 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19206), .B1(
        n19268), .B2(n19239), .ZN(n19197) );
  OAI211_X1 U22369 ( .C1(n19292), .C2(n19271), .A(n19198), .B(n19197), .ZN(
        P3_U2976) );
  AOI22_X1 U22370 ( .A1(n19231), .A2(n19201), .B1(n19272), .B2(n19204), .ZN(
        n19200) );
  AOI22_X1 U22371 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19206), .B1(
        n21306), .B2(n19274), .ZN(n19199) );
  OAI211_X1 U22372 ( .C1(n19234), .C2(n19220), .A(n19200), .B(n19199), .ZN(
        P3_U2977) );
  AOI22_X1 U22373 ( .A1(n19280), .A2(n19201), .B1(n19278), .B2(n19204), .ZN(
        n19203) );
  AOI22_X1 U22374 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19206), .B1(
        n19279), .B2(n19239), .ZN(n19202) );
  OAI211_X1 U22375 ( .C1(n19292), .C2(n19283), .A(n19203), .B(n19202), .ZN(
        P3_U2978) );
  AOI22_X1 U22376 ( .A1(n19205), .A2(n19239), .B1(n19284), .B2(n19204), .ZN(
        n19208) );
  AOI22_X1 U22377 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19206), .B1(
        n21306), .B2(n19287), .ZN(n19207) );
  OAI211_X1 U22378 ( .C1(n19210), .C2(n19209), .A(n19208), .B(n19207), .ZN(
        P3_U2979) );
  NOR2_X1 U22379 ( .A1(n19212), .A2(n19211), .ZN(n19238) );
  AOI22_X1 U22380 ( .A1(n19286), .A2(n19213), .B1(n19245), .B2(n19238), .ZN(
        n19219) );
  NOR2_X1 U22381 ( .A1(n19286), .A2(n19239), .ZN(n19215) );
  AOI221_X1 U22382 ( .B1(n19215), .B2(n19292), .C1(n19214), .C2(n19292), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19217) );
  OAI21_X1 U22383 ( .B1(n19240), .B2(n19217), .A(n19216), .ZN(n19241) );
  AOI22_X1 U22384 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19241), .B1(
        n19250), .B2(n19240), .ZN(n19218) );
  OAI211_X1 U22385 ( .C1(n19221), .C2(n19220), .A(n19219), .B(n19218), .ZN(
        P3_U2980) );
  AOI22_X1 U22386 ( .A1(n19286), .A2(n19256), .B1(n19254), .B2(n19238), .ZN(
        n19223) );
  AOI22_X1 U22387 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19241), .B1(
        n19255), .B2(n19239), .ZN(n19222) );
  OAI211_X1 U22388 ( .C1(n19237), .C2(n19259), .A(n19223), .B(n19222), .ZN(
        P3_U2981) );
  AOI22_X1 U22389 ( .A1(n19286), .A2(n21307), .B1(n21304), .B2(n19238), .ZN(
        n19226) );
  AOI22_X1 U22390 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19241), .B1(
        n19224), .B2(n19239), .ZN(n19225) );
  OAI211_X1 U22391 ( .C1(n21310), .C2(n19237), .A(n19226), .B(n19225), .ZN(
        P3_U2982) );
  AOI22_X1 U22392 ( .A1(n19286), .A2(n19261), .B1(n19260), .B2(n19238), .ZN(
        n19228) );
  AOI22_X1 U22393 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19241), .B1(
        n19262), .B2(n19239), .ZN(n19227) );
  OAI211_X1 U22394 ( .C1(n19237), .C2(n19265), .A(n19228), .B(n19227), .ZN(
        P3_U2983) );
  AOI22_X1 U22395 ( .A1(n19286), .A2(n19268), .B1(n19266), .B2(n19238), .ZN(
        n19230) );
  AOI22_X1 U22396 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19241), .B1(
        n19267), .B2(n19239), .ZN(n19229) );
  OAI211_X1 U22397 ( .C1(n19237), .C2(n19271), .A(n19230), .B(n19229), .ZN(
        P3_U2984) );
  AOI22_X1 U22398 ( .A1(n19231), .A2(n19239), .B1(n19272), .B2(n19238), .ZN(
        n19233) );
  AOI22_X1 U22399 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19274), .ZN(n19232) );
  OAI211_X1 U22400 ( .C1(n21312), .C2(n19234), .A(n19233), .B(n19232), .ZN(
        P3_U2985) );
  AOI22_X1 U22401 ( .A1(n19280), .A2(n19239), .B1(n19278), .B2(n19238), .ZN(
        n19236) );
  AOI22_X1 U22402 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19241), .B1(
        n19286), .B2(n19279), .ZN(n19235) );
  OAI211_X1 U22403 ( .C1(n19237), .C2(n19283), .A(n19236), .B(n19235), .ZN(
        P3_U2986) );
  AOI22_X1 U22404 ( .A1(n19285), .A2(n19239), .B1(n19284), .B2(n19238), .ZN(
        n19243) );
  AOI22_X1 U22405 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19287), .ZN(n19242) );
  OAI211_X1 U22406 ( .C1(n21312), .C2(n19291), .A(n19243), .B(n19242), .ZN(
        P3_U2987) );
  NOR2_X1 U22407 ( .A1(n19326), .A2(n19244), .ZN(n19248) );
  AND2_X1 U22408 ( .A1(n19248), .A2(n19350), .ZN(n21305) );
  AOI22_X1 U22409 ( .A1(n19286), .A2(n19246), .B1(n21305), .B2(n19245), .ZN(
        n19252) );
  AOI21_X1 U22410 ( .B1(n19249), .B2(n19248), .A(n19247), .ZN(n21315) );
  AOI22_X1 U22411 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21315), .B1(
        n19288), .B2(n19250), .ZN(n19251) );
  OAI211_X1 U22412 ( .C1(n19292), .C2(n19253), .A(n19252), .B(n19251), .ZN(
        P3_U2988) );
  AOI22_X1 U22413 ( .A1(n19286), .A2(n19255), .B1(n21305), .B2(n19254), .ZN(
        n19258) );
  AOI22_X1 U22414 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21315), .B1(
        n21306), .B2(n19256), .ZN(n19257) );
  OAI211_X1 U22415 ( .C1(n21309), .C2(n19259), .A(n19258), .B(n19257), .ZN(
        P3_U2989) );
  AOI22_X1 U22416 ( .A1(n21306), .A2(n19261), .B1(n21305), .B2(n19260), .ZN(
        n19264) );
  AOI22_X1 U22417 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21315), .B1(
        n19286), .B2(n19262), .ZN(n19263) );
  OAI211_X1 U22418 ( .C1(n21309), .C2(n19265), .A(n19264), .B(n19263), .ZN(
        P3_U2991) );
  AOI22_X1 U22419 ( .A1(n19286), .A2(n19267), .B1(n21305), .B2(n19266), .ZN(
        n19270) );
  AOI22_X1 U22420 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21315), .B1(
        n21306), .B2(n19268), .ZN(n19269) );
  OAI211_X1 U22421 ( .C1(n21309), .C2(n19271), .A(n19270), .B(n19269), .ZN(
        P3_U2992) );
  AOI22_X1 U22422 ( .A1(n21306), .A2(n19273), .B1(n21305), .B2(n19272), .ZN(
        n19276) );
  AOI22_X1 U22423 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21315), .B1(
        n19288), .B2(n19274), .ZN(n19275) );
  OAI211_X1 U22424 ( .C1(n21312), .C2(n19277), .A(n19276), .B(n19275), .ZN(
        P3_U2993) );
  AOI22_X1 U22425 ( .A1(n21306), .A2(n19279), .B1(n21305), .B2(n19278), .ZN(
        n19282) );
  AOI22_X1 U22426 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21315), .B1(
        n19286), .B2(n19280), .ZN(n19281) );
  OAI211_X1 U22427 ( .C1(n21309), .C2(n19283), .A(n19282), .B(n19281), .ZN(
        P3_U2994) );
  AOI22_X1 U22428 ( .A1(n19286), .A2(n19285), .B1(n21305), .B2(n19284), .ZN(
        n19290) );
  AOI22_X1 U22429 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21315), .B1(
        n19288), .B2(n19287), .ZN(n19289) );
  OAI211_X1 U22430 ( .C1(n19292), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P3_U2995) );
  OAI22_X1 U22431 ( .A1(n19296), .A2(n19295), .B1(n19294), .B2(n19293), .ZN(
        n19297) );
  AOI221_X1 U22432 ( .B1(n19300), .B2(n19299), .C1(n19298), .C2(n19299), .A(
        n19297), .ZN(n19464) );
  AOI211_X1 U22433 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19319), .A(
        n19302), .B(n19301), .ZN(n19336) );
  INV_X1 U22434 ( .A(n19319), .ZN(n19310) );
  NAND2_X1 U22435 ( .A1(n19310), .A2(n19303), .ZN(n19307) );
  INV_X1 U22436 ( .A(n19304), .ZN(n19305) );
  NOR2_X1 U22437 ( .A1(n19305), .A2(n19319), .ZN(n19306) );
  MUX2_X1 U22438 ( .A(n19307), .B(n19306), .S(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19329) );
  INV_X1 U22439 ( .A(n19329), .ZN(n19332) );
  INV_X1 U22440 ( .A(n19312), .ZN(n19308) );
  NOR2_X1 U22441 ( .A1(n19309), .A2(n19308), .ZN(n19315) );
  OAI21_X1 U22442 ( .B1(n19312), .B2(n19311), .A(n19310), .ZN(n19313) );
  INV_X1 U22443 ( .A(n19313), .ZN(n19314) );
  OAI21_X1 U22444 ( .B1(n19316), .B2(n19315), .A(n19314), .ZN(n19318) );
  AND2_X1 U22445 ( .A1(n19318), .A2(n19317), .ZN(n19321) );
  INV_X1 U22446 ( .A(n19321), .ZN(n19323) );
  MUX2_X1 U22447 ( .A(n19320), .B(n9896), .S(n19319), .Z(n19324) );
  AOI21_X1 U22448 ( .B1(n19321), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n19324), .ZN(n19322) );
  AOI21_X1 U22449 ( .B1(n18865), .B2(n19323), .A(n19322), .ZN(n19330) );
  INV_X1 U22450 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19327) );
  INV_X1 U22451 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19326) );
  INV_X1 U22452 ( .A(n19324), .ZN(n19325) );
  AOI21_X1 U22453 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19328) );
  OAI22_X1 U22454 ( .A1(n19330), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n19329), .B2(n19328), .ZN(n19331) );
  OAI21_X1 U22455 ( .B1(n19326), .B2(n19332), .A(n19331), .ZN(n19335) );
  OAI21_X1 U22456 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19333), .ZN(n19334) );
  NAND4_X1 U22457 ( .A1(n19464), .A2(n19336), .A3(n19335), .A4(n19334), .ZN(
        n19345) );
  AOI211_X1 U22458 ( .C1(n19339), .C2(n19338), .A(n19337), .B(n19345), .ZN(
        n19447) );
  AOI21_X1 U22459 ( .B1(n19473), .B2(n19472), .A(n19447), .ZN(n19351) );
  INV_X1 U22460 ( .A(n19340), .ZN(n19347) );
  NOR2_X1 U22461 ( .A1(n19349), .A2(n19350), .ZN(n19344) );
  NOR2_X1 U22462 ( .A1(n19466), .A2(n19341), .ZN(n19348) );
  AOI211_X1 U22463 ( .C1(n19342), .C2(n19478), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n19348), .ZN(n19343) );
  AOI211_X1 U22464 ( .C1(n19469), .C2(n19345), .A(n19344), .B(n19343), .ZN(
        n19346) );
  OAI221_X1 U22465 ( .B1(n19475), .B2(n19351), .C1(n19475), .C2(n19347), .A(
        n19346), .ZN(P3_U2996) );
  INV_X1 U22466 ( .A(n19348), .ZN(n19354) );
  NAND4_X1 U22467 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19473), .A4(n19472), .ZN(n19357) );
  INV_X1 U22468 ( .A(n19349), .ZN(n19352) );
  NAND3_X1 U22469 ( .A1(n19352), .A2(n19351), .A3(n19350), .ZN(n19353) );
  NAND4_X1 U22470 ( .A1(n19355), .A2(n19354), .A3(n19357), .A4(n19353), .ZN(
        P3_U2997) );
  OAI21_X1 U22471 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19356), .ZN(n19359) );
  INV_X1 U22472 ( .A(n19357), .ZN(n19358) );
  AOI21_X1 U22473 ( .B1(n19360), .B2(n19359), .A(n19358), .ZN(P3_U2998) );
  AND2_X1 U22474 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19443), .ZN(
        P3_U2999) );
  AND2_X1 U22475 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19443), .ZN(
        P3_U3000) );
  AND2_X1 U22476 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19443), .ZN(
        P3_U3001) );
  AND2_X1 U22477 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19443), .ZN(
        P3_U3002) );
  AND2_X1 U22478 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19443), .ZN(
        P3_U3003) );
  AND2_X1 U22479 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19443), .ZN(
        P3_U3004) );
  AND2_X1 U22480 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19443), .ZN(
        P3_U3005) );
  INV_X1 U22481 ( .A(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21376) );
  NOR2_X1 U22482 ( .A1(n21376), .A2(n19446), .ZN(P3_U3006) );
  AND2_X1 U22483 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19443), .ZN(
        P3_U3007) );
  AND2_X1 U22484 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19443), .ZN(
        P3_U3008) );
  AND2_X1 U22485 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19443), .ZN(
        P3_U3009) );
  AND2_X1 U22486 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19443), .ZN(
        P3_U3010) );
  AND2_X1 U22487 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19443), .ZN(
        P3_U3011) );
  AND2_X1 U22488 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19443), .ZN(
        P3_U3012) );
  AND2_X1 U22489 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19443), .ZN(
        P3_U3013) );
  AND2_X1 U22490 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19443), .ZN(
        P3_U3014) );
  AND2_X1 U22491 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19443), .ZN(
        P3_U3015) );
  AND2_X1 U22492 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19443), .ZN(
        P3_U3016) );
  AND2_X1 U22493 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19443), .ZN(
        P3_U3017) );
  AND2_X1 U22494 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19443), .ZN(
        P3_U3018) );
  AND2_X1 U22495 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19443), .ZN(
        P3_U3019) );
  AND2_X1 U22496 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19443), .ZN(
        P3_U3020) );
  AND2_X1 U22497 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19443), .ZN(P3_U3021) );
  AND2_X1 U22498 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19443), .ZN(P3_U3022) );
  AND2_X1 U22499 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19443), .ZN(P3_U3023) );
  AND2_X1 U22500 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19443), .ZN(P3_U3024) );
  AND2_X1 U22501 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19443), .ZN(P3_U3025) );
  AND2_X1 U22502 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19443), .ZN(P3_U3026) );
  AND2_X1 U22503 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19443), .ZN(P3_U3027) );
  AND2_X1 U22504 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19443), .ZN(P3_U3028) );
  OAI21_X1 U22505 ( .B1(n19361), .B2(n21254), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19362) );
  AOI22_X1 U22506 ( .A1(n19373), .A2(n19375), .B1(n19482), .B2(n19362), .ZN(
        n19363) );
  INV_X1 U22507 ( .A(NA), .ZN(n21248) );
  OR3_X1 U22508 ( .A1(n21248), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n19368) );
  OAI211_X1 U22509 ( .C1(n19466), .C2(n19364), .A(n19363), .B(n19368), .ZN(
        P3_U3029) );
  INV_X1 U22510 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19480) );
  NOR2_X1 U22511 ( .A1(n19375), .A2(n21254), .ZN(n19371) );
  OAI22_X1 U22512 ( .A1(n19480), .A2(n19371), .B1(n21254), .B2(n19364), .ZN(
        n19365) );
  INV_X1 U22513 ( .A(n19365), .ZN(n19367) );
  NAND2_X1 U22514 ( .A1(n19473), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19369) );
  OAI211_X1 U22515 ( .C1(n19367), .C2(n19373), .A(n19369), .B(n19366), .ZN(
        P3_U3030) );
  AOI22_X1 U22516 ( .A1(n19473), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n19373), 
        .B2(n19368), .ZN(n19374) );
  OAI22_X1 U22517 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19369), .ZN(n19370) );
  OAI22_X1 U22518 ( .A1(n19371), .A2(n19370), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19372) );
  OAI22_X1 U22519 ( .A1(n19374), .A2(n19375), .B1(n19373), .B2(n19372), .ZN(
        P3_U3031) );
  OAI222_X1 U22520 ( .A1(n18551), .A2(n9610), .B1(n19376), .B2(n19434), .C1(
        n19377), .C2(n19421), .ZN(P3_U3032) );
  OAI222_X1 U22521 ( .A1(n19421), .A2(n19380), .B1(n19378), .B2(n19434), .C1(
        n19377), .C2(n9610), .ZN(P3_U3033) );
  OAI222_X1 U22522 ( .A1(n19421), .A2(n19382), .B1(n19381), .B2(n19434), .C1(
        n19380), .C2(n9610), .ZN(P3_U3034) );
  OAI222_X1 U22523 ( .A1(n19421), .A2(n19385), .B1(n19383), .B2(n19434), .C1(
        n19382), .C2(n9610), .ZN(P3_U3035) );
  OAI222_X1 U22524 ( .A1(n19385), .A2(n9610), .B1(n19384), .B2(n19434), .C1(
        n19386), .C2(n19421), .ZN(P3_U3036) );
  OAI222_X1 U22525 ( .A1(n19421), .A2(n19388), .B1(n19387), .B2(n19434), .C1(
        n19386), .C2(n9610), .ZN(P3_U3037) );
  OAI222_X1 U22526 ( .A1(n19421), .A2(n19391), .B1(n19389), .B2(n19434), .C1(
        n19388), .C2(n9610), .ZN(P3_U3038) );
  OAI222_X1 U22527 ( .A1(n19391), .A2(n9610), .B1(n19390), .B2(n19434), .C1(
        n19392), .C2(n19421), .ZN(P3_U3039) );
  OAI222_X1 U22528 ( .A1(n19421), .A2(n19394), .B1(n19393), .B2(n19434), .C1(
        n19392), .C2(n9610), .ZN(P3_U3040) );
  OAI222_X1 U22529 ( .A1(n19421), .A2(n19396), .B1(n19395), .B2(n19434), .C1(
        n19394), .C2(n9610), .ZN(P3_U3041) );
  INV_X1 U22530 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19398) );
  OAI222_X1 U22531 ( .A1(n19421), .A2(n19398), .B1(n19397), .B2(n19434), .C1(
        n19396), .C2(n9610), .ZN(P3_U3042) );
  OAI222_X1 U22532 ( .A1(n19421), .A2(n19400), .B1(n19399), .B2(n19434), .C1(
        n19398), .C2(n9610), .ZN(P3_U3043) );
  OAI222_X1 U22533 ( .A1(n19421), .A2(n19402), .B1(n19401), .B2(n19434), .C1(
        n19400), .C2(n9610), .ZN(P3_U3044) );
  OAI222_X1 U22534 ( .A1(n19421), .A2(n19404), .B1(n19403), .B2(n19434), .C1(
        n19402), .C2(n9610), .ZN(P3_U3045) );
  OAI222_X1 U22535 ( .A1(n19421), .A2(n19406), .B1(n19405), .B2(n19434), .C1(
        n19404), .C2(n9610), .ZN(P3_U3046) );
  OAI222_X1 U22536 ( .A1(n19421), .A2(n19408), .B1(n19407), .B2(n19434), .C1(
        n19406), .C2(n9610), .ZN(P3_U3047) );
  OAI222_X1 U22537 ( .A1(n19421), .A2(n19410), .B1(n19409), .B2(n19434), .C1(
        n19408), .C2(n9610), .ZN(P3_U3048) );
  OAI222_X1 U22538 ( .A1(n19421), .A2(n19412), .B1(n19411), .B2(n19434), .C1(
        n19410), .C2(n9610), .ZN(P3_U3049) );
  INV_X1 U22539 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19415) );
  OAI222_X1 U22540 ( .A1(n19421), .A2(n19415), .B1(n19413), .B2(n19434), .C1(
        n19412), .C2(n9610), .ZN(P3_U3050) );
  OAI222_X1 U22541 ( .A1(n19415), .A2(n9610), .B1(n19414), .B2(n19434), .C1(
        n21391), .C2(n19421), .ZN(P3_U3051) );
  INV_X1 U22542 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19417) );
  OAI222_X1 U22543 ( .A1(n21391), .A2(n9610), .B1(n19416), .B2(n19434), .C1(
        n19417), .C2(n19421), .ZN(P3_U3052) );
  OAI222_X1 U22544 ( .A1(n19421), .A2(n19419), .B1(n19418), .B2(n19434), .C1(
        n19417), .C2(n9610), .ZN(P3_U3053) );
  OAI222_X1 U22545 ( .A1(n19421), .A2(n19423), .B1(n19420), .B2(n19434), .C1(
        n19419), .C2(n9610), .ZN(P3_U3054) );
  OAI222_X1 U22546 ( .A1(n19423), .A2(n9610), .B1(n19422), .B2(n19434), .C1(
        n21348), .C2(n19421), .ZN(P3_U3055) );
  OAI222_X1 U22547 ( .A1(n21348), .A2(n9610), .B1(n19424), .B2(n19434), .C1(
        n19426), .C2(n19421), .ZN(P3_U3056) );
  OAI222_X1 U22548 ( .A1(n19426), .A2(n9610), .B1(n19425), .B2(n19434), .C1(
        n19427), .C2(n19421), .ZN(P3_U3057) );
  INV_X1 U22549 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19430) );
  OAI222_X1 U22550 ( .A1(n19421), .A2(n19430), .B1(n19428), .B2(n19434), .C1(
        n19427), .C2(n9610), .ZN(P3_U3058) );
  OAI222_X1 U22551 ( .A1(n19430), .A2(n9610), .B1(n19429), .B2(n19434), .C1(
        n19431), .C2(n19421), .ZN(P3_U3059) );
  OAI222_X1 U22552 ( .A1(n19421), .A2(n19436), .B1(n19432), .B2(n19434), .C1(
        n19431), .C2(n9610), .ZN(P3_U3060) );
  OAI222_X1 U22553 ( .A1(n9610), .A2(n19436), .B1(n19435), .B2(n19434), .C1(
        n19433), .C2(n19421), .ZN(P3_U3061) );
  MUX2_X1 U22554 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n19434), .Z(P3_U3274) );
  INV_X1 U22555 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19437) );
  INV_X1 U22556 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n21335) );
  AOI22_X1 U22557 ( .A1(n19434), .A2(n19437), .B1(n21335), .B2(n19482), .ZN(
        P3_U3275) );
  INV_X1 U22558 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19438) );
  AOI22_X1 U22559 ( .A1(n19434), .A2(n19439), .B1(n19438), .B2(n19482), .ZN(
        P3_U3276) );
  INV_X1 U22560 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19460) );
  INV_X1 U22561 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19440) );
  AOI22_X1 U22562 ( .A1(n19434), .A2(n19460), .B1(n19440), .B2(n19482), .ZN(
        P3_U3277) );
  INV_X1 U22563 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19442) );
  INV_X1 U22564 ( .A(n19444), .ZN(n19441) );
  AOI21_X1 U22565 ( .B1(n19443), .B2(n19442), .A(n19441), .ZN(P3_U3280) );
  INV_X1 U22566 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22567 ( .B1(n19446), .B2(n19445), .A(n19444), .ZN(P3_U3281) );
  INV_X1 U22568 ( .A(n19447), .ZN(n19451) );
  NOR2_X1 U22569 ( .A1(n19449), .A2(n19448), .ZN(n19450) );
  OAI21_X1 U22570 ( .B1(n19452), .B2(n19451), .A(n19450), .ZN(P3_U3282) );
  INV_X1 U22571 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19458) );
  AOI211_X1 U22572 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_REIP_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19453) );
  INV_X1 U22573 ( .A(n19454), .ZN(n19459) );
  AOI22_X1 U22574 ( .A1(n19454), .A2(n19453), .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n19459), .ZN(n19455) );
  OAI21_X1 U22575 ( .B1(n19458), .B2(n19456), .A(n19455), .ZN(P3_U3292) );
  NOR2_X1 U22576 ( .A1(n19459), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19457) );
  AOI22_X1 U22577 ( .A1(n19460), .A2(n19459), .B1(n19458), .B2(n19457), .ZN(
        P3_U3293) );
  INV_X1 U22578 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19461) );
  AOI22_X1 U22579 ( .A1(n19434), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19461), 
        .B2(n19482), .ZN(P3_U3294) );
  INV_X1 U22580 ( .A(n19462), .ZN(n19465) );
  NAND2_X1 U22581 ( .A1(n19465), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19463) );
  OAI21_X1 U22582 ( .B1(n19465), .B2(n19464), .A(n19463), .ZN(P3_U3295) );
  AOI21_X1 U22583 ( .B1(n18184), .B2(n19466), .A(n19487), .ZN(n19467) );
  OAI21_X1 U22584 ( .B1(n19469), .B2(n19468), .A(n19467), .ZN(n19481) );
  OAI21_X1 U22585 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19471), .A(n19470), 
        .ZN(n19474) );
  AOI211_X1 U22586 ( .C1(n19485), .C2(n19474), .A(n19473), .B(n19472), .ZN(
        n19476) );
  NOR2_X1 U22587 ( .A1(n19476), .A2(n19475), .ZN(n19477) );
  OAI21_X1 U22588 ( .B1(n19478), .B2(n19477), .A(n19481), .ZN(n19479) );
  OAI21_X1 U22589 ( .B1(n19481), .B2(n19480), .A(n19479), .ZN(P3_U3296) );
  INV_X1 U22590 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n21410) );
  INV_X1 U22591 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19483) );
  AOI22_X1 U22592 ( .A1(n19434), .A2(n21410), .B1(n19483), .B2(n19482), .ZN(
        P3_U3297) );
  OAI21_X1 U22593 ( .B1(n19488), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19486), 
        .ZN(n19484) );
  OAI21_X1 U22594 ( .B1(n19486), .B2(n19485), .A(n19484), .ZN(P3_U3298) );
  NOR3_X1 U22595 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n19488), .A3(n19487), 
        .ZN(n19490) );
  NOR2_X1 U22596 ( .A1(n19490), .A2(n19489), .ZN(P3_U3299) );
  INV_X1 U22597 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20211) );
  INV_X1 U22598 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19491) );
  NAND2_X1 U22599 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20231), .ZN(n20221) );
  NAND2_X1 U22600 ( .A1(n20211), .A2(n19492), .ZN(n20218) );
  OAI21_X1 U22601 ( .B1(n20211), .B2(n20221), .A(n20218), .ZN(n20293) );
  OAI21_X1 U22602 ( .B1(n20211), .B2(n19491), .A(n20210), .ZN(P2_U2815) );
  INV_X2 U22603 ( .A(n20336), .ZN(n20347) );
  AOI22_X1 U22604 ( .A1(n20347), .A2(n19493), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20336), .ZN(n19494) );
  OAI21_X1 U22605 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20226), .A(n19494), 
        .ZN(P2_U2817) );
  OAI21_X1 U22606 ( .B1(n20213), .B2(BS16), .A(n20293), .ZN(n20291) );
  OAI21_X1 U22607 ( .B1(n20293), .B2(n16495), .A(n20291), .ZN(P2_U2818) );
  NOR4_X1 U22608 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19504) );
  NOR4_X1 U22609 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19503) );
  AOI211_X1 U22610 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_29__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19495) );
  INV_X1 U22611 ( .A(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21346) );
  INV_X1 U22612 ( .A(P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21352) );
  NAND3_X1 U22613 ( .A1(n19495), .A2(n21346), .A3(n21352), .ZN(n19501) );
  NOR4_X1 U22614 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(n19499) );
  NOR4_X1 U22615 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19498) );
  NOR4_X1 U22616 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19497) );
  NOR4_X1 U22617 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_22__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n19496) );
  NAND4_X1 U22618 ( .A1(n19499), .A2(n19498), .A3(n19497), .A4(n19496), .ZN(
        n19500) );
  NOR4_X1 U22619 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(n19501), .A4(n19500), .ZN(n19502)
         );
  NAND3_X1 U22620 ( .A1(n19504), .A2(n19503), .A3(n19502), .ZN(n19511) );
  NOR2_X1 U22621 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19511), .ZN(n19505) );
  INV_X1 U22622 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21398) );
  AOI22_X1 U22623 ( .A1(n19505), .A2(n19506), .B1(n21398), .B2(n19511), .ZN(
        P2_U2820) );
  OR3_X1 U22624 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19510) );
  INV_X1 U22625 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20288) );
  AOI22_X1 U22626 ( .A1(n19505), .A2(n19510), .B1(n19511), .B2(n20288), .ZN(
        P2_U2821) );
  INV_X1 U22627 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20292) );
  NAND2_X1 U22628 ( .A1(n19505), .A2(n20292), .ZN(n19509) );
  INV_X1 U22629 ( .A(n19511), .ZN(n19512) );
  OAI21_X1 U22630 ( .B1(n20232), .B2(n19506), .A(n19512), .ZN(n19507) );
  OAI21_X1 U22631 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19512), .A(n19507), 
        .ZN(n19508) );
  OAI221_X1 U22632 ( .B1(n19509), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19509), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19508), .ZN(P2_U2822) );
  INV_X1 U22633 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20286) );
  OAI221_X1 U22634 ( .B1(n19512), .B2(n20286), .C1(n19511), .C2(n19510), .A(
        n19509), .ZN(P2_U2823) );
  OAI21_X1 U22635 ( .B1(n19513), .B2(n16142), .A(n16032), .ZN(n19516) );
  NOR2_X1 U22636 ( .A1(n19514), .A2(n19549), .ZN(n19515) );
  AOI211_X1 U22637 ( .C1(n19547), .C2(P2_EBX_REG_12__SCAN_IN), .A(n19516), .B(
        n19515), .ZN(n19526) );
  NAND2_X1 U22638 ( .A1(n19559), .A2(n19517), .ZN(n19519) );
  XNOR2_X1 U22639 ( .A(n19519), .B(n19518), .ZN(n19524) );
  AND2_X1 U22640 ( .A1(n19520), .A2(n19542), .ZN(n19523) );
  NOR2_X1 U22641 ( .A1(n19521), .A2(n19555), .ZN(n19522) );
  AOI211_X1 U22642 ( .C1(n19524), .C2(n19563), .A(n19523), .B(n19522), .ZN(
        n19525) );
  OAI211_X1 U22643 ( .C1(n20250), .C2(n19546), .A(n19526), .B(n19525), .ZN(
        P2_U2843) );
  AOI21_X1 U22644 ( .B1(n19548), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19527), .ZN(n19528) );
  OAI21_X1 U22645 ( .B1(n12352), .B2(n19529), .A(n19528), .ZN(n19530) );
  AOI21_X1 U22646 ( .B1(n19532), .B2(n19531), .A(n19530), .ZN(n19545) );
  NOR2_X1 U22647 ( .A1(n19533), .A2(n19555), .ZN(n19541) );
  NOR2_X1 U22648 ( .A1(n19534), .A2(n19536), .ZN(n19535) );
  MUX2_X1 U22649 ( .A(n19536), .B(n19535), .S(n19559), .Z(n19539) );
  NOR3_X1 U22650 ( .A1(n19539), .A2(n19538), .A3(n19537), .ZN(n19540) );
  AOI211_X1 U22651 ( .C1(n19543), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        n19544) );
  OAI211_X1 U22652 ( .C1(n20239), .C2(n19546), .A(n19545), .B(n19544), .ZN(
        P2_U2849) );
  AOI22_X1 U22653 ( .A1(n19548), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19547), .ZN(n19568) );
  OAI22_X1 U22654 ( .A1(n19649), .A2(n19551), .B1(n19550), .B2(n19549), .ZN(
        n19552) );
  AOI211_X1 U22655 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19554), .A(n19553), .B(
        n19552), .ZN(n19567) );
  INV_X1 U22656 ( .A(n19651), .ZN(n19569) );
  OAI22_X1 U22657 ( .A1(n19580), .A2(n19556), .B1(n19555), .B2(n19569), .ZN(
        n19557) );
  INV_X1 U22658 ( .A(n19557), .ZN(n19566) );
  NAND2_X1 U22659 ( .A1(n19558), .A2(n19561), .ZN(n19560) );
  MUX2_X1 U22660 ( .A(n19561), .B(n19560), .S(n19559), .Z(n19564) );
  NAND3_X1 U22661 ( .A1(n19564), .A2(n19563), .A3(n19562), .ZN(n19565) );
  NAND4_X1 U22662 ( .A1(n19568), .A2(n19567), .A3(n19566), .A4(n19565), .ZN(
        P2_U2851) );
  OAI22_X1 U22663 ( .A1(n19580), .A2(n19571), .B1(n19570), .B2(n19569), .ZN(
        n19572) );
  INV_X1 U22664 ( .A(n19572), .ZN(n19573) );
  OAI21_X1 U22665 ( .B1(n19575), .B2(n19574), .A(n19573), .ZN(P2_U2883) );
  INV_X1 U22666 ( .A(n19649), .ZN(n19579) );
  AOI22_X1 U22667 ( .A1(n19579), .A2(n19578), .B1(n19577), .B2(n19576), .ZN(
        n19585) );
  XNOR2_X1 U22668 ( .A(n19581), .B(n19580), .ZN(n19583) );
  NAND2_X1 U22669 ( .A1(n19583), .A2(n19582), .ZN(n19584) );
  OAI211_X1 U22670 ( .C1(n19586), .C2(n19615), .A(n19585), .B(n19584), .ZN(
        P2_U2915) );
  NOR2_X1 U22671 ( .A1(n19592), .A2(n19587), .ZN(P2_U2920) );
  INV_X1 U22672 ( .A(n19588), .ZN(n19589) );
  AOI22_X1 U22673 ( .A1(n19589), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19623), .ZN(n19590) );
  OAI21_X1 U22674 ( .B1(n19592), .B2(n19591), .A(n19590), .ZN(P2_U2921) );
  AOI22_X1 U22675 ( .A1(n19623), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19593) );
  OAI21_X1 U22676 ( .B1(n13595), .B2(n19625), .A(n19593), .ZN(P2_U2936) );
  INV_X1 U22677 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19595) );
  AOI22_X1 U22678 ( .A1(n19623), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19594) );
  OAI21_X1 U22679 ( .B1(n19595), .B2(n19625), .A(n19594), .ZN(P2_U2937) );
  AOI22_X1 U22680 ( .A1(n19623), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19596) );
  OAI21_X1 U22681 ( .B1(n19597), .B2(n19625), .A(n19596), .ZN(P2_U2938) );
  AOI22_X1 U22682 ( .A1(n19623), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19598) );
  OAI21_X1 U22683 ( .B1(n19599), .B2(n19625), .A(n19598), .ZN(P2_U2939) );
  AOI22_X1 U22684 ( .A1(n19623), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19600) );
  OAI21_X1 U22685 ( .B1(n19601), .B2(n19625), .A(n19600), .ZN(P2_U2940) );
  AOI22_X1 U22686 ( .A1(n19623), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19602) );
  OAI21_X1 U22687 ( .B1(n19603), .B2(n19625), .A(n19602), .ZN(P2_U2941) );
  AOI22_X1 U22688 ( .A1(n19623), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19604) );
  OAI21_X1 U22689 ( .B1(n19605), .B2(n19625), .A(n19604), .ZN(P2_U2942) );
  AOI22_X1 U22690 ( .A1(n19623), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19606) );
  OAI21_X1 U22691 ( .B1(n19607), .B2(n19625), .A(n19606), .ZN(P2_U2943) );
  AOI22_X1 U22692 ( .A1(n19623), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19608) );
  OAI21_X1 U22693 ( .B1(n19609), .B2(n19625), .A(n19608), .ZN(P2_U2944) );
  AOI22_X1 U22694 ( .A1(n19623), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19610) );
  OAI21_X1 U22695 ( .B1(n19611), .B2(n19625), .A(n19610), .ZN(P2_U2945) );
  INV_X1 U22696 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19613) );
  AOI22_X1 U22697 ( .A1(n19623), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19612) );
  OAI21_X1 U22698 ( .B1(n19613), .B2(n19625), .A(n19612), .ZN(P2_U2946) );
  AOI22_X1 U22699 ( .A1(n19623), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19614) );
  OAI21_X1 U22700 ( .B1(n19615), .B2(n19625), .A(n19614), .ZN(P2_U2947) );
  INV_X1 U22701 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19617) );
  AOI22_X1 U22702 ( .A1(n19623), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19616) );
  OAI21_X1 U22703 ( .B1(n19617), .B2(n19625), .A(n19616), .ZN(P2_U2948) );
  AOI22_X1 U22704 ( .A1(n19623), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19618) );
  OAI21_X1 U22705 ( .B1(n19619), .B2(n19625), .A(n19618), .ZN(P2_U2949) );
  AOI22_X1 U22706 ( .A1(n19623), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19620) );
  OAI21_X1 U22707 ( .B1(n19621), .B2(n19625), .A(n19620), .ZN(P2_U2950) );
  AOI22_X1 U22708 ( .A1(n19623), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19622), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19624) );
  OAI21_X1 U22709 ( .B1(n12048), .B2(n19625), .A(n19624), .ZN(P2_U2951) );
  AOI22_X1 U22710 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19630), .B1(n19626), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19629) );
  NAND2_X1 U22711 ( .A1(n19628), .A2(n19627), .ZN(n19631) );
  NAND2_X1 U22712 ( .A1(n19629), .A2(n19631), .ZN(P2_U2966) );
  AOI22_X1 U22713 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19630), .B1(n13574), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19632) );
  NAND2_X1 U22714 ( .A1(n19632), .A2(n19631), .ZN(P2_U2981) );
  NOR2_X1 U22715 ( .A1(n19634), .A2(n19633), .ZN(n19646) );
  INV_X1 U22716 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19645) );
  NAND2_X1 U22717 ( .A1(n19636), .A2(n19635), .ZN(n19637) );
  OAI211_X1 U22718 ( .C1(n19640), .C2(n19639), .A(n19638), .B(n19637), .ZN(
        n19641) );
  AOI21_X1 U22719 ( .B1(n19643), .B2(n19642), .A(n19641), .ZN(n19644) );
  OAI21_X1 U22720 ( .B1(n19646), .B2(n19645), .A(n19644), .ZN(P2_U3014) );
  OAI21_X1 U22721 ( .B1(n19649), .B2(n19648), .A(n19647), .ZN(n19650) );
  AOI21_X1 U22722 ( .B1(n19651), .B2(n19669), .A(n19650), .ZN(n19652) );
  OAI21_X1 U22723 ( .B1(n19654), .B2(n19653), .A(n19652), .ZN(n19655) );
  AOI21_X1 U22724 ( .B1(n19657), .B2(n19656), .A(n19655), .ZN(n19658) );
  OAI221_X1 U22725 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19661), .C1(
        n19660), .C2(n19659), .A(n19658), .ZN(P2_U3042) );
  INV_X1 U22726 ( .A(n19662), .ZN(n19679) );
  AOI21_X1 U22727 ( .B1(n19665), .B2(n19664), .A(n19663), .ZN(n19666) );
  OAI21_X1 U22728 ( .B1(n19668), .B2(n19667), .A(n19666), .ZN(n19678) );
  NAND2_X1 U22729 ( .A1(n12404), .A2(n19669), .ZN(n19674) );
  NAND3_X1 U22730 ( .A1(n19672), .A2(n19671), .A3(n19670), .ZN(n19673) );
  OAI211_X1 U22731 ( .C1(n19676), .C2(n19675), .A(n19674), .B(n19673), .ZN(
        n19677) );
  AOI211_X1 U22732 ( .C1(n19679), .C2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n19678), .B(n19677), .ZN(n19681) );
  OAI211_X1 U22733 ( .C1(n19683), .C2(n19682), .A(n19681), .B(n19680), .ZN(
        P2_U3044) );
  INV_X1 U22734 ( .A(n19687), .ZN(n19686) );
  INV_X1 U22735 ( .A(n19684), .ZN(n19879) );
  NOR2_X1 U22736 ( .A1(n19808), .A2(n19746), .ZN(n19709) );
  NOR3_X1 U22737 ( .A1(n19685), .A2(n19709), .A3(n20145), .ZN(n19688) );
  AOI211_X2 U22738 ( .C1(n20145), .C2(n19686), .A(n19879), .B(n19688), .ZN(
        n19710) );
  AOI22_X1 U22739 ( .A1(n19710), .A2(n20150), .B1(n20149), .B2(n19709), .ZN(
        n19694) );
  INV_X1 U22740 ( .A(n19942), .ZN(n19933) );
  AOI21_X1 U22741 ( .B1(n19872), .B2(n19933), .A(n19687), .ZN(n19689) );
  NOR2_X1 U22742 ( .A1(n19689), .A2(n19688), .ZN(n19690) );
  OAI211_X1 U22743 ( .C1(n19709), .C2(n20318), .A(n19690), .B(n20152), .ZN(
        n19712) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20159), .ZN(n19693) );
  OAI211_X1 U22745 ( .C1(n20162), .C2(n19707), .A(n19694), .B(n19693), .ZN(
        P2_U3056) );
  AOI22_X1 U22746 ( .A1(n19710), .A2(n20164), .B1(n19709), .B2(n20163), .ZN(
        n19696) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20165), .ZN(n19695) );
  OAI211_X1 U22748 ( .C1(n20168), .C2(n19707), .A(n19696), .B(n19695), .ZN(
        P2_U3057) );
  AOI22_X1 U22749 ( .A1(n19710), .A2(n20170), .B1(n20169), .B2(n19709), .ZN(
        n19698) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20171), .ZN(n19697) );
  OAI211_X1 U22751 ( .C1(n20174), .C2(n19707), .A(n19698), .B(n19697), .ZN(
        P2_U3058) );
  AOI22_X1 U22752 ( .A1(n19710), .A2(n20176), .B1(n19709), .B2(n20175), .ZN(
        n19700) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20177), .ZN(n19699) );
  OAI211_X1 U22754 ( .C1(n20180), .C2(n19707), .A(n19700), .B(n19699), .ZN(
        P2_U3059) );
  AOI22_X1 U22755 ( .A1(n19710), .A2(n20182), .B1(n20181), .B2(n19709), .ZN(
        n19702) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20183), .ZN(n19701) );
  OAI211_X1 U22757 ( .C1(n20186), .C2(n19707), .A(n19702), .B(n19701), .ZN(
        P2_U3060) );
  AOI22_X1 U22758 ( .A1(n19710), .A2(n20188), .B1(n19709), .B2(n20187), .ZN(
        n19704) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20189), .ZN(n19703) );
  OAI211_X1 U22760 ( .C1(n20192), .C2(n19707), .A(n19704), .B(n19703), .ZN(
        P2_U3061) );
  AOI22_X1 U22761 ( .A1(n19710), .A2(n20194), .B1(n20193), .B2(n19709), .ZN(
        n19706) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19712), .B1(
        n19708), .B2(n20195), .ZN(n19705) );
  OAI211_X1 U22763 ( .C1(n20198), .C2(n19707), .A(n19706), .B(n19705), .ZN(
        P2_U3062) );
  INV_X1 U22764 ( .A(n20203), .ZN(n19870) );
  AOI22_X1 U22765 ( .A1(n19710), .A2(n20201), .B1(n20199), .B2(n19709), .ZN(
        n19714) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19712), .B1(
        n19711), .B2(n20136), .ZN(n19713) );
  OAI211_X1 U22767 ( .C1(n19870), .C2(n19743), .A(n19714), .B(n19713), .ZN(
        P2_U3063) );
  OR2_X1 U22768 ( .A1(n19971), .A2(n19746), .ZN(n19719) );
  INV_X1 U22769 ( .A(n19719), .ZN(n19738) );
  OAI21_X1 U22770 ( .B1(n19718), .B2(n19738), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19715) );
  NAND2_X1 U22771 ( .A1(n19838), .A2(n19745), .ZN(n19716) );
  NAND2_X1 U22772 ( .A1(n19715), .A2(n19716), .ZN(n19739) );
  AOI22_X1 U22773 ( .A1(n19739), .A2(n20150), .B1(n20149), .B2(n19738), .ZN(
        n19725) );
  INV_X1 U22774 ( .A(n19770), .ZN(n19717) );
  OAI221_X1 U22775 ( .B1(n16495), .B2(n19743), .C1(n16495), .C2(n19717), .A(
        n19716), .ZN(n19722) );
  INV_X1 U22776 ( .A(n19718), .ZN(n19720) );
  OAI21_X1 U22777 ( .B1(n19720), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19719), 
        .ZN(n19721) );
  MUX2_X1 U22778 ( .A(n19722), .B(n19721), .S(n20313), .Z(n19723) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20159), .ZN(n19724) );
  OAI211_X1 U22780 ( .C1(n20162), .C2(n19743), .A(n19725), .B(n19724), .ZN(
        P2_U3064) );
  AOI22_X1 U22781 ( .A1(n19739), .A2(n20164), .B1(n19738), .B2(n20163), .ZN(
        n19727) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20165), .ZN(n19726) );
  OAI211_X1 U22783 ( .C1(n20168), .C2(n19743), .A(n19727), .B(n19726), .ZN(
        P2_U3065) );
  AOI22_X1 U22784 ( .A1(n19739), .A2(n20170), .B1(n20169), .B2(n19738), .ZN(
        n19729) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20171), .ZN(n19728) );
  OAI211_X1 U22786 ( .C1(n20174), .C2(n19743), .A(n19729), .B(n19728), .ZN(
        P2_U3066) );
  AOI22_X1 U22787 ( .A1(n19739), .A2(n20176), .B1(n19738), .B2(n20175), .ZN(
        n19731) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20177), .ZN(n19730) );
  OAI211_X1 U22789 ( .C1(n20180), .C2(n19743), .A(n19731), .B(n19730), .ZN(
        P2_U3067) );
  AOI22_X1 U22790 ( .A1(n19739), .A2(n20182), .B1(n20181), .B2(n19738), .ZN(
        n19733) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20183), .ZN(n19732) );
  OAI211_X1 U22792 ( .C1(n20186), .C2(n19743), .A(n19733), .B(n19732), .ZN(
        P2_U3068) );
  AOI22_X1 U22793 ( .A1(n19739), .A2(n20188), .B1(n19738), .B2(n20187), .ZN(
        n19735) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20189), .ZN(n19734) );
  OAI211_X1 U22795 ( .C1(n20192), .C2(n19743), .A(n19735), .B(n19734), .ZN(
        P2_U3069) );
  AOI22_X1 U22796 ( .A1(n19739), .A2(n20194), .B1(n20193), .B2(n19738), .ZN(
        n19737) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20195), .ZN(n19736) );
  OAI211_X1 U22798 ( .C1(n20198), .C2(n19743), .A(n19737), .B(n19736), .ZN(
        P2_U3070) );
  AOI22_X1 U22799 ( .A1(n19739), .A2(n20201), .B1(n20199), .B2(n19738), .ZN(
        n19742) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19740), .B1(
        n19770), .B2(n20203), .ZN(n19741) );
  OAI211_X1 U22801 ( .C1(n20209), .C2(n19743), .A(n19742), .B(n19741), .ZN(
        P2_U3071) );
  INV_X1 U22802 ( .A(n20304), .ZN(n19744) );
  AOI21_X1 U22803 ( .B1(n19872), .B2(n19744), .A(n20313), .ZN(n19749) );
  AND2_X1 U22804 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19745), .ZN(
        n19753) );
  NOR2_X1 U22805 ( .A1(n19747), .A2(n19746), .ZN(n19769) );
  INV_X1 U22806 ( .A(n19769), .ZN(n19750) );
  AOI21_X1 U22807 ( .B1(n19751), .B2(n19750), .A(n20145), .ZN(n19748) );
  AOI22_X1 U22808 ( .A1(n20102), .A2(n19770), .B1(n20149), .B2(n19769), .ZN(
        n19756) );
  INV_X1 U22809 ( .A(n19749), .ZN(n19754) );
  OAI211_X1 U22810 ( .C1(n19751), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20313), 
        .B(n19750), .ZN(n19752) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19771), .B1(
        n19784), .B2(n20159), .ZN(n19755) );
  OAI211_X1 U22812 ( .C1(n19774), .C2(n19945), .A(n19756), .B(n19755), .ZN(
        P2_U3072) );
  AOI22_X1 U22813 ( .A1(n20165), .A2(n19784), .B1(n20163), .B2(n19769), .ZN(
        n19758) );
  AOI22_X1 U22814 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19771), .B1(
        n19770), .B2(n20111), .ZN(n19757) );
  OAI211_X1 U22815 ( .C1(n19774), .C2(n19948), .A(n19758), .B(n19757), .ZN(
        P2_U3073) );
  AOI22_X1 U22816 ( .A1(n20115), .A2(n19770), .B1(n20169), .B2(n19769), .ZN(
        n19760) );
  AOI22_X1 U22817 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19771), .B1(
        n19784), .B2(n20171), .ZN(n19759) );
  OAI211_X1 U22818 ( .C1(n19774), .C2(n19951), .A(n19760), .B(n19759), .ZN(
        P2_U3074) );
  AOI22_X1 U22819 ( .A1(n20177), .A2(n19784), .B1(n20175), .B2(n19769), .ZN(
        n19762) );
  AOI22_X1 U22820 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19771), .B1(
        n19770), .B2(n20119), .ZN(n19761) );
  OAI211_X1 U22821 ( .C1(n19774), .C2(n19954), .A(n19762), .B(n19761), .ZN(
        P2_U3075) );
  AOI22_X1 U22822 ( .A1(n20123), .A2(n19770), .B1(n20181), .B2(n19769), .ZN(
        n19764) );
  AOI22_X1 U22823 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19771), .B1(
        n19784), .B2(n20183), .ZN(n19763) );
  OAI211_X1 U22824 ( .C1(n19774), .C2(n19957), .A(n19764), .B(n19763), .ZN(
        P2_U3076) );
  AOI22_X1 U22825 ( .A1(n20189), .A2(n19784), .B1(n20187), .B2(n19769), .ZN(
        n19766) );
  AOI22_X1 U22826 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19771), .B1(
        n19770), .B2(n20127), .ZN(n19765) );
  OAI211_X1 U22827 ( .C1(n19774), .C2(n19960), .A(n19766), .B(n19765), .ZN(
        P2_U3077) );
  AOI22_X1 U22828 ( .A1(n20131), .A2(n19770), .B1(n20193), .B2(n19769), .ZN(
        n19768) );
  AOI22_X1 U22829 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19771), .B1(
        n19784), .B2(n20195), .ZN(n19767) );
  OAI211_X1 U22830 ( .C1(n19774), .C2(n19963), .A(n19768), .B(n19767), .ZN(
        P2_U3078) );
  AOI22_X1 U22831 ( .A1(n20136), .A2(n19770), .B1(n20199), .B2(n19769), .ZN(
        n19773) );
  AOI22_X1 U22832 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19771), .B1(
        n19784), .B2(n20203), .ZN(n19772) );
  OAI211_X1 U22833 ( .C1(n19774), .C2(n19969), .A(n19773), .B(n19772), .ZN(
        P2_U3079) );
  NOR2_X1 U22834 ( .A1(n19841), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19813) );
  INV_X1 U22835 ( .A(n19813), .ZN(n19815) );
  NOR2_X1 U22836 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19815), .ZN(
        n19802) );
  OAI21_X1 U22837 ( .B1(n12457), .B2(n19802), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19777) );
  INV_X1 U22838 ( .A(n19780), .ZN(n19842) );
  NAND3_X1 U22839 ( .A1(n19775), .A2(n19842), .A3(n20317), .ZN(n19776) );
  NAND2_X1 U22840 ( .A1(n19777), .A2(n19776), .ZN(n19803) );
  AOI22_X1 U22841 ( .A1(n19803), .A2(n20150), .B1(n20149), .B2(n19802), .ZN(
        n19789) );
  INV_X1 U22842 ( .A(n12457), .ZN(n19779) );
  INV_X1 U22843 ( .A(n19802), .ZN(n19778) );
  OAI211_X1 U22844 ( .C1(n19779), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20313), 
        .B(n19778), .ZN(n19787) );
  OR2_X1 U22845 ( .A1(n19781), .A2(n19780), .ZN(n20041) );
  OAI21_X1 U22846 ( .B1(n19784), .B2(n19833), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19785) );
  OAI21_X1 U22847 ( .B1(n20041), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19785), .ZN(n19786) );
  NAND3_X1 U22848 ( .A1(n19787), .A2(n20152), .A3(n19786), .ZN(n19804) );
  AOI22_X1 U22849 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20159), .ZN(n19788) );
  OAI211_X1 U22850 ( .C1(n20162), .C2(n19807), .A(n19789), .B(n19788), .ZN(
        P2_U3080) );
  AOI22_X1 U22851 ( .A1(n19803), .A2(n20164), .B1(n19802), .B2(n20163), .ZN(
        n19791) );
  AOI22_X1 U22852 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20165), .ZN(n19790) );
  OAI211_X1 U22853 ( .C1(n20168), .C2(n19807), .A(n19791), .B(n19790), .ZN(
        P2_U3081) );
  AOI22_X1 U22854 ( .A1(n19803), .A2(n20170), .B1(n20169), .B2(n19802), .ZN(
        n19793) );
  AOI22_X1 U22855 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20171), .ZN(n19792) );
  OAI211_X1 U22856 ( .C1(n20174), .C2(n19807), .A(n19793), .B(n19792), .ZN(
        P2_U3082) );
  AOI22_X1 U22857 ( .A1(n19803), .A2(n20176), .B1(n19802), .B2(n20175), .ZN(
        n19795) );
  AOI22_X1 U22858 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20177), .ZN(n19794) );
  OAI211_X1 U22859 ( .C1(n20180), .C2(n19807), .A(n19795), .B(n19794), .ZN(
        P2_U3083) );
  AOI22_X1 U22860 ( .A1(n19803), .A2(n20182), .B1(n20181), .B2(n19802), .ZN(
        n19797) );
  AOI22_X1 U22861 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20183), .ZN(n19796) );
  OAI211_X1 U22862 ( .C1(n20186), .C2(n19807), .A(n19797), .B(n19796), .ZN(
        P2_U3084) );
  AOI22_X1 U22863 ( .A1(n19803), .A2(n20188), .B1(n19802), .B2(n20187), .ZN(
        n19799) );
  AOI22_X1 U22864 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20189), .ZN(n19798) );
  OAI211_X1 U22865 ( .C1(n20192), .C2(n19807), .A(n19799), .B(n19798), .ZN(
        P2_U3085) );
  AOI22_X1 U22866 ( .A1(n19803), .A2(n20194), .B1(n20193), .B2(n19802), .ZN(
        n19801) );
  AOI22_X1 U22867 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20195), .ZN(n19800) );
  OAI211_X1 U22868 ( .C1(n20198), .C2(n19807), .A(n19801), .B(n19800), .ZN(
        P2_U3086) );
  AOI22_X1 U22869 ( .A1(n19803), .A2(n20201), .B1(n20199), .B2(n19802), .ZN(
        n19806) );
  AOI22_X1 U22870 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19804), .B1(
        n19833), .B2(n20203), .ZN(n19805) );
  OAI211_X1 U22871 ( .C1(n20209), .C2(n19807), .A(n19806), .B(n19805), .ZN(
        P2_U3087) );
  NOR2_X1 U22872 ( .A1(n19841), .A2(n19808), .ZN(n19832) );
  AOI22_X1 U22873 ( .A1(n20159), .A2(n19866), .B1(n20149), .B2(n19832), .ZN(
        n19818) );
  INV_X1 U22874 ( .A(n19872), .ZN(n19809) );
  OAI21_X1 U22875 ( .B1(n19809), .B2(n20072), .A(n20099), .ZN(n19816) );
  INV_X1 U22876 ( .A(n12454), .ZN(n19811) );
  INV_X1 U22877 ( .A(n19832), .ZN(n19810) );
  OAI211_X1 U22878 ( .C1(n19811), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20313), 
        .B(n19810), .ZN(n19812) );
  OAI211_X1 U22879 ( .C1(n19816), .C2(n19813), .A(n20152), .B(n19812), .ZN(
        n19835) );
  OAI21_X1 U22880 ( .B1(n12454), .B2(n19832), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19814) );
  AOI22_X1 U22881 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19835), .B1(
        n20150), .B2(n19834), .ZN(n19817) );
  OAI211_X1 U22882 ( .C1(n20162), .C2(n19783), .A(n19818), .B(n19817), .ZN(
        P2_U3088) );
  AOI22_X1 U22883 ( .A1(n20165), .A2(n19866), .B1(n20163), .B2(n19832), .ZN(
        n19820) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19835), .B1(
        n20164), .B2(n19834), .ZN(n19819) );
  OAI211_X1 U22885 ( .C1(n20168), .C2(n19783), .A(n19820), .B(n19819), .ZN(
        P2_U3089) );
  AOI22_X1 U22886 ( .A1(n20171), .A2(n19866), .B1(n20169), .B2(n19832), .ZN(
        n19822) );
  AOI22_X1 U22887 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19835), .B1(
        n20170), .B2(n19834), .ZN(n19821) );
  OAI211_X1 U22888 ( .C1(n20174), .C2(n19783), .A(n19822), .B(n19821), .ZN(
        P2_U3090) );
  AOI22_X1 U22889 ( .A1(n20177), .A2(n19866), .B1(n20175), .B2(n19832), .ZN(
        n19824) );
  AOI22_X1 U22890 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19835), .B1(
        n20176), .B2(n19834), .ZN(n19823) );
  OAI211_X1 U22891 ( .C1(n20180), .C2(n19783), .A(n19824), .B(n19823), .ZN(
        P2_U3091) );
  INV_X1 U22892 ( .A(n20183), .ZN(n20022) );
  AOI22_X1 U22893 ( .A1(n20123), .A2(n19833), .B1(n20181), .B2(n19832), .ZN(
        n19826) );
  AOI22_X1 U22894 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19835), .B1(
        n20182), .B2(n19834), .ZN(n19825) );
  OAI211_X1 U22895 ( .C1(n20022), .C2(n19863), .A(n19826), .B(n19825), .ZN(
        P2_U3092) );
  INV_X1 U22896 ( .A(n20189), .ZN(n19829) );
  AOI22_X1 U22897 ( .A1(n20127), .A2(n19833), .B1(n20187), .B2(n19832), .ZN(
        n19828) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19835), .B1(
        n20188), .B2(n19834), .ZN(n19827) );
  OAI211_X1 U22899 ( .C1(n19829), .C2(n19863), .A(n19828), .B(n19827), .ZN(
        P2_U3093) );
  AOI22_X1 U22900 ( .A1(n20195), .A2(n19866), .B1(n20193), .B2(n19832), .ZN(
        n19831) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19835), .B1(
        n20194), .B2(n19834), .ZN(n19830) );
  OAI211_X1 U22902 ( .C1(n20198), .C2(n19783), .A(n19831), .B(n19830), .ZN(
        P2_U3094) );
  AOI22_X1 U22903 ( .A1(n20136), .A2(n19833), .B1(n20199), .B2(n19832), .ZN(
        n19837) );
  AOI22_X1 U22904 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19835), .B1(
        n20201), .B2(n19834), .ZN(n19836) );
  OAI211_X1 U22905 ( .C1(n19870), .C2(n19863), .A(n19837), .B(n19836), .ZN(
        P2_U3095) );
  INV_X1 U22906 ( .A(n19838), .ZN(n19973) );
  OR2_X1 U22907 ( .A1(n19971), .A2(n19841), .ZN(n19844) );
  INV_X1 U22908 ( .A(n19844), .ZN(n19864) );
  OAI21_X1 U22909 ( .B1(n19843), .B2(n19864), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19839) );
  AOI22_X1 U22910 ( .A1(n19865), .A2(n20150), .B1(n20149), .B2(n19864), .ZN(
        n19850) );
  AOI21_X1 U22911 ( .B1(n19863), .B2(n19904), .A(n16495), .ZN(n19848) );
  NOR2_X1 U22912 ( .A1(n19842), .A2(n19841), .ZN(n19847) );
  INV_X1 U22913 ( .A(n19843), .ZN(n19845) );
  OAI211_X1 U22914 ( .C1(n19845), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20313), 
        .B(n19844), .ZN(n19846) );
  AOI22_X1 U22915 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20159), .ZN(n19849) );
  OAI211_X1 U22916 ( .C1(n20162), .C2(n19863), .A(n19850), .B(n19849), .ZN(
        P2_U3096) );
  AOI22_X1 U22917 ( .A1(n19865), .A2(n20164), .B1(n19864), .B2(n20163), .ZN(
        n19852) );
  AOI22_X1 U22918 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20165), .ZN(n19851) );
  OAI211_X1 U22919 ( .C1(n20168), .C2(n19863), .A(n19852), .B(n19851), .ZN(
        P2_U3097) );
  AOI22_X1 U22920 ( .A1(n19865), .A2(n20170), .B1(n20169), .B2(n19864), .ZN(
        n19854) );
  AOI22_X1 U22921 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20171), .ZN(n19853) );
  OAI211_X1 U22922 ( .C1(n20174), .C2(n19863), .A(n19854), .B(n19853), .ZN(
        P2_U3098) );
  AOI22_X1 U22923 ( .A1(n19865), .A2(n20176), .B1(n19864), .B2(n20175), .ZN(
        n19856) );
  AOI22_X1 U22924 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20177), .ZN(n19855) );
  OAI211_X1 U22925 ( .C1(n20180), .C2(n19863), .A(n19856), .B(n19855), .ZN(
        P2_U3099) );
  AOI22_X1 U22926 ( .A1(n19865), .A2(n20182), .B1(n20181), .B2(n19864), .ZN(
        n19858) );
  AOI22_X1 U22927 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20183), .ZN(n19857) );
  OAI211_X1 U22928 ( .C1(n20186), .C2(n19863), .A(n19858), .B(n19857), .ZN(
        P2_U3100) );
  AOI22_X1 U22929 ( .A1(n19865), .A2(n20188), .B1(n19864), .B2(n20187), .ZN(
        n19860) );
  AOI22_X1 U22930 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20189), .ZN(n19859) );
  OAI211_X1 U22931 ( .C1(n20192), .C2(n19863), .A(n19860), .B(n19859), .ZN(
        P2_U3101) );
  AOI22_X1 U22932 ( .A1(n19865), .A2(n20194), .B1(n20193), .B2(n19864), .ZN(
        n19862) );
  AOI22_X1 U22933 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19867), .B1(
        n19882), .B2(n20195), .ZN(n19861) );
  OAI211_X1 U22934 ( .C1(n20198), .C2(n19863), .A(n19862), .B(n19861), .ZN(
        P2_U3102) );
  AOI22_X1 U22935 ( .A1(n19865), .A2(n20201), .B1(n20199), .B2(n19864), .ZN(
        n19869) );
  AOI22_X1 U22936 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20136), .ZN(n19868) );
  OAI211_X1 U22937 ( .C1(n19870), .C2(n19904), .A(n19869), .B(n19868), .ZN(
        P2_U3103) );
  INV_X1 U22938 ( .A(n20156), .ZN(n19871) );
  NAND2_X1 U22939 ( .A1(n19872), .A2(n19871), .ZN(n20314) );
  OR2_X1 U22940 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20097), .ZN(
        n19880) );
  NAND2_X1 U22941 ( .A1(n20314), .A2(n19880), .ZN(n19876) );
  INV_X1 U22942 ( .A(n19911), .ZN(n19899) );
  NAND2_X1 U22943 ( .A1(n19911), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19873) );
  OAI211_X1 U22944 ( .C1(n19899), .C2(n20318), .A(n19877), .B(n20152), .ZN(
        n19874) );
  INV_X1 U22945 ( .A(n19874), .ZN(n19875) );
  INV_X1 U22946 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19885) );
  INV_X1 U22947 ( .A(n19877), .ZN(n19878) );
  AOI211_X2 U22948 ( .C1(n19880), .C2(n20145), .A(n19879), .B(n19878), .ZN(
        n19900) );
  AOI22_X1 U22949 ( .A1(n19900), .A2(n20150), .B1(n19899), .B2(n20149), .ZN(
        n19884) );
  AOI22_X1 U22950 ( .A1(n10291), .A2(n20159), .B1(n19882), .B2(n20102), .ZN(
        n19883) );
  OAI211_X1 U22951 ( .C1(n19886), .C2(n19885), .A(n19884), .B(n19883), .ZN(
        P2_U3104) );
  AOI22_X1 U22952 ( .A1(n19900), .A2(n20164), .B1(n19899), .B2(n20163), .ZN(
        n19888) );
  AOI22_X1 U22953 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20165), .ZN(n19887) );
  OAI211_X1 U22954 ( .C1(n20168), .C2(n19904), .A(n19888), .B(n19887), .ZN(
        P2_U3105) );
  AOI22_X1 U22955 ( .A1(n19900), .A2(n20170), .B1(n19899), .B2(n20169), .ZN(
        n19890) );
  AOI22_X1 U22956 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20171), .ZN(n19889) );
  OAI211_X1 U22957 ( .C1(n20174), .C2(n19904), .A(n19890), .B(n19889), .ZN(
        P2_U3106) );
  AOI22_X1 U22958 ( .A1(n19900), .A2(n20176), .B1(n19899), .B2(n20175), .ZN(
        n19892) );
  AOI22_X1 U22959 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20177), .ZN(n19891) );
  OAI211_X1 U22960 ( .C1(n20180), .C2(n19904), .A(n19892), .B(n19891), .ZN(
        P2_U3107) );
  AOI22_X1 U22961 ( .A1(n19900), .A2(n20182), .B1(n19899), .B2(n20181), .ZN(
        n19894) );
  AOI22_X1 U22962 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20183), .ZN(n19893) );
  OAI211_X1 U22963 ( .C1(n20186), .C2(n19904), .A(n19894), .B(n19893), .ZN(
        P2_U3108) );
  AOI22_X1 U22964 ( .A1(n19900), .A2(n20188), .B1(n19899), .B2(n20187), .ZN(
        n19896) );
  AOI22_X1 U22965 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20189), .ZN(n19895) );
  OAI211_X1 U22966 ( .C1(n20192), .C2(n19904), .A(n19896), .B(n19895), .ZN(
        P2_U3109) );
  AOI22_X1 U22967 ( .A1(n19900), .A2(n20194), .B1(n19899), .B2(n20193), .ZN(
        n19898) );
  AOI22_X1 U22968 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20195), .ZN(n19897) );
  OAI211_X1 U22969 ( .C1(n20198), .C2(n19904), .A(n19898), .B(n19897), .ZN(
        P2_U3110) );
  AOI22_X1 U22970 ( .A1(n19900), .A2(n20201), .B1(n19899), .B2(n20199), .ZN(
        n19903) );
  AOI22_X1 U22971 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19901), .B1(
        n10291), .B2(n20203), .ZN(n19902) );
  OAI211_X1 U22972 ( .C1(n20209), .C2(n19904), .A(n19903), .B(n19902), .ZN(
        P2_U3111) );
  NOR3_X1 U22973 ( .A1(n19965), .A2(n10291), .A3(n20313), .ZN(n19906) );
  INV_X1 U22974 ( .A(n20095), .ZN(n19905) );
  NOR2_X1 U22975 ( .A1(n19906), .A2(n19905), .ZN(n19908) );
  INV_X1 U22976 ( .A(n12460), .ZN(n19907) );
  AOI22_X1 U22977 ( .A1(n19908), .A2(n19907), .B1(n20145), .B2(n19911), .ZN(
        n19909) );
  NAND2_X1 U22978 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20325), .ZN(
        n20006) );
  NOR2_X1 U22979 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20006), .ZN(
        n19940) );
  AND2_X1 U22980 ( .A1(n19940), .A2(n20335), .ZN(n19928) );
  INV_X1 U22981 ( .A(n19908), .ZN(n19912) );
  AOI22_X1 U22982 ( .A1(n20102), .A2(n10291), .B1(n20149), .B2(n19928), .ZN(
        n19915) );
  OAI21_X1 U22983 ( .B1(n12460), .B2(n20145), .A(n20318), .ZN(n19910) );
  AOI21_X1 U22984 ( .B1(n19912), .B2(n19911), .A(n19910), .ZN(n19913) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19929), .B1(
        n19965), .B2(n20159), .ZN(n19914) );
  OAI211_X1 U22986 ( .C1(n19945), .C2(n19932), .A(n19915), .B(n19914), .ZN(
        P2_U3112) );
  AOI22_X1 U22987 ( .A1(n20111), .A2(n10291), .B1(n20163), .B2(n19928), .ZN(
        n19917) );
  AOI22_X1 U22988 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19929), .B1(
        n19965), .B2(n20165), .ZN(n19916) );
  OAI211_X1 U22989 ( .C1(n19948), .C2(n19932), .A(n19917), .B(n19916), .ZN(
        P2_U3113) );
  AOI22_X1 U22990 ( .A1(n20171), .A2(n19965), .B1(n20169), .B2(n19928), .ZN(
        n19919) );
  AOI22_X1 U22991 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19929), .B1(
        n10291), .B2(n20115), .ZN(n19918) );
  OAI211_X1 U22992 ( .C1(n19951), .C2(n19932), .A(n19919), .B(n19918), .ZN(
        P2_U3114) );
  AOI22_X1 U22993 ( .A1(n20177), .A2(n19965), .B1(n20175), .B2(n19928), .ZN(
        n19921) );
  AOI22_X1 U22994 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19929), .B1(
        n10291), .B2(n20119), .ZN(n19920) );
  OAI211_X1 U22995 ( .C1(n19954), .C2(n19932), .A(n19921), .B(n19920), .ZN(
        P2_U3115) );
  AOI22_X1 U22996 ( .A1(n20123), .A2(n10291), .B1(n20181), .B2(n19928), .ZN(
        n19923) );
  AOI22_X1 U22997 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19929), .B1(
        n19965), .B2(n20183), .ZN(n19922) );
  OAI211_X1 U22998 ( .C1(n19957), .C2(n19932), .A(n19923), .B(n19922), .ZN(
        P2_U3116) );
  AOI22_X1 U22999 ( .A1(n20127), .A2(n10291), .B1(n20187), .B2(n19928), .ZN(
        n19925) );
  AOI22_X1 U23000 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19929), .B1(
        n19965), .B2(n20189), .ZN(n19924) );
  OAI211_X1 U23001 ( .C1(n19960), .C2(n19932), .A(n19925), .B(n19924), .ZN(
        P2_U3117) );
  AOI22_X1 U23002 ( .A1(n20195), .A2(n19965), .B1(n20193), .B2(n19928), .ZN(
        n19927) );
  AOI22_X1 U23003 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19929), .B1(
        n10291), .B2(n20131), .ZN(n19926) );
  OAI211_X1 U23004 ( .C1(n19963), .C2(n19932), .A(n19927), .B(n19926), .ZN(
        P2_U3118) );
  AOI22_X1 U23005 ( .A1(n20136), .A2(n10291), .B1(n20199), .B2(n19928), .ZN(
        n19931) );
  AOI22_X1 U23006 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19929), .B1(
        n19965), .B2(n20203), .ZN(n19930) );
  OAI211_X1 U23007 ( .C1(n19969), .C2(n19932), .A(n19931), .B(n19930), .ZN(
        P2_U3119) );
  NAND2_X1 U23008 ( .A1(n20309), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20155) );
  INV_X1 U23009 ( .A(n20155), .ZN(n20068) );
  AOI21_X1 U23010 ( .B1(n20068), .B2(n19933), .A(n20313), .ZN(n19937) );
  INV_X1 U23011 ( .A(n19934), .ZN(n19938) );
  INV_X1 U23012 ( .A(n20006), .ZN(n20002) );
  NAND2_X1 U23013 ( .A1(n19935), .A2(n20002), .ZN(n19975) );
  AOI21_X1 U23014 ( .B1(n19938), .B2(n19975), .A(n20145), .ZN(n19936) );
  INV_X1 U23015 ( .A(n19975), .ZN(n19964) );
  AOI22_X1 U23016 ( .A1(n20102), .A2(n19965), .B1(n20149), .B2(n19964), .ZN(
        n19944) );
  INV_X1 U23017 ( .A(n19937), .ZN(n19941) );
  OAI211_X1 U23018 ( .C1(n19938), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19975), 
        .B(n20313), .ZN(n19939) );
  AOI22_X1 U23019 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19966), .B1(
        n19974), .B2(n20159), .ZN(n19943) );
  OAI211_X1 U23020 ( .C1(n19970), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        P2_U3120) );
  AOI22_X1 U23021 ( .A1(n20165), .A2(n19974), .B1(n20163), .B2(n19964), .ZN(
        n19947) );
  AOI22_X1 U23022 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19966), .B1(
        n19965), .B2(n20111), .ZN(n19946) );
  OAI211_X1 U23023 ( .C1(n19970), .C2(n19948), .A(n19947), .B(n19946), .ZN(
        P2_U3121) );
  AOI22_X1 U23024 ( .A1(n20115), .A2(n19965), .B1(n20169), .B2(n19964), .ZN(
        n19950) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19966), .B1(
        n19974), .B2(n20171), .ZN(n19949) );
  OAI211_X1 U23026 ( .C1(n19970), .C2(n19951), .A(n19950), .B(n19949), .ZN(
        P2_U3122) );
  AOI22_X1 U23027 ( .A1(n20177), .A2(n19974), .B1(n20175), .B2(n19964), .ZN(
        n19953) );
  AOI22_X1 U23028 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19966), .B1(
        n19965), .B2(n20119), .ZN(n19952) );
  OAI211_X1 U23029 ( .C1(n19970), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        P2_U3123) );
  AOI22_X1 U23030 ( .A1(n20183), .A2(n19974), .B1(n20181), .B2(n19964), .ZN(
        n19956) );
  AOI22_X1 U23031 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19966), .B1(
        n19965), .B2(n20123), .ZN(n19955) );
  OAI211_X1 U23032 ( .C1(n19970), .C2(n19957), .A(n19956), .B(n19955), .ZN(
        P2_U3124) );
  AOI22_X1 U23033 ( .A1(n20127), .A2(n19965), .B1(n20187), .B2(n19964), .ZN(
        n19959) );
  AOI22_X1 U23034 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19966), .B1(
        n19974), .B2(n20189), .ZN(n19958) );
  OAI211_X1 U23035 ( .C1(n19970), .C2(n19960), .A(n19959), .B(n19958), .ZN(
        P2_U3125) );
  AOI22_X1 U23036 ( .A1(n20195), .A2(n19974), .B1(n20193), .B2(n19964), .ZN(
        n19962) );
  AOI22_X1 U23037 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19966), .B1(
        n19965), .B2(n20131), .ZN(n19961) );
  OAI211_X1 U23038 ( .C1(n19970), .C2(n19963), .A(n19962), .B(n19961), .ZN(
        P2_U3126) );
  AOI22_X1 U23039 ( .A1(n20203), .A2(n19974), .B1(n20199), .B2(n19964), .ZN(
        n19968) );
  AOI22_X1 U23040 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19966), .B1(
        n19965), .B2(n20136), .ZN(n19967) );
  OAI211_X1 U23041 ( .C1(n19970), .C2(n19969), .A(n19968), .B(n19967), .ZN(
        P2_U3127) );
  OR2_X1 U23042 ( .A1(n19971), .A2(n20006), .ZN(n19978) );
  INV_X1 U23043 ( .A(n19978), .ZN(n19996) );
  OAI21_X1 U23044 ( .B1(n19977), .B2(n19996), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19972) );
  OAI21_X1 U23045 ( .B1(n20006), .B2(n19973), .A(n19972), .ZN(n19997) );
  AOI22_X1 U23046 ( .A1(n19997), .A2(n20150), .B1(n20149), .B2(n19996), .ZN(
        n19983) );
  OAI21_X1 U23047 ( .B1(n20019), .B2(n19974), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19976) );
  AOI21_X1 U23048 ( .B1(n19976), .B2(n19975), .A(n20313), .ZN(n19981) );
  NAND3_X1 U23049 ( .A1(n19977), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20318), 
        .ZN(n19979) );
  NAND2_X1 U23050 ( .A1(n19979), .A2(n19978), .ZN(n19980) );
  AOI22_X1 U23051 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20159), .ZN(n19982) );
  OAI211_X1 U23052 ( .C1(n20162), .C2(n20001), .A(n19983), .B(n19982), .ZN(
        P2_U3128) );
  AOI22_X1 U23053 ( .A1(n19997), .A2(n20164), .B1(n19996), .B2(n20163), .ZN(
        n19985) );
  AOI22_X1 U23054 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20165), .ZN(n19984) );
  OAI211_X1 U23055 ( .C1(n20168), .C2(n20001), .A(n19985), .B(n19984), .ZN(
        P2_U3129) );
  AOI22_X1 U23056 ( .A1(n19997), .A2(n20170), .B1(n20169), .B2(n19996), .ZN(
        n19987) );
  AOI22_X1 U23057 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20171), .ZN(n19986) );
  OAI211_X1 U23058 ( .C1(n20174), .C2(n20001), .A(n19987), .B(n19986), .ZN(
        P2_U3130) );
  AOI22_X1 U23059 ( .A1(n19997), .A2(n20176), .B1(n19996), .B2(n20175), .ZN(
        n19989) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20177), .ZN(n19988) );
  OAI211_X1 U23061 ( .C1(n20180), .C2(n20001), .A(n19989), .B(n19988), .ZN(
        P2_U3131) );
  AOI22_X1 U23062 ( .A1(n19997), .A2(n20182), .B1(n20181), .B2(n19996), .ZN(
        n19991) );
  AOI22_X1 U23063 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20183), .ZN(n19990) );
  OAI211_X1 U23064 ( .C1(n20186), .C2(n20001), .A(n19991), .B(n19990), .ZN(
        P2_U3132) );
  AOI22_X1 U23065 ( .A1(n19997), .A2(n20188), .B1(n19996), .B2(n20187), .ZN(
        n19993) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20189), .ZN(n19992) );
  OAI211_X1 U23067 ( .C1(n20192), .C2(n20001), .A(n19993), .B(n19992), .ZN(
        P2_U3133) );
  AOI22_X1 U23068 ( .A1(n19997), .A2(n20194), .B1(n20193), .B2(n19996), .ZN(
        n19995) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20195), .ZN(n19994) );
  OAI211_X1 U23070 ( .C1(n20198), .C2(n20001), .A(n19995), .B(n19994), .ZN(
        P2_U3134) );
  AOI22_X1 U23071 ( .A1(n19997), .A2(n20201), .B1(n20199), .B2(n19996), .ZN(
        n20000) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19998), .B1(
        n20019), .B2(n20203), .ZN(n19999) );
  OAI211_X1 U23073 ( .C1(n20209), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P2_U3135) );
  NAND2_X1 U23074 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20002), .ZN(
        n20005) );
  NAND2_X1 U23075 ( .A1(n20003), .A2(n20002), .ZN(n20007) );
  INV_X1 U23076 ( .A(n20007), .ZN(n20027) );
  OAI21_X1 U23077 ( .B1(n12452), .B2(n20027), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20004) );
  OAI21_X1 U23078 ( .B1(n20005), .B2(n20313), .A(n20004), .ZN(n20028) );
  AOI22_X1 U23079 ( .A1(n20028), .A2(n20150), .B1(n20149), .B2(n20027), .ZN(
        n20012) );
  OAI22_X1 U23080 ( .A1(n20155), .A2(n20304), .B1(n20006), .B2(n20034), .ZN(
        n20010) );
  INV_X1 U23081 ( .A(n12452), .ZN(n20008) );
  OAI211_X1 U23082 ( .C1(n20008), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20313), 
        .B(n20007), .ZN(n20009) );
  NAND3_X1 U23083 ( .A1(n20010), .A2(n20152), .A3(n20009), .ZN(n20029) );
  AOI22_X1 U23084 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20159), .ZN(n20011) );
  OAI211_X1 U23085 ( .C1(n20162), .C2(n20032), .A(n20012), .B(n20011), .ZN(
        P2_U3136) );
  AOI22_X1 U23086 ( .A1(n20028), .A2(n20164), .B1(n20027), .B2(n20163), .ZN(
        n20014) );
  AOI22_X1 U23087 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20165), .ZN(n20013) );
  OAI211_X1 U23088 ( .C1(n20168), .C2(n20032), .A(n20014), .B(n20013), .ZN(
        P2_U3137) );
  AOI22_X1 U23089 ( .A1(n20028), .A2(n20170), .B1(n20169), .B2(n20027), .ZN(
        n20016) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20171), .ZN(n20015) );
  OAI211_X1 U23091 ( .C1(n20174), .C2(n20032), .A(n20016), .B(n20015), .ZN(
        P2_U3138) );
  AOI22_X1 U23092 ( .A1(n20028), .A2(n20176), .B1(n20027), .B2(n20175), .ZN(
        n20018) );
  AOI22_X1 U23093 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20177), .ZN(n20017) );
  OAI211_X1 U23094 ( .C1(n20180), .C2(n20032), .A(n20018), .B(n20017), .ZN(
        P2_U3139) );
  AOI22_X1 U23095 ( .A1(n20028), .A2(n20182), .B1(n20181), .B2(n20027), .ZN(
        n20021) );
  AOI22_X1 U23096 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20029), .B1(
        n20019), .B2(n20123), .ZN(n20020) );
  OAI211_X1 U23097 ( .C1(n20022), .C2(n20063), .A(n20021), .B(n20020), .ZN(
        P2_U3140) );
  AOI22_X1 U23098 ( .A1(n20028), .A2(n20188), .B1(n20027), .B2(n20187), .ZN(
        n20024) );
  AOI22_X1 U23099 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20189), .ZN(n20023) );
  OAI211_X1 U23100 ( .C1(n20192), .C2(n20032), .A(n20024), .B(n20023), .ZN(
        P2_U3141) );
  AOI22_X1 U23101 ( .A1(n20028), .A2(n20194), .B1(n20193), .B2(n20027), .ZN(
        n20026) );
  AOI22_X1 U23102 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20195), .ZN(n20025) );
  OAI211_X1 U23103 ( .C1(n20198), .C2(n20032), .A(n20026), .B(n20025), .ZN(
        P2_U3142) );
  AOI22_X1 U23104 ( .A1(n20028), .A2(n20201), .B1(n20199), .B2(n20027), .ZN(
        n20031) );
  AOI22_X1 U23105 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20029), .B1(
        n20039), .B2(n20203), .ZN(n20030) );
  OAI211_X1 U23106 ( .C1(n20209), .C2(n20032), .A(n20031), .B(n20030), .ZN(
        P2_U3143) );
  INV_X1 U23107 ( .A(n20033), .ZN(n20036) );
  AND3_X1 U23108 ( .A1(n20034), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20066) );
  AND2_X1 U23109 ( .A1(n20066), .A2(n20335), .ZN(n20058) );
  OAI21_X1 U23110 ( .B1(n20037), .B2(n20058), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20035) );
  OAI21_X1 U23111 ( .B1(n20036), .B2(n20041), .A(n20035), .ZN(n20059) );
  AOI22_X1 U23112 ( .A1(n20059), .A2(n20150), .B1(n20149), .B2(n20058), .ZN(
        n20045) );
  INV_X1 U23113 ( .A(n20037), .ZN(n20038) );
  AOI21_X1 U23114 ( .B1(n20038), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20043) );
  OAI21_X1 U23115 ( .B1(n20039), .B2(n20064), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20040) );
  OAI21_X1 U23116 ( .B1(n20041), .B2(n20317), .A(n20040), .ZN(n20042) );
  AOI22_X1 U23117 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20159), .ZN(n20044) );
  OAI211_X1 U23118 ( .C1(n20162), .C2(n20063), .A(n20045), .B(n20044), .ZN(
        P2_U3144) );
  AOI22_X1 U23119 ( .A1(n20059), .A2(n20164), .B1(n20058), .B2(n20163), .ZN(
        n20047) );
  AOI22_X1 U23120 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20165), .ZN(n20046) );
  OAI211_X1 U23121 ( .C1(n20168), .C2(n20063), .A(n20047), .B(n20046), .ZN(
        P2_U3145) );
  AOI22_X1 U23122 ( .A1(n20059), .A2(n20170), .B1(n20169), .B2(n20058), .ZN(
        n20049) );
  AOI22_X1 U23123 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20171), .ZN(n20048) );
  OAI211_X1 U23124 ( .C1(n20174), .C2(n20063), .A(n20049), .B(n20048), .ZN(
        P2_U3146) );
  AOI22_X1 U23125 ( .A1(n20059), .A2(n20176), .B1(n20058), .B2(n20175), .ZN(
        n20051) );
  AOI22_X1 U23126 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20177), .ZN(n20050) );
  OAI211_X1 U23127 ( .C1(n20180), .C2(n20063), .A(n20051), .B(n20050), .ZN(
        P2_U3147) );
  AOI22_X1 U23128 ( .A1(n20059), .A2(n20182), .B1(n20181), .B2(n20058), .ZN(
        n20053) );
  AOI22_X1 U23129 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20183), .ZN(n20052) );
  OAI211_X1 U23130 ( .C1(n20186), .C2(n20063), .A(n20053), .B(n20052), .ZN(
        P2_U3148) );
  AOI22_X1 U23131 ( .A1(n20059), .A2(n20188), .B1(n20058), .B2(n20187), .ZN(
        n20055) );
  AOI22_X1 U23132 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20189), .ZN(n20054) );
  OAI211_X1 U23133 ( .C1(n20192), .C2(n20063), .A(n20055), .B(n20054), .ZN(
        P2_U3149) );
  AOI22_X1 U23134 ( .A1(n20059), .A2(n20194), .B1(n20193), .B2(n20058), .ZN(
        n20057) );
  AOI22_X1 U23135 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20195), .ZN(n20056) );
  OAI211_X1 U23136 ( .C1(n20198), .C2(n20063), .A(n20057), .B(n20056), .ZN(
        P2_U3150) );
  AOI22_X1 U23137 ( .A1(n20059), .A2(n20201), .B1(n20199), .B2(n20058), .ZN(
        n20062) );
  AOI22_X1 U23138 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20060), .B1(
        n20064), .B2(n20203), .ZN(n20061) );
  OAI211_X1 U23139 ( .C1(n20209), .C2(n20063), .A(n20062), .B(n20061), .ZN(
        P2_U3151) );
  AND2_X1 U23140 ( .A1(n20066), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20098) );
  NOR3_X1 U23141 ( .A1(n9641), .A2(n20098), .A3(n20145), .ZN(n20069) );
  AOI21_X1 U23142 ( .B1(n20066), .B2(n20318), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20065) );
  AOI22_X1 U23143 ( .A1(n20088), .A2(n20150), .B1(n20149), .B2(n20098), .ZN(
        n20075) );
  INV_X1 U23144 ( .A(n20072), .ZN(n20067) );
  AOI21_X1 U23145 ( .B1(n20068), .B2(n20067), .A(n20066), .ZN(n20070) );
  NOR2_X1 U23146 ( .A1(n20070), .A2(n20069), .ZN(n20071) );
  OAI211_X1 U23147 ( .C1(n20098), .C2(n20318), .A(n20071), .B(n20152), .ZN(
        n20089) );
  AOI22_X1 U23148 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20159), .ZN(n20074) );
  OAI211_X1 U23149 ( .C1(n20162), .C2(n20092), .A(n20075), .B(n20074), .ZN(
        P2_U3152) );
  AOI22_X1 U23150 ( .A1(n20088), .A2(n20164), .B1(n20098), .B2(n20163), .ZN(
        n20077) );
  AOI22_X1 U23151 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20165), .ZN(n20076) );
  OAI211_X1 U23152 ( .C1(n20168), .C2(n20092), .A(n20077), .B(n20076), .ZN(
        P2_U3153) );
  AOI22_X1 U23153 ( .A1(n20088), .A2(n20170), .B1(n20169), .B2(n20098), .ZN(
        n20079) );
  AOI22_X1 U23154 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20171), .ZN(n20078) );
  OAI211_X1 U23155 ( .C1(n20174), .C2(n20092), .A(n20079), .B(n20078), .ZN(
        P2_U3154) );
  AOI22_X1 U23156 ( .A1(n20088), .A2(n20176), .B1(n20098), .B2(n20175), .ZN(
        n20081) );
  AOI22_X1 U23157 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20177), .ZN(n20080) );
  OAI211_X1 U23158 ( .C1(n20180), .C2(n20092), .A(n20081), .B(n20080), .ZN(
        P2_U3155) );
  AOI22_X1 U23159 ( .A1(n20088), .A2(n20182), .B1(n20181), .B2(n20098), .ZN(
        n20083) );
  AOI22_X1 U23160 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20183), .ZN(n20082) );
  OAI211_X1 U23161 ( .C1(n20186), .C2(n20092), .A(n20083), .B(n20082), .ZN(
        P2_U3156) );
  AOI22_X1 U23162 ( .A1(n20088), .A2(n20188), .B1(n20098), .B2(n20187), .ZN(
        n20085) );
  AOI22_X1 U23163 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20189), .ZN(n20084) );
  OAI211_X1 U23164 ( .C1(n20192), .C2(n20092), .A(n20085), .B(n20084), .ZN(
        P2_U3157) );
  AOI22_X1 U23165 ( .A1(n20088), .A2(n20194), .B1(n20193), .B2(n20098), .ZN(
        n20087) );
  AOI22_X1 U23166 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20195), .ZN(n20086) );
  OAI211_X1 U23167 ( .C1(n20198), .C2(n20092), .A(n20087), .B(n20086), .ZN(
        P2_U3158) );
  AOI22_X1 U23168 ( .A1(n20088), .A2(n20201), .B1(n20199), .B2(n20098), .ZN(
        n20091) );
  AOI22_X1 U23169 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20089), .B1(
        n20137), .B2(n20203), .ZN(n20090) );
  OAI211_X1 U23170 ( .C1(n20209), .C2(n20092), .A(n20091), .B(n20090), .ZN(
        P2_U3159) );
  INV_X1 U23171 ( .A(n20137), .ZN(n20093) );
  NAND2_X1 U23172 ( .A1(n20093), .A2(n20099), .ZN(n20096) );
  OAI21_X1 U23173 ( .B1(n20096), .B2(n20143), .A(n20095), .ZN(n20103) );
  NOR3_X2 U23174 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20317), .A3(
        n20097), .ZN(n20135) );
  NOR2_X1 U23175 ( .A1(n20098), .A2(n20135), .ZN(n20106) );
  AOI211_X1 U23176 ( .C1(n20104), .C2(n20318), .A(n20099), .B(n20135), .ZN(
        n20100) );
  INV_X1 U23177 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U23178 ( .A1(n20102), .A2(n20137), .B1(n20149), .B2(n20135), .ZN(
        n20109) );
  INV_X1 U23179 ( .A(n20103), .ZN(n20107) );
  OAI21_X1 U23180 ( .B1(n20104), .B2(n20135), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20105) );
  AOI22_X1 U23181 ( .A1(n20150), .A2(n20138), .B1(n20143), .B2(n20159), .ZN(
        n20108) );
  OAI211_X1 U23182 ( .C1(n20142), .C2(n20110), .A(n20109), .B(n20108), .ZN(
        P2_U3160) );
  INV_X1 U23183 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U23184 ( .A1(n20165), .A2(n20143), .B1(n20163), .B2(n20135), .ZN(
        n20113) );
  AOI22_X1 U23185 ( .A1(n20164), .A2(n20138), .B1(n20137), .B2(n20111), .ZN(
        n20112) );
  OAI211_X1 U23186 ( .C1(n20142), .C2(n20114), .A(n20113), .B(n20112), .ZN(
        P2_U3161) );
  INV_X1 U23187 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20118) );
  AOI22_X1 U23188 ( .A1(n20171), .A2(n20143), .B1(n20169), .B2(n20135), .ZN(
        n20117) );
  AOI22_X1 U23189 ( .A1(n20170), .A2(n20138), .B1(n20137), .B2(n20115), .ZN(
        n20116) );
  OAI211_X1 U23190 ( .C1(n20142), .C2(n20118), .A(n20117), .B(n20116), .ZN(
        P2_U3162) );
  INV_X1 U23191 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U23192 ( .A1(n20119), .A2(n20137), .B1(n20175), .B2(n20135), .ZN(
        n20121) );
  AOI22_X1 U23193 ( .A1(n20176), .A2(n20138), .B1(n20143), .B2(n20177), .ZN(
        n20120) );
  OAI211_X1 U23194 ( .C1(n20142), .C2(n20122), .A(n20121), .B(n20120), .ZN(
        P2_U3163) );
  INV_X1 U23195 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U23196 ( .A1(n20183), .A2(n20143), .B1(n20181), .B2(n20135), .ZN(
        n20125) );
  AOI22_X1 U23197 ( .A1(n20182), .A2(n20138), .B1(n20137), .B2(n20123), .ZN(
        n20124) );
  OAI211_X1 U23198 ( .C1(n20142), .C2(n20126), .A(n20125), .B(n20124), .ZN(
        P2_U3164) );
  INV_X1 U23199 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U23200 ( .A1(n20189), .A2(n20143), .B1(n20187), .B2(n20135), .ZN(
        n20129) );
  AOI22_X1 U23201 ( .A1(n20188), .A2(n20138), .B1(n20137), .B2(n20127), .ZN(
        n20128) );
  OAI211_X1 U23202 ( .C1(n20142), .C2(n20130), .A(n20129), .B(n20128), .ZN(
        P2_U3165) );
  INV_X1 U23203 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U23204 ( .A1(n20195), .A2(n20143), .B1(n20193), .B2(n20135), .ZN(
        n20133) );
  AOI22_X1 U23205 ( .A1(n20194), .A2(n20138), .B1(n20137), .B2(n20131), .ZN(
        n20132) );
  OAI211_X1 U23206 ( .C1(n20142), .C2(n20134), .A(n20133), .B(n20132), .ZN(
        P2_U3166) );
  INV_X1 U23207 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U23208 ( .A1(n20203), .A2(n20143), .B1(n20199), .B2(n20135), .ZN(
        n20140) );
  AOI22_X1 U23209 ( .A1(n20201), .A2(n20138), .B1(n20137), .B2(n20136), .ZN(
        n20139) );
  OAI211_X1 U23210 ( .C1(n20142), .C2(n20141), .A(n20140), .B(n20139), .ZN(
        P2_U3167) );
  INV_X1 U23211 ( .A(n20144), .ZN(n20200) );
  NOR3_X1 U23212 ( .A1(n12453), .A2(n20200), .A3(n20145), .ZN(n20151) );
  NAND2_X1 U23213 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20146), .ZN(
        n20157) );
  INV_X1 U23214 ( .A(n20157), .ZN(n20147) );
  AOI21_X1 U23215 ( .B1(n20147), .B2(n20318), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20148) );
  AOI22_X1 U23216 ( .A1(n20202), .A2(n20150), .B1(n20200), .B2(n20149), .ZN(
        n20161) );
  INV_X1 U23217 ( .A(n20151), .ZN(n20153) );
  OAI211_X1 U23218 ( .C1(n20200), .C2(n20318), .A(n20153), .B(n20152), .ZN(
        n20154) );
  AOI221_X1 U23219 ( .B1(n20157), .B2(n20156), .C1(n20157), .C2(n20155), .A(
        n20154), .ZN(n20158) );
  AOI22_X1 U23220 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20159), .ZN(n20160) );
  OAI211_X1 U23221 ( .C1(n20162), .C2(n20208), .A(n20161), .B(n20160), .ZN(
        P2_U3168) );
  AOI22_X1 U23222 ( .A1(n20202), .A2(n20164), .B1(n20200), .B2(n20163), .ZN(
        n20167) );
  AOI22_X1 U23223 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20165), .ZN(n20166) );
  OAI211_X1 U23224 ( .C1(n20168), .C2(n20208), .A(n20167), .B(n20166), .ZN(
        P2_U3169) );
  AOI22_X1 U23225 ( .A1(n20202), .A2(n20170), .B1(n20200), .B2(n20169), .ZN(
        n20173) );
  AOI22_X1 U23226 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20171), .ZN(n20172) );
  OAI211_X1 U23227 ( .C1(n20174), .C2(n20208), .A(n20173), .B(n20172), .ZN(
        P2_U3170) );
  AOI22_X1 U23228 ( .A1(n20202), .A2(n20176), .B1(n20200), .B2(n20175), .ZN(
        n20179) );
  AOI22_X1 U23229 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20177), .ZN(n20178) );
  OAI211_X1 U23230 ( .C1(n20180), .C2(n20208), .A(n20179), .B(n20178), .ZN(
        P2_U3171) );
  AOI22_X1 U23231 ( .A1(n20202), .A2(n20182), .B1(n20200), .B2(n20181), .ZN(
        n20185) );
  AOI22_X1 U23232 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20183), .ZN(n20184) );
  OAI211_X1 U23233 ( .C1(n20186), .C2(n20208), .A(n20185), .B(n20184), .ZN(
        P2_U3172) );
  AOI22_X1 U23234 ( .A1(n20202), .A2(n20188), .B1(n20200), .B2(n20187), .ZN(
        n20191) );
  AOI22_X1 U23235 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20189), .ZN(n20190) );
  OAI211_X1 U23236 ( .C1(n20192), .C2(n20208), .A(n20191), .B(n20190), .ZN(
        P2_U3173) );
  AOI22_X1 U23237 ( .A1(n20202), .A2(n20194), .B1(n20200), .B2(n20193), .ZN(
        n20197) );
  AOI22_X1 U23238 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20195), .ZN(n20196) );
  OAI211_X1 U23239 ( .C1(n20198), .C2(n20208), .A(n20197), .B(n20196), .ZN(
        P2_U3174) );
  AOI22_X1 U23240 ( .A1(n20202), .A2(n20201), .B1(n20200), .B2(n20199), .ZN(
        n20207) );
  AOI22_X1 U23241 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20205), .B1(
        n20204), .B2(n20203), .ZN(n20206) );
  OAI211_X1 U23242 ( .C1(n20209), .C2(n20208), .A(n20207), .B(n20206), .ZN(
        P2_U3175) );
  AND2_X1 U23243 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20210), .ZN(
        P2_U3179) );
  AND2_X1 U23244 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20210), .ZN(
        P2_U3180) );
  INV_X1 U23245 ( .A(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n21351) );
  NOR2_X1 U23246 ( .A1(n21351), .A2(n20293), .ZN(P2_U3181) );
  AND2_X1 U23247 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20210), .ZN(
        P2_U3182) );
  NOR2_X1 U23248 ( .A1(n21346), .A2(n20293), .ZN(P2_U3183) );
  AND2_X1 U23249 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20210), .ZN(
        P2_U3184) );
  INV_X1 U23250 ( .A(P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21333) );
  NOR2_X1 U23251 ( .A1(n21333), .A2(n20293), .ZN(P2_U3185) );
  AND2_X1 U23252 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20210), .ZN(
        P2_U3186) );
  AND2_X1 U23253 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20210), .ZN(
        P2_U3187) );
  AND2_X1 U23254 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20210), .ZN(
        P2_U3188) );
  AND2_X1 U23255 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20210), .ZN(
        P2_U3189) );
  AND2_X1 U23256 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20210), .ZN(
        P2_U3190) );
  AND2_X1 U23257 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20210), .ZN(
        P2_U3191) );
  NOR2_X1 U23258 ( .A1(n21352), .A2(n20293), .ZN(P2_U3192) );
  AND2_X1 U23259 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20210), .ZN(
        P2_U3193) );
  AND2_X1 U23260 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20210), .ZN(
        P2_U3194) );
  AND2_X1 U23261 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20210), .ZN(
        P2_U3195) );
  AND2_X1 U23262 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20210), .ZN(
        P2_U3196) );
  AND2_X1 U23263 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20210), .ZN(
        P2_U3197) );
  AND2_X1 U23264 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20210), .ZN(
        P2_U3198) );
  AND2_X1 U23265 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20210), .ZN(
        P2_U3199) );
  AND2_X1 U23266 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20210), .ZN(
        P2_U3200) );
  AND2_X1 U23267 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20210), .ZN(P2_U3201) );
  AND2_X1 U23268 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20210), .ZN(P2_U3202) );
  AND2_X1 U23269 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20210), .ZN(P2_U3203) );
  AND2_X1 U23270 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20210), .ZN(P2_U3204) );
  AND2_X1 U23271 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20210), .ZN(P2_U3205) );
  INV_X1 U23272 ( .A(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21379) );
  NOR2_X1 U23273 ( .A1(n21379), .A2(n20293), .ZN(P2_U3206) );
  AND2_X1 U23274 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20210), .ZN(P2_U3207) );
  AND2_X1 U23275 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20210), .ZN(P2_U3208) );
  NOR2_X1 U23276 ( .A1(n21248), .A2(n20218), .ZN(n20230) );
  INV_X1 U23277 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20216) );
  NOR2_X1 U23278 ( .A1(n20211), .A2(n20216), .ZN(n20212) );
  NAND2_X1 U23279 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20224), .ZN(n20225) );
  AOI21_X1 U23280 ( .B1(n20212), .B2(n20225), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20215) );
  AOI211_X1 U23281 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21254), .A(
        n20213), .B(n20347), .ZN(n20214) );
  OR3_X1 U23282 ( .A1(n20230), .A2(n20215), .A3(n20214), .ZN(P2_U3209) );
  AOI21_X1 U23283 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21254), .A(n20231), 
        .ZN(n20222) );
  NOR2_X1 U23284 ( .A1(n20216), .A2(n20222), .ZN(n20219) );
  AOI21_X1 U23285 ( .B1(n20219), .B2(n20218), .A(n20217), .ZN(n20220) );
  OAI211_X1 U23286 ( .C1(n21254), .C2(n20221), .A(n20220), .B(n20225), .ZN(
        P2_U3210) );
  AOI21_X1 U23287 ( .B1(n20224), .B2(n20223), .A(n20222), .ZN(n20229) );
  OAI22_X1 U23288 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20226), .B1(NA), 
        .B2(n20225), .ZN(n20227) );
  OAI211_X1 U23289 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20227), .ZN(n20228) );
  OAI21_X1 U23290 ( .B1(n20230), .B2(n20229), .A(n20228), .ZN(P2_U3211) );
  OAI222_X1 U23291 ( .A1(n20284), .A2(n20234), .B1(n20233), .B2(n20347), .C1(
        n20232), .C2(n20281), .ZN(P2_U3212) );
  INV_X1 U23292 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20235) );
  OAI222_X1 U23293 ( .A1(n20284), .A2(n20235), .B1(n21345), .B2(n20347), .C1(
        n20234), .C2(n20281), .ZN(P2_U3213) );
  OAI222_X1 U23294 ( .A1(n20284), .A2(n11820), .B1(n20236), .B2(n20347), .C1(
        n20235), .C2(n20281), .ZN(P2_U3214) );
  OAI222_X1 U23295 ( .A1(n20284), .A2(n11827), .B1(n20237), .B2(n20347), .C1(
        n11820), .C2(n20281), .ZN(P2_U3215) );
  OAI222_X1 U23296 ( .A1(n20284), .A2(n20239), .B1(n20238), .B2(n20347), .C1(
        n11827), .C2(n20281), .ZN(P2_U3216) );
  OAI222_X1 U23297 ( .A1(n20284), .A2(n20241), .B1(n20240), .B2(n20347), .C1(
        n20239), .C2(n20281), .ZN(P2_U3217) );
  OAI222_X1 U23298 ( .A1(n20284), .A2(n20243), .B1(n20242), .B2(n20347), .C1(
        n20241), .C2(n20281), .ZN(P2_U3218) );
  OAI222_X1 U23299 ( .A1(n20284), .A2(n20245), .B1(n20244), .B2(n20347), .C1(
        n20243), .C2(n20281), .ZN(P2_U3219) );
  OAI222_X1 U23300 ( .A1(n20284), .A2(n20247), .B1(n20246), .B2(n20347), .C1(
        n20245), .C2(n20281), .ZN(P2_U3220) );
  OAI222_X1 U23301 ( .A1(n20284), .A2(n13488), .B1(n20248), .B2(n20347), .C1(
        n20247), .C2(n20281), .ZN(P2_U3221) );
  OAI222_X1 U23302 ( .A1(n20284), .A2(n20250), .B1(n20249), .B2(n20347), .C1(
        n13488), .C2(n20281), .ZN(P2_U3222) );
  OAI222_X1 U23303 ( .A1(n20284), .A2(n16131), .B1(n20251), .B2(n20347), .C1(
        n20250), .C2(n20281), .ZN(P2_U3223) );
  OAI222_X1 U23304 ( .A1(n20284), .A2(n16119), .B1(n20252), .B2(n20347), .C1(
        n16131), .C2(n20281), .ZN(P2_U3224) );
  OAI222_X1 U23305 ( .A1(n20284), .A2(n20254), .B1(n20253), .B2(n20347), .C1(
        n16119), .C2(n20281), .ZN(P2_U3225) );
  OAI222_X1 U23306 ( .A1(n20284), .A2(n16091), .B1(n20255), .B2(n20347), .C1(
        n20254), .C2(n20281), .ZN(P2_U3226) );
  OAI222_X1 U23307 ( .A1(n20284), .A2(n20257), .B1(n20256), .B2(n20347), .C1(
        n16091), .C2(n20281), .ZN(P2_U3227) );
  OAI222_X1 U23308 ( .A1(n20284), .A2(n16074), .B1(n20258), .B2(n20347), .C1(
        n20257), .C2(n20281), .ZN(P2_U3228) );
  OAI222_X1 U23309 ( .A1(n20284), .A2(n20260), .B1(n20259), .B2(n20347), .C1(
        n16074), .C2(n20281), .ZN(P2_U3229) );
  OAI222_X1 U23310 ( .A1(n20284), .A2(n20262), .B1(n20261), .B2(n20347), .C1(
        n20260), .C2(n20281), .ZN(P2_U3230) );
  OAI222_X1 U23311 ( .A1(n20284), .A2(n20264), .B1(n20263), .B2(n20347), .C1(
        n20262), .C2(n20281), .ZN(P2_U3231) );
  INV_X1 U23312 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20266) );
  OAI222_X1 U23313 ( .A1(n20284), .A2(n20266), .B1(n20265), .B2(n20347), .C1(
        n20264), .C2(n20281), .ZN(P2_U3232) );
  OAI222_X1 U23314 ( .A1(n20284), .A2(n20268), .B1(n20267), .B2(n20347), .C1(
        n20266), .C2(n20281), .ZN(P2_U3233) );
  OAI222_X1 U23315 ( .A1(n20284), .A2(n20270), .B1(n20269), .B2(n20347), .C1(
        n20268), .C2(n20281), .ZN(P2_U3234) );
  OAI222_X1 U23316 ( .A1(n20284), .A2(n20272), .B1(n20271), .B2(n20347), .C1(
        n20270), .C2(n20281), .ZN(P2_U3235) );
  INV_X1 U23317 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20274) );
  OAI222_X1 U23318 ( .A1(n20284), .A2(n20274), .B1(n20273), .B2(n20347), .C1(
        n20272), .C2(n20281), .ZN(P2_U3236) );
  OAI222_X1 U23319 ( .A1(n20284), .A2(n20276), .B1(n20275), .B2(n20347), .C1(
        n20274), .C2(n20281), .ZN(P2_U3237) );
  OAI222_X1 U23320 ( .A1(n20281), .A2(n20276), .B1(n21349), .B2(n20347), .C1(
        n20277), .C2(n20284), .ZN(P2_U3238) );
  OAI222_X1 U23321 ( .A1(n20284), .A2(n20279), .B1(n20278), .B2(n20347), .C1(
        n20277), .C2(n20281), .ZN(P2_U3239) );
  INV_X1 U23322 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20282) );
  OAI222_X1 U23323 ( .A1(n20284), .A2(n20282), .B1(n20280), .B2(n20347), .C1(
        n20279), .C2(n20281), .ZN(P2_U3240) );
  OAI222_X1 U23324 ( .A1(n20284), .A2(n12326), .B1(n20283), .B2(n20347), .C1(
        n20282), .C2(n20281), .ZN(P2_U3241) );
  INV_X1 U23325 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20285) );
  AOI22_X1 U23326 ( .A1(n20347), .A2(n20286), .B1(n20285), .B2(n20336), .ZN(
        P2_U3585) );
  MUX2_X1 U23327 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20347), .Z(P2_U3586) );
  INV_X1 U23328 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20287) );
  AOI22_X1 U23329 ( .A1(n20347), .A2(n20288), .B1(n20287), .B2(n20336), .ZN(
        P2_U3587) );
  INV_X1 U23330 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20289) );
  AOI22_X1 U23331 ( .A1(n20347), .A2(n21398), .B1(n20289), .B2(n20336), .ZN(
        P2_U3588) );
  OAI21_X1 U23332 ( .B1(n20293), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20291), 
        .ZN(n20290) );
  INV_X1 U23333 ( .A(n20290), .ZN(P2_U3591) );
  OAI21_X1 U23334 ( .B1(n20293), .B2(n20292), .A(n20291), .ZN(P2_U3592) );
  INV_X1 U23335 ( .A(n20294), .ZN(n20295) );
  OAI222_X1 U23336 ( .A1(n20300), .A2(n20299), .B1(n20298), .B2(n20297), .C1(
        n20296), .C2(n20295), .ZN(n20302) );
  MUX2_X1 U23337 ( .A(n20302), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n20301), .Z(P2_U3599) );
  NOR2_X1 U23338 ( .A1(n20304), .A2(n20303), .ZN(n20320) );
  NOR2_X1 U23339 ( .A1(n20305), .A2(n16495), .ZN(n20307) );
  INV_X1 U23340 ( .A(n20306), .ZN(n20329) );
  AOI21_X1 U23341 ( .B1(n20308), .B2(n20307), .A(n20329), .ZN(n20322) );
  OAI21_X1 U23342 ( .B1(n20320), .B2(n20322), .A(n20309), .ZN(n20312) );
  OR2_X1 U23343 ( .A1(n20310), .A2(n20318), .ZN(n20311) );
  OAI211_X1 U23344 ( .C1(n20314), .C2(n20313), .A(n20312), .B(n20311), .ZN(
        n20315) );
  INV_X1 U23345 ( .A(n20315), .ZN(n20316) );
  AOI22_X1 U23346 ( .A1(n20333), .A2(n20317), .B1(n20316), .B2(n20334), .ZN(
        P2_U3602) );
  NOR2_X1 U23347 ( .A1(n20319), .A2(n20318), .ZN(n20321) );
  AOI211_X1 U23348 ( .C1(n20323), .C2(n20322), .A(n20321), .B(n20320), .ZN(
        n20324) );
  AOI22_X1 U23349 ( .A1(n20333), .A2(n20325), .B1(n20324), .B2(n20334), .ZN(
        P2_U3603) );
  INV_X1 U23350 ( .A(n20326), .ZN(n20328) );
  OAI22_X1 U23351 ( .A1(n20330), .A2(n20329), .B1(n20328), .B2(n20327), .ZN(
        n20331) );
  AOI21_X1 U23352 ( .B1(n20335), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20331), 
        .ZN(n20332) );
  OAI22_X1 U23353 ( .A1(n20335), .A2(n20334), .B1(n20333), .B2(n20332), .ZN(
        P2_U3605) );
  INV_X1 U23354 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20337) );
  AOI22_X1 U23355 ( .A1(n20347), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20337), 
        .B2(n20336), .ZN(P2_U3608) );
  INV_X1 U23356 ( .A(n20338), .ZN(n20340) );
  AOI22_X1 U23357 ( .A1(n20342), .A2(n20341), .B1(n20340), .B2(n20339), .ZN(
        n20343) );
  NAND2_X1 U23358 ( .A1(n20344), .A2(n20343), .ZN(n20346) );
  MUX2_X1 U23359 ( .A(P2_MORE_REG_SCAN_IN), .B(n20346), .S(n20345), .Z(
        P2_U3609) );
  MUX2_X1 U23360 ( .A(P2_M_IO_N_REG_SCAN_IN), .B(P2_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20347), .Z(P2_U3611) );
  OAI21_X1 U23361 ( .B1(n20349), .B2(n20348), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20350) );
  OAI21_X1 U23362 ( .B1(n20352), .B2(n20351), .A(n20350), .ZN(P1_U2803) );
  INV_X1 U23363 ( .A(n21271), .ZN(n21275) );
  OAI21_X1 U23364 ( .B1(BS16), .B2(n20353), .A(n21275), .ZN(n21273) );
  OAI21_X1 U23365 ( .B1(n21275), .B2(n20900), .A(n21273), .ZN(P1_U2805) );
  OAI21_X1 U23366 ( .B1(n20355), .B2(n20354), .A(n15151), .ZN(P1_U2806) );
  NOR4_X1 U23367 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20359) );
  NOR4_X1 U23368 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20358) );
  NOR4_X1 U23369 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20357) );
  NOR4_X1 U23370 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20356) );
  NAND4_X1 U23371 ( .A1(n20359), .A2(n20358), .A3(n20357), .A4(n20356), .ZN(
        n20365) );
  NOR4_X1 U23372 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20363) );
  AOI211_X1 U23373 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20362) );
  NOR4_X1 U23374 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20361) );
  NOR4_X1 U23375 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20360) );
  NAND4_X1 U23376 ( .A1(n20363), .A2(n20362), .A3(n20361), .A4(n20360), .ZN(
        n20364) );
  NOR2_X1 U23377 ( .A1(n20365), .A2(n20364), .ZN(n21290) );
  NOR3_X1 U23378 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20368) );
  OAI21_X1 U23379 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20368), .A(n21290), .ZN(
        n20366) );
  OAI21_X1 U23380 ( .B1(n21290), .B2(n20367), .A(n20366), .ZN(P1_U2807) );
  INV_X1 U23381 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21274) );
  AOI21_X1 U23382 ( .B1(n21284), .B2(n21274), .A(n20368), .ZN(n20371) );
  INV_X1 U23383 ( .A(n21290), .ZN(n20369) );
  AOI22_X1 U23384 ( .A1(n21290), .A2(n20371), .B1(n20370), .B2(n20369), .ZN(
        P1_U2808) );
  OAI21_X1 U23385 ( .B1(n20399), .B2(n20372), .A(n20397), .ZN(n20384) );
  OAI22_X1 U23386 ( .A1(n20374), .A2(n20402), .B1(n20408), .B2(n20373), .ZN(
        n20375) );
  AOI21_X1 U23387 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n20411), .A(n20375), .ZN(
        n20379) );
  NAND2_X1 U23388 ( .A1(n20376), .A2(n13435), .ZN(n20378) );
  NAND2_X1 U23389 ( .A1(n20430), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20377) );
  OAI221_X1 U23390 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20382), .C1(n20381), 
        .C2(n20384), .A(n20380), .ZN(P1_U2833) );
  NAND2_X1 U23391 ( .A1(n20433), .A2(n20383), .ZN(n20385) );
  AOI21_X1 U23392 ( .B1(n20386), .B2(n20385), .A(n20384), .ZN(n20389) );
  INV_X1 U23393 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20447) );
  AOI22_X1 U23394 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20430), .B1(
        n20425), .B2(n20444), .ZN(n20387) );
  OAI211_X1 U23395 ( .C1(n20442), .C2(n20447), .A(n20387), .B(n20416), .ZN(
        n20388) );
  AOI211_X1 U23396 ( .C1(n20445), .C2(n13435), .A(n20389), .B(n20388), .ZN(
        n20390) );
  OAI21_X1 U23397 ( .B1(n20391), .B2(n20402), .A(n20390), .ZN(P1_U2834) );
  NOR3_X1 U23398 ( .A1(n20392), .A2(P1_REIP_REG_5__SCAN_IN), .A3(n20398), .ZN(
        n20396) );
  OAI21_X1 U23399 ( .B1(n20394), .B2(n20393), .A(n20416), .ZN(n20395) );
  AOI211_X1 U23400 ( .C1(n20411), .C2(P1_EBX_REG_5__SCAN_IN), .A(n20396), .B(
        n20395), .ZN(n20406) );
  OAI21_X1 U23401 ( .B1(n20399), .B2(n20398), .A(n20397), .ZN(n20422) );
  OAI22_X1 U23402 ( .A1(n20402), .A2(n20401), .B1(n20400), .B2(n20422), .ZN(
        n20403) );
  AOI21_X1 U23403 ( .B1(n20404), .B2(n20419), .A(n20403), .ZN(n20405) );
  OAI211_X1 U23404 ( .C1(n20408), .C2(n20407), .A(n20406), .B(n20405), .ZN(
        P1_U2835) );
  NOR3_X1 U23405 ( .A1(n21284), .A2(n21258), .A3(n20432), .ZN(n20409) );
  AOI21_X1 U23406 ( .B1(n20433), .B2(n20409), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n20423) );
  AOI21_X1 U23407 ( .B1(n20410), .B2(n13886), .A(n10125), .ZN(n20527) );
  AOI22_X1 U23408 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(n20411), .B1(n20425), .B2(
        n20527), .ZN(n20417) );
  OR2_X1 U23409 ( .A1(n20413), .A2(n20412), .ZN(n20415) );
  NAND2_X1 U23410 ( .A1(n20430), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20414) );
  AND4_X1 U23411 ( .A1(n20417), .A2(n20416), .A3(n20415), .A4(n20414), .ZN(
        n20421) );
  INV_X1 U23412 ( .A(n20523), .ZN(n20418) );
  AOI22_X1 U23413 ( .A1(n20520), .A2(n20419), .B1(n20418), .B2(n20426), .ZN(
        n20420) );
  OAI211_X1 U23414 ( .C1(n20423), .C2(n20422), .A(n20421), .B(n20420), .ZN(
        P1_U2836) );
  INV_X1 U23415 ( .A(n20424), .ZN(n20543) );
  AOI22_X1 U23416 ( .A1(n20427), .A2(n20426), .B1(n20425), .B2(n20543), .ZN(
        n20441) );
  NAND2_X1 U23417 ( .A1(n20429), .A2(n20428), .ZN(n20439) );
  AOI22_X1 U23418 ( .A1(n20431), .A2(n21031), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20430), .ZN(n20435) );
  NAND3_X1 U23419 ( .A1(n20433), .A2(n20432), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n20434) );
  OAI211_X1 U23420 ( .C1(n20437), .C2(n20436), .A(n20435), .B(n20434), .ZN(
        n20438) );
  AOI21_X1 U23421 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n20439), .A(n20438), .ZN(
        n20440) );
  OAI211_X1 U23422 ( .C1(n20443), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P1_U2838) );
  AOI22_X1 U23423 ( .A1(n20445), .A2(n20449), .B1(n20448), .B2(n20444), .ZN(
        n20446) );
  OAI21_X1 U23424 ( .B1(n20452), .B2(n20447), .A(n20446), .ZN(P1_U2866) );
  INV_X1 U23425 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20451) );
  AOI22_X1 U23426 ( .A1(n20520), .A2(n20449), .B1(n20448), .B2(n20527), .ZN(
        n20450) );
  OAI21_X1 U23427 ( .B1(n20452), .B2(n20451), .A(n20450), .ZN(P1_U2868) );
  AOI22_X1 U23428 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20453), .B1(n20471), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20454) );
  OAI21_X1 U23429 ( .B1(n20456), .B2(n20455), .A(n20454), .ZN(P1_U2921) );
  INV_X1 U23430 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20458) );
  AOI22_X1 U23431 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20457) );
  OAI21_X1 U23432 ( .B1(n20458), .B2(n20484), .A(n20457), .ZN(P1_U2922) );
  INV_X1 U23433 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20460) );
  AOI22_X1 U23434 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20459) );
  OAI21_X1 U23435 ( .B1(n20460), .B2(n20484), .A(n20459), .ZN(P1_U2923) );
  INV_X1 U23436 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20462) );
  AOI22_X1 U23437 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20461) );
  OAI21_X1 U23438 ( .B1(n20462), .B2(n20484), .A(n20461), .ZN(P1_U2924) );
  INV_X1 U23439 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20464) );
  AOI22_X1 U23440 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20463) );
  OAI21_X1 U23441 ( .B1(n20464), .B2(n20484), .A(n20463), .ZN(P1_U2925) );
  AOI22_X1 U23442 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20465) );
  OAI21_X1 U23443 ( .B1(n14933), .B2(n20484), .A(n20465), .ZN(P1_U2926) );
  INV_X1 U23444 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20467) );
  AOI22_X1 U23445 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20466) );
  OAI21_X1 U23446 ( .B1(n20467), .B2(n20484), .A(n20466), .ZN(P1_U2927) );
  INV_X1 U23447 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20469) );
  AOI22_X1 U23448 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20468) );
  OAI21_X1 U23449 ( .B1(n20469), .B2(n20484), .A(n20468), .ZN(P1_U2928) );
  AOI22_X1 U23450 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20470) );
  OAI21_X1 U23451 ( .B1(n10829), .B2(n20484), .A(n20470), .ZN(P1_U2929) );
  AOI22_X1 U23452 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20472) );
  OAI21_X1 U23453 ( .B1(n10823), .B2(n20484), .A(n20472), .ZN(P1_U2930) );
  AOI22_X1 U23454 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20473) );
  OAI21_X1 U23455 ( .B1(n20474), .B2(n20484), .A(n20473), .ZN(P1_U2931) );
  AOI22_X1 U23456 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20475) );
  OAI21_X1 U23457 ( .B1(n20476), .B2(n20484), .A(n20475), .ZN(P1_U2932) );
  AOI22_X1 U23458 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20477) );
  OAI21_X1 U23459 ( .B1(n20478), .B2(n20484), .A(n20477), .ZN(P1_U2933) );
  AOI22_X1 U23460 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20479) );
  OAI21_X1 U23461 ( .B1(n20480), .B2(n20484), .A(n20479), .ZN(P1_U2934) );
  AOI22_X1 U23462 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20481) );
  OAI21_X1 U23463 ( .B1(n20482), .B2(n20484), .A(n20481), .ZN(P1_U2935) );
  AOI22_X1 U23464 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21292), .B1(n20471), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20483) );
  OAI21_X1 U23465 ( .B1(n20485), .B2(n20484), .A(n20483), .ZN(P1_U2936) );
  AOI22_X1 U23466 ( .A1(n20509), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20512), .ZN(n20487) );
  NAND2_X1 U23467 ( .A1(n20497), .A2(n20486), .ZN(n20499) );
  NAND2_X1 U23468 ( .A1(n20487), .A2(n20499), .ZN(P1_U2945) );
  AOI22_X1 U23469 ( .A1(n20509), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20489) );
  NAND2_X1 U23470 ( .A1(n20497), .A2(n20488), .ZN(n20501) );
  NAND2_X1 U23471 ( .A1(n20489), .A2(n20501), .ZN(P1_U2946) );
  AOI22_X1 U23472 ( .A1(n20509), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20491) );
  NAND2_X1 U23473 ( .A1(n20497), .A2(n20490), .ZN(n20503) );
  NAND2_X1 U23474 ( .A1(n20491), .A2(n20503), .ZN(P1_U2947) );
  AOI22_X1 U23475 ( .A1(n20509), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20493) );
  NAND2_X1 U23476 ( .A1(n20497), .A2(n20492), .ZN(n20505) );
  NAND2_X1 U23477 ( .A1(n20493), .A2(n20505), .ZN(P1_U2948) );
  AOI22_X1 U23478 ( .A1(n20509), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20495) );
  NAND2_X1 U23479 ( .A1(n20497), .A2(n20494), .ZN(n20507) );
  NAND2_X1 U23480 ( .A1(n20495), .A2(n20507), .ZN(P1_U2949) );
  AOI22_X1 U23481 ( .A1(n20509), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20512), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20498) );
  NAND2_X1 U23482 ( .A1(n20497), .A2(n20496), .ZN(n20513) );
  NAND2_X1 U23483 ( .A1(n20498), .A2(n20513), .ZN(P1_U2951) );
  AOI22_X1 U23484 ( .A1(n20509), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20500) );
  NAND2_X1 U23485 ( .A1(n20500), .A2(n20499), .ZN(P1_U2960) );
  AOI22_X1 U23486 ( .A1(n20509), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20512), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20502) );
  NAND2_X1 U23487 ( .A1(n20502), .A2(n20501), .ZN(P1_U2961) );
  AOI22_X1 U23488 ( .A1(n20509), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20512), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20504) );
  NAND2_X1 U23489 ( .A1(n20504), .A2(n20503), .ZN(P1_U2962) );
  AOI22_X1 U23490 ( .A1(n20509), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20512), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20506) );
  NAND2_X1 U23491 ( .A1(n20506), .A2(n20505), .ZN(P1_U2963) );
  AOI22_X1 U23492 ( .A1(n20509), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20512), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20508) );
  NAND2_X1 U23493 ( .A1(n20508), .A2(n20507), .ZN(P1_U2964) );
  AOI22_X1 U23494 ( .A1(n20509), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20512), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20511) );
  NAND2_X1 U23495 ( .A1(n20511), .A2(n20510), .ZN(P1_U2965) );
  AOI22_X1 U23496 ( .A1(n20509), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20512), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20514) );
  NAND2_X1 U23497 ( .A1(n20514), .A2(n20513), .ZN(P1_U2966) );
  AOI22_X1 U23498 ( .A1(n17105), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20580), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20522) );
  XNOR2_X1 U23499 ( .A(n20515), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20516) );
  XNOR2_X1 U23500 ( .A(n20517), .B(n20516), .ZN(n20530) );
  AOI22_X1 U23501 ( .A1(n20520), .A2(n20519), .B1(n20530), .B2(n20518), .ZN(
        n20521) );
  OAI211_X1 U23502 ( .C1(n20524), .C2(n20523), .A(n20522), .B(n20521), .ZN(
        P1_U2995) );
  AOI21_X1 U23503 ( .B1(n20573), .B2(n20526), .A(n20525), .ZN(n20538) );
  AOI22_X1 U23504 ( .A1(n20544), .A2(n20527), .B1(n20580), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20532) );
  AOI211_X1 U23505 ( .C1(n20539), .C2(n20533), .A(n20528), .B(n20540), .ZN(
        n20529) );
  AOI21_X1 U23506 ( .B1(n20530), .B2(n20550), .A(n20529), .ZN(n20531) );
  OAI211_X1 U23507 ( .C1(n20538), .C2(n20533), .A(n20532), .B(n20531), .ZN(
        P1_U3027) );
  OAI222_X1 U23508 ( .A1(n20535), .A2(n20578), .B1(n20416), .B2(n21258), .C1(
        n20576), .C2(n20534), .ZN(n20536) );
  INV_X1 U23509 ( .A(n20536), .ZN(n20537) );
  OAI221_X1 U23510 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20540), .C1(
        n20539), .C2(n20538), .A(n20537), .ZN(P1_U3028) );
  NAND2_X1 U23511 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20542) );
  OAI21_X1 U23512 ( .B1(n20542), .B2(n20552), .A(n20541), .ZN(n20545) );
  AOI22_X1 U23513 ( .A1(n20573), .A2(n20545), .B1(n20544), .B2(n20543), .ZN(
        n20557) );
  INV_X1 U23514 ( .A(n20546), .ZN(n20548) );
  OAI21_X1 U23515 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20548), .A(
        n20547), .ZN(n20549) );
  AOI22_X1 U23516 ( .A1(n20551), .A2(n20550), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20549), .ZN(n20556) );
  NAND2_X1 U23517 ( .A1(n20580), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20555) );
  NAND3_X1 U23518 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20553), .A3(
        n20552), .ZN(n20554) );
  NAND4_X1 U23519 ( .A1(n20557), .A2(n20556), .A3(n20555), .A4(n20554), .ZN(
        P1_U3029) );
  AOI21_X1 U23520 ( .B1(n20573), .B2(n20559), .A(n20558), .ZN(n20583) );
  OAI21_X1 U23521 ( .B1(n20578), .B2(n20561), .A(n20560), .ZN(n20562) );
  INV_X1 U23522 ( .A(n20562), .ZN(n20570) );
  NOR3_X1 U23523 ( .A1(n20564), .A2(n20563), .A3(n20576), .ZN(n20568) );
  NOR3_X1 U23524 ( .A1(n20566), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20565), .ZN(n20567) );
  NOR2_X1 U23525 ( .A1(n20568), .A2(n20567), .ZN(n20569) );
  OAI211_X1 U23526 ( .C1(n20583), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3030) );
  INV_X1 U23527 ( .A(n20572), .ZN(n20574) );
  NOR3_X1 U23528 ( .A1(n20574), .A2(n20573), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20584) );
  OAI22_X1 U23529 ( .A1(n20578), .A2(n20577), .B1(n20576), .B2(n20575), .ZN(
        n20579) );
  AOI21_X1 U23530 ( .B1(n20580), .B2(P1_REIP_REG_0__SCAN_IN), .A(n20579), .ZN(
        n20581) );
  OAI221_X1 U23531 ( .B1(n20584), .B2(n20583), .C1(n20584), .C2(n20582), .A(
        n20581), .ZN(P1_U3031) );
  NOR2_X1 U23532 ( .A1(n20586), .A2(n20585), .ZN(P1_U3032) );
  INV_X1 U23533 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20596) );
  INV_X1 U23534 ( .A(DATAI_24_), .ZN(n20587) );
  OAI22_X2 U23535 ( .A1(n20588), .A2(n20644), .B1(n20587), .B2(n20646), .ZN(
        n21187) );
  OR2_X1 U23536 ( .A1(n10432), .A2(n20589), .ZN(n21034) );
  AOI22_X1 U23537 ( .A1(n21221), .A2(n21187), .B1(n20590), .B2(n21176), .ZN(
        n20595) );
  INV_X1 U23538 ( .A(n20690), .ZN(n20603) );
  INV_X1 U23539 ( .A(DATAI_16_), .ZN(n20592) );
  OAI22_X1 U23540 ( .A1(n20593), .A2(n20644), .B1(n20592), .B2(n20646), .ZN(
        n21095) );
  AOI22_X1 U23541 ( .A1(n21177), .A2(n20654), .B1(n20603), .B2(n21095), .ZN(
        n20594) );
  OAI211_X1 U23542 ( .C1(n20613), .C2(n20596), .A(n20595), .B(n20594), .ZN(
        P1_U3033) );
  INV_X1 U23543 ( .A(DATAI_25_), .ZN(n20597) );
  INV_X1 U23544 ( .A(n21142), .ZN(n21196) );
  INV_X1 U23545 ( .A(n21191), .ZN(n21047) );
  OAI22_X1 U23546 ( .A1(n21241), .A2(n21196), .B1(n20650), .B2(n21047), .ZN(
        n20599) );
  INV_X1 U23547 ( .A(n20599), .ZN(n20605) );
  INV_X1 U23548 ( .A(DATAI_17_), .ZN(n20602) );
  OAI22_X1 U23549 ( .A1(n20602), .A2(n20646), .B1(n20601), .B2(n20644), .ZN(
        n21193) );
  AOI22_X1 U23550 ( .A1(n21192), .A2(n20654), .B1(n20603), .B2(n21193), .ZN(
        n20604) );
  OAI211_X1 U23551 ( .C1(n20613), .C2(n20606), .A(n20605), .B(n20604), .ZN(
        P1_U3034) );
  INV_X1 U23552 ( .A(DATAI_19_), .ZN(n20607) );
  OAI22_X1 U23553 ( .A1(n20608), .A2(n20644), .B1(n20607), .B2(n20646), .ZN(
        n21208) );
  INV_X1 U23554 ( .A(n21208), .ZN(n21154) );
  INV_X1 U23555 ( .A(DATAI_27_), .ZN(n20609) );
  OAI22_X1 U23556 ( .A1(n20610), .A2(n20644), .B1(n20609), .B2(n20646), .ZN(
        n21151) );
  INV_X1 U23557 ( .A(n21151), .ZN(n21211) );
  INV_X1 U23558 ( .A(n21206), .ZN(n21055) );
  OAI22_X1 U23559 ( .A1(n21241), .A2(n21211), .B1(n20650), .B2(n21055), .ZN(
        n20612) );
  INV_X1 U23560 ( .A(n20612), .ZN(n20616) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20655), .B1(
        n21207), .B2(n20654), .ZN(n20615) );
  OAI211_X1 U23562 ( .C1(n21154), .C2(n20690), .A(n20616), .B(n20615), .ZN(
        P1_U3036) );
  INV_X1 U23563 ( .A(DATAI_20_), .ZN(n20617) );
  OAI22_X1 U23564 ( .A1(n20618), .A2(n20644), .B1(n20617), .B2(n20646), .ZN(
        n21214) );
  INV_X1 U23565 ( .A(n21214), .ZN(n21158) );
  INV_X1 U23566 ( .A(DATAI_28_), .ZN(n20619) );
  INV_X1 U23567 ( .A(n21155), .ZN(n21217) );
  INV_X1 U23568 ( .A(n21212), .ZN(n21060) );
  OAI22_X1 U23569 ( .A1(n21241), .A2(n21217), .B1(n20650), .B2(n21060), .ZN(
        n20621) );
  INV_X1 U23570 ( .A(n20621), .ZN(n20624) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20655), .B1(
        n21213), .B2(n20654), .ZN(n20623) );
  OAI211_X1 U23572 ( .C1(n21158), .C2(n20690), .A(n20624), .B(n20623), .ZN(
        P1_U3037) );
  INV_X1 U23573 ( .A(DATAI_21_), .ZN(n20626) );
  OAI22_X1 U23574 ( .A1(n20626), .A2(n20646), .B1(n20625), .B2(n20644), .ZN(
        n21220) );
  INV_X1 U23575 ( .A(n21220), .ZN(n21162) );
  INV_X1 U23576 ( .A(DATAI_29_), .ZN(n20627) );
  OAI22_X1 U23577 ( .A1(n20628), .A2(n20644), .B1(n20627), .B2(n20646), .ZN(
        n21159) );
  INV_X1 U23578 ( .A(n21159), .ZN(n21225) );
  INV_X1 U23579 ( .A(n21218), .ZN(n21065) );
  OAI22_X1 U23580 ( .A1(n21241), .A2(n21225), .B1(n20650), .B2(n21065), .ZN(
        n20630) );
  INV_X1 U23581 ( .A(n20630), .ZN(n20633) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20655), .B1(
        n21219), .B2(n20654), .ZN(n20632) );
  OAI211_X1 U23583 ( .C1(n21162), .C2(n20690), .A(n20633), .B(n20632), .ZN(
        P1_U3038) );
  INV_X1 U23584 ( .A(DATAI_22_), .ZN(n20634) );
  OAI22_X1 U23585 ( .A1(n20635), .A2(n20644), .B1(n20634), .B2(n20646), .ZN(
        n21114) );
  INV_X1 U23586 ( .A(n21114), .ZN(n21231) );
  INV_X1 U23587 ( .A(DATAI_30_), .ZN(n20636) );
  OAI22_X2 U23588 ( .A1(n20637), .A2(n20644), .B1(n20636), .B2(n20646), .ZN(
        n21228) );
  INV_X1 U23589 ( .A(n21228), .ZN(n21117) );
  INV_X1 U23590 ( .A(n21226), .ZN(n21070) );
  OAI22_X1 U23591 ( .A1(n21241), .A2(n21117), .B1(n20650), .B2(n21070), .ZN(
        n20638) );
  INV_X1 U23592 ( .A(n20638), .ZN(n20641) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20655), .B1(
        n21227), .B2(n20654), .ZN(n20640) );
  OAI211_X1 U23594 ( .C1(n21231), .C2(n20690), .A(n20641), .B(n20640), .ZN(
        P1_U3039) );
  INV_X1 U23595 ( .A(DATAI_23_), .ZN(n20643) );
  OAI22_X1 U23596 ( .A1(n20643), .A2(n20646), .B1(n20642), .B2(n20644), .ZN(
        n21120) );
  INV_X1 U23597 ( .A(DATAI_31_), .ZN(n20647) );
  OAI22_X2 U23598 ( .A1(n20647), .A2(n20646), .B1(n20645), .B2(n20644), .ZN(
        n21236) );
  INV_X1 U23599 ( .A(n21236), .ZN(n21125) );
  INV_X1 U23600 ( .A(n21232), .ZN(n21076) );
  OAI22_X1 U23601 ( .A1(n21241), .A2(n21125), .B1(n20650), .B2(n21076), .ZN(
        n20651) );
  INV_X1 U23602 ( .A(n20651), .ZN(n20657) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20655), .B1(
        n21235), .B2(n20654), .ZN(n20656) );
  OAI211_X1 U23604 ( .C1(n21242), .C2(n20690), .A(n20657), .B(n20656), .ZN(
        P1_U3040) );
  INV_X1 U23605 ( .A(n21187), .ZN(n21098) );
  NOR2_X1 U23606 ( .A1(n21084), .A2(n20659), .ZN(n20685) );
  INV_X1 U23607 ( .A(n20685), .ZN(n20672) );
  OAI21_X1 U23608 ( .B1(n20721), .B2(n20658), .A(n20672), .ZN(n20662) );
  NAND2_X1 U23609 ( .A1(n20662), .A2(n21186), .ZN(n20661) );
  INV_X1 U23610 ( .A(n20659), .ZN(n20666) );
  NAND2_X1 U23611 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20666), .ZN(n20660) );
  NAND2_X1 U23612 ( .A1(n20661), .A2(n20660), .ZN(n20686) );
  AOI22_X1 U23613 ( .A1(n21177), .A2(n20686), .B1(n21176), .B2(n20685), .ZN(
        n20669) );
  INV_X1 U23614 ( .A(n20727), .ZN(n20664) );
  INV_X1 U23615 ( .A(n20662), .ZN(n20663) );
  OAI21_X1 U23616 ( .B1(n20664), .B2(n20900), .A(n20663), .ZN(n20665) );
  OAI221_X1 U23617 ( .B1(n21186), .B2(n20666), .C1(n21184), .C2(n20665), .A(
        n21182), .ZN(n20687) );
  INV_X1 U23618 ( .A(n20936), .ZN(n20667) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21095), .ZN(n20668) );
  OAI211_X1 U23620 ( .C1(n21098), .C2(n20690), .A(n20669), .B(n20668), .ZN(
        P1_U3041) );
  AOI22_X1 U23621 ( .A1(n21192), .A2(n20686), .B1(n21191), .B2(n20685), .ZN(
        n20671) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21193), .ZN(n20670) );
  OAI211_X1 U23623 ( .C1(n21196), .C2(n20690), .A(n20671), .B(n20670), .ZN(
        P1_U3042) );
  INV_X1 U23624 ( .A(n21202), .ZN(n21107) );
  INV_X1 U23625 ( .A(n20686), .ZN(n20673) );
  OAI22_X1 U23626 ( .A1(n21200), .A2(n20673), .B1(n21197), .B2(n20672), .ZN(
        n20674) );
  INV_X1 U23627 ( .A(n20674), .ZN(n20676) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21104), .ZN(n20675) );
  OAI211_X1 U23629 ( .C1(n21107), .C2(n20690), .A(n20676), .B(n20675), .ZN(
        P1_U3043) );
  AOI22_X1 U23630 ( .A1(n21207), .A2(n20686), .B1(n21206), .B2(n20685), .ZN(
        n20678) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21208), .ZN(n20677) );
  OAI211_X1 U23632 ( .C1(n21211), .C2(n20690), .A(n20678), .B(n20677), .ZN(
        P1_U3044) );
  AOI22_X1 U23633 ( .A1(n21213), .A2(n20686), .B1(n21212), .B2(n20685), .ZN(
        n20680) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21214), .ZN(n20679) );
  OAI211_X1 U23635 ( .C1(n21217), .C2(n20690), .A(n20680), .B(n20679), .ZN(
        P1_U3045) );
  AOI22_X1 U23636 ( .A1(n21219), .A2(n20686), .B1(n21218), .B2(n20685), .ZN(
        n20682) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21220), .ZN(n20681) );
  OAI211_X1 U23638 ( .C1(n21225), .C2(n20690), .A(n20682), .B(n20681), .ZN(
        P1_U3046) );
  AOI22_X1 U23639 ( .A1(n21227), .A2(n20686), .B1(n21226), .B2(n20685), .ZN(
        n20684) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21114), .ZN(n20683) );
  OAI211_X1 U23641 ( .C1(n21117), .C2(n20690), .A(n20684), .B(n20683), .ZN(
        P1_U3047) );
  AOI22_X1 U23642 ( .A1(n21235), .A2(n20686), .B1(n21232), .B2(n20685), .ZN(
        n20689) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20687), .B1(
        n20714), .B2(n21120), .ZN(n20688) );
  OAI211_X1 U23644 ( .C1(n21125), .C2(n20690), .A(n20689), .B(n20688), .ZN(
        P1_U3048) );
  NOR3_X1 U23645 ( .A1(n20748), .A2(n20714), .A3(n21184), .ZN(n20692) );
  NOR2_X1 U23646 ( .A1(n20692), .A2(n20961), .ZN(n20698) );
  INV_X1 U23647 ( .A(n20698), .ZN(n20693) );
  NOR2_X1 U23648 ( .A1(n20721), .A2(n14172), .ZN(n20697) );
  NOR3_X1 U23649 ( .A1(n21033), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20728) );
  NAND2_X1 U23650 ( .A1(n21084), .A2(n20728), .ZN(n20695) );
  INV_X1 U23651 ( .A(n20695), .ZN(n20713) );
  AOI22_X1 U23652 ( .A1(n20748), .A2(n21095), .B1(n21176), .B2(n20713), .ZN(
        n20700) );
  NOR2_X1 U23653 ( .A1(n10290), .A2(n21246), .ZN(n20825) );
  AOI211_X1 U23654 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20695), .A(n20825), 
        .B(n20694), .ZN(n20696) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n21187), .ZN(n20699) );
  OAI211_X1 U23656 ( .C1(n20718), .C2(n21046), .A(n20700), .B(n20699), .ZN(
        P1_U3049) );
  INV_X1 U23657 ( .A(n21192), .ZN(n21051) );
  AOI22_X1 U23658 ( .A1(n20714), .A2(n21142), .B1(n21191), .B2(n20713), .ZN(
        n20702) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20715), .B1(
        n20748), .B2(n21193), .ZN(n20701) );
  OAI211_X1 U23660 ( .C1(n20718), .C2(n21051), .A(n20702), .B(n20701), .ZN(
        P1_U3050) );
  AOI22_X1 U23661 ( .A1(n20714), .A2(n21202), .B1(n20976), .B2(n20713), .ZN(
        n20704) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20715), .B1(
        n20748), .B2(n21104), .ZN(n20703) );
  OAI211_X1 U23663 ( .C1(n20718), .C2(n21200), .A(n20704), .B(n20703), .ZN(
        P1_U3051) );
  INV_X1 U23664 ( .A(n21207), .ZN(n21059) );
  AOI22_X1 U23665 ( .A1(n20748), .A2(n21208), .B1(n21206), .B2(n20713), .ZN(
        n20706) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n21151), .ZN(n20705) );
  OAI211_X1 U23667 ( .C1(n20718), .C2(n21059), .A(n20706), .B(n20705), .ZN(
        P1_U3052) );
  INV_X1 U23668 ( .A(n21213), .ZN(n21064) );
  AOI22_X1 U23669 ( .A1(n20748), .A2(n21214), .B1(n21212), .B2(n20713), .ZN(
        n20708) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n21155), .ZN(n20707) );
  OAI211_X1 U23671 ( .C1(n20718), .C2(n21064), .A(n20708), .B(n20707), .ZN(
        P1_U3053) );
  AOI22_X1 U23672 ( .A1(n20748), .A2(n21220), .B1(n21218), .B2(n20713), .ZN(
        n20710) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n21159), .ZN(n20709) );
  OAI211_X1 U23674 ( .C1(n20718), .C2(n21069), .A(n20710), .B(n20709), .ZN(
        P1_U3054) );
  INV_X1 U23675 ( .A(n21227), .ZN(n21074) );
  AOI22_X1 U23676 ( .A1(n20748), .A2(n21114), .B1(n21226), .B2(n20713), .ZN(
        n20712) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n21228), .ZN(n20711) );
  OAI211_X1 U23678 ( .C1(n20718), .C2(n21074), .A(n20712), .B(n20711), .ZN(
        P1_U3055) );
  INV_X1 U23679 ( .A(n21235), .ZN(n21082) );
  AOI22_X1 U23680 ( .A1(n20714), .A2(n21236), .B1(n21232), .B2(n20713), .ZN(
        n20717) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20715), .B1(
        n20748), .B2(n21120), .ZN(n20716) );
  OAI211_X1 U23682 ( .C1(n20718), .C2(n21082), .A(n20717), .B(n20716), .ZN(
        P1_U3056) );
  INV_X1 U23683 ( .A(n20719), .ZN(n20720) );
  OAI21_X1 U23684 ( .B1(n21184), .B2(n20727), .A(n20720), .ZN(n20730) );
  INV_X1 U23685 ( .A(n20721), .ZN(n20725) );
  INV_X1 U23686 ( .A(n20722), .ZN(n20723) );
  NAND2_X1 U23687 ( .A1(n20723), .A2(n10782), .ZN(n21171) );
  INV_X1 U23688 ( .A(n21171), .ZN(n20724) );
  NOR2_X1 U23689 ( .A1(n20995), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20747) );
  AOI21_X1 U23690 ( .B1(n20725), .B2(n20724), .A(n20747), .ZN(n20731) );
  INV_X1 U23691 ( .A(n20731), .ZN(n20726) );
  AOI22_X1 U23692 ( .A1(n20784), .A2(n21095), .B1(n21176), .B2(n20747), .ZN(
        n20734) );
  OAI21_X1 U23693 ( .B1(n21186), .B2(n20728), .A(n21182), .ZN(n20729) );
  AOI21_X1 U23694 ( .B1(n20731), .B2(n20730), .A(n20729), .ZN(n20732) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20749), .B1(
        n20748), .B2(n21187), .ZN(n20733) );
  OAI211_X1 U23696 ( .C1(n20752), .C2(n21046), .A(n20734), .B(n20733), .ZN(
        P1_U3057) );
  AOI22_X1 U23697 ( .A1(n20748), .A2(n21142), .B1(n21191), .B2(n20747), .ZN(
        n20736) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20749), .B1(
        n20784), .B2(n21193), .ZN(n20735) );
  OAI211_X1 U23699 ( .C1(n20752), .C2(n21051), .A(n20736), .B(n20735), .ZN(
        P1_U3058) );
  AOI22_X1 U23700 ( .A1(n20748), .A2(n21202), .B1(n20976), .B2(n20747), .ZN(
        n20738) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20749), .B1(
        n20784), .B2(n21104), .ZN(n20737) );
  OAI211_X1 U23702 ( .C1(n20752), .C2(n21200), .A(n20738), .B(n20737), .ZN(
        P1_U3059) );
  AOI22_X1 U23703 ( .A1(n20784), .A2(n21208), .B1(n21206), .B2(n20747), .ZN(
        n20740) );
  AOI22_X1 U23704 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20749), .B1(
        n20748), .B2(n21151), .ZN(n20739) );
  OAI211_X1 U23705 ( .C1(n20752), .C2(n21059), .A(n20740), .B(n20739), .ZN(
        P1_U3060) );
  AOI22_X1 U23706 ( .A1(n20748), .A2(n21155), .B1(n21212), .B2(n20747), .ZN(
        n20742) );
  AOI22_X1 U23707 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20749), .B1(
        n20784), .B2(n21214), .ZN(n20741) );
  OAI211_X1 U23708 ( .C1(n20752), .C2(n21064), .A(n20742), .B(n20741), .ZN(
        P1_U3061) );
  AOI22_X1 U23709 ( .A1(n20784), .A2(n21220), .B1(n21218), .B2(n20747), .ZN(
        n20744) );
  AOI22_X1 U23710 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20749), .B1(
        n20748), .B2(n21159), .ZN(n20743) );
  OAI211_X1 U23711 ( .C1(n20752), .C2(n21069), .A(n20744), .B(n20743), .ZN(
        P1_U3062) );
  AOI22_X1 U23712 ( .A1(n20748), .A2(n21228), .B1(n21226), .B2(n20747), .ZN(
        n20746) );
  AOI22_X1 U23713 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20749), .B1(
        n20784), .B2(n21114), .ZN(n20745) );
  OAI211_X1 U23714 ( .C1(n20752), .C2(n21074), .A(n20746), .B(n20745), .ZN(
        P1_U3063) );
  AOI22_X1 U23715 ( .A1(n20748), .A2(n21236), .B1(n21232), .B2(n20747), .ZN(
        n20751) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20749), .B1(
        n20784), .B2(n21120), .ZN(n20750) );
  OAI211_X1 U23717 ( .C1(n20752), .C2(n21082), .A(n20751), .B(n20750), .ZN(
        P1_U3064) );
  INV_X1 U23718 ( .A(n21095), .ZN(n21190) );
  NAND2_X1 U23719 ( .A1(n21031), .A2(n20754), .ZN(n20860) );
  NAND2_X1 U23720 ( .A1(n14172), .A2(n21186), .ZN(n20755) );
  OR2_X1 U23721 ( .A1(n20860), .A2(n20755), .ZN(n20758) );
  OR2_X1 U23722 ( .A1(n20821), .A2(n20756), .ZN(n20757) );
  NAND2_X1 U23723 ( .A1(n20758), .A2(n20757), .ZN(n20783) );
  NAND3_X1 U23724 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17071), .A3(
        n21033), .ZN(n20789) );
  NOR2_X1 U23725 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20789), .ZN(
        n20782) );
  AOI22_X1 U23726 ( .A1(n21177), .A2(n20783), .B1(n21176), .B2(n20782), .ZN(
        n20766) );
  INV_X1 U23727 ( .A(n20860), .ZN(n20761) );
  INV_X1 U23728 ( .A(n20784), .ZN(n20759) );
  AOI21_X1 U23729 ( .B1(n20759), .B2(n20818), .A(n20900), .ZN(n20760) );
  AOI21_X1 U23730 ( .B1(n20761), .B2(n14172), .A(n20760), .ZN(n20762) );
  NOR2_X1 U23731 ( .A1(n20762), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20764) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21187), .ZN(n20765) );
  OAI211_X1 U23733 ( .C1(n21190), .C2(n20818), .A(n20766), .B(n20765), .ZN(
        P1_U3065) );
  INV_X1 U23734 ( .A(n21193), .ZN(n21145) );
  AOI22_X1 U23735 ( .A1(n21192), .A2(n20783), .B1(n21191), .B2(n20782), .ZN(
        n20768) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21142), .ZN(n20767) );
  OAI211_X1 U23737 ( .C1(n21145), .C2(n20818), .A(n20768), .B(n20767), .ZN(
        P1_U3066) );
  INV_X1 U23738 ( .A(n20783), .ZN(n20770) );
  INV_X1 U23739 ( .A(n20782), .ZN(n20769) );
  OAI22_X1 U23740 ( .A1(n21200), .A2(n20770), .B1(n21197), .B2(n20769), .ZN(
        n20771) );
  INV_X1 U23741 ( .A(n20771), .ZN(n20773) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21202), .ZN(n20772) );
  OAI211_X1 U23743 ( .C1(n21205), .C2(n20818), .A(n20773), .B(n20772), .ZN(
        P1_U3067) );
  AOI22_X1 U23744 ( .A1(n21207), .A2(n20783), .B1(n21206), .B2(n20782), .ZN(
        n20775) );
  AOI22_X1 U23745 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21151), .ZN(n20774) );
  OAI211_X1 U23746 ( .C1(n21154), .C2(n20818), .A(n20775), .B(n20774), .ZN(
        P1_U3068) );
  AOI22_X1 U23747 ( .A1(n21213), .A2(n20783), .B1(n21212), .B2(n20782), .ZN(
        n20777) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21155), .ZN(n20776) );
  OAI211_X1 U23749 ( .C1(n21158), .C2(n20818), .A(n20777), .B(n20776), .ZN(
        P1_U3069) );
  AOI22_X1 U23750 ( .A1(n21219), .A2(n20783), .B1(n21218), .B2(n20782), .ZN(
        n20779) );
  AOI22_X1 U23751 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21159), .ZN(n20778) );
  OAI211_X1 U23752 ( .C1(n21162), .C2(n20818), .A(n20779), .B(n20778), .ZN(
        P1_U3070) );
  AOI22_X1 U23753 ( .A1(n21227), .A2(n20783), .B1(n21226), .B2(n20782), .ZN(
        n20781) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21228), .ZN(n20780) );
  OAI211_X1 U23755 ( .C1(n21231), .C2(n20818), .A(n20781), .B(n20780), .ZN(
        P1_U3071) );
  AOI22_X1 U23756 ( .A1(n21235), .A2(n20783), .B1(n21232), .B2(n20782), .ZN(
        n20787) );
  AOI22_X1 U23757 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20785), .B1(
        n20784), .B2(n21236), .ZN(n20786) );
  OAI211_X1 U23758 ( .C1(n21242), .C2(n20818), .A(n20787), .B(n20786), .ZN(
        P1_U3072) );
  OR2_X1 U23759 ( .A1(n20860), .A2(n20658), .ZN(n20788) );
  NOR2_X1 U23760 ( .A1(n21084), .A2(n20789), .ZN(n20813) );
  INV_X1 U23761 ( .A(n20813), .ZN(n20800) );
  NAND2_X1 U23762 ( .A1(n20788), .A2(n20800), .ZN(n20792) );
  NAND2_X1 U23763 ( .A1(n20792), .A2(n21186), .ZN(n20791) );
  INV_X1 U23764 ( .A(n20789), .ZN(n20795) );
  NAND2_X1 U23765 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20795), .ZN(n20790) );
  NAND2_X1 U23766 ( .A1(n20791), .A2(n20790), .ZN(n20814) );
  AOI22_X1 U23767 ( .A1(n21177), .A2(n20814), .B1(n21176), .B2(n20813), .ZN(
        n20797) );
  INV_X1 U23768 ( .A(n20792), .ZN(n20793) );
  OAI21_X1 U23769 ( .B1(n20866), .B2(n20900), .A(n20793), .ZN(n20794) );
  OAI221_X1 U23770 ( .B1(n21186), .B2(n20795), .C1(n21184), .C2(n20794), .A(
        n21182), .ZN(n20815) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21095), .ZN(n20796) );
  OAI211_X1 U23772 ( .C1(n21098), .C2(n20818), .A(n20797), .B(n20796), .ZN(
        P1_U3073) );
  AOI22_X1 U23773 ( .A1(n21192), .A2(n20814), .B1(n21191), .B2(n20813), .ZN(
        n20799) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21193), .ZN(n20798) );
  OAI211_X1 U23775 ( .C1(n21196), .C2(n20818), .A(n20799), .B(n20798), .ZN(
        P1_U3074) );
  INV_X1 U23776 ( .A(n20814), .ZN(n20801) );
  OAI22_X1 U23777 ( .A1(n21200), .A2(n20801), .B1(n21197), .B2(n20800), .ZN(
        n20802) );
  INV_X1 U23778 ( .A(n20802), .ZN(n20804) );
  AOI22_X1 U23779 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21104), .ZN(n20803) );
  OAI211_X1 U23780 ( .C1(n21107), .C2(n20818), .A(n20804), .B(n20803), .ZN(
        P1_U3075) );
  AOI22_X1 U23781 ( .A1(n21207), .A2(n20814), .B1(n21206), .B2(n20813), .ZN(
        n20806) );
  AOI22_X1 U23782 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21208), .ZN(n20805) );
  OAI211_X1 U23783 ( .C1(n21211), .C2(n20818), .A(n20806), .B(n20805), .ZN(
        P1_U3076) );
  AOI22_X1 U23784 ( .A1(n21213), .A2(n20814), .B1(n21212), .B2(n20813), .ZN(
        n20808) );
  AOI22_X1 U23785 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21214), .ZN(n20807) );
  OAI211_X1 U23786 ( .C1(n21217), .C2(n20818), .A(n20808), .B(n20807), .ZN(
        P1_U3077) );
  AOI22_X1 U23787 ( .A1(n21219), .A2(n20814), .B1(n21218), .B2(n20813), .ZN(
        n20810) );
  AOI22_X1 U23788 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21220), .ZN(n20809) );
  OAI211_X1 U23789 ( .C1(n21225), .C2(n20818), .A(n20810), .B(n20809), .ZN(
        P1_U3078) );
  AOI22_X1 U23790 ( .A1(n21227), .A2(n20814), .B1(n21226), .B2(n20813), .ZN(
        n20812) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21114), .ZN(n20811) );
  OAI211_X1 U23792 ( .C1(n21117), .C2(n20818), .A(n20812), .B(n20811), .ZN(
        P1_U3079) );
  AOI22_X1 U23793 ( .A1(n21235), .A2(n20814), .B1(n21232), .B2(n20813), .ZN(
        n20817) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20815), .B1(
        n20854), .B2(n21120), .ZN(n20816) );
  OAI211_X1 U23795 ( .C1(n21125), .C2(n20818), .A(n20817), .B(n20816), .ZN(
        P1_U3080) );
  NAND3_X1 U23796 ( .A1(n20852), .A2(n20844), .A3(n21186), .ZN(n20820) );
  NAND2_X1 U23797 ( .A1(n20820), .A2(n20819), .ZN(n20827) );
  NOR2_X1 U23798 ( .A1(n20860), .A2(n14172), .ZN(n20824) );
  INV_X1 U23799 ( .A(n20821), .ZN(n21129) );
  INV_X1 U23800 ( .A(n20869), .ZN(n20822) );
  NOR2_X1 U23801 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20822), .ZN(
        n20829) );
  INV_X1 U23802 ( .A(n20829), .ZN(n20851) );
  OAI22_X1 U23803 ( .A1(n20852), .A2(n21190), .B1(n21034), .B2(n20851), .ZN(
        n20823) );
  INV_X1 U23804 ( .A(n20823), .ZN(n20831) );
  INV_X1 U23805 ( .A(n20824), .ZN(n20826) );
  AOI21_X1 U23806 ( .B1(n20827), .B2(n20826), .A(n20825), .ZN(n20828) );
  OAI211_X1 U23807 ( .C1(n20829), .C2(n21041), .A(n21138), .B(n20828), .ZN(
        n20855) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n21187), .ZN(n20830) );
  OAI211_X1 U23809 ( .C1(n20858), .C2(n21046), .A(n20831), .B(n20830), .ZN(
        P1_U3081) );
  OAI22_X1 U23810 ( .A1(n20852), .A2(n21145), .B1(n21047), .B2(n20851), .ZN(
        n20832) );
  INV_X1 U23811 ( .A(n20832), .ZN(n20834) );
  AOI22_X1 U23812 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n21142), .ZN(n20833) );
  OAI211_X1 U23813 ( .C1(n20858), .C2(n21051), .A(n20834), .B(n20833), .ZN(
        P1_U3082) );
  OAI22_X1 U23814 ( .A1(n20852), .A2(n21205), .B1(n21197), .B2(n20851), .ZN(
        n20835) );
  INV_X1 U23815 ( .A(n20835), .ZN(n20837) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n21202), .ZN(n20836) );
  OAI211_X1 U23817 ( .C1(n20858), .C2(n21200), .A(n20837), .B(n20836), .ZN(
        P1_U3083) );
  OAI22_X1 U23818 ( .A1(n20844), .A2(n21211), .B1(n21055), .B2(n20851), .ZN(
        n20838) );
  INV_X1 U23819 ( .A(n20838), .ZN(n20840) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20855), .B1(
        n20889), .B2(n21208), .ZN(n20839) );
  OAI211_X1 U23821 ( .C1(n20858), .C2(n21059), .A(n20840), .B(n20839), .ZN(
        P1_U3084) );
  OAI22_X1 U23822 ( .A1(n20852), .A2(n21158), .B1(n21060), .B2(n20851), .ZN(
        n20841) );
  INV_X1 U23823 ( .A(n20841), .ZN(n20843) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n21155), .ZN(n20842) );
  OAI211_X1 U23825 ( .C1(n20858), .C2(n21064), .A(n20843), .B(n20842), .ZN(
        P1_U3085) );
  OAI22_X1 U23826 ( .A1(n20844), .A2(n21225), .B1(n21065), .B2(n20851), .ZN(
        n20845) );
  INV_X1 U23827 ( .A(n20845), .ZN(n20847) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20855), .B1(
        n20889), .B2(n21220), .ZN(n20846) );
  OAI211_X1 U23829 ( .C1(n20858), .C2(n21069), .A(n20847), .B(n20846), .ZN(
        P1_U3086) );
  OAI22_X1 U23830 ( .A1(n20852), .A2(n21231), .B1(n21070), .B2(n20851), .ZN(
        n20848) );
  INV_X1 U23831 ( .A(n20848), .ZN(n20850) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n21228), .ZN(n20849) );
  OAI211_X1 U23833 ( .C1(n20858), .C2(n21074), .A(n20850), .B(n20849), .ZN(
        P1_U3087) );
  OAI22_X1 U23834 ( .A1(n20852), .A2(n21242), .B1(n21076), .B2(n20851), .ZN(
        n20853) );
  INV_X1 U23835 ( .A(n20853), .ZN(n20857) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n21236), .ZN(n20856) );
  OAI211_X1 U23837 ( .C1(n20858), .C2(n21082), .A(n20857), .B(n20856), .ZN(
        P1_U3088) );
  INV_X1 U23838 ( .A(n20993), .ZN(n20859) );
  OR2_X1 U23839 ( .A1(n20860), .A2(n21171), .ZN(n20861) );
  NAND2_X1 U23840 ( .A1(n20861), .A2(n20874), .ZN(n20864) );
  NAND2_X1 U23841 ( .A1(n20864), .A2(n21186), .ZN(n20863) );
  NAND2_X1 U23842 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20869), .ZN(n20862) );
  NAND2_X1 U23843 ( .A1(n20863), .A2(n20862), .ZN(n20888) );
  INV_X1 U23844 ( .A(n20874), .ZN(n20887) );
  AOI22_X1 U23845 ( .A1(n21177), .A2(n20888), .B1(n20887), .B2(n21176), .ZN(
        n20871) );
  INV_X1 U23846 ( .A(n21179), .ZN(n20867) );
  INV_X1 U23847 ( .A(n20864), .ZN(n20865) );
  OAI21_X1 U23848 ( .B1(n20867), .B2(n20866), .A(n20865), .ZN(n20868) );
  OAI221_X1 U23849 ( .B1(n21186), .B2(n20869), .C1(n21184), .C2(n20868), .A(
        n21182), .ZN(n20890) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21187), .ZN(n20870) );
  OAI211_X1 U23851 ( .C1(n21190), .C2(n20904), .A(n20871), .B(n20870), .ZN(
        P1_U3089) );
  AOI22_X1 U23852 ( .A1(n21192), .A2(n20888), .B1(n20887), .B2(n21191), .ZN(
        n20873) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21142), .ZN(n20872) );
  OAI211_X1 U23854 ( .C1(n21145), .C2(n20904), .A(n20873), .B(n20872), .ZN(
        P1_U3090) );
  INV_X1 U23855 ( .A(n20888), .ZN(n20875) );
  OAI22_X1 U23856 ( .A1(n21200), .A2(n20875), .B1(n20874), .B2(n21197), .ZN(
        n20876) );
  INV_X1 U23857 ( .A(n20876), .ZN(n20878) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21202), .ZN(n20877) );
  OAI211_X1 U23859 ( .C1(n21205), .C2(n20904), .A(n20878), .B(n20877), .ZN(
        P1_U3091) );
  AOI22_X1 U23860 ( .A1(n21207), .A2(n20888), .B1(n20887), .B2(n21206), .ZN(
        n20880) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21151), .ZN(n20879) );
  OAI211_X1 U23862 ( .C1(n21154), .C2(n20904), .A(n20880), .B(n20879), .ZN(
        P1_U3092) );
  AOI22_X1 U23863 ( .A1(n21213), .A2(n20888), .B1(n20887), .B2(n21212), .ZN(
        n20882) );
  AOI22_X1 U23864 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21155), .ZN(n20881) );
  OAI211_X1 U23865 ( .C1(n21158), .C2(n20904), .A(n20882), .B(n20881), .ZN(
        P1_U3093) );
  AOI22_X1 U23866 ( .A1(n21219), .A2(n20888), .B1(n20887), .B2(n21218), .ZN(
        n20884) );
  AOI22_X1 U23867 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21159), .ZN(n20883) );
  OAI211_X1 U23868 ( .C1(n21162), .C2(n20904), .A(n20884), .B(n20883), .ZN(
        P1_U3094) );
  AOI22_X1 U23869 ( .A1(n21227), .A2(n20888), .B1(n20887), .B2(n21226), .ZN(
        n20886) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21228), .ZN(n20885) );
  OAI211_X1 U23871 ( .C1(n21231), .C2(n20904), .A(n20886), .B(n20885), .ZN(
        P1_U3095) );
  AOI22_X1 U23872 ( .A1(n21235), .A2(n20888), .B1(n20887), .B2(n21232), .ZN(
        n20892) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20890), .B1(
        n20889), .B2(n21236), .ZN(n20891) );
  OAI211_X1 U23874 ( .C1(n21242), .C2(n20904), .A(n20892), .B(n20891), .ZN(
        P1_U3096) );
  NAND2_X1 U23875 ( .A1(n20894), .A2(n20893), .ZN(n20997) );
  OR2_X1 U23876 ( .A1(n20997), .A2(n21133), .ZN(n20895) );
  NAND3_X1 U23877 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10743), .A3(
        n21033), .ZN(n20929) );
  NOR2_X1 U23878 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20929), .ZN(
        n20922) );
  INV_X1 U23879 ( .A(n20922), .ZN(n20909) );
  NAND2_X1 U23880 ( .A1(n20895), .A2(n20909), .ZN(n20901) );
  NAND2_X1 U23881 ( .A1(n20901), .A2(n21186), .ZN(n20899) );
  INV_X1 U23882 ( .A(n20896), .ZN(n20897) );
  AND2_X1 U23883 ( .A1(n20897), .A2(n20963), .ZN(n21036) );
  NAND2_X1 U23884 ( .A1(n20964), .A2(n21036), .ZN(n20898) );
  NAND2_X1 U23885 ( .A1(n20899), .A2(n20898), .ZN(n20923) );
  AOI22_X1 U23886 ( .A1(n21177), .A2(n20923), .B1(n21176), .B2(n20922), .ZN(
        n20906) );
  AOI21_X1 U23887 ( .B1(n20959), .B2(n20904), .A(n20900), .ZN(n20902) );
  AOI22_X1 U23888 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21187), .ZN(n20905) );
  OAI211_X1 U23889 ( .C1(n21190), .C2(n20959), .A(n20906), .B(n20905), .ZN(
        P1_U3097) );
  AOI22_X1 U23890 ( .A1(n21192), .A2(n20923), .B1(n21191), .B2(n20922), .ZN(
        n20908) );
  AOI22_X1 U23891 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21142), .ZN(n20907) );
  OAI211_X1 U23892 ( .C1(n21145), .C2(n20959), .A(n20908), .B(n20907), .ZN(
        P1_U3098) );
  INV_X1 U23893 ( .A(n20923), .ZN(n20910) );
  OAI22_X1 U23894 ( .A1(n21200), .A2(n20910), .B1(n21197), .B2(n20909), .ZN(
        n20911) );
  INV_X1 U23895 ( .A(n20911), .ZN(n20913) );
  AOI22_X1 U23896 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21202), .ZN(n20912) );
  OAI211_X1 U23897 ( .C1(n21205), .C2(n20959), .A(n20913), .B(n20912), .ZN(
        P1_U3099) );
  AOI22_X1 U23898 ( .A1(n21207), .A2(n20923), .B1(n21206), .B2(n20922), .ZN(
        n20915) );
  AOI22_X1 U23899 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21151), .ZN(n20914) );
  OAI211_X1 U23900 ( .C1(n21154), .C2(n20959), .A(n20915), .B(n20914), .ZN(
        P1_U3100) );
  AOI22_X1 U23901 ( .A1(n21213), .A2(n20923), .B1(n21212), .B2(n20922), .ZN(
        n20917) );
  AOI22_X1 U23902 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21155), .ZN(n20916) );
  OAI211_X1 U23903 ( .C1(n21158), .C2(n20959), .A(n20917), .B(n20916), .ZN(
        P1_U3101) );
  AOI22_X1 U23904 ( .A1(n21219), .A2(n20923), .B1(n21218), .B2(n20922), .ZN(
        n20919) );
  AOI22_X1 U23905 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21159), .ZN(n20918) );
  OAI211_X1 U23906 ( .C1(n21162), .C2(n20959), .A(n20919), .B(n20918), .ZN(
        P1_U3102) );
  AOI22_X1 U23907 ( .A1(n21227), .A2(n20923), .B1(n21226), .B2(n20922), .ZN(
        n20921) );
  AOI22_X1 U23908 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21228), .ZN(n20920) );
  OAI211_X1 U23909 ( .C1(n21231), .C2(n20959), .A(n20921), .B(n20920), .ZN(
        P1_U3103) );
  AOI22_X1 U23910 ( .A1(n21235), .A2(n20923), .B1(n21232), .B2(n20922), .ZN(
        n20927) );
  AOI22_X1 U23911 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20925), .B1(
        n20924), .B2(n21236), .ZN(n20926) );
  OAI211_X1 U23912 ( .C1(n21242), .C2(n20959), .A(n20927), .B(n20926), .ZN(
        P1_U3104) );
  NOR2_X1 U23913 ( .A1(n21084), .A2(n20929), .ZN(n20954) );
  INV_X1 U23914 ( .A(n20954), .ZN(n20941) );
  OAI21_X1 U23915 ( .B1(n20997), .B2(n20658), .A(n20941), .ZN(n20928) );
  NAND2_X1 U23916 ( .A1(n20928), .A2(n21186), .ZN(n20931) );
  INV_X1 U23917 ( .A(n20929), .ZN(n20935) );
  NAND2_X1 U23918 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20935), .ZN(n20930) );
  NAND2_X1 U23919 ( .A1(n20931), .A2(n20930), .ZN(n20955) );
  AOI22_X1 U23920 ( .A1(n21177), .A2(n20955), .B1(n21176), .B2(n20954), .ZN(
        n20938) );
  NOR2_X1 U23921 ( .A1(n20933), .A2(n20932), .ZN(n20934) );
  AOI22_X1 U23922 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21095), .ZN(n20937) );
  OAI211_X1 U23923 ( .C1(n21098), .C2(n20959), .A(n20938), .B(n20937), .ZN(
        P1_U3105) );
  AOI22_X1 U23924 ( .A1(n21192), .A2(n20955), .B1(n21191), .B2(n20954), .ZN(
        n20940) );
  AOI22_X1 U23925 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21193), .ZN(n20939) );
  OAI211_X1 U23926 ( .C1(n21196), .C2(n20959), .A(n20940), .B(n20939), .ZN(
        P1_U3106) );
  INV_X1 U23927 ( .A(n20955), .ZN(n20942) );
  OAI22_X1 U23928 ( .A1(n21200), .A2(n20942), .B1(n21197), .B2(n20941), .ZN(
        n20943) );
  INV_X1 U23929 ( .A(n20943), .ZN(n20945) );
  AOI22_X1 U23930 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21104), .ZN(n20944) );
  OAI211_X1 U23931 ( .C1(n21107), .C2(n20959), .A(n20945), .B(n20944), .ZN(
        P1_U3107) );
  AOI22_X1 U23932 ( .A1(n21207), .A2(n20955), .B1(n21206), .B2(n20954), .ZN(
        n20947) );
  AOI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21208), .ZN(n20946) );
  OAI211_X1 U23934 ( .C1(n21211), .C2(n20959), .A(n20947), .B(n20946), .ZN(
        P1_U3108) );
  AOI22_X1 U23935 ( .A1(n21213), .A2(n20955), .B1(n21212), .B2(n20954), .ZN(
        n20949) );
  AOI22_X1 U23936 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21214), .ZN(n20948) );
  OAI211_X1 U23937 ( .C1(n21217), .C2(n20959), .A(n20949), .B(n20948), .ZN(
        P1_U3109) );
  AOI22_X1 U23938 ( .A1(n21219), .A2(n20955), .B1(n21218), .B2(n20954), .ZN(
        n20951) );
  AOI22_X1 U23939 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21220), .ZN(n20950) );
  OAI211_X1 U23940 ( .C1(n21225), .C2(n20959), .A(n20951), .B(n20950), .ZN(
        P1_U3110) );
  AOI22_X1 U23941 ( .A1(n21227), .A2(n20955), .B1(n21226), .B2(n20954), .ZN(
        n20953) );
  AOI22_X1 U23942 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21114), .ZN(n20952) );
  OAI211_X1 U23943 ( .C1(n21117), .C2(n20959), .A(n20953), .B(n20952), .ZN(
        P1_U3111) );
  AOI22_X1 U23944 ( .A1(n21235), .A2(n20955), .B1(n21232), .B2(n20954), .ZN(
        n20958) );
  AOI22_X1 U23945 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20956), .B1(
        n20988), .B2(n21120), .ZN(n20957) );
  OAI211_X1 U23946 ( .C1(n21125), .C2(n20959), .A(n20958), .B(n20957), .ZN(
        P1_U3112) );
  NOR3_X1 U23947 ( .A1(n21025), .A2(n20988), .A3(n21184), .ZN(n20962) );
  NOR2_X1 U23948 ( .A1(n20962), .A2(n20961), .ZN(n20971) );
  INV_X1 U23949 ( .A(n20971), .ZN(n20965) );
  NOR2_X1 U23950 ( .A1(n20997), .A2(n14172), .ZN(n20970) );
  OR2_X1 U23951 ( .A1(n20963), .A2(n17071), .ZN(n20966) );
  INV_X1 U23952 ( .A(n20966), .ZN(n21128) );
  NAND3_X1 U23953 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n10743), .ZN(n21002) );
  NOR2_X1 U23954 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21002), .ZN(
        n20987) );
  AOI22_X1 U23955 ( .A1(n20988), .A2(n21187), .B1(n21176), .B2(n20987), .ZN(
        n20973) );
  NAND2_X1 U23956 ( .A1(n20966), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21137) );
  OAI211_X1 U23957 ( .C1(n21041), .C2(n20987), .A(n21137), .B(n20967), .ZN(
        n20968) );
  INV_X1 U23958 ( .A(n20968), .ZN(n20969) );
  AOI22_X1 U23959 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20989), .B1(
        n21025), .B2(n21095), .ZN(n20972) );
  OAI211_X1 U23960 ( .C1(n20992), .C2(n21046), .A(n20973), .B(n20972), .ZN(
        P1_U3113) );
  AOI22_X1 U23961 ( .A1(n21025), .A2(n21193), .B1(n21191), .B2(n20987), .ZN(
        n20975) );
  AOI22_X1 U23962 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20989), .B1(
        n20988), .B2(n21142), .ZN(n20974) );
  OAI211_X1 U23963 ( .C1(n20992), .C2(n21051), .A(n20975), .B(n20974), .ZN(
        P1_U3114) );
  AOI22_X1 U23964 ( .A1(n21025), .A2(n21104), .B1(n20976), .B2(n20987), .ZN(
        n20978) );
  AOI22_X1 U23965 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20989), .B1(
        n20988), .B2(n21202), .ZN(n20977) );
  OAI211_X1 U23966 ( .C1(n20992), .C2(n21200), .A(n20978), .B(n20977), .ZN(
        P1_U3115) );
  AOI22_X1 U23967 ( .A1(n20988), .A2(n21151), .B1(n21206), .B2(n20987), .ZN(
        n20980) );
  AOI22_X1 U23968 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20989), .B1(
        n21025), .B2(n21208), .ZN(n20979) );
  OAI211_X1 U23969 ( .C1(n20992), .C2(n21059), .A(n20980), .B(n20979), .ZN(
        P1_U3116) );
  AOI22_X1 U23970 ( .A1(n21025), .A2(n21214), .B1(n21212), .B2(n20987), .ZN(
        n20982) );
  AOI22_X1 U23971 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20989), .B1(
        n20988), .B2(n21155), .ZN(n20981) );
  OAI211_X1 U23972 ( .C1(n20992), .C2(n21064), .A(n20982), .B(n20981), .ZN(
        P1_U3117) );
  AOI22_X1 U23973 ( .A1(n20988), .A2(n21159), .B1(n21218), .B2(n20987), .ZN(
        n20984) );
  AOI22_X1 U23974 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20989), .B1(
        n21025), .B2(n21220), .ZN(n20983) );
  OAI211_X1 U23975 ( .C1(n20992), .C2(n21069), .A(n20984), .B(n20983), .ZN(
        P1_U3118) );
  AOI22_X1 U23976 ( .A1(n20988), .A2(n21228), .B1(n21226), .B2(n20987), .ZN(
        n20986) );
  AOI22_X1 U23977 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20989), .B1(
        n21025), .B2(n21114), .ZN(n20985) );
  OAI211_X1 U23978 ( .C1(n20992), .C2(n21074), .A(n20986), .B(n20985), .ZN(
        P1_U3119) );
  AOI22_X1 U23979 ( .A1(n21025), .A2(n21120), .B1(n21232), .B2(n20987), .ZN(
        n20991) );
  AOI22_X1 U23980 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20989), .B1(
        n20988), .B2(n21236), .ZN(n20990) );
  OAI211_X1 U23981 ( .C1(n20992), .C2(n21082), .A(n20991), .B(n20990), .ZN(
        P1_U3120) );
  INV_X1 U23982 ( .A(n20995), .ZN(n20996) );
  NAND2_X1 U23983 ( .A1(n20996), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21010) );
  OAI21_X1 U23984 ( .B1(n20997), .B2(n21171), .A(n21010), .ZN(n20998) );
  NAND2_X1 U23985 ( .A1(n20998), .A2(n21186), .ZN(n21001) );
  INV_X1 U23986 ( .A(n21002), .ZN(n20999) );
  NAND2_X1 U23987 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20999), .ZN(n21000) );
  NAND2_X1 U23988 ( .A1(n21001), .A2(n21000), .ZN(n21024) );
  INV_X1 U23989 ( .A(n21010), .ZN(n21023) );
  AOI22_X1 U23990 ( .A1(n21177), .A2(n21024), .B1(n21176), .B2(n21023), .ZN(
        n21007) );
  OAI21_X1 U23991 ( .B1(n21004), .B2(n21003), .A(n21002), .ZN(n21005) );
  NAND2_X1 U23992 ( .A1(n21005), .A2(n21182), .ZN(n21026) );
  AOI22_X1 U23993 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21187), .ZN(n21006) );
  OAI211_X1 U23994 ( .C1(n21190), .C2(n21043), .A(n21007), .B(n21006), .ZN(
        P1_U3121) );
  AOI22_X1 U23995 ( .A1(n21192), .A2(n21024), .B1(n21191), .B2(n21023), .ZN(
        n21009) );
  AOI22_X1 U23996 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21142), .ZN(n21008) );
  OAI211_X1 U23997 ( .C1(n21145), .C2(n21043), .A(n21009), .B(n21008), .ZN(
        P1_U3122) );
  INV_X1 U23998 ( .A(n21024), .ZN(n21011) );
  OAI22_X1 U23999 ( .A1(n21200), .A2(n21011), .B1(n21197), .B2(n21010), .ZN(
        n21012) );
  INV_X1 U24000 ( .A(n21012), .ZN(n21014) );
  AOI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21202), .ZN(n21013) );
  OAI211_X1 U24002 ( .C1(n21205), .C2(n21043), .A(n21014), .B(n21013), .ZN(
        P1_U3123) );
  AOI22_X1 U24003 ( .A1(n21207), .A2(n21024), .B1(n21206), .B2(n21023), .ZN(
        n21016) );
  AOI22_X1 U24004 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21151), .ZN(n21015) );
  OAI211_X1 U24005 ( .C1(n21154), .C2(n21043), .A(n21016), .B(n21015), .ZN(
        P1_U3124) );
  AOI22_X1 U24006 ( .A1(n21213), .A2(n21024), .B1(n21212), .B2(n21023), .ZN(
        n21018) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21155), .ZN(n21017) );
  OAI211_X1 U24008 ( .C1(n21158), .C2(n21043), .A(n21018), .B(n21017), .ZN(
        P1_U3125) );
  AOI22_X1 U24009 ( .A1(n21219), .A2(n21024), .B1(n21218), .B2(n21023), .ZN(
        n21020) );
  AOI22_X1 U24010 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21159), .ZN(n21019) );
  OAI211_X1 U24011 ( .C1(n21162), .C2(n21043), .A(n21020), .B(n21019), .ZN(
        P1_U3126) );
  AOI22_X1 U24012 ( .A1(n21227), .A2(n21024), .B1(n21226), .B2(n21023), .ZN(
        n21022) );
  AOI22_X1 U24013 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21228), .ZN(n21021) );
  OAI211_X1 U24014 ( .C1(n21231), .C2(n21043), .A(n21022), .B(n21021), .ZN(
        P1_U3127) );
  AOI22_X1 U24015 ( .A1(n21235), .A2(n21024), .B1(n21232), .B2(n21023), .ZN(
        n21028) );
  AOI22_X1 U24016 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21026), .B1(
        n21025), .B2(n21236), .ZN(n21027) );
  OAI211_X1 U24017 ( .C1(n21242), .C2(n21043), .A(n21028), .B(n21027), .ZN(
        P1_U3128) );
  NAND2_X1 U24018 ( .A1(n21043), .A2(n21124), .ZN(n21029) );
  AOI21_X1 U24019 ( .B1(n21029), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21184), 
        .ZN(n21039) );
  NAND2_X1 U24020 ( .A1(n21031), .A2(n21030), .ZN(n21172) );
  OR2_X1 U24021 ( .A1(n21172), .A2(n21133), .ZN(n21038) );
  INV_X1 U24022 ( .A(n21038), .ZN(n21032) );
  NAND3_X1 U24023 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21033), .ZN(n21090) );
  NOR2_X1 U24024 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21090), .ZN(
        n21042) );
  INV_X1 U24025 ( .A(n21042), .ZN(n21075) );
  OAI22_X1 U24026 ( .A1(n21124), .A2(n21190), .B1(n21034), .B2(n21075), .ZN(
        n21035) );
  INV_X1 U24027 ( .A(n21035), .ZN(n21045) );
  NOR2_X1 U24028 ( .A1(n21036), .A2(n21246), .ZN(n21037) );
  AOI21_X1 U24029 ( .B1(n21039), .B2(n21038), .A(n21037), .ZN(n21040) );
  AOI22_X1 U24030 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21187), .ZN(n21044) );
  OAI211_X1 U24031 ( .C1(n21083), .C2(n21046), .A(n21045), .B(n21044), .ZN(
        P1_U3129) );
  OAI22_X1 U24032 ( .A1(n21124), .A2(n21145), .B1(n21047), .B2(n21075), .ZN(
        n21048) );
  INV_X1 U24033 ( .A(n21048), .ZN(n21050) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21142), .ZN(n21049) );
  OAI211_X1 U24035 ( .C1(n21083), .C2(n21051), .A(n21050), .B(n21049), .ZN(
        P1_U3130) );
  OAI22_X1 U24036 ( .A1(n21124), .A2(n21205), .B1(n21197), .B2(n21075), .ZN(
        n21052) );
  INV_X1 U24037 ( .A(n21052), .ZN(n21054) );
  AOI22_X1 U24038 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21202), .ZN(n21053) );
  OAI211_X1 U24039 ( .C1(n21083), .C2(n21200), .A(n21054), .B(n21053), .ZN(
        P1_U3131) );
  OAI22_X1 U24040 ( .A1(n21124), .A2(n21154), .B1(n21055), .B2(n21075), .ZN(
        n21056) );
  INV_X1 U24041 ( .A(n21056), .ZN(n21058) );
  AOI22_X1 U24042 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21151), .ZN(n21057) );
  OAI211_X1 U24043 ( .C1(n21083), .C2(n21059), .A(n21058), .B(n21057), .ZN(
        P1_U3132) );
  OAI22_X1 U24044 ( .A1(n21124), .A2(n21158), .B1(n21060), .B2(n21075), .ZN(
        n21061) );
  INV_X1 U24045 ( .A(n21061), .ZN(n21063) );
  AOI22_X1 U24046 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21155), .ZN(n21062) );
  OAI211_X1 U24047 ( .C1(n21083), .C2(n21064), .A(n21063), .B(n21062), .ZN(
        P1_U3133) );
  OAI22_X1 U24048 ( .A1(n21124), .A2(n21162), .B1(n21065), .B2(n21075), .ZN(
        n21066) );
  INV_X1 U24049 ( .A(n21066), .ZN(n21068) );
  AOI22_X1 U24050 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21159), .ZN(n21067) );
  OAI211_X1 U24051 ( .C1(n21083), .C2(n21069), .A(n21068), .B(n21067), .ZN(
        P1_U3134) );
  OAI22_X1 U24052 ( .A1(n21124), .A2(n21231), .B1(n21070), .B2(n21075), .ZN(
        n21071) );
  INV_X1 U24053 ( .A(n21071), .ZN(n21073) );
  AOI22_X1 U24054 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21228), .ZN(n21072) );
  OAI211_X1 U24055 ( .C1(n21083), .C2(n21074), .A(n21073), .B(n21072), .ZN(
        P1_U3135) );
  OAI22_X1 U24056 ( .A1(n21124), .A2(n21242), .B1(n21076), .B2(n21075), .ZN(
        n21077) );
  INV_X1 U24057 ( .A(n21077), .ZN(n21081) );
  AOI22_X1 U24058 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21079), .B1(
        n21078), .B2(n21236), .ZN(n21080) );
  OAI211_X1 U24059 ( .C1(n21083), .C2(n21082), .A(n21081), .B(n21080), .ZN(
        P1_U3136) );
  NOR2_X1 U24060 ( .A1(n21084), .A2(n21090), .ZN(n21118) );
  INV_X1 U24061 ( .A(n21118), .ZN(n21101) );
  OAI21_X1 U24062 ( .B1(n21172), .B2(n20658), .A(n21101), .ZN(n21085) );
  NAND2_X1 U24063 ( .A1(n21085), .A2(n21186), .ZN(n21088) );
  INV_X1 U24064 ( .A(n21090), .ZN(n21086) );
  NAND2_X1 U24065 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21086), .ZN(n21087) );
  NAND2_X1 U24066 ( .A1(n21088), .A2(n21087), .ZN(n21119) );
  AOI22_X1 U24067 ( .A1(n21177), .A2(n21119), .B1(n21176), .B2(n21118), .ZN(
        n21097) );
  OAI21_X1 U24068 ( .B1(n21094), .B2(n21091), .A(n21090), .ZN(n21092) );
  NAND2_X1 U24069 ( .A1(n21092), .A2(n21182), .ZN(n21121) );
  AOI22_X1 U24070 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21095), .ZN(n21096) );
  OAI211_X1 U24071 ( .C1(n21098), .C2(n21124), .A(n21097), .B(n21096), .ZN(
        P1_U3137) );
  AOI22_X1 U24072 ( .A1(n21192), .A2(n21119), .B1(n21191), .B2(n21118), .ZN(
        n21100) );
  AOI22_X1 U24073 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21193), .ZN(n21099) );
  OAI211_X1 U24074 ( .C1(n21196), .C2(n21124), .A(n21100), .B(n21099), .ZN(
        P1_U3138) );
  INV_X1 U24075 ( .A(n21119), .ZN(n21102) );
  OAI22_X1 U24076 ( .A1(n21200), .A2(n21102), .B1(n21197), .B2(n21101), .ZN(
        n21103) );
  INV_X1 U24077 ( .A(n21103), .ZN(n21106) );
  AOI22_X1 U24078 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21104), .ZN(n21105) );
  OAI211_X1 U24079 ( .C1(n21107), .C2(n21124), .A(n21106), .B(n21105), .ZN(
        P1_U3139) );
  AOI22_X1 U24080 ( .A1(n21207), .A2(n21119), .B1(n21206), .B2(n21118), .ZN(
        n21109) );
  AOI22_X1 U24081 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21208), .ZN(n21108) );
  OAI211_X1 U24082 ( .C1(n21211), .C2(n21124), .A(n21109), .B(n21108), .ZN(
        P1_U3140) );
  AOI22_X1 U24083 ( .A1(n21213), .A2(n21119), .B1(n21212), .B2(n21118), .ZN(
        n21111) );
  AOI22_X1 U24084 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21214), .ZN(n21110) );
  OAI211_X1 U24085 ( .C1(n21217), .C2(n21124), .A(n21111), .B(n21110), .ZN(
        P1_U3141) );
  AOI22_X1 U24086 ( .A1(n21219), .A2(n21119), .B1(n21218), .B2(n21118), .ZN(
        n21113) );
  AOI22_X1 U24087 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21220), .ZN(n21112) );
  OAI211_X1 U24088 ( .C1(n21225), .C2(n21124), .A(n21113), .B(n21112), .ZN(
        P1_U3142) );
  AOI22_X1 U24089 ( .A1(n21227), .A2(n21119), .B1(n21226), .B2(n21118), .ZN(
        n21116) );
  AOI22_X1 U24090 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21114), .ZN(n21115) );
  OAI211_X1 U24091 ( .C1(n21117), .C2(n21124), .A(n21116), .B(n21115), .ZN(
        P1_U3143) );
  AOI22_X1 U24092 ( .A1(n21235), .A2(n21119), .B1(n21232), .B2(n21118), .ZN(
        n21123) );
  AOI22_X1 U24093 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21121), .B1(
        n21167), .B2(n21120), .ZN(n21122) );
  OAI211_X1 U24094 ( .C1(n21125), .C2(n21124), .A(n21123), .B(n21122), .ZN(
        P1_U3144) );
  NAND2_X1 U24095 ( .A1(n21133), .A2(n21186), .ZN(n21127) );
  OR2_X1 U24096 ( .A1(n21172), .A2(n21127), .ZN(n21131) );
  NAND2_X1 U24097 ( .A1(n21129), .A2(n21128), .ZN(n21130) );
  NAND2_X1 U24098 ( .A1(n21131), .A2(n21130), .ZN(n21166) );
  NOR2_X1 U24099 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21132), .ZN(
        n21165) );
  AOI22_X1 U24100 ( .A1(n21177), .A2(n21166), .B1(n21176), .B2(n21165), .ZN(
        n21141) );
  OAI21_X1 U24101 ( .B1(n21167), .B2(n21237), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21136) );
  INV_X1 U24102 ( .A(n21172), .ZN(n21134) );
  NAND2_X1 U24103 ( .A1(n21134), .A2(n21133), .ZN(n21135) );
  AOI21_X1 U24104 ( .B1(n21136), .B2(n21135), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21139) );
  AOI22_X1 U24105 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21187), .ZN(n21140) );
  OAI211_X1 U24106 ( .C1(n21190), .C2(n21224), .A(n21141), .B(n21140), .ZN(
        P1_U3145) );
  AOI22_X1 U24107 ( .A1(n21192), .A2(n21166), .B1(n21191), .B2(n21165), .ZN(
        n21144) );
  AOI22_X1 U24108 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21142), .ZN(n21143) );
  OAI211_X1 U24109 ( .C1(n21145), .C2(n21224), .A(n21144), .B(n21143), .ZN(
        P1_U3146) );
  INV_X1 U24110 ( .A(n21166), .ZN(n21147) );
  INV_X1 U24111 ( .A(n21165), .ZN(n21146) );
  OAI22_X1 U24112 ( .A1(n21200), .A2(n21147), .B1(n21197), .B2(n21146), .ZN(
        n21148) );
  INV_X1 U24113 ( .A(n21148), .ZN(n21150) );
  AOI22_X1 U24114 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21202), .ZN(n21149) );
  OAI211_X1 U24115 ( .C1(n21205), .C2(n21224), .A(n21150), .B(n21149), .ZN(
        P1_U3147) );
  AOI22_X1 U24116 ( .A1(n21207), .A2(n21166), .B1(n21206), .B2(n21165), .ZN(
        n21153) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21151), .ZN(n21152) );
  OAI211_X1 U24118 ( .C1(n21154), .C2(n21224), .A(n21153), .B(n21152), .ZN(
        P1_U3148) );
  AOI22_X1 U24119 ( .A1(n21213), .A2(n21166), .B1(n21212), .B2(n21165), .ZN(
        n21157) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21155), .ZN(n21156) );
  OAI211_X1 U24121 ( .C1(n21158), .C2(n21224), .A(n21157), .B(n21156), .ZN(
        P1_U3149) );
  AOI22_X1 U24122 ( .A1(n21219), .A2(n21166), .B1(n21218), .B2(n21165), .ZN(
        n21161) );
  AOI22_X1 U24123 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21159), .ZN(n21160) );
  OAI211_X1 U24124 ( .C1(n21162), .C2(n21224), .A(n21161), .B(n21160), .ZN(
        P1_U3150) );
  AOI22_X1 U24125 ( .A1(n21227), .A2(n21166), .B1(n21226), .B2(n21165), .ZN(
        n21164) );
  AOI22_X1 U24126 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21228), .ZN(n21163) );
  OAI211_X1 U24127 ( .C1(n21231), .C2(n21224), .A(n21164), .B(n21163), .ZN(
        P1_U3151) );
  AOI22_X1 U24128 ( .A1(n21235), .A2(n21166), .B1(n21232), .B2(n21165), .ZN(
        n21170) );
  AOI22_X1 U24129 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21236), .ZN(n21169) );
  OAI211_X1 U24130 ( .C1(n21242), .C2(n21224), .A(n21170), .B(n21169), .ZN(
        P1_U3152) );
  OR2_X1 U24131 ( .A1(n21172), .A2(n21171), .ZN(n21173) );
  NAND2_X1 U24132 ( .A1(n21173), .A2(n21198), .ZN(n21178) );
  NAND2_X1 U24133 ( .A1(n21178), .A2(n21186), .ZN(n21175) );
  NAND2_X1 U24134 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21185), .ZN(n21174) );
  NAND2_X1 U24135 ( .A1(n21175), .A2(n21174), .ZN(n21234) );
  INV_X1 U24136 ( .A(n21198), .ZN(n21233) );
  AOI22_X1 U24137 ( .A1(n21177), .A2(n21234), .B1(n21233), .B2(n21176), .ZN(
        n21189) );
  AOI21_X1 U24138 ( .B1(n21180), .B2(n21179), .A(n21178), .ZN(n21181) );
  INV_X1 U24139 ( .A(n21181), .ZN(n21183) );
  OAI221_X1 U24140 ( .B1(n21186), .B2(n21185), .C1(n21184), .C2(n21183), .A(
        n21182), .ZN(n21238) );
  AOI22_X1 U24141 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21238), .B1(
        n21237), .B2(n21187), .ZN(n21188) );
  OAI211_X1 U24142 ( .C1(n21190), .C2(n21241), .A(n21189), .B(n21188), .ZN(
        P1_U3153) );
  AOI22_X1 U24143 ( .A1(n21192), .A2(n21234), .B1(n21233), .B2(n21191), .ZN(
        n21195) );
  AOI22_X1 U24144 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21238), .B1(
        n21221), .B2(n21193), .ZN(n21194) );
  OAI211_X1 U24145 ( .C1(n21196), .C2(n21224), .A(n21195), .B(n21194), .ZN(
        P1_U3154) );
  INV_X1 U24146 ( .A(n21234), .ZN(n21199) );
  OAI22_X1 U24147 ( .A1(n21200), .A2(n21199), .B1(n21198), .B2(n21197), .ZN(
        n21201) );
  INV_X1 U24148 ( .A(n21201), .ZN(n21204) );
  AOI22_X1 U24149 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21238), .B1(
        n21237), .B2(n21202), .ZN(n21203) );
  OAI211_X1 U24150 ( .C1(n21205), .C2(n21241), .A(n21204), .B(n21203), .ZN(
        P1_U3155) );
  AOI22_X1 U24151 ( .A1(n21207), .A2(n21234), .B1(n21233), .B2(n21206), .ZN(
        n21210) );
  AOI22_X1 U24152 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21238), .B1(
        n21221), .B2(n21208), .ZN(n21209) );
  OAI211_X1 U24153 ( .C1(n21211), .C2(n21224), .A(n21210), .B(n21209), .ZN(
        P1_U3156) );
  AOI22_X1 U24154 ( .A1(n21213), .A2(n21234), .B1(n21233), .B2(n21212), .ZN(
        n21216) );
  AOI22_X1 U24155 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21238), .B1(
        n21221), .B2(n21214), .ZN(n21215) );
  OAI211_X1 U24156 ( .C1(n21217), .C2(n21224), .A(n21216), .B(n21215), .ZN(
        P1_U3157) );
  AOI22_X1 U24157 ( .A1(n21219), .A2(n21234), .B1(n21233), .B2(n21218), .ZN(
        n21223) );
  AOI22_X1 U24158 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21238), .B1(
        n21221), .B2(n21220), .ZN(n21222) );
  OAI211_X1 U24159 ( .C1(n21225), .C2(n21224), .A(n21223), .B(n21222), .ZN(
        P1_U3158) );
  AOI22_X1 U24160 ( .A1(n21227), .A2(n21234), .B1(n21233), .B2(n21226), .ZN(
        n21230) );
  AOI22_X1 U24161 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21238), .B1(
        n21237), .B2(n21228), .ZN(n21229) );
  OAI211_X1 U24162 ( .C1(n21231), .C2(n21241), .A(n21230), .B(n21229), .ZN(
        P1_U3159) );
  AOI22_X1 U24163 ( .A1(n21235), .A2(n21234), .B1(n21233), .B2(n21232), .ZN(
        n21240) );
  AOI22_X1 U24164 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21238), .B1(
        n21237), .B2(n21236), .ZN(n21239) );
  OAI211_X1 U24165 ( .C1(n21242), .C2(n21241), .A(n21240), .B(n21239), .ZN(
        P1_U3160) );
  INV_X1 U24166 ( .A(n21243), .ZN(n21245) );
  OAI211_X1 U24167 ( .C1(n21247), .C2(n21246), .A(n21245), .B(n21244), .ZN(
        P1_U3163) );
  AND2_X1 U24168 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21271), .ZN(
        P1_U3164) );
  AND2_X1 U24169 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21271), .ZN(
        P1_U3165) );
  AND2_X1 U24170 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21271), .ZN(
        P1_U3166) );
  AND2_X1 U24171 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21271), .ZN(
        P1_U3167) );
  AND2_X1 U24172 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21271), .ZN(
        P1_U3168) );
  AND2_X1 U24173 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21271), .ZN(
        P1_U3169) );
  AND2_X1 U24174 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21271), .ZN(
        P1_U3170) );
  AND2_X1 U24175 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21271), .ZN(
        P1_U3171) );
  AND2_X1 U24176 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21271), .ZN(
        P1_U3172) );
  AND2_X1 U24177 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21271), .ZN(
        P1_U3173) );
  AND2_X1 U24178 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21271), .ZN(
        P1_U3174) );
  AND2_X1 U24179 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21271), .ZN(
        P1_U3175) );
  AND2_X1 U24180 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21271), .ZN(
        P1_U3176) );
  AND2_X1 U24181 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21271), .ZN(
        P1_U3177) );
  AND2_X1 U24182 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21271), .ZN(
        P1_U3178) );
  AND2_X1 U24183 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21271), .ZN(
        P1_U3179) );
  AND2_X1 U24184 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21271), .ZN(
        P1_U3180) );
  AND2_X1 U24185 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21271), .ZN(
        P1_U3181) );
  AND2_X1 U24186 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21271), .ZN(
        P1_U3182) );
  AND2_X1 U24187 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21271), .ZN(
        P1_U3183) );
  AND2_X1 U24188 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21271), .ZN(
        P1_U3184) );
  AND2_X1 U24189 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21271), .ZN(
        P1_U3185) );
  AND2_X1 U24190 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21271), .ZN(P1_U3186) );
  AND2_X1 U24191 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21271), .ZN(P1_U3187) );
  AND2_X1 U24192 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21271), .ZN(P1_U3188) );
  AND2_X1 U24193 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21271), .ZN(P1_U3189) );
  AND2_X1 U24194 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21271), .ZN(P1_U3190) );
  AND2_X1 U24195 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21271), .ZN(P1_U3191) );
  AND2_X1 U24196 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21271), .ZN(P1_U3192) );
  AND2_X1 U24197 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21271), .ZN(P1_U3193) );
  NOR3_X1 U24198 ( .A1(n21302), .A2(NA), .A3(n21251), .ZN(n21249) );
  OAI22_X1 U24199 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21249), .B1(
        P1_STATE_REG_1__SCAN_IN), .B2(n21248), .ZN(n21255) );
  OAI21_X1 U24200 ( .B1(n21293), .B2(NA), .A(P1_STATE_REG_1__SCAN_IN), .ZN(
        n21250) );
  AOI21_X1 U24201 ( .B1(n21250), .B2(n21302), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21252) );
  OR2_X1 U24202 ( .A1(n21252), .A2(n21251), .ZN(n21253) );
  OAI22_X1 U24203 ( .A1(n21256), .A2(n21255), .B1(n21254), .B2(n21253), .ZN(
        P1_U3196) );
  AOI22_X1 U24204 ( .A1(n21266), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21265), .ZN(n21257) );
  OAI21_X1 U24205 ( .B1(n21258), .B2(n21268), .A(n21257), .ZN(P1_U3199) );
  AOI22_X1 U24206 ( .A1(n21266), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21265), .ZN(n21259) );
  OAI21_X1 U24207 ( .B1(n21260), .B2(n21268), .A(n21259), .ZN(P1_U3204) );
  AOI22_X1 U24208 ( .A1(n21266), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21265), .ZN(n21261) );
  OAI21_X1 U24209 ( .B1(n21262), .B2(n21268), .A(n21261), .ZN(P1_U3214) );
  AOI22_X1 U24210 ( .A1(n21266), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21265), .ZN(n21263) );
  OAI21_X1 U24211 ( .B1(n21264), .B2(n21268), .A(n21263), .ZN(P1_U3218) );
  AOI22_X1 U24212 ( .A1(n21266), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21265), .ZN(n21267) );
  OAI21_X1 U24213 ( .B1(n21269), .B2(n21268), .A(n21267), .ZN(P1_U3223) );
  INV_X1 U24214 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21272) );
  INV_X1 U24215 ( .A(n21273), .ZN(n21270) );
  AOI21_X1 U24216 ( .B1(n21272), .B2(n21271), .A(n21270), .ZN(P1_U3464) );
  OAI21_X1 U24217 ( .B1(n21275), .B2(n21274), .A(n21273), .ZN(P1_U3465) );
  AOI22_X1 U24218 ( .A1(n21279), .A2(n21278), .B1(n21277), .B2(n21276), .ZN(
        n21280) );
  INV_X1 U24219 ( .A(n21280), .ZN(n21283) );
  MUX2_X1 U24220 ( .A(n21283), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21281), .Z(P1_U3469) );
  AOI21_X1 U24221 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21285) );
  OAI221_X1 U24222 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21285), .C1(n21284), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n21290), .ZN(n21286) );
  OAI21_X1 U24223 ( .B1(n21290), .B2(n21287), .A(n21286), .ZN(P1_U3481) );
  OAI21_X1 U24224 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21290), .ZN(n21288) );
  OAI21_X1 U24225 ( .B1(n21290), .B2(n21289), .A(n21288), .ZN(P1_U3482) );
  AOI21_X1 U24226 ( .B1(n21293), .B2(n21292), .A(n21291), .ZN(n21295) );
  NAND3_X1 U24227 ( .A1(n9667), .A2(n21295), .A3(n21294), .ZN(n21303) );
  NOR2_X1 U24228 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21296), .ZN(n21301) );
  OAI211_X1 U24229 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21298), .A(n21297), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21299) );
  NAND2_X1 U24230 ( .A1(n21303), .A2(n21299), .ZN(n21300) );
  OAI22_X1 U24231 ( .A1(n21303), .A2(n21302), .B1(n21301), .B2(n21300), .ZN(
        P1_U3485) );
  AOI22_X1 U24232 ( .A1(n21307), .A2(n21306), .B1(n21305), .B2(n21304), .ZN(
        n21308) );
  INV_X1 U24233 ( .A(n21308), .ZN(n21314) );
  OAI22_X1 U24234 ( .A1(n21312), .A2(n21311), .B1(n21310), .B2(n21309), .ZN(
        n21313) );
  AOI211_X1 U24235 ( .C1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .C2(n21315), .A(
        n21314), .B(n21313), .ZN(n21470) );
  INV_X1 U24236 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n21317) );
  AOI22_X1 U24237 ( .A1(n21318), .A2(keyinput49), .B1(n21317), .B2(keyinput46), 
        .ZN(n21316) );
  OAI221_X1 U24238 ( .B1(n21318), .B2(keyinput49), .C1(n21317), .C2(keyinput46), .A(n21316), .ZN(n21328) );
  AOI22_X1 U24239 ( .A1(n17720), .A2(keyinput25), .B1(n21452), .B2(keyinput20), 
        .ZN(n21319) );
  OAI221_X1 U24240 ( .B1(n17720), .B2(keyinput25), .C1(n21452), .C2(keyinput20), .A(n21319), .ZN(n21327) );
  AOI22_X1 U24241 ( .A1(n21321), .A2(keyinput28), .B1(n17721), .B2(keyinput62), 
        .ZN(n21320) );
  OAI221_X1 U24242 ( .B1(n21321), .B2(keyinput28), .C1(n17721), .C2(keyinput62), .A(n21320), .ZN(n21326) );
  AOI22_X1 U24243 ( .A1(n21324), .A2(keyinput7), .B1(keyinput27), .B2(n21323), 
        .ZN(n21322) );
  OAI221_X1 U24244 ( .B1(n21324), .B2(keyinput7), .C1(n21323), .C2(keyinput27), 
        .A(n21322), .ZN(n21325) );
  NOR4_X1 U24245 ( .A1(n21328), .A2(n21327), .A3(n21326), .A4(n21325), .ZN(
        n21468) );
  INV_X1 U24246 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n21330) );
  AOI22_X1 U24247 ( .A1(n21451), .A2(keyinput50), .B1(keyinput45), .B2(n21330), 
        .ZN(n21329) );
  OAI221_X1 U24248 ( .B1(n21451), .B2(keyinput50), .C1(n21330), .C2(keyinput45), .A(n21329), .ZN(n21341) );
  AOI22_X1 U24249 ( .A1(n21333), .A2(keyinput47), .B1(n21332), .B2(keyinput6), 
        .ZN(n21331) );
  OAI221_X1 U24250 ( .B1(n21333), .B2(keyinput47), .C1(n21332), .C2(keyinput6), 
        .A(n21331), .ZN(n21340) );
  AOI22_X1 U24251 ( .A1(n21335), .A2(keyinput44), .B1(n16236), .B2(keyinput40), 
        .ZN(n21334) );
  OAI221_X1 U24252 ( .B1(n21335), .B2(keyinput44), .C1(n16236), .C2(keyinput40), .A(n21334), .ZN(n21339) );
  XNOR2_X1 U24253 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B(keyinput34), .ZN(
        n21337) );
  XNOR2_X1 U24254 ( .A(keyinput48), .B(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n21336) );
  NAND2_X1 U24255 ( .A1(n21337), .A2(n21336), .ZN(n21338) );
  NOR4_X1 U24256 ( .A1(n21341), .A2(n21340), .A3(n21339), .A4(n21338), .ZN(
        n21467) );
  AOI22_X1 U24257 ( .A1(n21343), .A2(keyinput24), .B1(n12363), .B2(keyinput13), 
        .ZN(n21342) );
  OAI221_X1 U24258 ( .B1(n21343), .B2(keyinput24), .C1(n12363), .C2(keyinput13), .A(n21342), .ZN(n21427) );
  AOI22_X1 U24259 ( .A1(n21346), .A2(keyinput30), .B1(n21345), .B2(keyinput38), 
        .ZN(n21344) );
  OAI221_X1 U24260 ( .B1(n21346), .B2(keyinput30), .C1(n21345), .C2(keyinput38), .A(n21344), .ZN(n21426) );
  OAI22_X1 U24261 ( .A1(n21349), .A2(keyinput33), .B1(n21348), .B2(keyinput36), 
        .ZN(n21347) );
  AOI221_X1 U24262 ( .B1(n21349), .B2(keyinput33), .C1(keyinput36), .C2(n21348), .A(n21347), .ZN(n21369) );
  OAI22_X1 U24263 ( .A1(n21352), .A2(keyinput55), .B1(n21351), .B2(keyinput51), 
        .ZN(n21350) );
  AOI221_X1 U24264 ( .B1(n21352), .B2(keyinput55), .C1(keyinput51), .C2(n21351), .A(n21350), .ZN(n21368) );
  AOI22_X1 U24265 ( .A1(n21437), .A2(keyinput3), .B1(keyinput17), .B2(n21354), 
        .ZN(n21353) );
  OAI221_X1 U24266 ( .B1(n21437), .B2(keyinput3), .C1(n21354), .C2(keyinput17), 
        .A(n21353), .ZN(n21366) );
  INV_X1 U24267 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n21356) );
  AOI22_X1 U24268 ( .A1(n21357), .A2(keyinput60), .B1(keyinput39), .B2(n21356), 
        .ZN(n21355) );
  OAI221_X1 U24269 ( .B1(n21357), .B2(keyinput60), .C1(n21356), .C2(keyinput39), .A(n21355), .ZN(n21365) );
  INV_X1 U24270 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n21436) );
  INV_X1 U24271 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21359) );
  AOI22_X1 U24272 ( .A1(n21436), .A2(keyinput59), .B1(n21359), .B2(keyinput1), 
        .ZN(n21358) );
  OAI221_X1 U24273 ( .B1(n21436), .B2(keyinput59), .C1(n21359), .C2(keyinput1), 
        .A(n21358), .ZN(n21364) );
  INV_X1 U24274 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n21360) );
  XOR2_X1 U24275 ( .A(n21360), .B(keyinput43), .Z(n21362) );
  XNOR2_X1 U24276 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B(keyinput15), .ZN(
        n21361) );
  NAND2_X1 U24277 ( .A1(n21362), .A2(n21361), .ZN(n21363) );
  NOR4_X1 U24278 ( .A1(n21366), .A2(n21365), .A3(n21364), .A4(n21363), .ZN(
        n21367) );
  NAND3_X1 U24279 ( .A1(n21369), .A2(n21368), .A3(n21367), .ZN(n21425) );
  INV_X1 U24280 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21372) );
  INV_X1 U24281 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21371) );
  AOI22_X1 U24282 ( .A1(n21372), .A2(keyinput4), .B1(keyinput5), .B2(n21371), 
        .ZN(n21370) );
  OAI221_X1 U24283 ( .B1(n21372), .B2(keyinput4), .C1(n21371), .C2(keyinput5), 
        .A(n21370), .ZN(n21383) );
  AOI22_X1 U24284 ( .A1(n21374), .A2(keyinput23), .B1(keyinput18), .B2(n21446), 
        .ZN(n21373) );
  OAI221_X1 U24285 ( .B1(n21374), .B2(keyinput23), .C1(n21446), .C2(keyinput18), .A(n21373), .ZN(n21382) );
  AOI22_X1 U24286 ( .A1(n21377), .A2(keyinput56), .B1(keyinput63), .B2(n21376), 
        .ZN(n21375) );
  OAI221_X1 U24287 ( .B1(n21377), .B2(keyinput56), .C1(n21376), .C2(keyinput63), .A(n21375), .ZN(n21381) );
  INV_X1 U24288 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n21442) );
  AOI22_X1 U24289 ( .A1(n21442), .A2(keyinput54), .B1(keyinput21), .B2(n21379), 
        .ZN(n21378) );
  OAI221_X1 U24290 ( .B1(n21442), .B2(keyinput54), .C1(n21379), .C2(keyinput21), .A(n21378), .ZN(n21380) );
  NOR4_X1 U24291 ( .A1(n21383), .A2(n21382), .A3(n21381), .A4(n21380), .ZN(
        n21423) );
  INV_X1 U24292 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n21447) );
  AOI22_X1 U24293 ( .A1(n21447), .A2(keyinput52), .B1(n21443), .B2(keyinput10), 
        .ZN(n21384) );
  OAI221_X1 U24294 ( .B1(n21447), .B2(keyinput52), .C1(n21443), .C2(keyinput10), .A(n21384), .ZN(n21395) );
  INV_X1 U24295 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21445) );
  AOI22_X1 U24296 ( .A1(n21386), .A2(keyinput2), .B1(keyinput26), .B2(n21445), 
        .ZN(n21385) );
  OAI221_X1 U24297 ( .B1(n21386), .B2(keyinput2), .C1(n21445), .C2(keyinput26), 
        .A(n21385), .ZN(n21394) );
  AOI22_X1 U24298 ( .A1(n21388), .A2(keyinput53), .B1(n21444), .B2(keyinput58), 
        .ZN(n21387) );
  OAI221_X1 U24299 ( .B1(n21388), .B2(keyinput53), .C1(n21444), .C2(keyinput58), .A(n21387), .ZN(n21393) );
  AOI22_X1 U24300 ( .A1(n21391), .A2(keyinput12), .B1(n21390), .B2(keyinput61), 
        .ZN(n21389) );
  OAI221_X1 U24301 ( .B1(n21391), .B2(keyinput12), .C1(n21390), .C2(keyinput61), .A(n21389), .ZN(n21392) );
  NOR4_X1 U24302 ( .A1(n21395), .A2(n21394), .A3(n21393), .A4(n21392), .ZN(
        n21422) );
  AOI22_X1 U24303 ( .A1(n21397), .A2(keyinput29), .B1(n10708), .B2(keyinput35), 
        .ZN(n21396) );
  OAI221_X1 U24304 ( .B1(n21397), .B2(keyinput29), .C1(n10708), .C2(keyinput35), .A(n21396), .ZN(n21401) );
  XNOR2_X1 U24305 ( .A(n21398), .B(keyinput19), .ZN(n21400) );
  XOR2_X1 U24306 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B(keyinput8), .Z(
        n21399) );
  OR3_X1 U24307 ( .A1(n21401), .A2(n21400), .A3(n21399), .ZN(n21408) );
  AOI22_X1 U24308 ( .A1(n12350), .A2(keyinput32), .B1(keyinput42), .B2(n21429), 
        .ZN(n21402) );
  OAI221_X1 U24309 ( .B1(n12350), .B2(keyinput32), .C1(n21429), .C2(keyinput42), .A(n21402), .ZN(n21407) );
  AOI22_X1 U24310 ( .A1(n21405), .A2(keyinput16), .B1(n21404), .B2(keyinput0), 
        .ZN(n21403) );
  OAI221_X1 U24311 ( .B1(n21405), .B2(keyinput16), .C1(n21404), .C2(keyinput0), 
        .A(n21403), .ZN(n21406) );
  NOR3_X1 U24312 ( .A1(n21408), .A2(n21407), .A3(n21406), .ZN(n21421) );
  AOI22_X1 U24313 ( .A1(n21410), .A2(keyinput11), .B1(n21450), .B2(keyinput37), 
        .ZN(n21409) );
  OAI221_X1 U24314 ( .B1(n21410), .B2(keyinput11), .C1(n21450), .C2(keyinput37), .A(n21409), .ZN(n21419) );
  AOI22_X1 U24315 ( .A1(n21428), .A2(keyinput41), .B1(n11232), .B2(keyinput9), 
        .ZN(n21411) );
  OAI221_X1 U24316 ( .B1(n21428), .B2(keyinput41), .C1(n11232), .C2(keyinput9), 
        .A(n21411), .ZN(n21418) );
  AOI22_X1 U24317 ( .A1(n9918), .A2(keyinput57), .B1(n13620), .B2(keyinput31), 
        .ZN(n21412) );
  OAI221_X1 U24318 ( .B1(n9918), .B2(keyinput57), .C1(n13620), .C2(keyinput31), 
        .A(n21412), .ZN(n21417) );
  INV_X1 U24319 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n21413) );
  XOR2_X1 U24320 ( .A(n21413), .B(keyinput14), .Z(n21415) );
  XNOR2_X1 U24321 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B(keyinput22), .ZN(
        n21414) );
  NAND2_X1 U24322 ( .A1(n21415), .A2(n21414), .ZN(n21416) );
  NOR4_X1 U24323 ( .A1(n21419), .A2(n21418), .A3(n21417), .A4(n21416), .ZN(
        n21420) );
  NAND4_X1 U24324 ( .A1(n21423), .A2(n21422), .A3(n21421), .A4(n21420), .ZN(
        n21424) );
  NOR4_X1 U24325 ( .A1(n21427), .A2(n21426), .A3(n21425), .A4(n21424), .ZN(
        n21466) );
  NAND4_X1 U24326 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(
        P3_MEMORYFETCH_REG_SCAN_IN), .A3(n21428), .A4(n11232), .ZN(n21435) );
  NAND4_X1 U24327 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_13__3__SCAN_IN), .A3(P2_BYTEENABLE_REG_0__SCAN_IN), 
        .A4(n10708), .ZN(n21434) );
  NOR2_X1 U24328 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(
        P1_REIP_REG_25__SCAN_IN), .ZN(n21432) );
  NAND2_X1 U24329 ( .A1(n21429), .A2(n13620), .ZN(n21430) );
  NOR2_X1 U24330 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21430), .ZN(
        n21431) );
  NAND4_X1 U24331 ( .A1(n21432), .A2(n21431), .A3(P2_DATAO_REG_8__SCAN_IN), 
        .A4(n9918), .ZN(n21433) );
  NOR4_X1 U24332 ( .A1(n21435), .A2(P3_REIP_REG_21__SCAN_IN), .A3(n21434), 
        .A4(n21433), .ZN(n21464) );
  NOR4_X1 U24333 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .A3(P1_UWORD_REG_7__SCAN_IN), .A4(
        n21436), .ZN(n21463) );
  NAND4_X1 U24334 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(P2_EBX_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(n17721), .ZN(n21441) );
  NAND4_X1 U24335 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P3_REIP_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n21440) );
  INV_X1 U24336 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n21438) );
  NAND4_X1 U24337 ( .A1(n21438), .A2(n21437), .A3(P3_LWORD_REG_14__SCAN_IN), 
        .A4(P3_LWORD_REG_7__SCAN_IN), .ZN(n21439) );
  NOR3_X1 U24338 ( .A1(n21441), .A2(n21440), .A3(n21439), .ZN(n21462) );
  NAND4_X1 U24339 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(n21443), .A4(n21442), .ZN(n21460) );
  NAND4_X1 U24340 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(DATAI_2_), .A3(n21445), 
        .A4(n21444), .ZN(n21459) );
  NOR4_X1 U24341 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(
        BUF1_REG_26__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A4(n21446), .ZN(n21448) );
  NAND4_X1 U24342 ( .A1(n21449), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A3(
        n21448), .A4(n21447), .ZN(n21458) );
  NOR4_X1 U24343 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(n16949), .A4(n21450), .ZN(n21456)
         );
  NOR4_X1 U24344 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(n21451), .A4(n16236), .ZN(n21455) );
  NOR4_X1 U24345 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_LWORD_REG_2__SCAN_IN), .A3(n17720), .A4(n21452), .ZN(n21454) );
  NOR4_X1 U24346 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        BUF2_REG_27__SCAN_IN), .A3(P1_DATAO_REG_13__SCAN_IN), .A4(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n21453) );
  NAND4_X1 U24347 ( .A1(n21456), .A2(n21455), .A3(n21454), .A4(n21453), .ZN(
        n21457) );
  NOR4_X1 U24348 ( .A1(n21460), .A2(n21459), .A3(n21458), .A4(n21457), .ZN(
        n21461) );
  NAND4_X1 U24349 ( .A1(n21464), .A2(n21463), .A3(n21462), .A4(n21461), .ZN(
        n21465) );
  NAND4_X1 U24350 ( .A1(n21468), .A2(n21467), .A3(n21466), .A4(n21465), .ZN(
        n21469) );
  XOR2_X1 U24351 ( .A(n21470), .B(n21469), .Z(P3_U2990) );
  INV_X1 U11096 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13862) );
  NAND2_X2 U11437 ( .A1(n10340), .A2(n10339), .ZN(n10414) );
  BUF_X1 U11432 ( .A(n11754), .Z(n12066) );
  CLKBUF_X1 U11384 ( .A(n10418), .Z(n20649) );
  XNOR2_X1 U11459 ( .A(n10509), .B(n10508), .ZN(n10775) );
  AND4_X1 U13425 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10340) );
  AND2_X2 U15094 ( .A1(n11908), .A2(n13875), .ZN(n11930) );
  AND2_X2 U15104 ( .A1(n13078), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11975) );
  CLKBUF_X1 U11048 ( .A(n13414), .Z(n11184) );
  CLKBUF_X2 U11082 ( .A(n10555), .Z(n9612) );
  XNOR2_X1 U11085 ( .A(n10691), .B(n10680), .ZN(n10831) );
  AND3_X1 U11106 ( .A1(n14122), .A2(n10444), .A3(n9815), .ZN(n9820) );
  CLKBUF_X1 U11109 ( .A(n14166), .Z(n20893) );
  CLKBUF_X1 U11111 ( .A(n12090), .Z(n12285) );
  CLKBUF_X1 U11116 ( .A(n12065), .Z(n12342) );
  CLKBUF_X1 U11130 ( .A(n12461), .Z(n19977) );
  CLKBUF_X1 U11135 ( .A(n11252), .Z(n17793) );
  CLKBUF_X1 U11148 ( .A(n10597), .Z(n20629) );
  CLKBUF_X1 U11156 ( .A(n9606), .Z(n20104) );
  CLKBUF_X1 U11167 ( .A(n14507), .Z(n14629) );
  NAND2_X1 U11173 ( .A1(n12478), .A2(n12004), .ZN(n21471) );
  AND2_X1 U11404 ( .A1(n10243), .A2(n10430), .ZN(n21472) );
endmodule

