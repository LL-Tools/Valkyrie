

module b20_C_AntiSAT_k_128_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10135;

  OAI222_X1 U4824 ( .A1(n7826), .A2(n7825), .B1(P1_U3086), .B2(n7858), .C1(
        n9807), .C2(n7823), .ZN(P1_U3328) );
  INV_X2 U4825 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4827 ( .A(n9383), .ZN(n9369) );
  CLKBUF_X1 U4828 ( .A(n5021), .Z(n7859) );
  BUF_X2 U4829 ( .A(n5824), .Z(n6132) );
  CLKBUF_X2 U4830 ( .A(n5049), .Z(n7862) );
  AND2_X1 U4831 ( .A1(n5778), .A2(n5769), .ZN(n5824) );
  NAND2_X2 U4832 ( .A1(n4463), .A2(n4390), .ZN(n4462) );
  NAND2_X1 U4833 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5768) );
  NAND4_X2 U4834 ( .A1(n5027), .A2(n5026), .A3(n5025), .A4(n5024), .ZN(n9411)
         );
  INV_X1 U4835 ( .A(n5021), .ZN(n5075) );
  CLKBUF_X2 U4836 ( .A(n6499), .Z(n4320) );
  CLKBUF_X1 U4837 ( .A(n10135), .Z(P2_U3893) );
  NOR2_X1 U4838 ( .A1(n6570), .A2(n6512), .ZN(n10135) );
  AND3_X1 U4839 ( .A1(n4873), .A2(n4870), .A3(n4869), .ZN(n8186) );
  INV_X1 U4840 ( .A(n5060), .ZN(n5394) );
  XNOR2_X1 U4841 ( .A(n8384), .B(n8073), .ZN(n8069) );
  NAND2_X1 U4842 ( .A1(n8614), .A2(n8589), .ZN(n8605) );
  AND2_X1 U4843 ( .A1(n8617), .A2(n8616), .ZN(n8633) );
  INV_X1 U4844 ( .A(n5694), .ZN(n6482) );
  INV_X1 U4845 ( .A(n4937), .ZN(n4938) );
  AND2_X2 U4846 ( .A1(n6631), .A2(n6650), .ZN(n5060) );
  OAI211_X1 U4847 ( .C1(n6653), .C2(n5217), .A(n4970), .B(n4969), .ZN(n6242)
         );
  AND3_X1 U4848 ( .A1(n5833), .A2(n5832), .A3(n5831), .ZN(n7088) );
  INV_X1 U4849 ( .A(n8606), .ZN(n8577) );
  AND3_X1 U4850 ( .A1(n5844), .A2(n5843), .A3(n5842), .ZN(n7346) );
  NAND2_X1 U4851 ( .A1(n8949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U4852 ( .A1(n6631), .A2(n7969), .ZN(n5217) );
  AND2_X1 U4853 ( .A1(n5460), .A2(n5459), .ZN(n9101) );
  CLKBUF_X3 U4854 ( .A(n6499), .Z(n4319) );
  INV_X1 U4855 ( .A(n9614), .ZN(n6260) );
  INV_X1 U4856 ( .A(n7240), .ZN(n9921) );
  OAI22_X1 U4857 ( .A1(n9554), .A2(n9553), .B1(n9560), .B2(n9544), .ZN(n9536)
         );
  XNOR2_X1 U4858 ( .A(n5315), .B(n5313), .ZN(n6783) );
  NAND4_X1 U4859 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n8388)
         );
  AOI21_X1 U4860 ( .B1(n8540), .B2(n8755), .A(n8539), .ZN(n8795) );
  AND3_X1 U4861 ( .A1(n5855), .A2(n5854), .A3(n5853), .ZN(n7875) );
  NAND3_X2 U4862 ( .A1(n4942), .A2(n4940), .A3(n4941), .ZN(n9413) );
  OAI222_X1 U4863 ( .A1(n7825), .A2(n6678), .B1(n9807), .B2(n6677), .C1(
        P1_U3086), .C2(n6820), .ZN(P1_U3347) );
  NAND2_X1 U4864 ( .A1(n9805), .A2(n4937), .ZN(n6499) );
  NOR2_X2 U4865 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4953) );
  NAND2_X2 U4866 ( .A1(n4441), .A2(n4880), .ZN(n6141) );
  OAI22_X2 U4868 ( .A1(n7614), .A2(n4586), .B1(n4585), .B2(n4587), .ZN(n8773)
         );
  NAND2_X2 U4871 ( .A1(n9688), .A2(n9687), .ZN(n9686) );
  OAI21_X2 U4872 ( .B1(n9700), .B2(n9228), .A(n9304), .ZN(n9688) );
  OAI222_X4 U4873 ( .A1(n8953), .A2(n6676), .B1(n8955), .B2(n6677), .C1(
        P2_U3151), .C2(n6675), .ZN(P2_U3287) );
  XNOR2_X2 U4874 ( .A(n5087), .B(SI_3_), .ZN(n5085) );
  NOR2_X2 U4875 ( .A1(n9108), .A2(n5703), .ZN(n6493) );
  INV_X1 U4876 ( .A(n6242), .ZN(n9205) );
  AOI22_X2 U4877 ( .A1(n7888), .A2(n7887), .B1(n7886), .B2(n8382), .ZN(n7890)
         );
  AOI22_X2 U4878 ( .A1(n9570), .A2(n9571), .B1(n9752), .B2(n9399), .ZN(n9554)
         );
  XNOR2_X2 U4879 ( .A(n5765), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5778) );
  XNOR2_X2 U4880 ( .A(n5768), .B(n5767), .ZN(n5777) );
  AOI21_X1 U4881 ( .B1(n9739), .B2(n10004), .A(n6306), .ZN(n6477) );
  AND2_X1 U4882 ( .A1(n4672), .A2(n4359), .ZN(n9188) );
  OR2_X1 U4883 ( .A1(n7453), .A2(n9145), .ZN(n7452) );
  OAI21_X2 U4884 ( .B1(n9214), .B2(n9859), .A(n9213), .ZN(n7453) );
  INV_X2 U4885 ( .A(n7936), .ZN(n7438) );
  NAND4_X1 U4886 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8384)
         );
  AND4_X1 U4887 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n8777)
         );
  NOR2_X1 U4888 ( .A1(n8392), .A2(n7054), .ZN(n8037) );
  AND3_X1 U4889 ( .A1(n5813), .A2(n5812), .A3(n5814), .ZN(n4560) );
  AND2_X1 U4891 ( .A1(n6628), .A2(n4997), .ZN(n6484) );
  NAND2_X2 U4892 ( .A1(n4846), .A2(n6177), .ZN(n5821) );
  NAND2_X1 U4893 ( .A1(n5711), .A2(n4950), .ZN(n6628) );
  NAND2_X1 U4894 ( .A1(n4957), .A2(n4956), .ZN(n9197) );
  NOR2_X1 U4895 ( .A1(n6141), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6138) );
  BUF_X2 U4896 ( .A(n7969), .Z(n9136) );
  CLKBUF_X3 U4897 ( .A(n5035), .Z(n7969) );
  INV_X4 U4899 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6993) );
  OAI21_X1 U4900 ( .B1(n4620), .B2(n4344), .A(n9113), .ZN(n4614) );
  AND2_X1 U4901 ( .A1(n9074), .A2(n4623), .ZN(n4622) );
  AND2_X1 U4902 ( .A1(n4325), .A2(n4623), .ZN(n4619) );
  AND2_X1 U4903 ( .A1(n4895), .A2(n4896), .ZN(n4325) );
  NOR2_X1 U4904 ( .A1(n9532), .A2(n9531), .ZN(n9737) );
  NAND2_X1 U4905 ( .A1(n7925), .A2(n7924), .ZN(n8324) );
  NOR2_X1 U4906 ( .A1(n9539), .A2(n9350), .ZN(n7853) );
  NAND2_X1 U4907 ( .A1(n4733), .A2(n4731), .ZN(n8247) );
  AOI21_X1 U4908 ( .B1(n4721), .B2(n4724), .A(n4719), .ZN(n4718) );
  AND2_X1 U4909 ( .A1(n8332), .A2(n8334), .ZN(n7891) );
  NAND2_X1 U4910 ( .A1(n4424), .A2(n4370), .ZN(n4672) );
  NAND2_X1 U4911 ( .A1(n8756), .A2(n4365), .ZN(n8744) );
  AOI21_X1 U4912 ( .B1(n4354), .B2(n4330), .A(n4728), .ZN(n4727) );
  OAI21_X1 U4913 ( .B1(n7571), .B2(n9158), .A(n6253), .ZN(n7625) );
  AOI21_X1 U4914 ( .B1(n4662), .B2(n4668), .A(n4660), .ZN(n4659) );
  NAND2_X1 U4915 ( .A1(n7452), .A2(n6284), .ZN(n7575) );
  NAND2_X1 U4916 ( .A1(n7205), .A2(n7204), .ZN(n7416) );
  NAND2_X2 U4917 ( .A1(n5748), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9129) );
  OR2_X1 U4918 ( .A1(n8968), .A2(n9127), .ZN(n9299) );
  INV_X2 U4919 ( .A(n9713), .ZN(n4321) );
  AND2_X1 U4920 ( .A1(n9278), .A2(n9281), .ZN(n9158) );
  OR2_X1 U4921 ( .A1(n7586), .A2(n8989), .ZN(n9278) );
  NAND2_X1 U4922 ( .A1(n5294), .A2(n5293), .ZN(n7631) );
  INV_X1 U4923 ( .A(n8777), .ZN(n8382) );
  OR2_X1 U4924 ( .A1(n7590), .A2(n7295), .ZN(n9843) );
  NAND4_X1 U4925 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(n8383)
         );
  NAND2_X1 U4926 ( .A1(n5191), .A2(n5190), .ZN(n7590) );
  NAND4_X1 U4927 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n8392)
         );
  NAND2_X1 U4929 ( .A1(n5237), .A2(n5236), .ZN(n5259) );
  CLKBUF_X1 U4930 ( .A(n5728), .Z(n9384) );
  NAND2_X1 U4931 ( .A1(n5163), .A2(n5162), .ZN(n9945) );
  AND3_X1 U4932 ( .A1(n4562), .A2(n4561), .A3(n5815), .ZN(n6976) );
  INV_X2 U4933 ( .A(n7984), .ZN(n7975) );
  INV_X4 U4934 ( .A(n5014), .ZN(n5697) );
  NAND4_X1 U4935 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n9410)
         );
  NOR2_X1 U4936 ( .A1(n5445), .A2(n4982), .ZN(n4988) );
  INV_X1 U4937 ( .A(n6484), .ZN(n5014) );
  NAND4_X1 U4938 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n9880)
         );
  NAND4_X1 U4939 ( .A1(n5199), .A2(n5198), .A3(n5197), .A4(n5196), .ZN(n9408)
         );
  NAND2_X1 U4940 ( .A1(n5160), .A2(n5159), .ZN(n5176) );
  NAND2_X1 U4941 ( .A1(n5426), .A2(n4981), .ZN(n5445) );
  MUX2_X1 U4942 ( .A(n6199), .B(n5865), .S(n5762), .Z(n6201) );
  XNOR2_X1 U4943 ( .A(n5784), .B(n5783), .ZN(n6177) );
  OR2_X1 U4944 ( .A1(n5921), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5968) );
  AND2_X1 U4945 ( .A1(n5707), .A2(n5708), .ZN(n4950) );
  AND2_X1 U4946 ( .A1(n9197), .A2(n9375), .ZN(n4997) );
  AOI21_X1 U4947 ( .B1(n4549), .B2(n4547), .A(n4546), .ZN(n4545) );
  MUX2_X1 U4948 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4947), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n4949) );
  NOR2_X1 U4949 ( .A1(n6141), .A2(n4606), .ZN(n6200) );
  NOR2_X1 U4950 ( .A1(n5896), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5908) );
  AND2_X1 U4951 ( .A1(n4965), .A2(n4964), .ZN(n4656) );
  OAI211_X2 U4952 ( .C1(n4769), .C2(n4655), .A(n4654), .B(n4652), .ZN(n7858)
         );
  NAND2_X1 U4953 ( .A1(n4493), .A2(n4420), .ZN(n4657) );
  NAND2_X1 U4954 ( .A1(n4769), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U4955 ( .A1(n5261), .A2(n5260), .ZN(n5285) );
  NAND2_X2 U4956 ( .A1(n4817), .A2(n4815), .ZN(n5035) );
  INV_X1 U4957 ( .A(n4743), .ZN(n4440) );
  AND3_X1 U4958 ( .A1(n5289), .A2(n4976), .A3(n4920), .ZN(n4923) );
  NOR2_X2 U4959 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5289) );
  INV_X4 U4960 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4961 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5829) );
  INV_X1 U4962 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4921) );
  INV_X1 U4963 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4952) );
  INV_X1 U4964 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8504) );
  INV_X1 U4965 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4476) );
  INV_X1 U4966 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4655) );
  INV_X2 U4967 ( .A(n8622), .ZN(n8327) );
  NAND2_X1 U4968 ( .A1(n4985), .A2(n4921), .ZN(n4982) );
  OAI221_X1 U4969 ( .B1(n8203), .B2(keyinput58), .C1(n4921), .C2(keyinput39), 
        .A(n6453), .ZN(n6461) );
  NOR2_X2 U4970 ( .A1(n9563), .A2(n9562), .ZN(n9561) );
  NAND3_X1 U4971 ( .A1(n4998), .A2(n6628), .A3(n7237), .ZN(n6486) );
  NOR3_X4 U4972 ( .A1(n9111), .A2(n9110), .A3(n9109), .ZN(n9108) );
  NAND2_X2 U4973 ( .A1(n4890), .A2(n4891), .ZN(n9111) );
  NOR2_X2 U4974 ( .A1(n9528), .A2(n9529), .ZN(n9527) );
  AND2_X2 U4975 ( .A1(n5728), .A2(n9197), .ZN(n6267) );
  AND2_X1 U4976 ( .A1(n6631), .A2(n6650), .ZN(n4322) );
  AOI21_X1 U4977 ( .B1(n4545), .B2(n4548), .A(n4544), .ZN(n4543) );
  NAND2_X1 U4978 ( .A1(n4506), .A2(n4858), .ZN(n4857) );
  NAND2_X1 U4979 ( .A1(n8034), .A2(n8171), .ZN(n4506) );
  NAND2_X1 U4980 ( .A1(n5214), .A2(n5213), .ZN(n5236) );
  AOI21_X1 U4981 ( .B1(n4574), .B2(n4572), .A(n4379), .ZN(n4571) );
  INV_X1 U4982 ( .A(n4353), .ZN(n4572) );
  INV_X1 U4983 ( .A(n5209), .ZN(n4546) );
  INV_X1 U4984 ( .A(n5175), .ZN(n4547) );
  NAND2_X1 U4985 ( .A1(n7120), .A2(n7121), .ZN(n7119) );
  NAND2_X1 U4986 ( .A1(n4855), .A2(n4371), .ZN(n8044) );
  NAND2_X1 U4987 ( .A1(n4856), .A2(n8039), .ZN(n4855) );
  NAND2_X1 U4988 ( .A1(n4857), .A2(n8038), .ZN(n4856) );
  NAND2_X1 U4989 ( .A1(n8098), .A2(n8097), .ZN(n8102) );
  NAND2_X1 U4990 ( .A1(n4862), .A2(n4860), .ZN(n4859) );
  AND2_X1 U4991 ( .A1(n8126), .A2(n4864), .ZN(n8112) );
  NOR2_X1 U4992 ( .A1(n8695), .A2(n8110), .ZN(n4864) );
  NAND2_X1 U4993 ( .A1(n4814), .A2(n8113), .ZN(n6163) );
  INV_X1 U4994 ( .A(n8658), .ZN(n4814) );
  AND2_X1 U4995 ( .A1(n5355), .A2(n4887), .ZN(n4886) );
  NAND2_X1 U4996 ( .A1(n9066), .A2(n4888), .ZN(n4887) );
  INV_X1 U4997 ( .A(n5312), .ZN(n4888) );
  AND2_X1 U4998 ( .A1(n4324), .A2(n4927), .ZN(n4492) );
  INV_X1 U4999 ( .A(n5492), .ZN(n4535) );
  INV_X1 U5000 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U5001 ( .A1(n5210), .A2(n4550), .ZN(n4549) );
  INV_X1 U5002 ( .A(n5179), .ZN(n4550) );
  OR2_X1 U5003 ( .A1(n8791), .A2(n7993), .ZN(n8176) );
  NAND2_X1 U5004 ( .A1(n4878), .A2(n4607), .ZN(n4606) );
  INV_X1 U5005 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4607) );
  NOR2_X1 U5006 ( .A1(n5761), .A2(n4879), .ZN(n4878) );
  NAND2_X1 U5007 ( .A1(n5762), .A2(n5759), .ZN(n4879) );
  OAI21_X1 U5008 ( .B1(n6172), .B2(n4460), .A(n4459), .ZN(n7992) );
  AOI21_X1 U5009 ( .B1(n4788), .B2(n8159), .A(n4789), .ZN(n4459) );
  INV_X1 U5010 ( .A(n4788), .ZN(n4460) );
  OR2_X1 U5011 ( .A1(n8178), .A2(n8208), .ZN(n7943) );
  INV_X1 U5012 ( .A(n8106), .ZN(n4458) );
  OR2_X2 U5013 ( .A1(n6976), .A2(n8390), .ZN(n8039) );
  OR2_X1 U5014 ( .A1(n8530), .A2(n8538), .ZN(n8175) );
  OR2_X1 U5015 ( .A1(n8268), .A2(n8358), .ZN(n8155) );
  OR2_X1 U5016 ( .A1(n8650), .A2(n8251), .ZN(n8132) );
  OR2_X1 U5017 ( .A1(n8907), .A2(n8645), .ZN(n8130) );
  OR2_X1 U5018 ( .A1(n8925), .A2(n8710), .ZN(n8654) );
  OR2_X1 U5019 ( .A1(n8941), .A2(n8759), .ZN(n4578) );
  INV_X1 U5020 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U5021 ( .A1(n4341), .A2(n4897), .ZN(n4896) );
  OR2_X1 U5022 ( .A1(n9728), .A2(n9530), .ZN(n9363) );
  NAND2_X1 U5023 ( .A1(n7958), .A2(n9543), .ZN(n4699) );
  NAND2_X1 U5024 ( .A1(n6298), .A2(n9543), .ZN(n9182) );
  OR2_X1 U5025 ( .A1(n6298), .A2(n9543), .ZN(n9354) );
  OR2_X1 U5026 ( .A1(n9742), .A2(n9564), .ZN(n9349) );
  NOR2_X1 U5027 ( .A1(n4339), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4900) );
  AND2_X1 U5028 ( .A1(n4927), .A2(n4928), .ZN(n4773) );
  NAND2_X1 U5029 ( .A1(n4540), .A2(n5622), .ZN(n5645) );
  OAI21_X1 U5030 ( .B1(n5544), .B2(n5543), .A(n5542), .ZN(n5567) );
  INV_X1 U5031 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4981) );
  AND2_X1 U5032 ( .A1(n5515), .A2(n5497), .ZN(n5513) );
  NOR2_X1 U5033 ( .A1(n5464), .A2(n4539), .ZN(n4538) );
  INV_X1 U5034 ( .A(n5444), .ZN(n4539) );
  NAND2_X1 U5035 ( .A1(n5285), .A2(n5263), .ZN(n5286) );
  INV_X1 U5036 ( .A(n5255), .ZN(n4808) );
  NAND2_X1 U5037 ( .A1(n5181), .A2(n5180), .ZN(n5209) );
  INV_X1 U5038 ( .A(n7667), .ZN(n4730) );
  INV_X1 U5039 ( .A(n6118), .ZN(n6181) );
  INV_X1 U5040 ( .A(n5857), .ZN(n6054) );
  OAI211_X1 U5041 ( .C1(n7119), .C2(n4831), .A(n4825), .B(n4826), .ZN(n7192)
         );
  NOR2_X1 U5042 ( .A1(n4827), .A2(n7065), .ZN(n4826) );
  XNOR2_X1 U5043 ( .A(n7992), .B(n8024), .ZN(n6188) );
  AOI21_X1 U5044 ( .B1(n8773), .B2(n5925), .A(n4902), .ZN(n8758) );
  NOR2_X1 U5045 ( .A1(n4356), .A2(n4583), .ZN(n4582) );
  INV_X1 U5046 ( .A(n5874), .ZN(n4583) );
  INV_X1 U5047 ( .A(n4571), .ZN(n4567) );
  NAND2_X1 U5048 ( .A1(n4576), .A2(n4569), .ZN(n4566) );
  OAI22_X1 U5049 ( .A1(n9801), .A2(n7984), .B1(n7983), .B2(n6700), .ZN(n7999)
         );
  AND2_X1 U5050 ( .A1(n8095), .A2(n4387), .ZN(n4457) );
  INV_X1 U5051 ( .A(n7983), .ZN(n6013) );
  INV_X1 U5052 ( .A(n5821), .ZN(n6012) );
  NAND2_X1 U5053 ( .A1(n4462), .A2(n6177), .ZN(n4461) );
  INV_X1 U5054 ( .A(n5035), .ZN(n6650) );
  NAND2_X1 U5055 ( .A1(n9458), .A2(n9457), .ZN(n9472) );
  AND2_X1 U5056 ( .A1(n9762), .A2(n9400), .ZN(n6263) );
  INV_X2 U5057 ( .A(n5217), .ZN(n9137) );
  AND2_X1 U5058 ( .A1(n4771), .A2(n4655), .ZN(n4653) );
  XNOR2_X1 U5059 ( .A(n5645), .B(n5644), .ZN(n7796) );
  OAI21_X1 U5060 ( .B1(n5259), .B2(n4802), .A(n4800), .ZN(n5332) );
  XNOR2_X1 U5061 ( .A(n5057), .B(n5036), .ZN(n5055) );
  NAND2_X1 U5062 ( .A1(n9250), .A2(n4497), .ZN(n4496) );
  OR2_X1 U5063 ( .A1(n9259), .A2(n9383), .ZN(n4495) );
  NOR2_X1 U5064 ( .A1(n9369), .A2(n4498), .ZN(n4497) );
  NAND2_X1 U5065 ( .A1(n8092), .A2(n8091), .ZN(n4862) );
  NAND2_X1 U5066 ( .A1(n9707), .A2(n4332), .ZN(n4487) );
  INV_X1 U5067 ( .A(n9324), .ZN(n4486) );
  AOI21_X1 U5068 ( .B1(n8129), .B2(n8133), .A(n8128), .ZN(n4854) );
  NAND2_X1 U5069 ( .A1(n8117), .A2(n8684), .ZN(n4851) );
  NAND2_X1 U5070 ( .A1(n4865), .A2(n8707), .ZN(n8126) );
  OAI21_X1 U5071 ( .B1(n8103), .B2(n4867), .A(n4866), .ZN(n4865) );
  INV_X1 U5072 ( .A(n8108), .ZN(n4866) );
  INV_X1 U5073 ( .A(n8140), .ZN(n4853) );
  NAND2_X1 U5074 ( .A1(n4489), .A2(n9253), .ZN(n9249) );
  INV_X1 U5075 ( .A(n9252), .ZN(n4489) );
  INV_X1 U5076 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4915) );
  OR4_X1 U5077 ( .A1(n8025), .A2(n8024), .A3(n8541), .A4(n8023), .ZN(n8026) );
  OR3_X1 U5078 ( .A1(n8558), .A2(n8548), .A3(n8022), .ZN(n8023) );
  NOR2_X1 U5079 ( .A1(n7546), .A2(n6613), .ZN(n6615) );
  AOI21_X1 U5080 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7745), .A(n7739), .ZN(
        n6617) );
  AND3_X1 U5081 ( .A1(n4840), .A2(n4839), .A3(n4417), .ZN(n8425) );
  NOR2_X1 U5082 ( .A1(n6050), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U5083 ( .A1(n6027), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4433) );
  NOR2_X1 U5084 ( .A1(n5972), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4432) );
  NOR2_X1 U5085 ( .A1(n5916), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4431) );
  OAI21_X1 U5086 ( .B1(n7613), .B2(n4589), .A(n5913), .ZN(n4588) );
  NAND2_X1 U5087 ( .A1(n7775), .A2(n8382), .ZN(n4590) );
  NAND2_X1 U5088 ( .A1(n4810), .A2(n4809), .ZN(n6172) );
  NOR2_X1 U5089 ( .A1(n8157), .A2(n8160), .ZN(n4809) );
  AND2_X1 U5090 ( .A1(n6082), .A2(n6081), .ZN(n8568) );
  AND2_X1 U5091 ( .A1(n8597), .A2(n8606), .ZN(n8148) );
  AND2_X1 U5092 ( .A1(n6170), .A2(n8622), .ZN(n8145) );
  INV_X1 U5093 ( .A(n8896), .ZN(n7919) );
  OR2_X1 U5094 ( .A1(n8896), .A2(n8646), .ZN(n8138) );
  NAND2_X1 U5095 ( .A1(n8352), .A2(n8686), .ZN(n8120) );
  INV_X1 U5096 ( .A(n8125), .ZN(n4451) );
  OR2_X1 U5097 ( .A1(n6200), .A2(n5865), .ZN(n5785) );
  NOR2_X1 U5098 ( .A1(n4596), .A2(n4593), .ZN(n4882) );
  NOR2_X1 U5099 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4594) );
  INV_X1 U5100 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U5101 ( .A1(n4633), .A2(n4355), .ZN(n4898) );
  AOI21_X1 U5102 ( .B1(n7292), .B2(n7293), .A(n4635), .ZN(n4634) );
  AOI21_X1 U5103 ( .B1(n4886), .B2(n4889), .A(n4405), .ZN(n4885) );
  INV_X1 U5104 ( .A(n9066), .ZN(n4889) );
  OR2_X1 U5105 ( .A1(n9735), .A2(n7866), .ZN(n9358) );
  NOR2_X1 U5106 ( .A1(n9752), .A2(n9757), .ZN(n4783) );
  NOR2_X1 U5107 ( .A1(n9746), .A2(n4782), .ZN(n4781) );
  INV_X1 U5108 ( .A(n4783), .ZN(n4782) );
  NOR2_X1 U5109 ( .A1(n9586), .A2(n4707), .ZN(n4706) );
  NOR2_X1 U5110 ( .A1(n4708), .A2(n6263), .ZN(n4707) );
  OR2_X1 U5111 ( .A1(n9752), .A2(n9592), .ZN(n9340) );
  OR2_X1 U5112 ( .A1(n9757), .A2(n9079), .ZN(n9336) );
  NOR2_X1 U5113 ( .A1(n6288), .A2(n6287), .ZN(n4671) );
  OR2_X1 U5114 ( .A1(n9772), .A2(n9663), .ZN(n9321) );
  OR2_X1 U5115 ( .A1(n9719), .A2(n9046), .ZN(n9304) );
  OR2_X1 U5116 ( .A1(n7817), .A2(n9037), .ZN(n9300) );
  INV_X1 U5117 ( .A(n7622), .ZN(n4665) );
  AND2_X1 U5118 ( .A1(n7303), .A2(n4323), .ZN(n4680) );
  INV_X1 U5119 ( .A(n4348), .ZN(n4684) );
  INV_X1 U5120 ( .A(n6249), .ZN(n4702) );
  INV_X1 U5121 ( .A(n6276), .ZN(n4647) );
  INV_X1 U5122 ( .A(n9207), .ZN(n4650) );
  NOR2_X1 U5123 ( .A1(n9653), .A2(n9772), .ZN(n9644) );
  OR2_X1 U5124 ( .A1(n7631), .A2(n8968), .ZN(n4775) );
  NOR2_X1 U5125 ( .A1(n7813), .A2(n7817), .ZN(n9716) );
  OR2_X1 U5126 ( .A1(n9869), .A2(n9945), .ZN(n9852) );
  AOI21_X1 U5127 ( .B1(n5647), .B2(n4525), .A(n4523), .ZN(n4522) );
  NAND2_X1 U5128 ( .A1(n4524), .A2(n5677), .ZN(n4523) );
  NAND2_X1 U5129 ( .A1(n4525), .A2(n4527), .ZN(n4524) );
  NAND2_X1 U5130 ( .A1(n4541), .A2(n5596), .ZN(n5621) );
  NAND2_X1 U5131 ( .A1(n5516), .A2(n5515), .ZN(n5544) );
  AOI21_X1 U5132 ( .B1(n4531), .B2(n4534), .A(n4530), .ZN(n4529) );
  INV_X1 U5133 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4978) );
  INV_X1 U5134 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4979) );
  AOI21_X1 U5135 ( .B1(n4800), .B2(n4802), .A(n5331), .ZN(n4799) );
  NAND2_X1 U5136 ( .A1(n5257), .A2(SI_10_), .ZN(n5258) );
  INV_X1 U5137 ( .A(n4549), .ZN(n4548) );
  INV_X1 U5138 ( .A(n5114), .ZN(n4520) );
  INV_X1 U5139 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4816) );
  NAND2_X1 U5140 ( .A1(n4430), .A2(n4429), .ZN(n5902) );
  INV_X1 U5141 ( .A(n5890), .ZN(n4430) );
  NOR2_X1 U5142 ( .A1(n8308), .A2(n4735), .ZN(n4734) );
  INV_X1 U5143 ( .A(n4736), .ZN(n4735) );
  NOR2_X1 U5144 ( .A1(n4739), .A2(n8308), .ZN(n4732) );
  XNOR2_X1 U5145 ( .A(n8872), .B(n7438), .ZN(n7935) );
  NAND2_X1 U5146 ( .A1(n7440), .A2(n7441), .ZN(n4716) );
  INV_X1 U5147 ( .A(n7282), .ZN(n4715) );
  OR2_X1 U5148 ( .A1(n7280), .A2(n7341), .ZN(n4717) );
  NOR2_X1 U5149 ( .A1(n7767), .A2(n7768), .ZN(n4728) );
  AOI21_X1 U5150 ( .B1(n4739), .B2(n4738), .A(n4737), .ZN(n4736) );
  INV_X1 U5151 ( .A(n8238), .ZN(n4737) );
  INV_X1 U5152 ( .A(n7913), .ZN(n4738) );
  AND2_X1 U5153 ( .A1(n7912), .A2(n8341), .ZN(n7913) );
  OR2_X1 U5154 ( .A1(n8342), .A2(n8288), .ZN(n7912) );
  AND2_X1 U5155 ( .A1(n6047), .A2(n6046), .ZN(n7927) );
  OAI21_X1 U5156 ( .B1(n7038), .B2(n6597), .A(n4823), .ZN(n7041) );
  AOI22_X1 U5157 ( .A1(n7036), .A2(n7037), .B1(n7038), .B2(n6519), .ZN(n6935)
         );
  INV_X1 U5158 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6928) );
  INV_X1 U5159 ( .A(n6604), .ZN(n4830) );
  NAND2_X1 U5160 ( .A1(n4765), .A2(n7185), .ZN(n7187) );
  INV_X1 U5161 ( .A(n4766), .ZN(n4765) );
  OR2_X1 U5162 ( .A1(n6607), .A2(n7329), .ZN(n4474) );
  NAND2_X1 U5163 ( .A1(n6581), .A2(n7329), .ZN(n7367) );
  NAND2_X1 U5164 ( .A1(n4750), .A2(n7367), .ZN(n7369) );
  INV_X1 U5165 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U5166 ( .A1(n4474), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5167 ( .A1(n6607), .A2(n7329), .ZN(n7354) );
  AND2_X1 U5168 ( .A1(n6585), .A2(n7474), .ZN(n6587) );
  NOR2_X1 U5169 ( .A1(n7548), .A2(n7547), .ZN(n7546) );
  NAND2_X1 U5170 ( .A1(n4758), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4757) );
  INV_X1 U5171 ( .A(n6587), .ZN(n4756) );
  XNOR2_X1 U5172 ( .A(n6615), .B(n6614), .ZN(n7655) );
  NAND2_X1 U5173 ( .A1(n4475), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4822) );
  INV_X1 U5174 ( .A(n7655), .ZN(n4475) );
  NOR2_X1 U5175 ( .A1(n7543), .A2(n6589), .ZN(n6590) );
  AOI21_X1 U5176 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7745), .A(n7732), .ZN(
        n6592) );
  OR2_X1 U5177 ( .A1(n7787), .A2(n4841), .ZN(n4839) );
  OR2_X1 U5178 ( .A1(n6620), .A2(n6555), .ZN(n4841) );
  OR2_X1 U5179 ( .A1(n4346), .A2(n6620), .ZN(n4840) );
  OR2_X1 U5180 ( .A1(n7787), .A2(n6555), .ZN(n4842) );
  XNOR2_X1 U5181 ( .A(n8425), .B(n8426), .ZN(n8403) );
  NOR2_X1 U5182 ( .A1(n8393), .A2(n4426), .ZN(n8414) );
  NOR2_X1 U5183 ( .A1(n6619), .A2(n7883), .ZN(n4426) );
  NOR2_X1 U5184 ( .A1(n8403), .A2(n8404), .ZN(n8427) );
  AOI21_X1 U5185 ( .B1(n6188), .B2(n7757), .A(n6185), .ZN(n6186) );
  AND2_X1 U5186 ( .A1(n6110), .A2(n6109), .ZN(n8537) );
  NAND2_X1 U5187 ( .A1(n4575), .A2(n4351), .ZN(n4574) );
  INV_X1 U5188 ( .A(n8548), .ZN(n4575) );
  AND2_X1 U5189 ( .A1(n7944), .A2(n7943), .ZN(n8535) );
  OR2_X1 U5190 ( .A1(n6088), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U5191 ( .A1(n4427), .A2(n8301), .ZN(n6066) );
  INV_X1 U5192 ( .A(n4427), .ZN(n6057) );
  OR2_X1 U5193 ( .A1(n6044), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6050) );
  OR2_X1 U5194 ( .A1(n5999), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6018) );
  AND4_X1 U5195 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8710)
         );
  NAND2_X1 U5196 ( .A1(n4455), .A2(n4458), .ZN(n4452) );
  NAND2_X1 U5197 ( .A1(n4458), .A2(n6157), .ZN(n4453) );
  OR2_X1 U5198 ( .A1(n5943), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5957) );
  INV_X1 U5199 ( .A(n4431), .ZN(n5792) );
  NAND2_X1 U5200 ( .A1(n4385), .A2(n8080), .ZN(n4446) );
  NAND2_X1 U5201 ( .A1(n8080), .A2(n8079), .ZN(n4447) );
  NAND2_X1 U5202 ( .A1(n4448), .A2(n8072), .ZN(n7754) );
  OR2_X1 U5203 ( .A1(n7611), .A2(n6153), .ZN(n4448) );
  NAND2_X1 U5204 ( .A1(n7559), .A2(n8078), .ZN(n7611) );
  OR2_X1 U5205 ( .A1(n7666), .A2(n8073), .ZN(n5901) );
  NAND2_X1 U5206 ( .A1(n7614), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U5207 ( .A1(n4581), .A2(n4579), .ZN(n7561) );
  NOR2_X1 U5208 ( .A1(n5887), .A2(n4580), .ZN(n4579) );
  OAI21_X1 U5209 ( .B1(n7481), .B2(n7480), .A(n8063), .ZN(n7558) );
  OR2_X1 U5210 ( .A1(n7558), .A2(n8069), .ZN(n7559) );
  NAND2_X1 U5211 ( .A1(n5772), .A2(n5771), .ZN(n5876) );
  INV_X1 U5212 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5771) );
  INV_X1 U5213 ( .A(n5859), .ZN(n5772) );
  OR2_X1 U5214 ( .A1(n7983), .A2(n6654), .ZN(n4562) );
  OR2_X1 U5215 ( .A1(n7984), .A2(n6653), .ZN(n4561) );
  INV_X1 U5216 ( .A(n8535), .ZN(n8541) );
  NAND2_X1 U5217 ( .A1(n6172), .A2(n8000), .ZN(n8547) );
  OR2_X1 U5218 ( .A1(n8159), .A2(n8160), .ZN(n8558) );
  NAND2_X1 U5219 ( .A1(n8581), .A2(n8155), .ZN(n4810) );
  AOI21_X1 U5220 ( .B1(n8586), .B2(n8149), .A(n8148), .ZN(n8581) );
  NAND2_X1 U5221 ( .A1(n4611), .A2(n4609), .ZN(n8573) );
  NOR2_X1 U5222 ( .A1(n6075), .A2(n4610), .ZN(n4609) );
  INV_X1 U5223 ( .A(n6024), .ZN(n4610) );
  OR2_X1 U5224 ( .A1(n8890), .A2(n7927), .ZN(n8143) );
  NAND2_X1 U5225 ( .A1(n8612), .A2(n8141), .ZN(n4812) );
  NAND2_X1 U5226 ( .A1(n6165), .A2(n4914), .ZN(n6166) );
  OR2_X1 U5227 ( .A1(n8919), .A2(n8698), .ZN(n8670) );
  AND4_X1 U5228 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n8699)
         );
  NAND2_X1 U5229 ( .A1(n8744), .A2(n4578), .ZN(n4577) );
  INV_X1 U5230 ( .A(n8780), .ZN(n8760) );
  INV_X1 U5231 ( .A(n8778), .ZN(n8761) );
  AND2_X1 U5232 ( .A1(n8095), .A2(n8096), .ZN(n8743) );
  NAND2_X1 U5233 ( .A1(n4441), .A2(n4397), .ZN(n5896) );
  NOR2_X1 U5234 ( .A1(n5591), .A2(n5590), .ZN(n9052) );
  NAND2_X1 U5235 ( .A1(n6265), .A2(n9204), .ZN(n4642) );
  NAND2_X1 U5236 ( .A1(n5279), .A2(n5280), .ZN(n9012) );
  INV_X1 U5237 ( .A(n9024), .ZN(n4892) );
  NAND2_X1 U5238 ( .A1(n8972), .A2(n4335), .ZN(n4895) );
  INV_X1 U5239 ( .A(n9052), .ZN(n4625) );
  NAND2_X1 U5240 ( .A1(n4899), .A2(n7593), .ZN(n4631) );
  NOR2_X1 U5241 ( .A1(n5133), .A2(n5132), .ZN(n5164) );
  OR2_X1 U5242 ( .A1(n5075), .A2(n5076), .ZN(n5083) );
  NOR2_X1 U5243 ( .A1(n4977), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n4637) );
  NOR2_X1 U5244 ( .A1(n7677), .A2(n4411), .ZN(n9438) );
  NAND2_X1 U5245 ( .A1(n9472), .A2(n9471), .ZN(n9475) );
  OR2_X1 U5246 ( .A1(n9475), .A2(n9474), .ZN(n4509) );
  NAND2_X1 U5247 ( .A1(n9140), .A2(n9139), .ZN(n9503) );
  NAND2_X1 U5248 ( .A1(n7846), .A2(n7845), .ZN(n9728) );
  NOR2_X1 U5249 ( .A1(n9728), .A2(n9520), .ZN(n9512) );
  NOR2_X1 U5250 ( .A1(n9545), .A2(n6298), .ZN(n9519) );
  NAND2_X1 U5251 ( .A1(n9358), .A2(n9359), .ZN(n9529) );
  NAND2_X1 U5252 ( .A1(n4386), .A2(n4699), .ZN(n4695) );
  AND2_X1 U5253 ( .A1(n4693), .A2(n9529), .ZN(n4692) );
  NAND2_X1 U5254 ( .A1(n4695), .A2(n4697), .ZN(n4693) );
  INV_X1 U5255 ( .A(n4695), .ZN(n4694) );
  NAND2_X1 U5256 ( .A1(n6291), .A2(n9537), .ZN(n6292) );
  AND2_X1 U5257 ( .A1(n9537), .A2(n9347), .ZN(n9553) );
  AND2_X1 U5258 ( .A1(n4709), .A2(n6261), .ZN(n4708) );
  NAND2_X1 U5259 ( .A1(n9606), .A2(n9626), .ZN(n4709) );
  AND2_X1 U5260 ( .A1(n9336), .A2(n9335), .ZN(n9586) );
  NAND2_X1 U5261 ( .A1(n9772), .A2(n9663), .ZN(n9621) );
  NAND2_X1 U5262 ( .A1(n9636), .A2(n6258), .ZN(n9620) );
  OR2_X1 U5263 ( .A1(n9772), .A2(n9401), .ZN(n6258) );
  AOI22_X1 U5264 ( .A1(n9165), .A2(n9667), .B1(n9664), .B2(n4786), .ZN(n9652)
         );
  OR2_X1 U5265 ( .A1(n6271), .A2(n6256), .ZN(n9674) );
  NAND2_X1 U5266 ( .A1(n9686), .A2(n4349), .ZN(n9675) );
  NAND2_X1 U5267 ( .A1(n9674), .A2(n9308), .ZN(n9684) );
  OR2_X1 U5268 ( .A1(n9708), .A2(n9707), .ZN(n9706) );
  OAI22_X1 U5269 ( .A1(n7811), .A2(n9298), .B1(n7817), .B2(n9702), .ZN(n9708)
         );
  OAI21_X1 U5270 ( .B1(n7689), .B2(n9160), .A(n6254), .ZN(n7720) );
  NAND2_X1 U5271 ( .A1(n4425), .A2(n9159), .ZN(n4670) );
  AOI22_X1 U5272 ( .A1(n7625), .A2(n7624), .B1(n9985), .B2(n9091), .ZN(n7689)
         );
  CLKBUF_X1 U5273 ( .A(n7622), .Z(n4425) );
  AOI22_X1 U5274 ( .A1(n7451), .A2(n9145), .B1(n9970), .B2(n7701), .ZN(n7571)
         );
  NAND2_X1 U5275 ( .A1(n4687), .A2(n4334), .ZN(n4686) );
  NAND2_X1 U5276 ( .A1(n7301), .A2(n7303), .ZN(n4688) );
  OAI211_X1 U5277 ( .C1(n6657), .C2(n5217), .A(n5065), .B(n5064), .ZN(n7240)
         );
  INV_X1 U5278 ( .A(n9835), .ZN(n9879) );
  NAND2_X1 U5279 ( .A1(n5220), .A2(n5219), .ZN(n9960) );
  NAND2_X1 U5280 ( .A1(n7968), .A2(n7967), .ZN(n7980) );
  OR2_X1 U5281 ( .A1(n7964), .A2(n7963), .ZN(n7968) );
  XNOR2_X1 U5282 ( .A(n7980), .B(n7979), .ZN(n9138) );
  NOR2_X1 U5283 ( .A1(n4963), .A2(n5288), .ZN(n4420) );
  INV_X1 U5284 ( .A(n4772), .ZN(n4771) );
  OAI21_X1 U5285 ( .B1(n4773), .B2(n5288), .A(n4966), .ZN(n4772) );
  NAND2_X1 U5286 ( .A1(n6112), .A2(n5679), .ZN(n7820) );
  OR2_X1 U5287 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  OAI21_X1 U5288 ( .B1(n5647), .B2(n4527), .A(n4525), .ZN(n5678) );
  XNOR2_X1 U5289 ( .A(n5671), .B(n5670), .ZN(n7802) );
  NAND2_X1 U5290 ( .A1(n5647), .A2(n5646), .ZN(n5671) );
  OAI21_X1 U5291 ( .B1(n5442), .B2(n4534), .A(n4531), .ZN(n5514) );
  NAND3_X1 U5292 ( .A1(n5445), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U5293 ( .A1(n4536), .A2(n4537), .ZN(n5493) );
  NAND2_X1 U5294 ( .A1(n5442), .A2(n4538), .ZN(n4536) );
  NAND2_X1 U5295 ( .A1(n4803), .A2(n4804), .ZN(n5315) );
  NAND2_X1 U5296 ( .A1(n5259), .A2(n4806), .ZN(n4803) );
  NAND2_X1 U5297 ( .A1(n5209), .A2(n5183), .ZN(n5210) );
  NAND2_X1 U5298 ( .A1(n5059), .A2(n4796), .ZN(n4795) );
  NOR2_X1 U5299 ( .A1(n4345), .A2(n4797), .ZN(n4796) );
  OAI21_X1 U5300 ( .B1(n5085), .B2(n4345), .A(n5110), .ZN(n4794) );
  AND2_X1 U5301 ( .A1(n5118), .A2(n5117), .ZN(n6720) );
  INV_X1 U5302 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4677) );
  INV_X1 U5303 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4678) );
  XNOR2_X1 U5304 ( .A(n7084), .B(n8390), .ZN(n7085) );
  AND4_X1 U5305 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n8251)
         );
  NAND2_X1 U5306 ( .A1(n6063), .A2(n6062), .ZN(n8268) );
  AND4_X1 U5307 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n7889)
         );
  INV_X1 U5308 ( .A(n8759), .ZN(n8735) );
  AOI211_X1 U5309 ( .C1(n8181), .C2(n7999), .A(n8028), .B(n7998), .ZN(n8032)
         );
  NAND2_X1 U5310 ( .A1(n4608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5784) );
  NAND4_X1 U5311 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n8385)
         );
  AND3_X1 U5312 ( .A1(n4745), .A2(n4744), .A3(n8510), .ZN(n8513) );
  INV_X1 U5313 ( .A(n6986), .ZN(n4847) );
  XNOR2_X1 U5314 ( .A(n4470), .B(n8502), .ZN(n4469) );
  NAND2_X1 U5315 ( .A1(n8500), .A2(n8499), .ZN(n4470) );
  NAND2_X1 U5316 ( .A1(n6131), .A2(n6130), .ZN(n8530) );
  INV_X1 U5317 ( .A(n4601), .ZN(n4600) );
  OAI21_X1 U5318 ( .B1(n4602), .B2(n10090), .A(n4603), .ZN(n4601) );
  OR2_X1 U5319 ( .A1(n10092), .A2(n4604), .ZN(n4603) );
  INV_X1 U5320 ( .A(n4467), .ZN(n4602) );
  NAND2_X1 U5321 ( .A1(n8024), .A2(n4569), .ZN(n4568) );
  OAI21_X1 U5322 ( .B1(n4576), .B2(n4361), .A(n4566), .ZN(n4565) );
  NAND2_X1 U5323 ( .A1(n5930), .A2(n5929), .ZN(n8841) );
  INV_X1 U5324 ( .A(n8530), .ZN(n8164) );
  INV_X1 U5325 ( .A(n9689), .ZN(n9664) );
  OR2_X1 U5326 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NAND2_X1 U5327 ( .A1(n6788), .A2(n6787), .ZN(n4884) );
  AOI21_X1 U5328 ( .B1(n5206), .B2(n9880), .A(n5125), .ZN(n7158) );
  NAND2_X1 U5329 ( .A1(n5550), .A2(n5549), .ZN(n9762) );
  INV_X1 U5330 ( .A(n9404), .ZN(n9091) );
  AND2_X2 U5331 ( .A1(n4357), .A2(n4491), .ZN(n9917) );
  NOR2_X1 U5332 ( .A1(n4910), .A2(n4350), .ZN(n4491) );
  AND2_X1 U5333 ( .A1(n5061), .A2(n9417), .ZN(n4910) );
  INV_X1 U5334 ( .A(n9574), .ZN(n9544) );
  NAND4_X1 U5335 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n9878)
         );
  NAND4_X2 U5336 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n6272)
         );
  OR2_X1 U5337 ( .A1(n5075), .A2(n7250), .ZN(n5006) );
  OR2_X1 U5338 ( .A1(n5738), .A2(n6629), .ZN(n5004) );
  OR2_X1 U5339 ( .A1(n6748), .A2(n6747), .ZN(n4513) );
  OR2_X1 U5340 ( .A1(n6737), .A2(n6736), .ZN(n4511) );
  AND2_X1 U5341 ( .A1(n4513), .A2(n4512), .ZN(n6737) );
  NAND2_X1 U5342 ( .A1(n6720), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4512) );
  NOR2_X1 U5343 ( .A1(n6758), .A2(n4401), .ZN(n6715) );
  NOR2_X1 U5344 ( .A1(n6715), .A2(n6714), .ZN(n6827) );
  INV_X1 U5345 ( .A(n5728), .ZN(n9496) );
  NAND2_X1 U5346 ( .A1(n4554), .A2(n4552), .ZN(n9724) );
  NOR2_X1 U5347 ( .A1(n5061), .A2(n4553), .ZN(n4552) );
  NAND2_X1 U5348 ( .A1(n9801), .A2(n9136), .ZN(n4554) );
  NOR2_X1 U5349 ( .A1(n9136), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U5350 ( .A1(n7869), .A2(n7868), .ZN(n9731) );
  NAND2_X1 U5351 ( .A1(n7856), .A2(n9876), .ZN(n7869) );
  NAND2_X1 U5352 ( .A1(n4505), .A2(n8059), .ZN(n4504) );
  NAND2_X1 U5353 ( .A1(n8050), .A2(n6148), .ZN(n4505) );
  INV_X1 U5354 ( .A(n9254), .ZN(n4498) );
  NAND2_X1 U5355 ( .A1(n4494), .A2(n9263), .ZN(n9269) );
  NOR2_X1 U5356 ( .A1(n4861), .A2(n8171), .ZN(n4860) );
  OR2_X1 U5357 ( .A1(n8094), .A2(n8185), .ZN(n4863) );
  OAI21_X1 U5358 ( .B1(n8102), .B2(n5939), .A(n4868), .ZN(n4867) );
  INV_X1 U5359 ( .A(n8104), .ZN(n4868) );
  AOI21_X1 U5360 ( .B1(n4347), .B2(n4488), .A(n4486), .ZN(n4485) );
  NAND2_X1 U5361 ( .A1(n4853), .A2(n4364), .ZN(n4849) );
  AOI21_X1 U5362 ( .B1(n4853), .B2(n8131), .A(n4852), .ZN(n4850) );
  NAND2_X1 U5363 ( .A1(n6077), .A2(n8139), .ZN(n4852) );
  AOI22_X1 U5364 ( .A1(n8175), .A2(n8165), .B1(n8164), .B2(n8185), .ZN(n8172)
         );
  OR2_X1 U5365 ( .A1(n8161), .A2(n8548), .ZN(n4909) );
  NAND2_X1 U5366 ( .A1(n9351), .A2(n9383), .ZN(n4478) );
  NAND2_X1 U5367 ( .A1(n8449), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4838) );
  NOR2_X1 U5368 ( .A1(n7942), .A2(n8168), .ZN(n4788) );
  NOR2_X1 U5369 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4597) );
  AND2_X1 U5370 ( .A1(n5756), .A2(n5755), .ZN(n4595) );
  AND2_X1 U5371 ( .A1(n4599), .A2(n4598), .ZN(n5966) );
  INV_X1 U5372 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4599) );
  INV_X1 U5373 ( .A(n7268), .ZN(n4635) );
  NOR2_X1 U5374 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  INV_X1 U5375 ( .A(n7593), .ZN(n4628) );
  OR2_X1 U5376 ( .A1(n9265), .A2(n9262), .ZN(n6281) );
  INV_X1 U5377 ( .A(n5513), .ZN(n4530) );
  INV_X1 U5378 ( .A(n4908), .ZN(n4544) );
  INV_X1 U5379 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4818) );
  INV_X1 U5380 ( .A(n5777), .ZN(n5769) );
  NAND2_X1 U5381 ( .A1(n4767), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5382 ( .A1(n4752), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4751) );
  NAND2_X1 U5383 ( .A1(n8430), .A2(n4838), .ZN(n4835) );
  OR2_X1 U5384 ( .A1(n4836), .A2(n8427), .ZN(n4834) );
  NAND2_X1 U5385 ( .A1(n4837), .A2(n4838), .ZN(n4836) );
  INV_X1 U5386 ( .A(n8428), .ZN(n4837) );
  AND2_X1 U5387 ( .A1(n8178), .A2(n8208), .ZN(n7942) );
  OR2_X1 U5388 ( .A1(n8383), .A2(n10056), .ZN(n8072) );
  INV_X1 U5389 ( .A(n8145), .ZN(n6171) );
  INV_X1 U5390 ( .A(n8001), .ZN(n8146) );
  AND2_X1 U5391 ( .A1(n6078), .A2(n8613), .ZN(n8589) );
  OR2_X1 U5392 ( .A1(n8615), .A2(n6077), .ZN(n8588) );
  OR2_X1 U5393 ( .A1(n8643), .A2(n8631), .ZN(n8615) );
  OR2_X1 U5394 ( .A1(n8631), .A2(n8630), .ZN(n8616) );
  NAND2_X1 U5395 ( .A1(n6163), .A2(n4813), .ZN(n6165) );
  NOR2_X1 U5396 ( .A1(n6160), .A2(n6161), .ZN(n4813) );
  INV_X1 U5397 ( .A(n8120), .ZN(n8124) );
  NAND2_X1 U5398 ( .A1(n4907), .A2(n5760), .ZN(n5761) );
  INV_X1 U5399 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5760) );
  INV_X1 U5400 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U5401 ( .A1(n5908), .A2(n5909), .ZN(n5921) );
  INV_X1 U5402 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4883) );
  AOI21_X1 U5403 ( .B1(n5206), .B2(n9413), .A(n4999), .ZN(n5002) );
  AND2_X1 U5404 ( .A1(n5501), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U5405 ( .A1(n4500), .A2(n9365), .ZN(n9366) );
  AND2_X1 U5406 ( .A1(n6289), .A2(n9319), .ZN(n9247) );
  NAND2_X1 U5407 ( .A1(n4674), .A2(n4676), .ZN(n4673) );
  OAI21_X1 U5408 ( .B1(n4349), .B2(n4675), .A(n9144), .ZN(n4674) );
  AND2_X1 U5409 ( .A1(n5472), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5501) );
  AND2_X1 U5410 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(n5449), .ZN(n5472) );
  NOR2_X1 U5411 ( .A1(n6271), .A2(n9719), .ZN(n4787) );
  AND2_X1 U5412 ( .A1(n4666), .A2(n4663), .ZN(n4662) );
  INV_X1 U5413 ( .A(n9299), .ZN(n4660) );
  NAND2_X1 U5414 ( .A1(n9991), .A2(n9977), .ZN(n4776) );
  AOI21_X1 U5415 ( .B1(n4658), .B2(n9160), .A(n4667), .ZN(n4666) );
  INV_X1 U5416 ( .A(n9288), .ZN(n4667) );
  NOR2_X1 U5417 ( .A1(n9159), .A2(n6285), .ZN(n4658) );
  AND2_X1 U5418 ( .A1(n9921), .A2(n9927), .ZN(n4778) );
  NAND2_X1 U5419 ( .A1(n5728), .A2(n9388), .ZN(n6265) );
  NAND2_X1 U5420 ( .A1(n9604), .A2(n4338), .ZN(n9545) );
  NAND2_X1 U5421 ( .A1(n9604), .A2(n9600), .ZN(n9593) );
  AND2_X1 U5422 ( .A1(n9716), .A2(n9819), .ZN(n9714) );
  NOR3_X1 U5423 ( .A1(n7581), .A2(n7631), .A3(n7586), .ZN(n7691) );
  NOR2_X1 U5424 ( .A1(n7581), .A2(n7586), .ZN(n7628) );
  NAND3_X1 U5425 ( .A1(n7239), .A2(n9933), .A3(n4336), .ZN(n9869) );
  NAND2_X1 U5426 ( .A1(n4517), .A2(n6128), .ZN(n7966) );
  AND2_X1 U5427 ( .A1(n4333), .A2(n4927), .ZN(n4712) );
  XNOR2_X1 U5428 ( .A(n7966), .B(n7965), .ZN(n7964) );
  NAND2_X1 U5429 ( .A1(n4963), .A2(n5288), .ZN(n4964) );
  NAND2_X1 U5430 ( .A1(n4943), .A2(n4900), .ZN(n4493) );
  INV_X1 U5431 ( .A(n4526), .ZN(n4525) );
  OAI21_X1 U5432 ( .B1(n4527), .B2(n5646), .A(n5672), .ZN(n4526) );
  NAND2_X1 U5433 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  INV_X1 U5434 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5705) );
  AOI21_X1 U5435 ( .B1(n4352), .B2(n4533), .A(n4532), .ZN(n4531) );
  INV_X1 U5436 ( .A(n5491), .ZN(n4532) );
  INV_X1 U5437 ( .A(n4538), .ZN(n4533) );
  INV_X1 U5438 ( .A(n4352), .ZN(n4534) );
  AOI21_X1 U5439 ( .B1(n5443), .B2(n4538), .A(n4382), .ZN(n4537) );
  AND2_X1 U5440 ( .A1(n4637), .A2(n4978), .ZN(n4636) );
  AOI21_X1 U5441 ( .B1(n4327), .B2(n4801), .A(n4378), .ZN(n4800) );
  INV_X1 U5442 ( .A(n4806), .ZN(n4801) );
  INV_X1 U5443 ( .A(n4327), .ZN(n4802) );
  NOR2_X1 U5444 ( .A1(n5286), .A2(n4807), .ZN(n4806) );
  INV_X1 U5445 ( .A(n5258), .ZN(n4807) );
  AOI21_X1 U5446 ( .B1(n4808), .B2(n4806), .A(n4805), .ZN(n4804) );
  INV_X1 U5447 ( .A(n5285), .ZN(n4805) );
  NAND2_X1 U5448 ( .A1(n4952), .A2(n4639), .ZN(n4638) );
  NOR2_X1 U5449 ( .A1(n4951), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5142) );
  INV_X1 U5450 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5089) );
  CLKBUF_X1 U5451 ( .A(n5062), .Z(n5063) );
  OAI21_X1 U5452 ( .B1(n5035), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n4959), .ZN(
        n5031) );
  NAND2_X1 U5453 ( .A1(n5035), .A2(n6647), .ZN(n4959) );
  INV_X1 U5454 ( .A(n8353), .ZN(n4719) );
  NAND2_X1 U5455 ( .A1(n4428), .A2(n5775), .ZN(n5914) );
  INV_X1 U5456 ( .A(n5902), .ZN(n4428) );
  AOI21_X1 U5457 ( .B1(n4328), .B2(n7913), .A(n4372), .ZN(n4742) );
  OR2_X1 U5458 ( .A1(n7665), .A2(n4354), .ZN(n7711) );
  AND2_X1 U5459 ( .A1(n7906), .A2(n7904), .ZN(n8284) );
  OR2_X1 U5460 ( .A1(n5914), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5916) );
  AOI21_X1 U5461 ( .B1(n4723), .B2(n4722), .A(n4406), .ZN(n4721) );
  INV_X1 U5462 ( .A(n7933), .ZN(n4722) );
  AND2_X1 U5463 ( .A1(n6981), .A2(n6980), .ZN(n8347) );
  AOI211_X1 U5464 ( .C1(n7997), .C2(n8175), .A(n7996), .B(n7995), .ZN(n7998)
         );
  AND2_X1 U5465 ( .A1(n6209), .A2(n8030), .ZN(n8031) );
  NAND2_X1 U5466 ( .A1(n7040), .A2(n7041), .ZN(n7039) );
  NAND2_X1 U5467 ( .A1(n4762), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4761) );
  NAND2_X1 U5468 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  INV_X1 U5469 ( .A(n6939), .ZN(n4763) );
  INV_X1 U5470 ( .A(n6575), .ZN(n4764) );
  NAND2_X1 U5471 ( .A1(n6575), .A2(n6939), .ZN(n7123) );
  OR2_X1 U5472 ( .A1(n6926), .A2(n6927), .ZN(n6924) );
  NAND2_X1 U5473 ( .A1(n4473), .A2(n7354), .ZN(n6608) );
  NAND2_X1 U5474 ( .A1(n4845), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4843) );
  OR2_X1 U5475 ( .A1(n6610), .A2(n7474), .ZN(n4845) );
  AND2_X1 U5476 ( .A1(n6610), .A2(n7474), .ZN(n6611) );
  AND2_X1 U5477 ( .A1(n4843), .A2(n4471), .ZN(n7548) );
  INV_X1 U5478 ( .A(n6611), .ZN(n4471) );
  AND2_X1 U5479 ( .A1(n4822), .A2(n4388), .ZN(n7741) );
  NOR2_X1 U5480 ( .A1(n7741), .A2(n7740), .ZN(n7739) );
  NOR2_X1 U5481 ( .A1(n6593), .A2(n7778), .ZN(n6595) );
  NOR2_X1 U5482 ( .A1(n8399), .A2(n8398), .ZN(n8420) );
  NAND2_X1 U5483 ( .A1(n5980), .A2(n5979), .ZN(n5992) );
  OAI21_X1 U5484 ( .B1(n8446), .B2(n8445), .A(n8444), .ZN(n8470) );
  OR2_X1 U5485 ( .A1(n8443), .A2(n8827), .ZN(n4749) );
  AND2_X1 U5486 ( .A1(n4834), .A2(n4832), .ZN(n8481) );
  NOR2_X1 U5487 ( .A1(n4833), .A2(n8468), .ZN(n4832) );
  INV_X1 U5488 ( .A(n4835), .ZN(n4833) );
  OR2_X1 U5489 ( .A1(n8443), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5490 ( .A1(n4747), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U5491 ( .A1(n8463), .A2(n4747), .ZN(n4744) );
  OR2_X1 U5492 ( .A1(n6116), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U5493 ( .A1(n6065), .A2(n6064), .ZN(n6088) );
  INV_X1 U5494 ( .A(n6066), .ZN(n6065) );
  NAND2_X1 U5495 ( .A1(n4433), .A2(n6035), .ZN(n6044) );
  INV_X1 U5496 ( .A(n4433), .ZN(n6036) );
  NAND2_X1 U5497 ( .A1(n6017), .A2(n6016), .ZN(n6027) );
  INV_X1 U5498 ( .A(n6018), .ZN(n6017) );
  NAND2_X1 U5499 ( .A1(n4432), .A2(n5984), .ZN(n5999) );
  NAND2_X1 U5500 ( .A1(n5956), .A2(n5955), .ZN(n5972) );
  INV_X1 U5501 ( .A(n5957), .ZN(n5956) );
  INV_X1 U5502 ( .A(n4432), .ZN(n5985) );
  NAND2_X1 U5503 ( .A1(n5932), .A2(n5931), .ZN(n5943) );
  INV_X1 U5504 ( .A(n5933), .ZN(n5932) );
  NAND2_X1 U5505 ( .A1(n4431), .A2(n7743), .ZN(n5933) );
  NAND2_X1 U5506 ( .A1(n4445), .A2(n4443), .ZN(n8753) );
  AOI21_X1 U5507 ( .B1(n4446), .B2(n4447), .A(n4444), .ZN(n4443) );
  INV_X1 U5508 ( .A(n8089), .ZN(n4444) );
  INV_X1 U5509 ( .A(n4590), .ZN(n4585) );
  NAND2_X1 U5510 ( .A1(n4591), .A2(n4590), .ZN(n4586) );
  INV_X1 U5511 ( .A(n4588), .ZN(n4587) );
  NAND2_X1 U5512 ( .A1(n5774), .A2(n5773), .ZN(n5890) );
  INV_X1 U5513 ( .A(n5888), .ZN(n5774) );
  NAND2_X1 U5514 ( .A1(n5875), .A2(n5874), .ZN(n7482) );
  AOI21_X1 U5515 ( .B1(n7336), .B2(n4437), .A(n4435), .ZN(n7481) );
  NOR2_X1 U5516 ( .A1(n7334), .A2(n6152), .ZN(n4437) );
  NOR2_X1 U5517 ( .A1(n8059), .A2(n6152), .ZN(n4435) );
  OR2_X1 U5518 ( .A1(n5876), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5888) );
  OR2_X1 U5519 ( .A1(n8387), .A2(n7875), .ZN(n7412) );
  NAND2_X1 U5520 ( .A1(n6928), .A2(n5770), .ZN(n5859) );
  INV_X1 U5521 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4604) );
  AOI21_X1 U5522 ( .B1(n4571), .B2(n4573), .A(n4383), .ZN(n4569) );
  INV_X1 U5523 ( .A(n4574), .ZN(n4573) );
  NAND2_X1 U5524 ( .A1(n4906), .A2(n6186), .ZN(n4467) );
  NAND2_X1 U5525 ( .A1(n6173), .A2(n8166), .ZN(n8548) );
  AND2_X1 U5526 ( .A1(n8155), .A2(n8154), .ZN(n8580) );
  OR2_X1 U5527 ( .A1(n6083), .A2(n8568), .ZN(n8572) );
  NAND2_X1 U5528 ( .A1(n4812), .A2(n4811), .ZN(n8586) );
  AND2_X1 U5529 ( .A1(n6171), .A2(n8143), .ZN(n4811) );
  NOR2_X1 U5530 ( .A1(n8148), .A2(n8146), .ZN(n8594) );
  OR2_X1 U5531 ( .A1(n6077), .A2(n6076), .ZN(n8613) );
  AND2_X1 U5532 ( .A1(n8618), .A2(n8616), .ZN(n6076) );
  INV_X1 U5533 ( .A(n8628), .ZN(n8631) );
  OAI21_X1 U5534 ( .B1(n8640), .B2(n6168), .A(n8133), .ZN(n8629) );
  AND4_X1 U5535 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n8646)
         );
  AND2_X1 U5536 ( .A1(n8132), .A2(n8133), .ZN(n8643) );
  OR2_X1 U5537 ( .A1(n8003), .A2(n6159), .ZN(n8658) );
  AND4_X1 U5538 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n8698)
         );
  AOI21_X1 U5539 ( .B1(n4452), .B2(n4453), .A(n4451), .ZN(n4450) );
  NOR2_X1 U5540 ( .A1(n8730), .A2(n8105), .ZN(n7878) );
  INV_X1 U5541 ( .A(n7635), .ZN(n10051) );
  INV_X1 U5542 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6192) );
  INV_X1 U5543 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6194) );
  INV_X1 U5544 ( .A(n4882), .ZN(n4881) );
  AND2_X1 U5545 ( .A1(n4882), .A2(n5758), .ZN(n4880) );
  INV_X1 U5546 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5909) );
  INV_X1 U5547 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5802) );
  INV_X1 U5548 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5867) );
  NOR2_X1 U5549 ( .A1(n5850), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U5550 ( .A1(n4877), .A2(n4440), .ZN(n5850) );
  AND2_X1 U5551 ( .A1(n5829), .A2(n5753), .ZN(n4877) );
  INV_X1 U5552 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5753) );
  XNOR2_X1 U5553 ( .A(n5068), .B(n6482), .ZN(n5070) );
  AND2_X1 U5554 ( .A1(n5669), .A2(n5668), .ZN(n5701) );
  AND2_X1 U5555 ( .A1(n5312), .A2(n5310), .ZN(n9013) );
  NAND2_X1 U5556 ( .A1(n5398), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5429) );
  NOR2_X1 U5557 ( .A1(n8978), .A2(n5587), .ZN(n4621) );
  INV_X1 U5558 ( .A(n7077), .ZN(n4632) );
  AND2_X1 U5559 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5105) );
  NAND2_X1 U5560 ( .A1(n9015), .A2(n5312), .ZN(n9065) );
  AND2_X1 U5561 ( .A1(n9012), .A2(n5283), .ZN(n9086) );
  NAND2_X1 U5562 ( .A1(n5253), .A2(n5252), .ZN(n9085) );
  NOR2_X1 U5563 ( .A1(n5429), .A2(n9045), .ZN(n5449) );
  NAND2_X1 U5564 ( .A1(n5105), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5133) );
  NOR2_X1 U5565 ( .A1(n5643), .A2(n5642), .ZN(n9110) );
  AND2_X1 U5566 ( .A1(n4885), .A2(n5380), .ZN(n4640) );
  NAND2_X1 U5567 ( .A1(n9366), .A2(n4499), .ZN(n9367) );
  AND2_X1 U5568 ( .A1(n9503), .A2(n9396), .ZN(n4499) );
  OR2_X1 U5569 ( .A1(n9444), .A2(n9443), .ZN(n9456) );
  AND2_X1 U5570 ( .A1(n9456), .A2(n9455), .ZN(n9458) );
  NAND2_X1 U5571 ( .A1(n4509), .A2(n4418), .ZN(n9483) );
  NAND2_X1 U5572 ( .A1(n9354), .A2(n9182), .ZN(n9356) );
  INV_X1 U5573 ( .A(n9397), .ZN(n9543) );
  NAND2_X1 U5574 ( .A1(n9349), .A2(n9180), .ZN(n9541) );
  INV_X1 U5575 ( .A(n9398), .ZN(n9564) );
  NAND2_X1 U5576 ( .A1(n9604), .A2(n4781), .ZN(n9555) );
  NOR2_X1 U5577 ( .A1(n9588), .A2(n4643), .ZN(n9577) );
  NAND2_X1 U5578 ( .A1(n4644), .A2(n9335), .ZN(n4643) );
  AOI21_X1 U5579 ( .B1(n4706), .B2(n6263), .A(n4374), .ZN(n4705) );
  NAND2_X1 U5580 ( .A1(n9611), .A2(n9142), .ZN(n9589) );
  AND2_X1 U5581 ( .A1(n9644), .A2(n9633), .ZN(n9627) );
  AND2_X1 U5582 ( .A1(n9627), .A2(n9606), .ZN(n9604) );
  NAND2_X1 U5583 ( .A1(n4672), .A2(n4673), .ZN(n9641) );
  AOI22_X1 U5584 ( .A1(n9652), .A2(n6257), .B1(n9777), .B2(n9678), .ZN(n9637)
         );
  NAND2_X1 U5585 ( .A1(n9321), .A2(n9621), .ZN(n9640) );
  NAND2_X1 U5586 ( .A1(n9637), .A2(n9640), .ZN(n9636) );
  NAND2_X1 U5587 ( .A1(n9716), .A2(n4785), .ZN(n9653) );
  AND2_X1 U5588 ( .A1(n4331), .A2(n9655), .ZN(n4785) );
  NAND2_X1 U5589 ( .A1(n9716), .A2(n4787), .ZN(n9693) );
  NAND2_X1 U5590 ( .A1(n9716), .A2(n4331), .ZN(n9668) );
  NAND2_X1 U5591 ( .A1(n4711), .A2(n4710), .ZN(n9667) );
  AOI21_X1 U5592 ( .B1(n4326), .B2(n9707), .A(n4380), .ZN(n4710) );
  AND2_X1 U5593 ( .A1(n5369), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5398) );
  NOR2_X1 U5594 ( .A1(n5342), .A2(n5341), .ZN(n5369) );
  AOI22_X1 U5595 ( .A1(n7720), .A2(n9162), .B1(n9997), .B2(n9127), .ZN(n7811)
         );
  AND2_X1 U5596 ( .A1(n9300), .A2(n9301), .ZN(n9298) );
  NAND2_X1 U5597 ( .A1(n4664), .A2(n4666), .ZN(n7721) );
  NAND2_X1 U5598 ( .A1(n4665), .A2(n4669), .ZN(n4664) );
  OR2_X1 U5599 ( .A1(n5321), .A2(n5320), .ZN(n5342) );
  OR2_X1 U5600 ( .A1(n7586), .A2(n9405), .ZN(n6253) );
  NAND2_X1 U5601 ( .A1(n5269), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5296) );
  NOR2_X1 U5602 ( .A1(n7572), .A2(n7573), .ZN(n6284) );
  NAND2_X1 U5603 ( .A1(n5240), .A2(n5239), .ZN(n7459) );
  OR2_X1 U5604 ( .A1(n7455), .A2(n7459), .ZN(n7581) );
  AOI21_X1 U5605 ( .B1(n4323), .B2(n4684), .A(n4381), .ZN(n4683) );
  NOR2_X1 U5606 ( .A1(n5221), .A2(n6824), .ZN(n5241) );
  OR2_X1 U5607 ( .A1(n5193), .A2(n5192), .ZN(n5221) );
  NOR2_X1 U5608 ( .A1(n9852), .A2(n7590), .ZN(n9853) );
  AOI21_X1 U5609 ( .B1(n9151), .B2(n4702), .A(n4373), .ZN(n4700) );
  OAI21_X1 U5610 ( .B1(n4650), .B2(n9206), .A(n4648), .ZN(n4646) );
  AND2_X1 U5611 ( .A1(n7227), .A2(n9917), .ZN(n7239) );
  NAND2_X1 U5612 ( .A1(n7239), .A2(n9921), .ZN(n9888) );
  XNOR2_X1 U5613 ( .A(n9917), .B(n9411), .ZN(n9147) );
  CLKBUF_X1 U5614 ( .A(n6242), .Z(n9900) );
  AND2_X1 U5615 ( .A1(n9728), .A2(n9959), .ZN(n9729) );
  NAND2_X1 U5616 ( .A1(n5681), .A2(n5680), .ZN(n6298) );
  NAND2_X1 U5617 ( .A1(n7820), .A2(n9137), .ZN(n5681) );
  NAND2_X1 U5618 ( .A1(n7802), .A2(n9137), .ZN(n5652) );
  NAND2_X1 U5619 ( .A1(n5602), .A2(n5601), .ZN(n9752) );
  NAND2_X1 U5620 ( .A1(n5518), .A2(n5517), .ZN(n9767) );
  NAND2_X1 U5621 ( .A1(n5499), .A2(n5498), .ZN(n9772) );
  INV_X1 U5622 ( .A(n7252), .ZN(n6943) );
  INV_X1 U5623 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4931) );
  XNOR2_X1 U5624 ( .A(n6125), .B(n6124), .ZN(n7827) );
  NAND2_X1 U5625 ( .A1(n4770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U5626 ( .A1(n4945), .A2(n4773), .ZN(n4770) );
  INV_X1 U5627 ( .A(n4982), .ZN(n4922) );
  INV_X1 U5628 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5392) );
  OAI21_X1 U5629 ( .B1(n5259), .B2(n4808), .A(n5258), .ZN(n5287) );
  OAI21_X1 U5630 ( .B1(n5176), .B2(n4548), .A(n4545), .ZN(n5235) );
  AOI21_X1 U5631 ( .B1(n5139), .B2(n4520), .A(n4377), .ZN(n4519) );
  XNOR2_X1 U5632 ( .A(n5157), .B(SI_6_), .ZN(n5155) );
  XNOR2_X1 U5633 ( .A(n5112), .B(SI_4_), .ZN(n5110) );
  XNOR2_X1 U5634 ( .A(n5031), .B(SI_1_), .ZN(n5030) );
  XNOR2_X1 U5635 ( .A(n4968), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6723) );
  AND2_X1 U5636 ( .A1(n5942), .A2(n5941), .ZN(n8222) );
  INV_X1 U5637 ( .A(n8786), .ZN(n10067) );
  NAND2_X1 U5638 ( .A1(n7109), .A2(n7110), .ZN(n7279) );
  NAND2_X1 U5639 ( .A1(n4741), .A2(n4742), .ZN(n8240) );
  NAND2_X1 U5640 ( .A1(n8271), .A2(n7913), .ZN(n4741) );
  NAND2_X1 U5641 ( .A1(n7711), .A2(n7710), .ZN(n7769) );
  AOI21_X1 U5642 ( .B1(n4732), .B2(n4736), .A(n4404), .ZN(n4731) );
  AND4_X1 U5643 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n8779)
         );
  INV_X1 U5644 ( .A(n4716), .ZN(n4714) );
  NAND2_X1 U5645 ( .A1(n7279), .A2(n4717), .ZN(n7281) );
  NAND2_X1 U5646 ( .A1(n4729), .A2(n4727), .ZN(n7888) );
  OAI21_X1 U5647 ( .B1(n8271), .B2(n4740), .A(n4736), .ZN(n8307) );
  INV_X1 U5648 ( .A(n8322), .ZN(n7924) );
  AND2_X1 U5649 ( .A1(n5998), .A2(n5997), .ZN(n8352) );
  AND4_X1 U5650 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n8645)
         );
  OAI21_X1 U5651 ( .B1(n8271), .B2(n4328), .A(n7913), .ZN(n8343) );
  OAI21_X1 U5652 ( .B1(n8223), .B2(n4724), .A(n4721), .ZN(n8356) );
  INV_X1 U5653 ( .A(n8362), .ZN(n8378) );
  AND4_X1 U5654 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n8734)
         );
  NAND2_X1 U5655 ( .A1(n6094), .A2(n6093), .ZN(n8550) );
  OAI211_X1 U5656 ( .C1(n6181), .C2(n6061), .A(n6060), .B(n6059), .ZN(n8606)
         );
  OAI211_X1 U5657 ( .C1(n6054), .C2(n8810), .A(n6053), .B(n6052), .ZN(n8622)
         );
  INV_X1 U5658 ( .A(n8645), .ZN(n8676) );
  INV_X1 U5659 ( .A(n7889), .ZN(n8762) );
  NAND2_X1 U5660 ( .A1(n5858), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4563) );
  XNOR2_X1 U5661 ( .A(n6519), .B(n4434), .ZN(n7036) );
  NAND2_X1 U5662 ( .A1(n4760), .A2(n7123), .ZN(n7125) );
  INV_X1 U5663 ( .A(n4761), .ZN(n4760) );
  NAND2_X1 U5664 ( .A1(n4828), .A2(n4825), .ZN(n7064) );
  NAND2_X1 U5665 ( .A1(n4767), .A2(n7185), .ZN(n7067) );
  AOI21_X1 U5666 ( .B1(n6521), .B2(n7118), .A(n7132), .ZN(n7062) );
  NAND2_X1 U5667 ( .A1(n4474), .A2(n7354), .ZN(n7328) );
  NAND2_X1 U5668 ( .A1(n4752), .A2(n7367), .ZN(n7324) );
  AOI21_X1 U5669 ( .B1(n7363), .B2(n7362), .A(n7361), .ZN(n7468) );
  NAND2_X1 U5670 ( .A1(n4472), .A2(n7354), .ZN(n7359) );
  INV_X1 U5671 ( .A(n4473), .ZN(n4472) );
  NAND2_X1 U5672 ( .A1(n4758), .A2(n4756), .ZN(n7472) );
  NOR2_X1 U5673 ( .A1(n4757), .A2(n6587), .ZN(n7471) );
  NOR2_X1 U5674 ( .A1(n4843), .A2(n6611), .ZN(n7464) );
  OR2_X1 U5675 ( .A1(n4844), .A2(n6611), .ZN(n7465) );
  INV_X1 U5676 ( .A(n4845), .ZN(n4844) );
  INV_X1 U5677 ( .A(n4822), .ZN(n7654) );
  AOI21_X1 U5678 ( .B1(n7737), .B2(n7736), .A(n7735), .ZN(n7783) );
  NOR2_X1 U5679 ( .A1(n6591), .A2(n7647), .ZN(n7734) );
  NAND2_X1 U5680 ( .A1(n4840), .A2(n4839), .ZN(n8401) );
  NOR2_X1 U5681 ( .A1(n8416), .A2(n8415), .ZN(n8418) );
  NOR2_X1 U5682 ( .A1(n8427), .A2(n8428), .ZN(n8431) );
  NAND2_X1 U5683 ( .A1(n4570), .A2(n4574), .ZN(n8536) );
  NAND2_X1 U5684 ( .A1(n6026), .A2(n6025), .ZN(n8650) );
  OAI21_X1 U5685 ( .B1(n6156), .B2(n4453), .A(n4452), .ZN(n8712) );
  NAND2_X1 U5686 ( .A1(n4442), .A2(n4446), .ZN(n8772) );
  OR2_X1 U5687 ( .A1(n7611), .A2(n4447), .ZN(n4442) );
  INV_X1 U5688 ( .A(n10061), .ZN(n7775) );
  NAND2_X1 U5689 ( .A1(n7612), .A2(n4591), .ZN(n7755) );
  AND2_X1 U5690 ( .A1(n4581), .A2(n4584), .ZN(n7562) );
  INV_X1 U5691 ( .A(n8782), .ZN(n10033) );
  INV_X1 U5692 ( .A(n8715), .ZN(n10031) );
  NAND2_X1 U5693 ( .A1(n7977), .A2(n7976), .ZN(n8791) );
  INV_X1 U5694 ( .A(n7346), .ZN(n7212) );
  INV_X1 U5695 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4464) );
  OAI21_X1 U5696 ( .B1(n4467), .B2(n4466), .A(n10078), .ZN(n4465) );
  INV_X1 U5697 ( .A(n6187), .ZN(n4466) );
  NAND2_X1 U5698 ( .A1(n8547), .A2(n8166), .ZN(n4790) );
  NAND2_X1 U5699 ( .A1(n6101), .A2(n6100), .ZN(n8861) );
  NAND2_X1 U5700 ( .A1(n6087), .A2(n6086), .ZN(n8867) );
  NAND2_X1 U5701 ( .A1(n4810), .A2(n8154), .ZN(n8557) );
  INV_X1 U5702 ( .A(n8268), .ZN(n8872) );
  NAND2_X1 U5703 ( .A1(n6056), .A2(n6055), .ZN(n8878) );
  NAND2_X1 U5704 ( .A1(n6049), .A2(n6048), .ZN(n8884) );
  NAND2_X1 U5705 ( .A1(n4812), .A2(n8143), .ZN(n8603) );
  NAND2_X1 U5706 ( .A1(n6043), .A2(n6042), .ZN(n8890) );
  NAND2_X1 U5707 ( .A1(n6034), .A2(n6033), .ZN(n8896) );
  NAND2_X1 U5708 ( .A1(n6015), .A2(n6014), .ZN(n8907) );
  INV_X1 U5709 ( .A(n8352), .ZN(n8913) );
  NAND2_X1 U5710 ( .A1(n5983), .A2(n5982), .ZN(n8919) );
  AND2_X1 U5711 ( .A1(n8689), .A2(n8688), .ZN(n8917) );
  NAND2_X1 U5712 ( .A1(n5971), .A2(n5970), .ZN(n8925) );
  INV_X1 U5713 ( .A(n7901), .ZN(n8932) );
  INV_X1 U5714 ( .A(n8222), .ZN(n8722) );
  NAND2_X1 U5715 ( .A1(n4454), .A2(n6157), .ZN(n7877) );
  NAND2_X1 U5716 ( .A1(n6156), .A2(n4457), .ZN(n4454) );
  NAND2_X1 U5717 ( .A1(n6156), .A2(n8095), .ZN(n8729) );
  NAND2_X1 U5718 ( .A1(n5789), .A2(n5788), .ZN(n8941) );
  INV_X1 U5719 ( .A(n8934), .ZN(n8942) );
  AND3_X1 U5720 ( .A1(n5900), .A2(n5899), .A3(n5898), .ZN(n8073) );
  INV_X1 U5721 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U5722 ( .A1(n4743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U5723 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4477) );
  NAND2_X1 U5724 ( .A1(n5340), .A2(n5339), .ZN(n8968) );
  CLKBUF_X1 U5725 ( .A(n6954), .Z(n6955) );
  INV_X1 U5726 ( .A(n4631), .ZN(n4630) );
  INV_X1 U5727 ( .A(n9399), .ZN(n9592) );
  NAND2_X1 U5728 ( .A1(n4894), .A2(n4892), .ZN(n4891) );
  NAND2_X1 U5729 ( .A1(n7796), .A2(n9137), .ZN(n5628) );
  INV_X1 U5730 ( .A(n4614), .ZN(n4613) );
  INV_X1 U5731 ( .A(n9406), .ZN(n7701) );
  OR2_X1 U5732 ( .A1(n5733), .A2(n7828), .ZN(n9115) );
  AND2_X1 U5733 ( .A1(n5130), .A2(n7157), .ZN(n7266) );
  NAND2_X1 U5734 ( .A1(n9196), .A2(n9374), .ZN(n4556) );
  AOI21_X1 U5735 ( .B1(n9193), .B2(n4558), .A(n9387), .ZN(n4557) );
  AOI21_X1 U5736 ( .B1(n9195), .B2(n9194), .A(n4559), .ZN(n4558) );
  NAND2_X1 U5737 ( .A1(n9384), .A2(n9192), .ZN(n4559) );
  INV_X1 U5738 ( .A(n9376), .ZN(n9388) );
  AND4_X1 U5739 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n7866)
         );
  NAND4_X1 U5740 ( .A1(n5138), .A2(n5137), .A3(n5136), .A4(n5135), .ZN(n9409)
         );
  OR2_X1 U5741 ( .A1(n4320), .A2(n9862), .ZN(n5136) );
  OR2_X1 U5742 ( .A1(n5075), .A2(n5131), .ZN(n5137) );
  AND2_X1 U5743 ( .A1(n4511), .A2(n4510), .ZN(n6760) );
  NAND2_X1 U5744 ( .A1(n6718), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4510) );
  NOR2_X1 U5745 ( .A1(n6827), .A2(n4402), .ZN(n6831) );
  NAND2_X1 U5746 ( .A1(n6831), .A2(n6830), .ZN(n6839) );
  OAI21_X1 U5747 ( .B1(n6842), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6839), .ZN(
        n6840) );
  NOR2_X1 U5748 ( .A1(n6908), .A2(n4516), .ZN(n6912) );
  AND2_X1 U5749 ( .A1(n6909), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4516) );
  NOR2_X1 U5750 ( .A1(n6912), .A2(n6911), .ZN(n7148) );
  NOR2_X1 U5751 ( .A1(n7148), .A2(n4515), .ZN(n7152) );
  AND2_X1 U5752 ( .A1(n7149), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5753 ( .A1(n7152), .A2(n7151), .ZN(n7169) );
  OAI21_X1 U5754 ( .B1(n7170), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7169), .ZN(
        n7171) );
  NOR2_X1 U5755 ( .A1(n7402), .A2(n4514), .ZN(n7406) );
  AND2_X1 U5756 ( .A1(n7403), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U5757 ( .A1(n7406), .A2(n7405), .ZN(n7677) );
  AND2_X1 U5758 ( .A1(n4975), .A2(n4637), .ZN(n5336) );
  XNOR2_X1 U5759 ( .A(n9438), .B(n9437), .ZN(n7679) );
  INV_X1 U5760 ( .A(n4509), .ZN(n9482) );
  INV_X1 U5761 ( .A(n9503), .ZN(n9727) );
  XNOR2_X1 U5762 ( .A(n7847), .B(n9362), .ZN(n9733) );
  NAND2_X1 U5763 ( .A1(n4690), .A2(n4689), .ZN(n7847) );
  AOI21_X1 U5764 ( .B1(n4692), .B2(n4694), .A(n4384), .ZN(n4689) );
  OAI21_X1 U5765 ( .B1(n9536), .B2(n4694), .A(n4692), .ZN(n9517) );
  NAND2_X1 U5766 ( .A1(n4691), .A2(n4695), .ZN(n9518) );
  INV_X1 U5767 ( .A(n6298), .ZN(n7958) );
  AOI21_X1 U5768 ( .B1(n6262), .B2(n4708), .A(n6263), .ZN(n9587) );
  NAND2_X1 U5769 ( .A1(n6262), .A2(n6261), .ZN(n9603) );
  NAND2_X1 U5770 ( .A1(n9675), .A2(n9312), .ZN(n9661) );
  NAND2_X1 U5771 ( .A1(n9706), .A2(n4326), .ZN(n9683) );
  AND2_X1 U5772 ( .A1(n9706), .A2(n6255), .ZN(n9685) );
  NAND2_X1 U5773 ( .A1(n5368), .A2(n5367), .ZN(n7817) );
  NAND2_X1 U5774 ( .A1(n4670), .A2(n4669), .ZN(n7687) );
  NAND2_X1 U5775 ( .A1(n5319), .A2(n5318), .ZN(n7694) );
  NAND2_X1 U5776 ( .A1(n4685), .A2(n4686), .ZN(n7424) );
  NAND2_X1 U5777 ( .A1(n4688), .A2(n4348), .ZN(n4685) );
  OR2_X1 U5778 ( .A1(n4321), .A2(n7238), .ZN(n9709) );
  NAND2_X1 U5779 ( .A1(n4688), .A2(n6252), .ZN(n9832) );
  NAND2_X1 U5780 ( .A1(n4703), .A2(n6249), .ZN(n7257) );
  OR2_X1 U5781 ( .A1(n4321), .A2(n7228), .ZN(n9884) );
  NAND2_X1 U5782 ( .A1(n4651), .A2(n9207), .ZN(n9874) );
  NAND2_X1 U5783 ( .A1(n6277), .A2(n6276), .ZN(n7233) );
  INV_X1 U5784 ( .A(n9897), .ZN(n9710) );
  INV_X1 U5785 ( .A(n9884), .ZN(n9901) );
  INV_X1 U5786 ( .A(n10019), .ZN(n10017) );
  NAND2_X1 U5787 ( .A1(n4423), .A2(n4421), .ZN(n9787) );
  INV_X1 U5788 ( .A(n4422), .ZN(n4421) );
  INV_X1 U5789 ( .A(n9731), .ZN(n4423) );
  OAI21_X1 U5790 ( .B1(n9733), .B2(n9963), .A(n9732), .ZN(n4422) );
  NOR2_X1 U5791 ( .A1(n10004), .A2(n6305), .ZN(n6306) );
  XNOR2_X1 U5792 ( .A(n4555), .B(n7982), .ZN(n9801) );
  OAI21_X1 U5793 ( .B1(n7980), .B2(n7979), .A(n7978), .ZN(n4555) );
  NAND2_X1 U5794 ( .A1(n9798), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4930) );
  OR2_X1 U5795 ( .A1(n4771), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U5796 ( .A1(n4551), .A2(n5179), .ZN(n5211) );
  NAND2_X1 U5797 ( .A1(n5176), .A2(n5175), .ZN(n4551) );
  INV_X1 U5798 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U5799 ( .A1(n4521), .A2(n5114), .ZN(n5140) );
  NAND2_X1 U5800 ( .A1(n4795), .A2(n4793), .ZN(n4521) );
  INV_X1 U5801 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U5802 ( .A1(n5059), .A2(n5058), .ZN(n5086) );
  XNOR2_X1 U5803 ( .A(n5028), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U5804 ( .A1(n4678), .A2(n4677), .ZN(n4679) );
  AOI211_X1 U5805 ( .C1(n8488), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8487), .B(
        n8486), .ZN(n8489) );
  NAND2_X1 U5806 ( .A1(n4821), .A2(n8514), .ZN(n4820) );
  NAND2_X1 U5807 ( .A1(n4469), .A2(n8509), .ZN(n4468) );
  OAI21_X1 U5808 ( .B1(n6187), .B2(n10090), .A(n4600), .ZN(n6231) );
  NAND2_X1 U5809 ( .A1(n4884), .A2(n5019), .ZN(n6855) );
  INV_X1 U5810 ( .A(n4513), .ZN(n6746) );
  INV_X1 U5811 ( .A(n4511), .ZN(n6735) );
  AND2_X1 U5812 ( .A1(n9289), .A2(n9288), .ZN(n9160) );
  AND2_X1 U5813 ( .A1(n4686), .A2(n4409), .ZN(n4323) );
  AND2_X1 U5814 ( .A1(n4926), .A2(n4367), .ZN(n4324) );
  AND3_X1 U5815 ( .A1(n5743), .A2(n9380), .A3(n5731), .ZN(n9113) );
  AND2_X1 U5816 ( .A1(n9684), .A2(n6255), .ZN(n4326) );
  NAND2_X1 U5817 ( .A1(n4925), .A2(n4924), .ZN(n4956) );
  AND2_X1 U5818 ( .A1(n4804), .A2(n5313), .ZN(n4327) );
  OR2_X1 U5819 ( .A1(n8287), .A2(n8342), .ZN(n4328) );
  OAI211_X1 U5820 ( .C1(n6651), .C2(n5217), .A(n5094), .B(n5093), .ZN(n7079)
         );
  NAND2_X1 U5821 ( .A1(n4759), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4329) );
  AND3_X1 U5822 ( .A1(n4925), .A2(n4924), .A3(n4492), .ZN(n4943) );
  AND2_X1 U5823 ( .A1(n7710), .A2(n4358), .ZN(n4330) );
  AND2_X1 U5824 ( .A1(n4787), .A2(n4786), .ZN(n4331) );
  AND3_X1 U5825 ( .A1(n9302), .A2(n9383), .A3(n9301), .ZN(n4332) );
  AND2_X1 U5826 ( .A1(n4900), .A2(n4963), .ZN(n4333) );
  OR2_X1 U5827 ( .A1(n7590), .A2(n9408), .ZN(n4334) );
  AND2_X1 U5828 ( .A1(n4897), .A2(n5593), .ZN(n4335) );
  AND3_X1 U5829 ( .A1(n9927), .A2(n9921), .A3(n9939), .ZN(n4336) );
  AND4_X1 U5830 ( .A1(n4981), .A2(n4979), .A3(n5392), .A4(n4978), .ZN(n4337)
         );
  OR2_X1 U5831 ( .A1(n8867), .A2(n8576), .ZN(n8000) );
  NAND2_X1 U5832 ( .A1(n9340), .A2(n9341), .ZN(n9571) );
  INV_X1 U5833 ( .A(n9571), .ZN(n4644) );
  OR2_X1 U5834 ( .A1(n8769), .A2(n8779), .ZN(n8093) );
  INV_X1 U5835 ( .A(n8093), .ZN(n4861) );
  NAND2_X1 U5836 ( .A1(n5428), .A2(n5427), .ZN(n6271) );
  AND2_X1 U5837 ( .A1(n4781), .A2(n4780), .ZN(n4338) );
  NAND2_X1 U5838 ( .A1(n4655), .A2(n4929), .ZN(n4339) );
  AND2_X1 U5839 ( .A1(n4465), .A2(n4410), .ZN(n4340) );
  OR2_X1 U5840 ( .A1(n5592), .A2(n9052), .ZN(n4341) );
  OR2_X1 U5841 ( .A1(n8518), .A2(n8517), .ZN(n4342) );
  INV_X1 U5842 ( .A(n8383), .ZN(n7768) );
  INV_X1 U5843 ( .A(n9312), .ZN(n4675) );
  AND2_X1 U5844 ( .A1(n4333), .A2(n4362), .ZN(n4343) );
  AND2_X1 U5845 ( .A1(n9051), .A2(n4625), .ZN(n4344) );
  NAND2_X1 U5846 ( .A1(n6955), .A2(n5073), .ZN(n7074) );
  INV_X1 U5847 ( .A(n8465), .ZN(n4747) );
  INV_X1 U5848 ( .A(n4846), .ZN(n8493) );
  AND2_X1 U5849 ( .A1(n5088), .A2(SI_3_), .ZN(n4345) );
  NAND2_X1 U5850 ( .A1(n5448), .A2(n5447), .ZN(n9781) );
  INV_X1 U5851 ( .A(n5858), .ZN(n5790) );
  OR2_X1 U5852 ( .A1(n6618), .A2(n6617), .ZN(n4346) );
  NAND2_X1 U5853 ( .A1(n5421), .A2(n5420), .ZN(n5442) );
  NAND2_X1 U5854 ( .A1(n6112), .A2(n6111), .ZN(n6125) );
  OR2_X1 U5855 ( .A1(n7631), .A2(n9091), .ZN(n9283) );
  NAND2_X1 U5856 ( .A1(n9058), .A2(n9059), .ZN(n9002) );
  AND2_X1 U5857 ( .A1(n9307), .A2(n4487), .ZN(n4347) );
  OR2_X1 U5858 ( .A1(n9878), .A2(n9921), .ZN(n6278) );
  INV_X1 U5859 ( .A(n4724), .ZN(n4723) );
  NAND2_X1 U5860 ( .A1(n8264), .A2(n4725), .ZN(n4724) );
  AND2_X1 U5861 ( .A1(n6252), .A2(n4334), .ZN(n4348) );
  INV_X1 U5862 ( .A(n6173), .ZN(n8167) );
  OR2_X1 U5863 ( .A1(n8861), .A2(n8537), .ZN(n6173) );
  AND2_X1 U5864 ( .A1(n9676), .A2(n9674), .ZN(n4349) );
  NAND2_X1 U5865 ( .A1(n4742), .A2(n4412), .ZN(n4740) );
  AND2_X1 U5866 ( .A1(n4322), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4350) );
  OR2_X1 U5867 ( .A1(n8861), .A2(n8560), .ZN(n4351) );
  AND2_X1 U5868 ( .A1(n4537), .A2(n4535), .ZN(n4352) );
  XNOR2_X1 U5869 ( .A(n5256), .B(SI_10_), .ZN(n5255) );
  INV_X1 U5870 ( .A(n9735), .ZN(n9526) );
  NAND2_X1 U5871 ( .A1(n6479), .A2(n6478), .ZN(n9735) );
  AND2_X1 U5872 ( .A1(n4351), .A2(n6097), .ZN(n4353) );
  OR2_X1 U5873 ( .A1(n4730), .A2(n4911), .ZN(n4354) );
  OAI211_X1 U5874 ( .C1(n6661), .C2(n5217), .A(n5120), .B(n5119), .ZN(n7261)
         );
  NAND2_X1 U5875 ( .A1(n4938), .A2(n4936), .ZN(n5049) );
  OR2_X1 U5876 ( .A1(n7292), .A2(n7293), .ZN(n4355) );
  AND2_X1 U5877 ( .A1(n8385), .A2(n7635), .ZN(n4356) );
  XNOR2_X1 U5878 ( .A(n7964), .B(SI_29_), .ZN(n7844) );
  OR2_X1 U5879 ( .A1(n5217), .A2(n6655), .ZN(n4357) );
  OR2_X1 U5880 ( .A1(n7766), .A2(n8383), .ZN(n4358) );
  INV_X1 U5881 ( .A(n4824), .ZN(n4828) );
  AND2_X1 U5882 ( .A1(n4673), .A2(n4671), .ZN(n4359) );
  OR2_X1 U5883 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4360) );
  NAND2_X1 U5884 ( .A1(n5866), .A2(n5867), .ZN(n5882) );
  AND2_X1 U5885 ( .A1(n4569), .A2(n4567), .ZN(n4361) );
  NAND2_X1 U5886 ( .A1(n4975), .A2(n4920), .ZN(n5238) );
  AND2_X1 U5887 ( .A1(n4927), .A2(n4931), .ZN(n4362) );
  INV_X1 U5888 ( .A(n9311), .ZN(n4676) );
  OR2_X1 U5889 ( .A1(n5882), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4363) );
  AND2_X1 U5890 ( .A1(n4854), .A2(n4851), .ZN(n4364) );
  OR2_X1 U5891 ( .A1(n10073), .A2(n8779), .ZN(n4365) );
  XNOR2_X1 U5892 ( .A(n5314), .B(n6431), .ZN(n5313) );
  INV_X1 U5893 ( .A(n6157), .ZN(n4456) );
  INV_X1 U5894 ( .A(n9757), .ZN(n9600) );
  NAND2_X1 U5895 ( .A1(n5573), .A2(n5572), .ZN(n9757) );
  AND2_X1 U5896 ( .A1(n4834), .A2(n4835), .ZN(n4366) );
  AND2_X1 U5897 ( .A1(n4993), .A2(n5705), .ZN(n4367) );
  NAND2_X1 U5898 ( .A1(n9757), .A2(n9079), .ZN(n9335) );
  INV_X1 U5899 ( .A(n9746), .ZN(n9560) );
  NAND2_X1 U5900 ( .A1(n5628), .A2(n5627), .ZN(n9746) );
  AND2_X1 U5901 ( .A1(n4749), .A2(n4748), .ZN(n4368) );
  AND2_X1 U5902 ( .A1(n5089), .A2(n4916), .ZN(n4369) );
  AND2_X1 U5903 ( .A1(n4676), .A2(n9312), .ZN(n4370) );
  OR2_X1 U5904 ( .A1(n8039), .A2(n8185), .ZN(n4371) );
  INV_X1 U5905 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4963) );
  OR2_X1 U5906 ( .A1(n9880), .A2(n9933), .ZN(n9253) );
  NOR2_X1 U5907 ( .A1(n7915), .A2(n8686), .ZN(n4372) );
  NOR2_X1 U5908 ( .A1(n9880), .A2(n7261), .ZN(n4373) );
  NOR2_X1 U5909 ( .A1(n9600), .A2(n9079), .ZN(n4374) );
  NOR2_X1 U5910 ( .A1(n5872), .A2(n7417), .ZN(n4375) );
  INV_X1 U5911 ( .A(n4740), .ZN(n4739) );
  OR2_X1 U5912 ( .A1(n4881), .A2(n5882), .ZN(n4376) );
  INV_X1 U5913 ( .A(n4697), .ZN(n4696) );
  NAND2_X1 U5914 ( .A1(n4699), .A2(n9541), .ZN(n4697) );
  INV_X1 U5915 ( .A(n8024), .ZN(n4576) );
  AND2_X1 U5916 ( .A1(n5141), .A2(SI_5_), .ZN(n4377) );
  AND2_X1 U5917 ( .A1(n5314), .A2(SI_12_), .ZN(n4378) );
  AND2_X1 U5918 ( .A1(n8796), .A2(n8208), .ZN(n4379) );
  NOR2_X1 U5919 ( .A1(n6271), .A2(n9703), .ZN(n4380) );
  NOR2_X1 U5920 ( .A1(n9960), .A2(n9407), .ZN(n4381) );
  AND2_X1 U5921 ( .A1(n8867), .A2(n8576), .ZN(n8160) );
  INV_X1 U5922 ( .A(n8463), .ZN(n4748) );
  AND2_X1 U5923 ( .A1(n5463), .A2(SI_18_), .ZN(n4382) );
  INV_X1 U5924 ( .A(n9707), .ZN(n4488) );
  AND2_X1 U5925 ( .A1(n9304), .A2(n9306), .ZN(n9707) );
  OAI21_X1 U5926 ( .B1(n7942), .B2(n6173), .A(n7943), .ZN(n4789) );
  AND2_X1 U5927 ( .A1(n8178), .A2(n8551), .ZN(n4383) );
  AND2_X1 U5928 ( .A1(n9735), .A2(n7843), .ZN(n4384) );
  NAND2_X1 U5929 ( .A1(n8861), .A2(n8537), .ZN(n8166) );
  OAI21_X1 U5930 ( .B1(n4457), .B2(n4456), .A(n7876), .ZN(n4455) );
  INV_X1 U5931 ( .A(n4591), .ZN(n4589) );
  NAND2_X1 U5932 ( .A1(n8383), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5933 ( .A1(n6154), .A2(n8072), .ZN(n4385) );
  NAND2_X1 U5934 ( .A1(n9356), .A2(n4698), .ZN(n4386) );
  INV_X1 U5935 ( .A(n4894), .ZN(n4893) );
  NAND2_X1 U5936 ( .A1(n4896), .A2(n5619), .ZN(n4894) );
  NAND2_X1 U5937 ( .A1(n9363), .A2(n9364), .ZN(n9362) );
  INV_X1 U5938 ( .A(n9362), .ZN(n4501) );
  OR2_X1 U5939 ( .A1(n8841), .A2(n8218), .ZN(n4387) );
  OR2_X1 U5940 ( .A1(n6614), .A2(n6615), .ZN(n4388) );
  AND2_X1 U5941 ( .A1(n4790), .A2(n6173), .ZN(n4389) );
  AND2_X1 U5942 ( .A1(n4608), .A2(n4360), .ZN(n4390) );
  AND2_X1 U5943 ( .A1(n4576), .A2(n4571), .ZN(n4391) );
  NAND2_X1 U5944 ( .A1(n5146), .A2(n5145), .ZN(n6270) );
  XNOR2_X1 U5945 ( .A(n5141), .B(n5115), .ZN(n5139) );
  NOR2_X1 U5946 ( .A1(n8431), .A2(n8430), .ZN(n4392) );
  OR2_X1 U5947 ( .A1(n6190), .A2(n5761), .ZN(n4393) );
  INV_X1 U5948 ( .A(n8208), .ZN(n8551) );
  AND2_X1 U5949 ( .A1(n6123), .A2(n6122), .ZN(n8208) );
  INV_X1 U5950 ( .A(n4649), .ZN(n4648) );
  NOR2_X1 U5951 ( .A1(n9927), .A2(n9410), .ZN(n4649) );
  NAND2_X1 U5952 ( .A1(n9742), .A2(n9564), .ZN(n9180) );
  INV_X1 U5953 ( .A(n8796), .ZN(n8178) );
  AND2_X1 U5954 ( .A1(n6115), .A2(n6114), .ZN(n8796) );
  AND2_X1 U5955 ( .A1(n4895), .A2(n4893), .ZN(n4394) );
  OR2_X1 U5956 ( .A1(n9746), .A2(n9544), .ZN(n9537) );
  INV_X1 U5957 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5865) );
  AND2_X1 U5958 ( .A1(n4892), .A2(n4335), .ZN(n4395) );
  AND2_X1 U5959 ( .A1(n8144), .A2(n6171), .ZN(n4396) );
  AND2_X1 U5960 ( .A1(n5754), .A2(n4883), .ZN(n4397) );
  NOR2_X1 U5961 ( .A1(n4606), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4398) );
  INV_X1 U5962 ( .A(n4436), .ZN(n8059) );
  NAND2_X1 U5963 ( .A1(n8055), .A2(n7412), .ZN(n4436) );
  OR2_X1 U5964 ( .A1(n4714), .A2(n4717), .ZN(n4399) );
  INV_X1 U5965 ( .A(n7544), .ZN(n4759) );
  INV_X1 U5966 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4639) );
  AND2_X1 U5967 ( .A1(n8173), .A2(n8179), .ZN(n4400) );
  INV_X1 U5968 ( .A(n9781), .ZN(n4786) );
  INV_X1 U5969 ( .A(n7631), .ZN(n9985) );
  NAND2_X1 U5970 ( .A1(n9299), .A2(n9223), .ZN(n9162) );
  INV_X1 U5971 ( .A(n9162), .ZN(n4663) );
  INV_X1 U5972 ( .A(n7329), .ZN(n4753) );
  NAND2_X1 U5973 ( .A1(n9065), .A2(n9066), .ZN(n8957) );
  NAND2_X1 U5974 ( .A1(n5652), .A2(n5651), .ZN(n9742) );
  INV_X1 U5975 ( .A(n9742), .ZN(n4780) );
  AND2_X1 U5976 ( .A1(n6716), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4401) );
  AND2_X1 U5977 ( .A1(n6828), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U5978 ( .A1(n5471), .A2(n5470), .ZN(n9777) );
  NAND2_X1 U5979 ( .A1(n5397), .A2(n5396), .ZN(n9719) );
  NAND2_X1 U5980 ( .A1(n4975), .A2(n4636), .ZN(n5364) );
  INV_X1 U5981 ( .A(n8358), .ZN(n8595) );
  AND2_X1 U5982 ( .A1(n6073), .A2(n6072), .ZN(n8358) );
  NAND2_X1 U5983 ( .A1(n9604), .A2(n4783), .ZN(n4784) );
  OR2_X1 U5984 ( .A1(n5926), .A2(n8735), .ZN(n4403) );
  NOR2_X1 U5985 ( .A1(n7918), .A2(n8663), .ZN(n4404) );
  AND2_X1 U5986 ( .A1(n5357), .A2(n8960), .ZN(n4405) );
  INV_X1 U5987 ( .A(n5939), .ZN(n8105) );
  OR2_X1 U5988 ( .A1(n8841), .A2(n8746), .ZN(n5939) );
  AND2_X1 U5989 ( .A1(n4726), .A2(n8358), .ZN(n4406) );
  INV_X1 U5990 ( .A(n9051), .ZN(n4897) );
  AND2_X1 U5991 ( .A1(n4670), .A2(n9283), .ZN(n4407) );
  AND2_X1 U5992 ( .A1(n4842), .A2(n4346), .ZN(n4408) );
  INV_X1 U5993 ( .A(n6264), .ZN(n4698) );
  AND2_X1 U5994 ( .A1(n9742), .A2(n9398), .ZN(n6264) );
  INV_X1 U5995 ( .A(n10092), .ZN(n10090) );
  NAND2_X1 U5996 ( .A1(n5268), .A2(n5267), .ZN(n7586) );
  NAND2_X1 U5997 ( .A1(n9274), .A2(n9270), .ZN(n4409) );
  INV_X1 U5998 ( .A(n8069), .ZN(n4580) );
  OR2_X1 U5999 ( .A1(n10078), .A2(n4464), .ZN(n4410) );
  AND2_X1 U6000 ( .A1(n7678), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4411) );
  INV_X1 U6001 ( .A(n7303), .ZN(n4682) );
  NAND2_X1 U6002 ( .A1(n5154), .A2(n7268), .ZN(n7291) );
  OR2_X1 U6003 ( .A1(n7916), .A2(n8676), .ZN(n4412) );
  INV_X1 U6004 ( .A(n4669), .ZN(n4668) );
  AND2_X1 U6005 ( .A1(n9160), .A2(n9283), .ZN(n4669) );
  INV_X1 U6006 ( .A(n9838), .ZN(n4687) );
  NAND2_X1 U6007 ( .A1(n4630), .A2(n5208), .ZN(n7592) );
  NOR2_X1 U6008 ( .A1(n7665), .A2(n4911), .ZN(n4413) );
  AND3_X1 U6009 ( .A1(n4715), .A2(n4717), .A3(n7279), .ZN(n4414) );
  INV_X1 U6010 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4598) );
  AND2_X1 U6011 ( .A1(n4757), .A2(n4756), .ZN(n4415) );
  INV_X1 U6012 ( .A(n4774), .ZN(n7725) );
  NOR3_X1 U6013 ( .A1(n7581), .A2(n4776), .A3(n7631), .ZN(n4774) );
  NOR3_X1 U6014 ( .A1(n7581), .A2(n4776), .A3(n4775), .ZN(n4777) );
  NAND2_X1 U6015 ( .A1(n7239), .A2(n4778), .ZN(n4779) );
  NAND2_X1 U6016 ( .A1(n4898), .A2(n5203), .ZN(n5208) );
  NOR2_X1 U6017 ( .A1(n8507), .A2(n8508), .ZN(n4416) );
  OR2_X1 U6018 ( .A1(n6619), .A2(n8725), .ZN(n4417) );
  INV_X1 U6019 ( .A(n5887), .ZN(n4584) );
  NAND2_X1 U6020 ( .A1(n4612), .A2(n5020), .ZN(n6852) );
  AND3_X1 U6021 ( .A1(n5806), .A2(n5805), .A3(n5804), .ZN(n10056) );
  INV_X1 U6022 ( .A(n10056), .ZN(n4592) );
  NAND2_X1 U6023 ( .A1(n9486), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U6024 ( .A1(n7119), .A2(n4829), .ZN(n4825) );
  XNOR2_X1 U6025 ( .A(n4930), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4937) );
  AND2_X1 U6026 ( .A1(n4762), .A2(n7123), .ZN(n4419) );
  INV_X1 U6027 ( .A(n7038), .ZN(n4434) );
  INV_X1 U6028 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4429) );
  INV_X1 U6029 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n4439) );
  INV_X1 U6030 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4819) );
  INV_X1 U6031 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n4438) );
  INV_X1 U6032 ( .A(n6659), .ZN(n4831) );
  NAND2_X1 U6033 ( .A1(n6578), .A2(n6659), .ZN(n7185) );
  NOR2_X1 U6034 ( .A1(n4830), .A2(n6659), .ZN(n4829) );
  INV_X1 U6035 ( .A(P2_U3893), .ZN(n8391) );
  NAND2_X2 U6036 ( .A1(n7113), .A2(n8200), .ZN(n8375) );
  NOR2_X1 U6037 ( .A1(n9577), .A2(n6290), .ZN(n9563) );
  NOR2_X1 U6038 ( .A1(n9561), .A2(n6292), .ZN(n9539) );
  NOR2_X1 U6039 ( .A1(n9589), .A2(n9590), .ZN(n9588) );
  OAI21_X1 U6040 ( .B1(n7853), .B2(n9356), .A(n9182), .ZN(n9528) );
  INV_X1 U6041 ( .A(n9686), .ZN(n4424) );
  NAND2_X1 U6042 ( .A1(n7809), .A2(n9298), .ZN(n7808) );
  OAI21_X1 U6043 ( .B1(n4665), .B2(n4661), .A(n4659), .ZN(n6286) );
  NOR2_X1 U6044 ( .A1(n9188), .A2(n9247), .ZN(n9613) );
  NAND2_X4 U6045 ( .A1(n6679), .A2(n7858), .ZN(n6631) );
  NAND2_X1 U6046 ( .A1(n9613), .A2(n9612), .ZN(n9611) );
  NAND2_X1 U6047 ( .A1(n4768), .A2(n4831), .ZN(n4767) );
  NAND2_X1 U6048 ( .A1(n4754), .A2(n4753), .ZN(n4752) );
  INV_X1 U6049 ( .A(n8492), .ZN(n4821) );
  OAI21_X1 U6050 ( .B1(n8032), .B2(n8036), .A(n8031), .ZN(n8193) );
  OR2_X1 U6051 ( .A1(n8029), .A2(n8033), .ZN(n8030) );
  NAND2_X4 U6052 ( .A1(n4657), .A2(n4656), .ZN(n6679) );
  NAND2_X2 U6053 ( .A1(n5205), .A2(n5204), .ZN(n4899) );
  INV_X1 U6054 ( .A(n5043), .ZN(n5041) );
  NAND2_X1 U6055 ( .A1(n6953), .A2(n6956), .ZN(n6954) );
  AOI21_X1 U6056 ( .B1(n8978), .B2(n8977), .A(n9053), .ZN(n8983) );
  NAND2_X1 U6057 ( .A1(n4325), .A2(n4621), .ZN(n4618) );
  NAND3_X1 U6058 ( .A1(n9031), .A2(n9033), .A3(n9032), .ZN(n9030) );
  OAI211_X1 U6059 ( .C1(n5208), .C2(n4629), .A(n5234), .B(n4626), .ZN(n5253)
         );
  OR2_X2 U6060 ( .A1(n9073), .A2(n9076), .ZN(n4624) );
  NAND2_X1 U6061 ( .A1(n9015), .A2(n4886), .ZN(n4641) );
  NOR2_X2 U6062 ( .A1(n4951), .A2(n4919), .ZN(n4925) );
  NAND4_X1 U6063 ( .A1(n4884), .A2(n4612), .A3(n5020), .A4(n5019), .ZN(n6853)
         );
  INV_X1 U6064 ( .A(n7334), .ZN(n8050) );
  OR2_X1 U6065 ( .A1(n4743), .A2(n4438), .ZN(n6573) );
  NAND2_X1 U6066 ( .A1(n4440), .A2(n5829), .ZN(n5840) );
  OR2_X1 U6067 ( .A1(n4743), .A2(n4439), .ZN(n6599) );
  NAND2_X1 U6068 ( .A1(n7611), .A2(n4446), .ZN(n4445) );
  NAND2_X1 U6069 ( .A1(n4449), .A2(n4450), .ZN(n6158) );
  NAND2_X1 U6070 ( .A1(n6156), .A2(n4452), .ZN(n4449) );
  NAND2_X1 U6071 ( .A1(n4463), .A2(n4390), .ZN(n4846) );
  NAND2_X4 U6072 ( .A1(n4461), .A2(n9136), .ZN(n7983) );
  NAND4_X1 U6073 ( .A1(n4342), .A2(n8516), .A3(n4416), .A4(n4468), .ZN(
        P2_U3201) );
  XNOR2_X1 U6074 ( .A(n4477), .B(n4476), .ZN(n7010) );
  NAND2_X1 U6075 ( .A1(n4479), .A2(n4478), .ZN(n9357) );
  NAND2_X1 U6076 ( .A1(n4480), .A2(n9369), .ZN(n4479) );
  NAND2_X1 U6077 ( .A1(n4481), .A2(n9349), .ZN(n4480) );
  NAND2_X1 U6078 ( .A1(n4482), .A2(n9180), .ZN(n4481) );
  NAND2_X1 U6079 ( .A1(n4483), .A2(n9537), .ZN(n4482) );
  NAND2_X1 U6080 ( .A1(n9348), .A2(n9347), .ZN(n4483) );
  NAND2_X1 U6081 ( .A1(n9343), .A2(n9342), .ZN(n9348) );
  NAND2_X1 U6082 ( .A1(n9303), .A2(n4347), .ZN(n4484) );
  OAI21_X1 U6083 ( .B1(n9303), .B2(n4488), .A(n4347), .ZN(n9325) );
  NAND2_X1 U6084 ( .A1(n4484), .A2(n4485), .ZN(n9327) );
  AND2_X2 U6085 ( .A1(n4490), .A2(n4646), .ZN(n9252) );
  NAND3_X1 U6086 ( .A1(n4645), .A2(n6278), .A3(n6277), .ZN(n4490) );
  NAND2_X1 U6087 ( .A1(n7217), .A2(n7216), .ZN(n6277) );
  INV_X2 U6088 ( .A(n9917), .ZN(n9201) );
  AND3_X2 U6089 ( .A1(n4925), .A2(n4924), .A3(n4324), .ZN(n4945) );
  NAND3_X1 U6090 ( .A1(n4496), .A2(n9260), .A3(n4495), .ZN(n4494) );
  NAND3_X1 U6091 ( .A1(n9361), .A2(n9360), .A3(n4501), .ZN(n4500) );
  NAND3_X1 U6092 ( .A1(n8051), .A2(n4504), .A3(n8062), .ZN(n4503) );
  NAND3_X1 U6093 ( .A1(n4503), .A2(n8063), .A3(n4502), .ZN(n8065) );
  NAND3_X1 U6094 ( .A1(n4504), .A2(n8062), .A3(n4436), .ZN(n4502) );
  NAND2_X1 U6095 ( .A1(n8051), .A2(n8050), .ZN(n8061) );
  NAND2_X2 U6096 ( .A1(n8197), .A2(n8033), .ZN(n8171) );
  NAND2_X1 U6097 ( .A1(n4848), .A2(n4850), .ZN(n4507) );
  NAND3_X1 U6098 ( .A1(n8118), .A2(n8117), .A3(n4850), .ZN(n4508) );
  NAND3_X1 U6099 ( .A1(n4508), .A2(n4396), .A3(n4507), .ZN(n8150) );
  NAND2_X1 U6100 ( .A1(n6125), .A2(n6124), .ZN(n4517) );
  NAND2_X1 U6101 ( .A1(n4518), .A2(n4519), .ZN(n5156) );
  NAND3_X1 U6102 ( .A1(n4795), .A2(n4793), .A3(n5139), .ZN(n4518) );
  INV_X1 U6103 ( .A(n4522), .ZN(n6112) );
  INV_X1 U6104 ( .A(n5670), .ZN(n4527) );
  NAND2_X1 U6105 ( .A1(n5442), .A2(n4531), .ZN(n4528) );
  NAND2_X1 U6106 ( .A1(n4528), .A2(n4529), .ZN(n5516) );
  OAI21_X1 U6107 ( .B1(n5442), .B2(n5443), .A(n5444), .ZN(n5465) );
  NAND2_X1 U6108 ( .A1(n5621), .A2(n5620), .ZN(n4540) );
  NAND2_X1 U6109 ( .A1(n5595), .A2(n5594), .ZN(n4541) );
  NAND2_X1 U6110 ( .A1(n5176), .A2(n4545), .ZN(n4542) );
  NAND2_X1 U6111 ( .A1(n4542), .A2(n4543), .ZN(n5237) );
  NAND4_X1 U6112 ( .A1(n9377), .A2(n9378), .A3(n4557), .A4(n4556), .ZN(n9395)
         );
  NAND2_X4 U6113 ( .A1(n4560), .A2(n4563), .ZN(n8390) );
  NAND2_X1 U6114 ( .A1(n8040), .A2(n8039), .ZN(n7097) );
  NAND2_X1 U6115 ( .A1(n6098), .A2(n4391), .ZN(n4564) );
  OAI211_X1 U6116 ( .C1(n6098), .C2(n4568), .A(n4565), .B(n4564), .ZN(n6146)
         );
  NAND2_X1 U6117 ( .A1(n6098), .A2(n4353), .ZN(n4570) );
  NAND2_X1 U6118 ( .A1(n6098), .A2(n6097), .ZN(n8549) );
  NAND2_X1 U6121 ( .A1(n5875), .A2(n4582), .ZN(n4581) );
  NAND4_X1 U6122 ( .A1(n4595), .A2(n5757), .A3(n5994), .A4(n4594), .ZN(n4593)
         );
  NAND4_X1 U6123 ( .A1(n4397), .A2(n5966), .A3(n4597), .A4(n5802), .ZN(n4596)
         );
  NAND2_X1 U6124 ( .A1(n6187), .A2(n6186), .ZN(n8526) );
  INV_X1 U6125 ( .A(n6141), .ZN(n4605) );
  NAND2_X1 U6126 ( .A1(n4605), .A2(n4398), .ZN(n4608) );
  INV_X1 U6127 ( .A(n4608), .ZN(n5786) );
  NAND2_X1 U6128 ( .A1(n8662), .A2(n8659), .ZN(n4611) );
  NAND2_X1 U6129 ( .A1(n8573), .A2(n6085), .ZN(n8559) );
  NAND2_X2 U6130 ( .A1(n4611), .A2(n6024), .ZN(n8566) );
  NAND2_X1 U6131 ( .A1(n5001), .A2(n5000), .ZN(n4612) );
  NAND2_X1 U6132 ( .A1(n4615), .A2(n4613), .ZN(n9057) );
  NAND2_X1 U6133 ( .A1(n4616), .A2(n9074), .ZN(n4615) );
  NAND2_X1 U6134 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U6135 ( .A1(n4619), .A2(n9073), .ZN(n4617) );
  INV_X1 U6136 ( .A(n4325), .ZN(n4620) );
  NAND2_X1 U6137 ( .A1(n4624), .A2(n9074), .ZN(n8977) );
  AND2_X1 U6138 ( .A1(n4624), .A2(n4622), .ZN(n9053) );
  INV_X1 U6139 ( .A(n8978), .ZN(n4623) );
  NAND2_X1 U6140 ( .A1(n4899), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U6141 ( .A1(n7697), .A2(n7699), .ZN(n7698) );
  NAND2_X1 U6142 ( .A1(n4631), .A2(n5208), .ZN(n7697) );
  INV_X1 U6143 ( .A(n7699), .ZN(n4629) );
  NAND3_X1 U6144 ( .A1(n6954), .A2(n4632), .A3(n5073), .ZN(n7075) );
  NAND2_X1 U6145 ( .A1(n5154), .A2(n4634), .ZN(n4633) );
  INV_X1 U6146 ( .A(n4898), .ZN(n5205) );
  INV_X1 U6147 ( .A(n5364), .ZN(n4980) );
  NOR2_X1 U6148 ( .A1(n4951), .A2(n4638), .ZN(n5161) );
  NAND2_X1 U6149 ( .A1(n4641), .A2(n4885), .ZN(n5384) );
  NAND2_X1 U6150 ( .A1(n4641), .A2(n4640), .ZN(n9121) );
  INV_X2 U6151 ( .A(n8972), .ZN(n9006) );
  NAND2_X2 U6152 ( .A1(n9002), .A2(n5535), .ZN(n8972) );
  NAND2_X4 U6153 ( .A1(n4642), .A2(n9386), .ZN(n5694) );
  NAND2_X2 U6154 ( .A1(n4989), .A2(n4990), .ZN(n5728) );
  NOR2_X1 U6155 ( .A1(n4649), .A2(n4647), .ZN(n4645) );
  NAND2_X1 U6156 ( .A1(n9252), .A2(n6279), .ZN(n6280) );
  NAND3_X1 U6157 ( .A1(n6277), .A2(n6278), .A3(n6276), .ZN(n4651) );
  INV_X1 U6158 ( .A(n4662), .ZN(n4661) );
  NAND3_X1 U6159 ( .A1(n4677), .A2(n4678), .A3(n4915), .ZN(n5062) );
  NAND2_X1 U6160 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4679), .ZN(n5028) );
  NAND2_X1 U6161 ( .A1(n6484), .A2(n9413), .ZN(n4973) );
  NAND2_X1 U6162 ( .A1(n7301), .A2(n4680), .ZN(n4681) );
  NAND2_X1 U6163 ( .A1(n4681), .A2(n4683), .ZN(n7451) );
  NAND2_X1 U6164 ( .A1(n9536), .A2(n4692), .ZN(n4690) );
  NAND2_X1 U6165 ( .A1(n9536), .A2(n4696), .ZN(n4691) );
  AOI21_X1 U6166 ( .B1(n9536), .B2(n9541), .A(n6264), .ZN(n7842) );
  NAND2_X1 U6167 ( .A1(n4701), .A2(n4700), .ZN(n9866) );
  NAND3_X1 U6168 ( .A1(n9886), .A2(n9151), .A3(n9887), .ZN(n4701) );
  NAND2_X1 U6169 ( .A1(n9886), .A2(n9887), .ZN(n4703) );
  NAND2_X1 U6170 ( .A1(n6262), .A2(n4706), .ZN(n4704) );
  NAND2_X1 U6171 ( .A1(n4704), .A2(n4705), .ZN(n9570) );
  NAND2_X1 U6172 ( .A1(n9708), .A2(n4326), .ZN(n4711) );
  NAND2_X1 U6173 ( .A1(n4945), .A2(n4343), .ZN(n9798) );
  AND2_X1 U6174 ( .A1(n4945), .A2(n4712), .ZN(n4962) );
  AOI211_X2 U6175 ( .C1(n9959), .C2(n6298), .A(n7953), .B(n7960), .ZN(n6299)
         );
  INV_X2 U6176 ( .A(n4954), .ZN(n4924) );
  MUX2_X1 U6177 ( .A(n6681), .B(n9809), .S(n6631), .Z(n7252) );
  NOR2_X1 U6178 ( .A1(n9527), .A2(n7854), .ZN(n7855) );
  XNOR2_X1 U6179 ( .A(n7936), .B(n6977), .ZN(n7084) );
  AND3_X2 U6180 ( .A1(n6975), .A2(n6974), .A3(n6973), .ZN(n7936) );
  OAI21_X2 U6181 ( .B1(n5992), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5995) );
  NOR2_X2 U6182 ( .A1(n5968), .A2(n5967), .ZN(n5980) );
  OAI211_X1 U6183 ( .C1(n4715), .C2(n4714), .A(n4399), .B(n4713), .ZN(n7640)
         );
  NAND3_X1 U6184 ( .A1(n7109), .A2(n4716), .A3(n7110), .ZN(n4713) );
  NAND2_X1 U6185 ( .A1(n8223), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U6186 ( .A1(n4720), .A2(n4718), .ZN(n7939) );
  OAI21_X1 U6187 ( .B1(n8223), .B2(n7934), .A(n7933), .ZN(n8263) );
  NAND2_X1 U6188 ( .A1(n7933), .A2(n7934), .ZN(n4725) );
  INV_X1 U6189 ( .A(n7935), .ZN(n4726) );
  NAND2_X1 U6190 ( .A1(n7665), .A2(n4330), .ZN(n4729) );
  NAND2_X1 U6191 ( .A1(n8271), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6192 ( .A1(n4744), .A2(n4745), .ZN(n8511) );
  INV_X1 U6193 ( .A(n4749), .ZN(n8462) );
  NAND2_X1 U6194 ( .A1(n4751), .A2(n7367), .ZN(n6583) );
  INV_X1 U6195 ( .A(n6581), .ZN(n4754) );
  NAND2_X1 U6196 ( .A1(n6587), .A2(n4759), .ZN(n4755) );
  OAI21_X1 U6197 ( .B1(n6586), .B2(n4329), .A(n4755), .ZN(n7543) );
  INV_X1 U6198 ( .A(n6586), .ZN(n4758) );
  NAND2_X1 U6199 ( .A1(n4761), .A2(n7123), .ZN(n6576) );
  NAND2_X1 U6200 ( .A1(n4766), .A2(n7185), .ZN(n6579) );
  INV_X1 U6201 ( .A(n6578), .ZN(n4768) );
  NAND2_X1 U6202 ( .A1(n4322), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4970) );
  OR2_X2 U6203 ( .A1(n4945), .A2(n5288), .ZN(n4769) );
  INV_X1 U6204 ( .A(n4777), .ZN(n7813) );
  NAND3_X1 U6205 ( .A1(n7239), .A2(n9933), .A3(n4778), .ZN(n9868) );
  INV_X1 U6206 ( .A(n4779), .ZN(n9889) );
  INV_X1 U6207 ( .A(n4784), .ZN(n9578) );
  INV_X1 U6208 ( .A(n5058), .ZN(n4797) );
  OAI21_X1 U6209 ( .B1(n5059), .B2(n4792), .A(n4791), .ZN(n5111) );
  AOI21_X1 U6210 ( .B1(n4797), .B2(n5085), .A(n4345), .ZN(n4791) );
  INV_X1 U6211 ( .A(n5085), .ZN(n4792) );
  INV_X1 U6212 ( .A(n4794), .ZN(n4793) );
  NAND2_X1 U6213 ( .A1(n5259), .A2(n4800), .ZN(n4798) );
  NAND2_X1 U6214 ( .A1(n4798), .A2(n4799), .ZN(n5335) );
  NAND3_X1 U6215 ( .A1(n4816), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4815) );
  NAND3_X1 U6216 ( .A1(n8504), .A2(n4819), .A3(n4818), .ZN(n4817) );
  NAND3_X1 U6217 ( .A1(n8489), .A2(n8490), .A3(n4820), .ZN(P2_U3200) );
  NAND2_X1 U6218 ( .A1(n7038), .A2(n6597), .ZN(n4823) );
  XNOR2_X2 U6219 ( .A(n5830), .B(n5829), .ZN(n7038) );
  NAND2_X1 U6220 ( .A1(n7039), .A2(n6600), .ZN(n6601) );
  AOI21_X1 U6221 ( .B1(n7119), .B2(n6604), .A(n4831), .ZN(n4824) );
  NOR2_X1 U6222 ( .A1(n4831), .A2(n6604), .ZN(n4827) );
  INV_X1 U6223 ( .A(n4842), .ZN(n7786) );
  MUX2_X1 U6224 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n8493), .Z(n6516) );
  MUX2_X1 U6225 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n8493), .Z(n6987) );
  MUX2_X1 U6226 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n8493), .Z(n6520) );
  MUX2_X1 U6227 ( .A(P2_REG1_REG_5__SCAN_IN), .B(P2_REG2_REG_5__SCAN_IN), .S(
        n8493), .Z(n6522) );
  MUX2_X1 U6228 ( .A(n6547), .B(n8767), .S(n8493), .Z(n6548) );
  NOR2_X1 U6229 ( .A1(n4847), .A2(n8493), .ZN(n8514) );
  OR2_X1 U6230 ( .A1(n8127), .A2(n4849), .ZN(n4848) );
  NAND3_X1 U6231 ( .A1(n8040), .A2(n8035), .A3(n8197), .ZN(n4858) );
  NAND3_X1 U6232 ( .A1(n4863), .A2(n8743), .A3(n4859), .ZN(n8098) );
  NAND2_X1 U6233 ( .A1(n8180), .A2(n8179), .ZN(n4869) );
  NAND2_X1 U6234 ( .A1(n4871), .A2(n8171), .ZN(n4870) );
  NAND2_X1 U6235 ( .A1(n4872), .A2(n8174), .ZN(n4871) );
  NAND2_X1 U6236 ( .A1(n4876), .A2(n8208), .ZN(n4872) );
  NAND2_X1 U6237 ( .A1(n4874), .A2(n8185), .ZN(n4873) );
  NAND2_X1 U6238 ( .A1(n4875), .A2(n8177), .ZN(n4874) );
  NAND2_X1 U6239 ( .A1(n4876), .A2(n8796), .ZN(n4875) );
  OR2_X1 U6240 ( .A1(n8180), .A2(n4400), .ZN(n4876) );
  NAND2_X1 U6241 ( .A1(n6138), .A2(n5759), .ZN(n6190) );
  NAND2_X1 U6242 ( .A1(n5003), .A2(n5002), .ZN(n5020) );
  NAND3_X1 U6243 ( .A1(n4925), .A2(n4924), .A3(n4926), .ZN(n4991) );
  NAND2_X1 U6244 ( .A1(n8972), .A2(n4395), .ZN(n4890) );
  AND2_X1 U6245 ( .A1(n5208), .A2(n4899), .ZN(n7591) );
  AND2_X1 U6246 ( .A1(n4937), .A2(n4936), .ZN(n5021) );
  NAND3_X1 U6247 ( .A1(n5130), .A2(n7267), .A3(n7157), .ZN(n5154) );
  OAI21_X1 U6248 ( .B1(n8629), .B2(n6169), .A(n8138), .ZN(n8612) );
  NAND2_X1 U6249 ( .A1(n5835), .A2(n5834), .ZN(n7205) );
  INV_X1 U6250 ( .A(n6188), .ZN(n8534) );
  NAND2_X1 U6251 ( .A1(n8683), .A2(n5991), .ZN(n8673) );
  NAND2_X1 U6252 ( .A1(n9526), .A2(n9519), .ZN(n9520) );
  NAND2_X1 U6253 ( .A1(n8673), .A2(n6006), .ZN(n6008) );
  INV_X1 U6254 ( .A(n7097), .ZN(n8006) );
  NAND2_X1 U6255 ( .A1(n8758), .A2(n8757), .ZN(n8756) );
  NAND2_X1 U6256 ( .A1(n9620), .A2(n6259), .ZN(n6262) );
  NAND2_X1 U6257 ( .A1(n5786), .A2(n5783), .ZN(n5766) );
  NAND2_X1 U6258 ( .A1(n5786), .A2(n5764), .ZN(n8949) );
  NAND2_X1 U6259 ( .A1(n8333), .A2(n7892), .ZN(n8256) );
  NAND2_X1 U6260 ( .A1(n8229), .A2(n7891), .ZN(n8333) );
  NAND2_X1 U6261 ( .A1(n6251), .A2(n6250), .ZN(n7301) );
  OR2_X1 U6262 ( .A1(n5049), .A2(n4933), .ZN(n4934) );
  NAND2_X1 U6263 ( .A1(n5129), .A2(n5128), .ZN(n7157) );
  NOR2_X1 U6264 ( .A1(n6201), .A2(n6200), .ZN(n6203) );
  NAND2_X1 U6265 ( .A1(n7075), .A2(n5103), .ZN(n5126) );
  INV_X1 U6266 ( .A(n5126), .ZN(n5129) );
  AOI21_X1 U6267 ( .B1(n8163), .B2(n8162), .A(n4909), .ZN(n8170) );
  NAND2_X1 U6268 ( .A1(n8153), .A2(n8580), .ZN(n8163) );
  INV_X1 U6269 ( .A(n5778), .ZN(n8202) );
  NAND2_X1 U6270 ( .A1(n8390), .A2(n6976), .ZN(n8040) );
  INV_X1 U6271 ( .A(n4962), .ZN(n4965) );
  OR2_X1 U6272 ( .A1(n4962), .A2(n5288), .ZN(n4932) );
  OAI21_X1 U6273 ( .B1(n5567), .B2(n5566), .A(n5565), .ZN(n5595) );
  XNOR2_X1 U6274 ( .A(n5567), .B(n5566), .ZN(n7599) );
  NOR2_X1 U6275 ( .A1(n6272), .A2(n7252), .ZN(n6946) );
  AOI21_X1 U6276 ( .B1(n6272), .B2(n6484), .A(n5012), .ZN(n5018) );
  OAI22_X1 U6277 ( .A1(n7640), .A2(n7639), .B1(n7638), .B2(n8386), .ZN(n7641)
         );
  NAND2_X1 U6278 ( .A1(n8231), .A2(n8230), .ZN(n8229) );
  OAI21_X2 U6279 ( .B1(n9097), .B2(n9101), .A(n8996), .ZN(n8995) );
  XNOR2_X1 U6280 ( .A(n7890), .B(n8762), .ZN(n8231) );
  NOR2_X2 U6281 ( .A1(n9099), .A2(n9098), .ZN(n9097) );
  NOR2_X2 U6282 ( .A1(n5460), .A2(n5459), .ZN(n9099) );
  OAI21_X1 U6283 ( .B1(n5725), .B2(n6493), .A(n9113), .ZN(n5752) );
  INV_X1 U6284 ( .A(n9283), .ZN(n6285) );
  OR2_X1 U6285 ( .A1(n8164), .A2(n8838), .ZN(n4901) );
  INV_X1 U6286 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5762) );
  AND2_X1 U6287 ( .A1(n10067), .A2(n7889), .ZN(n4902) );
  OR2_X1 U6288 ( .A1(n7958), .A2(n9135), .ZN(n4903) );
  AND2_X1 U6289 ( .A1(n7897), .A2(n8746), .ZN(n4904) );
  OR2_X1 U6290 ( .A1(n8164), .A2(n8934), .ZN(n4905) );
  OR2_X1 U6291 ( .A1(n8534), .A2(n10062), .ZN(n4906) );
  AND2_X1 U6292 ( .A1(n6194), .A2(n6192), .ZN(n4907) );
  AND2_X1 U6293 ( .A1(n5236), .A2(n5216), .ZN(n4908) );
  INV_X1 U6294 ( .A(n8384), .ZN(n7666) );
  AND2_X1 U6295 ( .A1(n7664), .A2(n8385), .ZN(n4911) );
  INV_X2 U6296 ( .A(n6054), .ZN(n7985) );
  AND2_X1 U6297 ( .A1(n8289), .A2(n8288), .ZN(n4912) );
  NAND2_X1 U6298 ( .A1(n8573), .A2(n8572), .ZN(n4913) );
  NAND2_X1 U6299 ( .A1(n6164), .A2(n8130), .ZN(n4914) );
  AND2_X1 U6300 ( .A1(n8176), .A2(n8175), .ZN(n8177) );
  INV_X1 U6301 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4916) );
  INV_X1 U6302 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4920) );
  INV_X1 U6303 ( .A(n8686), .ZN(n6005) );
  INV_X1 U6304 ( .A(n5204), .ZN(n5203) );
  INV_X1 U6305 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4918) );
  OR2_X1 U6306 ( .A1(n8567), .A2(n6083), .ZN(n6075) );
  AND2_X1 U6307 ( .A1(n7443), .A2(n10051), .ZN(n5887) );
  NAND2_X1 U6308 ( .A1(n5102), .A2(n5101), .ZN(n5103) );
  NAND2_X1 U6309 ( .A1(n7899), .A2(n8734), .ZN(n7900) );
  NOR2_X1 U6310 ( .A1(n6585), .A2(n7474), .ZN(n6586) );
  AND2_X1 U6311 ( .A1(n6084), .A2(n8572), .ZN(n6085) );
  INV_X1 U6312 ( .A(n5252), .ZN(n5250) );
  AND2_X1 U6313 ( .A1(n9003), .A2(n9004), .ZN(n5535) );
  INV_X1 U6314 ( .A(n5383), .ZN(n5380) );
  AND2_X1 U6315 ( .A1(n5520), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5551) );
  INV_X1 U6316 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5132) );
  INV_X1 U6317 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4926) );
  OAI22_X1 U6318 ( .A1(n7878), .A2(n5949), .B1(n8722), .B2(n8381), .ZN(n8708)
         );
  INV_X1 U6319 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U6320 ( .A1(n8685), .A2(n8684), .ZN(n8683) );
  INV_X1 U6321 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U6322 ( .A1(n5384), .A2(n5383), .ZN(n9032) );
  AND2_X1 U6323 ( .A1(n5551), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5575) );
  AND2_X1 U6324 ( .A1(n5241), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5269) );
  OAI22_X1 U6325 ( .A1(n7866), .A2(n9835), .B1(n9833), .B2(n9564), .ZN(n6295)
         );
  OR2_X1 U6326 ( .A1(n5296), .A2(n5295), .ZN(n5321) );
  INV_X1 U6327 ( .A(n9553), .ZN(n9562) );
  OR2_X1 U6328 ( .A1(n7694), .A2(n9403), .ZN(n6254) );
  OR2_X1 U6329 ( .A1(n7966), .A2(n7965), .ZN(n7967) );
  NAND2_X1 U6330 ( .A1(n7709), .A2(n7666), .ZN(n7710) );
  AOI21_X1 U6331 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8449), .A(n8442), .ZN(
        n8461) );
  NAND2_X1 U6332 ( .A1(n8175), .A2(n7994), .ZN(n8024) );
  AND2_X1 U6333 ( .A1(n8194), .A2(n8190), .ZN(n7384) );
  INV_X1 U6334 ( .A(n8550), .ZN(n8576) );
  AND2_X1 U6335 ( .A1(n5912), .A2(n5911), .ZN(n10061) );
  OR2_X1 U6336 ( .A1(n6978), .A2(n8171), .ZN(n8778) );
  AND2_X1 U6337 ( .A1(n6896), .A2(n8947), .ZN(n6981) );
  INV_X1 U6338 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5767) );
  NOR2_X1 U6339 ( .A1(n9006), .A2(n8973), .ZN(n9073) );
  AND2_X1 U6340 ( .A1(n5490), .A2(n5489), .ZN(n8996) );
  INV_X1 U6341 ( .A(n9615), .ZN(n9079) );
  AND2_X1 U6342 ( .A1(n9433), .A2(n9432), .ZN(n9434) );
  INV_X1 U6343 ( .A(n7867), .ZN(n7868) );
  INV_X1 U6344 ( .A(n9762), .ZN(n9606) );
  INV_X1 U6345 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6305) );
  INV_X1 U6346 ( .A(n7261), .ZN(n9933) );
  OR2_X1 U6347 ( .A1(n6790), .A2(n6302), .ZN(n7220) );
  XNOR2_X1 U6348 ( .A(n5333), .B(SI_13_), .ZN(n5331) );
  NAND2_X1 U6349 ( .A1(n5113), .A2(SI_4_), .ZN(n5114) );
  INV_X1 U6350 ( .A(SI_2_), .ZN(n5036) );
  INV_X1 U6351 ( .A(n6174), .ZN(n8194) );
  OR2_X1 U6352 ( .A1(P2_U3150), .A2(n6571), .ZN(n8505) );
  NAND2_X1 U6353 ( .A1(n8093), .A2(n8091), .ZN(n8757) );
  AND2_X1 U6354 ( .A1(n10038), .A2(n10029), .ZN(n8717) );
  AND2_X1 U6355 ( .A1(n7601), .A2(n8036), .ZN(n7382) );
  INV_X1 U6356 ( .A(n8838), .ZN(n8845) );
  AND2_X1 U6357 ( .A1(n5561), .A2(n5560), .ZN(n9076) );
  OR2_X1 U6358 ( .A1(n5738), .A2(n6728), .ZN(n5198) );
  OR2_X1 U6359 ( .A1(n5049), .A2(n5080), .ZN(n5081) );
  NOR2_X1 U6360 ( .A1(n6841), .A2(n6840), .ZN(n6908) );
  NOR2_X1 U6361 ( .A1(n7172), .A2(n7171), .ZN(n7402) );
  AOI211_X1 U6362 ( .C1(n9735), .C2(n9522), .A(n9670), .B(n9521), .ZN(n9734)
         );
  AND2_X1 U6363 ( .A1(n9142), .A2(n9143), .ZN(n9612) );
  INV_X1 U6364 ( .A(n9833), .ZN(n9877) );
  AND2_X1 U6365 ( .A1(n6303), .A2(n9380), .ZN(n9897) );
  INV_X1 U6366 ( .A(n9904), .ZN(n9893) );
  NOR2_X1 U6367 ( .A1(n9730), .A2(n9729), .ZN(n9732) );
  AND2_X1 U6368 ( .A1(n7579), .A2(n6940), .ZN(n9963) );
  INV_X1 U6369 ( .A(n9963), .ZN(n10000) );
  AND2_X1 U6370 ( .A1(n6628), .A2(n6626), .ZN(n9380) );
  XNOR2_X1 U6371 ( .A(n5177), .B(SI_7_), .ZN(n5175) );
  INV_X1 U6372 ( .A(n8344), .ZN(n8366) );
  AND2_X1 U6373 ( .A1(n7991), .A2(n6137), .ZN(n8538) );
  INV_X1 U6374 ( .A(n8734), .ZN(n8381) );
  INV_X1 U6375 ( .A(n8509), .ZN(n8484) );
  INV_X1 U6376 ( .A(n8514), .ZN(n8491) );
  AND2_X1 U6377 ( .A1(n7028), .A2(n8782), .ZN(n8739) );
  INV_X1 U6378 ( .A(n8717), .ZN(n8789) );
  INV_X1 U6379 ( .A(n7999), .ZN(n8851) );
  XOR2_X1 U6380 ( .A(n8594), .B(n8587), .Z(n8881) );
  OR2_X1 U6381 ( .A1(n10080), .A2(n10072), .ZN(n8934) );
  OR2_X1 U6382 ( .A1(n10080), .A2(n10074), .ZN(n8945) );
  AND2_X1 U6383 ( .A1(n6241), .A2(n6240), .ZN(n10080) );
  AND2_X1 U6384 ( .A1(n6570), .A2(n6899), .ZN(n8947) );
  INV_X1 U6385 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6666) );
  AND2_X1 U6386 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  INV_X1 U6387 ( .A(n9767), .ZN(n9633) );
  INV_X1 U6388 ( .A(n9082), .ZN(n9135) );
  AND4_X1 U6389 ( .A1(n6504), .A2(n6503), .A3(n6502), .A4(n6501), .ZN(n9530)
         );
  OR2_X1 U6390 ( .A1(n4321), .A2(n9496), .ZN(n9904) );
  INV_X1 U6391 ( .A(n10004), .ZN(n10002) );
  INV_X1 U6392 ( .A(n9912), .ZN(n9913) );
  INV_X1 U6393 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6678) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6649) );
  INV_X1 U6395 ( .A(n5062), .ZN(n4917) );
  NAND2_X1 U6396 ( .A1(n4917), .A2(n4369), .ZN(n4951) );
  NAND4_X1 U6397 ( .A1(n4953), .A2(n4952), .A3(n4639), .A4(n4918), .ZN(n4919)
         );
  NOR2_X2 U6398 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4976) );
  NAND3_X1 U6399 ( .A1(n4923), .A2(n4922), .A3(n4337), .ZN(n4954) );
  INV_X1 U6400 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4993) );
  INV_X1 U6401 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4927) );
  INV_X1 U6402 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4928) );
  INV_X1 U6403 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4929) );
  XNOR2_X2 U6404 ( .A(n4932), .B(n4931), .ZN(n4936) );
  NAND2_X1 U6405 ( .A1(n5021), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4935) );
  INV_X1 U6406 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4933) );
  AND2_X1 U6407 ( .A1(n4935), .A2(n4934), .ZN(n4942) );
  INV_X2 U6408 ( .A(n4936), .ZN(n9805) );
  INV_X1 U6409 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6856) );
  OR2_X1 U6410 ( .A1(n6499), .A2(n6856), .ZN(n4941) );
  NAND2_X4 U6411 ( .A1(n4938), .A2(n9805), .ZN(n5738) );
  INV_X1 U6412 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U6414 ( .A(n4967), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5711) );
  INV_X1 U6415 ( .A(n4943), .ZN(n4948) );
  NAND2_X1 U6416 ( .A1(n4948), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4944) );
  XNOR2_X1 U6417 ( .A(n4944), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5707) );
  INV_X1 U6418 ( .A(n4945), .ZN(n4946) );
  NAND2_X1 U6419 ( .A1(n4946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4947) );
  AND2_X1 U6420 ( .A1(n4949), .A2(n4948), .ZN(n5708) );
  NAND2_X1 U6421 ( .A1(n5161), .A2(n4953), .ZN(n4974) );
  OAI21_X1 U6422 ( .B1(n4974), .B2(n4954), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4955) );
  MUX2_X1 U6423 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4955), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n4957) );
  NAND2_X1 U6424 ( .A1(n4956), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4958) );
  XNOR2_X1 U6425 ( .A(n4958), .B(n4926), .ZN(n9204) );
  INV_X1 U6426 ( .A(n9204), .ZN(n9375) );
  INV_X1 U6427 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6654) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6647) );
  AND2_X1 U6429 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U6430 ( .A1(n5035), .A2(n4960), .ZN(n5010) );
  NAND3_X1 U6431 ( .A1(n6650), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4961) );
  NAND2_X1 U6432 ( .A1(n5010), .A2(n4961), .ZN(n5029) );
  XNOR2_X1 U6433 ( .A(n5030), .B(n5029), .ZN(n6653) );
  NAND2_X1 U6434 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n4966) );
  INV_X4 U6435 ( .A(n6631), .ZN(n5061) );
  NAND2_X1 U6436 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4968) );
  NAND2_X1 U6437 ( .A1(n5061), .A2(n6723), .ZN(n4969) );
  INV_X1 U6438 ( .A(n4997), .ZN(n4971) );
  NAND2_X1 U6439 ( .A1(n6628), .A2(n4971), .ZN(n5121) );
  INV_X1 U6440 ( .A(n5121), .ZN(n5682) );
  NAND2_X1 U6441 ( .A1(n6242), .A2(n5682), .ZN(n4972) );
  NAND2_X1 U6442 ( .A1(n4973), .A2(n4972), .ZN(n4996) );
  INV_X1 U6443 ( .A(n4974), .ZN(n4975) );
  NAND2_X1 U6444 ( .A1(n5289), .A2(n4976), .ZN(n4977) );
  NAND2_X1 U6445 ( .A1(n4980), .A2(n4979), .ZN(n5391) );
  OAI21_X2 U6446 ( .B1(n5391), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6447 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n4983) );
  NAND2_X1 U6448 ( .A1(n4983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4984) );
  OAI21_X1 U6449 ( .B1(n4985), .B2(P1_IR_REG_31__SCAN_IN), .A(n4984), .ZN(
        n4986) );
  INV_X1 U6450 ( .A(n4986), .ZN(n4987) );
  NOR2_X1 U6451 ( .A1(n4988), .A2(n4987), .ZN(n4989) );
  AND2_X1 U6452 ( .A1(n4991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6453 ( .A1(n4992), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n4995) );
  INV_X1 U6454 ( .A(n4992), .ZN(n4994) );
  NAND2_X1 U6455 ( .A1(n4994), .A2(n4993), .ZN(n5704) );
  NAND2_X1 U6456 ( .A1(n4995), .A2(n5704), .ZN(n9376) );
  OR2_X1 U6457 ( .A1(n9197), .A2(n9204), .ZN(n9386) );
  XNOR2_X1 U6458 ( .A(n4996), .B(n5694), .ZN(n5003) );
  INV_X1 U6459 ( .A(n5003), .ZN(n5001) );
  NAND2_X1 U6460 ( .A1(n6267), .A2(n9376), .ZN(n4998) );
  NAND2_X1 U6461 ( .A1(n9496), .A2(n4997), .ZN(n7237) );
  INV_X4 U6462 ( .A(n6486), .ZN(n5206) );
  AND2_X1 U6463 ( .A1(n6242), .A2(n6484), .ZN(n4999) );
  INV_X1 U6464 ( .A(n5002), .ZN(n5000) );
  INV_X1 U6465 ( .A(n5049), .ZN(n5104) );
  NAND2_X1 U6466 ( .A1(n5104), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5007) );
  INV_X1 U6467 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7250) );
  INV_X1 U6468 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6792) );
  OR2_X1 U6469 ( .A1(n4320), .A2(n6792), .ZN(n5005) );
  INV_X1 U6470 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6629) );
  INV_X1 U6471 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U6472 ( .A1(n9136), .A2(SI_0_), .ZN(n5009) );
  INV_X1 U6473 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6474 ( .A1(n5009), .A2(n5008), .ZN(n5011) );
  NAND2_X1 U6475 ( .A1(n5011), .A2(n5010), .ZN(n9809) );
  NOR2_X1 U6476 ( .A1(n7252), .A2(n5121), .ZN(n5012) );
  INV_X1 U6477 ( .A(n6628), .ZN(n5015) );
  NAND2_X1 U6478 ( .A1(n5015), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6479 ( .A1(n5018), .A2(n5013), .ZN(n6788) );
  NAND2_X1 U6480 ( .A1(n5206), .A2(n6272), .ZN(n5017) );
  AOI22_X1 U6481 ( .A1(n6943), .A2(n6484), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5015), .ZN(n5016) );
  NAND2_X1 U6482 ( .A1(n5017), .A2(n5016), .ZN(n6787) );
  NAND2_X1 U6483 ( .A1(n5018), .A2(n5694), .ZN(n5019) );
  NAND2_X1 U6484 ( .A1(n6853), .A2(n5020), .ZN(n5046) );
  NAND2_X1 U6485 ( .A1(n5021), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5027) );
  INV_X1 U6486 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5022) );
  OR2_X1 U6487 ( .A1(n5738), .A2(n5022), .ZN(n5026) );
  INV_X1 U6488 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5023) );
  OR2_X1 U6489 ( .A1(n5049), .A2(n5023), .ZN(n5025) );
  INV_X1 U6490 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9414) );
  OR2_X1 U6491 ( .A1(n4319), .A2(n9414), .ZN(n5024) );
  NAND2_X1 U6492 ( .A1(n9411), .A2(n6484), .ZN(n5038) );
  NAND2_X1 U6493 ( .A1(n5030), .A2(n5029), .ZN(n5034) );
  INV_X1 U6494 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6495 ( .A1(n5032), .A2(SI_1_), .ZN(n5033) );
  NAND2_X1 U6496 ( .A1(n5034), .A2(n5033), .ZN(n5056) );
  MUX2_X1 U6497 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5035), .Z(n5057) );
  XNOR2_X1 U6498 ( .A(n5056), .B(n5055), .ZN(n6655) );
  INV_X1 U6499 ( .A(n5121), .ZN(n5639) );
  NAND2_X1 U6500 ( .A1(n9201), .A2(n5639), .ZN(n5037) );
  NAND2_X1 U6501 ( .A1(n5038), .A2(n5037), .ZN(n5039) );
  XNOR2_X1 U6502 ( .A(n5039), .B(n5694), .ZN(n5044) );
  INV_X1 U6503 ( .A(n5044), .ZN(n5042) );
  AND2_X1 U6504 ( .A1(n9201), .A2(n6484), .ZN(n5040) );
  AOI21_X2 U6505 ( .B1(n5206), .B2(n9411), .A(n5040), .ZN(n5043) );
  NAND2_X1 U6506 ( .A1(n5042), .A2(n5041), .ZN(n5045) );
  NAND2_X1 U6507 ( .A1(n5044), .A2(n5043), .ZN(n5047) );
  AND2_X1 U6508 ( .A1(n5045), .A2(n5047), .ZN(n6866) );
  NAND2_X1 U6509 ( .A1(n5046), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U6510 ( .A1(n6865), .A2(n5047), .ZN(n6953) );
  NAND2_X1 U6511 ( .A1(n5021), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6512 ( .A1(n4320), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5053) );
  INV_X1 U6513 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5048) );
  OR2_X1 U6514 ( .A1(n5738), .A2(n5048), .ZN(n5052) );
  INV_X1 U6515 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5050) );
  OR2_X1 U6516 ( .A1(n5049), .A2(n5050), .ZN(n5051) );
  NAND2_X1 U6517 ( .A1(n9878), .A2(n6484), .ZN(n5067) );
  NAND2_X1 U6518 ( .A1(n5056), .A2(n5055), .ZN(n5059) );
  NAND2_X1 U6519 ( .A1(n5057), .A2(SI_2_), .ZN(n5058) );
  MUX2_X1 U6520 ( .A(n6658), .B(n6648), .S(n5035), .Z(n5087) );
  XNOR2_X1 U6521 ( .A(n5086), .B(n5085), .ZN(n6657) );
  NAND2_X1 U6522 ( .A1(n5060), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6523 ( .A1(n5063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6524 ( .A(n5090), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U6525 ( .A1(n5061), .A2(n6724), .ZN(n5064) );
  NAND2_X1 U6526 ( .A1(n7240), .A2(n5639), .ZN(n5066) );
  NAND2_X1 U6527 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  AND2_X1 U6528 ( .A1(n7240), .A2(n5697), .ZN(n5069) );
  AOI21_X1 U6529 ( .B1(n5206), .B2(n9878), .A(n5069), .ZN(n5071) );
  XNOR2_X1 U6530 ( .A(n5070), .B(n5071), .ZN(n6956) );
  INV_X1 U6531 ( .A(n5070), .ZN(n5072) );
  NAND2_X1 U6532 ( .A1(n5072), .A2(n5071), .ZN(n5073) );
  INV_X1 U6533 ( .A(n5738), .ZN(n5074) );
  NAND2_X1 U6534 ( .A1(n5074), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5084) );
  INV_X1 U6535 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5076) );
  INV_X1 U6536 ( .A(n5105), .ZN(n5079) );
  INV_X1 U6537 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7241) );
  INV_X1 U6538 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6539 ( .A1(n7241), .A2(n5077), .ZN(n5078) );
  NAND2_X1 U6540 ( .A1(n5079), .A2(n5078), .ZN(n9881) );
  OR2_X1 U6541 ( .A1(n4320), .A2(n9881), .ZN(n5082) );
  INV_X1 U6542 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6543 ( .A1(n9410), .A2(n6484), .ZN(n5096) );
  INV_X1 U6544 ( .A(n5087), .ZN(n5088) );
  INV_X1 U6545 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6652) );
  MUX2_X1 U6546 ( .A(n6652), .B(n6649), .S(n5035), .Z(n5112) );
  XNOR2_X1 U6547 ( .A(n5111), .B(n5110), .ZN(n6651) );
  NAND2_X1 U6548 ( .A1(n5060), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6549 ( .A1(n5090), .A2(n5089), .ZN(n5091) );
  NAND2_X1 U6550 ( .A1(n5091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U6551 ( .A(n5092), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U6552 ( .A1(n5061), .A2(n6725), .ZN(n5093) );
  NAND2_X1 U6553 ( .A1(n7079), .A2(n5639), .ZN(n5095) );
  NAND2_X1 U6554 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  XNOR2_X1 U6555 ( .A(n5097), .B(n5694), .ZN(n5099) );
  AND2_X1 U6556 ( .A1(n7079), .A2(n6484), .ZN(n5098) );
  AOI21_X1 U6557 ( .B1(n5206), .B2(n9410), .A(n5098), .ZN(n5100) );
  XNOR2_X1 U6558 ( .A(n5099), .B(n5100), .ZN(n7077) );
  INV_X1 U6559 ( .A(n5099), .ZN(n5102) );
  INV_X1 U6560 ( .A(n5100), .ZN(n5101) );
  NAND2_X1 U6561 ( .A1(n5104), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5109) );
  INV_X1 U6562 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7259) );
  OR2_X1 U6563 ( .A1(n5075), .A2(n7259), .ZN(n5108) );
  OAI21_X1 U6564 ( .B1(n5105), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5133), .ZN(
        n7258) );
  OR2_X1 U6565 ( .A1(n4319), .A2(n7258), .ZN(n5107) );
  INV_X1 U6566 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6721) );
  OR2_X1 U6567 ( .A1(n5738), .A2(n6721), .ZN(n5106) );
  NAND2_X1 U6568 ( .A1(n9880), .A2(n5697), .ZN(n5123) );
  INV_X1 U6569 ( .A(n5112), .ZN(n5113) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5035), .Z(n5141) );
  INV_X1 U6571 ( .A(SI_5_), .ZN(n5115) );
  XNOR2_X1 U6572 ( .A(n5140), .B(n5139), .ZN(n6661) );
  NAND2_X1 U6573 ( .A1(n5060), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6574 ( .A1(n4951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6575 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5116), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5118) );
  INV_X1 U6576 ( .A(n5142), .ZN(n5117) );
  NAND2_X1 U6577 ( .A1(n5061), .A2(n6720), .ZN(n5119) );
  NAND2_X1 U6578 ( .A1(n7261), .A2(n5639), .ZN(n5122) );
  NAND2_X1 U6579 ( .A1(n5123), .A2(n5122), .ZN(n5124) );
  XNOR2_X1 U6580 ( .A(n5124), .B(n6482), .ZN(n5127) );
  NAND2_X1 U6581 ( .A1(n5126), .A2(n5127), .ZN(n7156) );
  AND2_X1 U6582 ( .A1(n7261), .A2(n5697), .ZN(n5125) );
  NAND2_X1 U6583 ( .A1(n7156), .A2(n7158), .ZN(n5130) );
  INV_X1 U6584 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6585 ( .A1(n5104), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5138) );
  INV_X1 U6586 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5131) );
  AND2_X1 U6587 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  OR2_X1 U6588 ( .A1(n5134), .A2(n5164), .ZN(n9862) );
  INV_X1 U6589 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6719) );
  OR2_X1 U6590 ( .A1(n5738), .A2(n6719), .ZN(n5135) );
  NAND2_X1 U6591 ( .A1(n9409), .A2(n6484), .ZN(n5148) );
  MUX2_X1 U6592 ( .A(n6666), .B(n6663), .S(n5035), .Z(n5157) );
  XNOR2_X1 U6593 ( .A(n5156), .B(n5155), .ZN(n6665) );
  OR2_X1 U6594 ( .A1(n5217), .A2(n6665), .ZN(n5146) );
  INV_X1 U6595 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5288) );
  OR2_X1 U6596 ( .A1(n5142), .A2(n5288), .ZN(n5143) );
  XNOR2_X1 U6597 ( .A(n5143), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6718) );
  INV_X1 U6598 ( .A(n6718), .ZN(n6743) );
  OAI22_X1 U6599 ( .A1(n5394), .A2(n6663), .B1(n6631), .B2(n6743), .ZN(n5144)
         );
  INV_X1 U6600 ( .A(n5144), .ZN(n5145) );
  NAND2_X1 U6601 ( .A1(n6270), .A2(n5639), .ZN(n5147) );
  NAND2_X1 U6602 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  XNOR2_X1 U6603 ( .A(n5149), .B(n5694), .ZN(n5150) );
  AOI22_X1 U6604 ( .A1(n5206), .A2(n9409), .B1(n6484), .B2(n6270), .ZN(n5151)
         );
  NAND2_X1 U6605 ( .A1(n5150), .A2(n5151), .ZN(n7267) );
  INV_X1 U6606 ( .A(n5150), .ZN(n5153) );
  INV_X1 U6607 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6608 ( .A1(n5153), .A2(n5152), .ZN(n7268) );
  NAND2_X1 U6609 ( .A1(n5156), .A2(n5155), .ZN(n5160) );
  INV_X1 U6610 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6611 ( .A1(n5158), .A2(SI_6_), .ZN(n5159) );
  INV_X1 U6612 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6667) );
  INV_X1 U6613 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6669) );
  MUX2_X1 U6614 ( .A(n6667), .B(n6669), .S(n7969), .Z(n5177) );
  XNOR2_X1 U6615 ( .A(n5176), .B(n5175), .ZN(n6668) );
  OR2_X1 U6616 ( .A1(n6668), .A2(n5217), .ZN(n5163) );
  OR2_X1 U6617 ( .A1(n5161), .A2(n5288), .ZN(n5186) );
  XNOR2_X1 U6618 ( .A(n5186), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U6619 ( .A1(n5060), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5061), .B2(
        n6716), .ZN(n5162) );
  NAND2_X1 U6620 ( .A1(n9945), .A2(n5697), .ZN(n5171) );
  NAND2_X1 U6621 ( .A1(n5104), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5169) );
  INV_X1 U6622 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7312) );
  OR2_X1 U6623 ( .A1(n5075), .A2(n7312), .ZN(n5168) );
  INV_X1 U6624 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6717) );
  OR2_X1 U6625 ( .A1(n5738), .A2(n6717), .ZN(n5167) );
  NAND2_X1 U6626 ( .A1(n5164), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5193) );
  OR2_X1 U6627 ( .A1(n5164), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6628 ( .A1(n5193), .A2(n5165), .ZN(n7311) );
  OR2_X1 U6629 ( .A1(n4319), .A2(n7311), .ZN(n5166) );
  NAND4_X1 U6630 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n9861)
         );
  NAND2_X1 U6631 ( .A1(n5206), .A2(n9861), .ZN(n5170) );
  NAND2_X1 U6632 ( .A1(n5171), .A2(n5170), .ZN(n7293) );
  NAND2_X1 U6633 ( .A1(n9945), .A2(n5639), .ZN(n5173) );
  NAND2_X1 U6634 ( .A1(n9861), .A2(n5697), .ZN(n5172) );
  NAND2_X1 U6635 ( .A1(n5173), .A2(n5172), .ZN(n5174) );
  XNOR2_X1 U6636 ( .A(n5174), .B(n6482), .ZN(n7292) );
  INV_X1 U6637 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6638 ( .A1(n5178), .A2(SI_7_), .ZN(n5179) );
  INV_X1 U6639 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U6640 ( .A(n6676), .B(n6678), .S(n7969), .Z(n5181) );
  INV_X1 U6641 ( .A(SI_8_), .ZN(n5180) );
  INV_X1 U6642 ( .A(n5181), .ZN(n5182) );
  NAND2_X1 U6643 ( .A1(n5182), .A2(SI_8_), .ZN(n5183) );
  INV_X1 U6644 ( .A(n5210), .ZN(n5184) );
  XNOR2_X1 U6645 ( .A(n5211), .B(n5184), .ZN(n6677) );
  OR2_X1 U6646 ( .A1(n6677), .A2(n5217), .ZN(n5191) );
  INV_X1 U6647 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6648 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6649 ( .A1(n5187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5188) );
  XNOR2_X1 U6650 ( .A(n5188), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6828) );
  INV_X1 U6651 ( .A(n6828), .ZN(n6820) );
  OAI22_X1 U6652 ( .A1(n5394), .A2(n6678), .B1(n6631), .B2(n6820), .ZN(n5189)
         );
  INV_X1 U6653 ( .A(n5189), .ZN(n5190) );
  NAND2_X1 U6654 ( .A1(n7590), .A2(n5639), .ZN(n5201) );
  NAND2_X1 U6655 ( .A1(n7859), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5199) );
  INV_X1 U6656 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6728) );
  INV_X1 U6657 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6658 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  NAND2_X1 U6659 ( .A1(n5221), .A2(n5194), .ZN(n9848) );
  OR2_X1 U6660 ( .A1(n4319), .A2(n9848), .ZN(n5197) );
  INV_X1 U6661 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5195) );
  OR2_X1 U6662 ( .A1(n7862), .A2(n5195), .ZN(n5196) );
  NAND2_X1 U6663 ( .A1(n9408), .A2(n5697), .ZN(n5200) );
  NAND2_X1 U6664 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  XNOR2_X1 U6665 ( .A(n5202), .B(n6482), .ZN(n5204) );
  AND2_X1 U6666 ( .A1(n5206), .A2(n9408), .ZN(n5207) );
  AOI21_X1 U6667 ( .B1(n7590), .B2(n5697), .A(n5207), .ZN(n7593) );
  INV_X1 U6668 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6689) );
  INV_X1 U6669 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5212) );
  MUX2_X1 U6670 ( .A(n6689), .B(n5212), .S(n7969), .Z(n5214) );
  INV_X1 U6671 ( .A(SI_9_), .ZN(n5213) );
  INV_X1 U6672 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6673 ( .A1(n5215), .A2(SI_9_), .ZN(n5216) );
  XNOR2_X1 U6674 ( .A(n5235), .B(n4908), .ZN(n6687) );
  NAND2_X1 U6675 ( .A1(n6687), .A2(n9137), .ZN(n5220) );
  NAND2_X1 U6676 ( .A1(n4974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6677 ( .A(n5218), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6842) );
  AOI22_X1 U6678 ( .A1(n5060), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5061), .B2(
        n6842), .ZN(n5219) );
  NAND2_X1 U6679 ( .A1(n9960), .A2(n5639), .ZN(n5228) );
  NAND2_X1 U6680 ( .A1(n5104), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5226) );
  INV_X1 U6681 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7432) );
  OR2_X1 U6682 ( .A1(n5075), .A2(n7432), .ZN(n5225) );
  INV_X1 U6683 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6824) );
  AND2_X1 U6684 ( .A1(n5221), .A2(n6824), .ZN(n5222) );
  OR2_X1 U6685 ( .A1(n5222), .A2(n5241), .ZN(n7702) );
  OR2_X1 U6686 ( .A1(n4320), .A2(n7702), .ZN(n5224) );
  INV_X1 U6687 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6821) );
  OR2_X1 U6688 ( .A1(n5738), .A2(n6821), .ZN(n5223) );
  NAND4_X1 U6689 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), .ZN(n9407)
         );
  NAND2_X1 U6690 ( .A1(n9407), .A2(n5697), .ZN(n5227) );
  NAND2_X1 U6691 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  XNOR2_X1 U6692 ( .A(n5229), .B(n6482), .ZN(n5231) );
  AND2_X1 U6693 ( .A1(n5206), .A2(n9407), .ZN(n5230) );
  AOI21_X1 U6694 ( .B1(n9960), .B2(n5697), .A(n5230), .ZN(n5232) );
  XNOR2_X1 U6695 ( .A(n5231), .B(n5232), .ZN(n7699) );
  INV_X1 U6696 ( .A(n5231), .ZN(n5233) );
  NAND2_X1 U6697 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  INV_X1 U6698 ( .A(n5253), .ZN(n5251) );
  INV_X1 U6699 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6692) );
  INV_X1 U6700 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6694) );
  MUX2_X1 U6701 ( .A(n6692), .B(n6694), .S(n7969), .Z(n5256) );
  XNOR2_X1 U6702 ( .A(n5259), .B(n5255), .ZN(n6691) );
  NAND2_X1 U6703 ( .A1(n6691), .A2(n9137), .ZN(n5240) );
  NAND2_X1 U6704 ( .A1(n5238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U6705 ( .A(n5291), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U6706 ( .A1(n5060), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5061), .B2(
        n6909), .ZN(n5239) );
  NAND2_X1 U6707 ( .A1(n7459), .A2(n5639), .ZN(n5248) );
  NAND2_X1 U6708 ( .A1(n5104), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5246) );
  INV_X1 U6709 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7457) );
  OR2_X1 U6710 ( .A1(n5075), .A2(n7457), .ZN(n5245) );
  INV_X1 U6711 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6845) );
  OR2_X1 U6712 ( .A1(n5738), .A2(n6845), .ZN(n5244) );
  NOR2_X1 U6713 ( .A1(n5241), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5242) );
  OR2_X1 U6714 ( .A1(n5269), .A2(n5242), .ZN(n8990) );
  OR2_X1 U6715 ( .A1(n4320), .A2(n8990), .ZN(n5243) );
  NAND4_X1 U6716 ( .A1(n5246), .A2(n5245), .A3(n5244), .A4(n5243), .ZN(n9406)
         );
  NAND2_X1 U6717 ( .A1(n9406), .A2(n5697), .ZN(n5247) );
  NAND2_X1 U6718 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  XNOR2_X1 U6719 ( .A(n5249), .B(n5694), .ZN(n5252) );
  NAND2_X1 U6720 ( .A1(n5251), .A2(n5250), .ZN(n8984) );
  AND2_X1 U6721 ( .A1(n5206), .A2(n9406), .ZN(n5254) );
  AOI21_X1 U6722 ( .B1(n7459), .B2(n5697), .A(n5254), .ZN(n8987) );
  NAND3_X1 U6723 ( .A1(n8984), .A2(n9085), .A3(n8987), .ZN(n8985) );
  NAND2_X1 U6724 ( .A1(n8985), .A2(n9085), .ZN(n5284) );
  INV_X1 U6725 ( .A(n5256), .ZN(n5257) );
  INV_X1 U6726 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6708) );
  INV_X1 U6727 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6706) );
  MUX2_X1 U6728 ( .A(n6708), .B(n6706), .S(n7969), .Z(n5261) );
  INV_X1 U6729 ( .A(SI_11_), .ZN(n5260) );
  INV_X1 U6730 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6731 ( .A1(n5262), .A2(SI_11_), .ZN(n5263) );
  XNOR2_X1 U6732 ( .A(n5287), .B(n5286), .ZN(n6705) );
  NAND2_X1 U6733 ( .A1(n6705), .A2(n9137), .ZN(n5268) );
  INV_X1 U6734 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6735 ( .A1(n5291), .A2(n5264), .ZN(n5265) );
  NAND2_X1 U6736 ( .A1(n5265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5266) );
  XNOR2_X1 U6737 ( .A(n5266), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7149) );
  AOI22_X1 U6738 ( .A1(n5060), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5061), .B2(
        n7149), .ZN(n5267) );
  NAND2_X1 U6739 ( .A1(n7586), .A2(n5639), .ZN(n5276) );
  NAND2_X1 U6740 ( .A1(n5104), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5274) );
  INV_X1 U6741 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7580) );
  OR2_X1 U6742 ( .A1(n5075), .A2(n7580), .ZN(n5273) );
  INV_X1 U6743 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6915) );
  OR2_X1 U6744 ( .A1(n5738), .A2(n6915), .ZN(n5272) );
  OR2_X1 U6745 ( .A1(n5269), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6746 ( .A1(n5296), .A2(n5270), .ZN(n9092) );
  OR2_X1 U6747 ( .A1(n4319), .A2(n9092), .ZN(n5271) );
  NAND4_X1 U6748 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n9405)
         );
  NAND2_X1 U6749 ( .A1(n9405), .A2(n5697), .ZN(n5275) );
  NAND2_X1 U6750 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  XNOR2_X1 U6751 ( .A(n5277), .B(n5694), .ZN(n5279) );
  AND2_X1 U6752 ( .A1(n5206), .A2(n9405), .ZN(n5278) );
  AOI21_X1 U6753 ( .B1(n7586), .B2(n5697), .A(n5278), .ZN(n5280) );
  INV_X1 U6754 ( .A(n5279), .ZN(n5282) );
  INV_X1 U6755 ( .A(n5280), .ZN(n5281) );
  NAND2_X1 U6756 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  NAND2_X1 U6757 ( .A1(n5284), .A2(n9086), .ZN(n9011) );
  NAND2_X1 U6758 ( .A1(n9011), .A2(n9012), .ZN(n5311) );
  MUX2_X1 U6759 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7969), .Z(n5314) );
  INV_X1 U6760 ( .A(SI_12_), .ZN(n6431) );
  NAND2_X1 U6761 ( .A1(n6783), .A2(n9137), .ZN(n5294) );
  OR2_X1 U6762 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6763 ( .A1(n5291), .A2(n5290), .ZN(n5316) );
  INV_X1 U6764 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5292) );
  XNOR2_X1 U6765 ( .A(n5316), .B(n5292), .ZN(n7170) );
  AOI22_X1 U6766 ( .A1(n5060), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5061), .B2(
        n7170), .ZN(n5293) );
  NAND2_X1 U6767 ( .A1(n7631), .A2(n5639), .ZN(n5303) );
  NAND2_X1 U6768 ( .A1(n5104), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5301) );
  INV_X1 U6769 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7626) );
  OR2_X1 U6770 ( .A1(n5075), .A2(n7626), .ZN(n5300) );
  INV_X1 U6771 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7143) );
  OR2_X1 U6772 ( .A1(n5738), .A2(n7143), .ZN(n5299) );
  INV_X1 U6773 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6774 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U6775 ( .A1(n5321), .A2(n5297), .ZN(n9019) );
  OR2_X1 U6776 ( .A1(n4319), .A2(n9019), .ZN(n5298) );
  NAND4_X1 U6777 ( .A1(n5301), .A2(n5300), .A3(n5299), .A4(n5298), .ZN(n9404)
         );
  NAND2_X1 U6778 ( .A1(n9404), .A2(n5697), .ZN(n5302) );
  NAND2_X1 U6779 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  XNOR2_X1 U6780 ( .A(n5304), .B(n5694), .ZN(n5306) );
  AND2_X1 U6781 ( .A1(n5206), .A2(n9404), .ZN(n5305) );
  AOI21_X1 U6782 ( .B1(n7631), .B2(n5697), .A(n5305), .ZN(n5307) );
  NAND2_X1 U6783 ( .A1(n5306), .A2(n5307), .ZN(n5312) );
  INV_X1 U6784 ( .A(n5306), .ZN(n5309) );
  INV_X1 U6785 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U6786 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U6787 ( .A1(n5311), .A2(n9013), .ZN(n9015) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7969), .Z(n5333) );
  XNOR2_X1 U6789 ( .A(n5332), .B(n5331), .ZN(n6796) );
  NAND2_X1 U6790 ( .A1(n6796), .A2(n9137), .ZN(n5319) );
  OAI21_X1 U6791 ( .B1(n5316), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  XNOR2_X1 U6792 ( .A(n5317), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7403) );
  AOI22_X1 U6793 ( .A1(n5060), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5061), .B2(
        n7403), .ZN(n5318) );
  NAND2_X1 U6794 ( .A1(n7694), .A2(n5639), .ZN(n5328) );
  NAND2_X1 U6795 ( .A1(n5104), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5326) );
  INV_X1 U6796 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7690) );
  OR2_X1 U6797 ( .A1(n5075), .A2(n7690), .ZN(n5325) );
  INV_X1 U6798 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6799 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  NAND2_X1 U6800 ( .A1(n5342), .A2(n5322), .ZN(n9068) );
  OR2_X1 U6801 ( .A1(n4319), .A2(n9068), .ZN(n5324) );
  INV_X1 U6802 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7175) );
  OR2_X1 U6803 ( .A1(n5738), .A2(n7175), .ZN(n5323) );
  NAND4_X1 U6804 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n9403)
         );
  NAND2_X1 U6805 ( .A1(n9403), .A2(n5697), .ZN(n5327) );
  NAND2_X1 U6806 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  XNOR2_X1 U6807 ( .A(n5329), .B(n6482), .ZN(n5352) );
  AND2_X1 U6808 ( .A1(n5206), .A2(n9403), .ZN(n5330) );
  AOI21_X1 U6809 ( .B1(n7694), .B2(n5697), .A(n5330), .ZN(n5353) );
  XNOR2_X1 U6810 ( .A(n5352), .B(n5353), .ZN(n9066) );
  NAND2_X1 U6811 ( .A1(n5333), .A2(SI_13_), .ZN(n5334) );
  NAND2_X1 U6812 ( .A1(n5335), .A2(n5334), .ZN(n5360) );
  MUX2_X1 U6813 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7969), .Z(n5361) );
  XNOR2_X1 U6814 ( .A(n5361), .B(SI_14_), .ZN(n5358) );
  XNOR2_X1 U6815 ( .A(n5360), .B(n5358), .ZN(n6861) );
  NAND2_X1 U6816 ( .A1(n6861), .A2(n9137), .ZN(n5340) );
  INV_X1 U6817 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6862) );
  OR2_X1 U6818 ( .A1(n5336), .A2(n5288), .ZN(n5337) );
  XNOR2_X1 U6819 ( .A(n5337), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7678) );
  INV_X1 U6820 ( .A(n7678), .ZN(n7681) );
  OAI22_X1 U6821 ( .A1(n5394), .A2(n6862), .B1(n6631), .B2(n7681), .ZN(n5338)
         );
  INV_X1 U6822 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U6823 ( .A1(n5104), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5347) );
  INV_X1 U6824 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7726) );
  OR2_X1 U6825 ( .A1(n5075), .A2(n7726), .ZN(n5346) );
  INV_X1 U6826 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5341) );
  AND2_X1 U6827 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  OR2_X1 U6828 ( .A1(n5343), .A2(n5369), .ZN(n8965) );
  OR2_X1 U6829 ( .A1(n4320), .A2(n8965), .ZN(n5345) );
  INV_X1 U6830 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7397) );
  OR2_X1 U6831 ( .A1(n5738), .A2(n7397), .ZN(n5344) );
  NAND4_X1 U6832 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n9402)
         );
  AND2_X1 U6833 ( .A1(n5206), .A2(n9402), .ZN(n5348) );
  AOI21_X1 U6834 ( .B1(n8968), .B2(n5697), .A(n5348), .ZN(n5356) );
  NAND2_X1 U6835 ( .A1(n8968), .A2(n5639), .ZN(n5350) );
  NAND2_X1 U6836 ( .A1(n9402), .A2(n5697), .ZN(n5349) );
  NAND2_X1 U6837 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  XNOR2_X1 U6838 ( .A(n5351), .B(n5694), .ZN(n8961) );
  INV_X1 U6839 ( .A(n5352), .ZN(n5354) );
  AND2_X1 U6840 ( .A1(n5354), .A2(n5353), .ZN(n8958) );
  AOI21_X1 U6841 ( .B1(n5356), .B2(n8961), .A(n8958), .ZN(n5355) );
  INV_X1 U6842 ( .A(n8961), .ZN(n5357) );
  INV_X1 U6843 ( .A(n5356), .ZN(n8960) );
  INV_X1 U6844 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U6845 ( .A1(n5360), .A2(n5359), .ZN(n5363) );
  NAND2_X1 U6846 ( .A1(n5361), .A2(SI_14_), .ZN(n5362) );
  NAND2_X1 U6847 ( .A1(n5363), .A2(n5362), .ZN(n5387) );
  MUX2_X1 U6848 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n9136), .Z(n5388) );
  XNOR2_X1 U6849 ( .A(n5388), .B(SI_15_), .ZN(n5385) );
  XNOR2_X1 U6850 ( .A(n5387), .B(n5385), .ZN(n6874) );
  NAND2_X1 U6851 ( .A1(n6874), .A2(n9137), .ZN(n5368) );
  INV_X1 U6852 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U6853 ( .A1(n5364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5365) );
  XNOR2_X1 U6854 ( .A(n5365), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9431) );
  INV_X1 U6855 ( .A(n9431), .ZN(n9437) );
  OAI22_X1 U6856 ( .A1(n5394), .A2(n6875), .B1(n6631), .B2(n9437), .ZN(n5366)
         );
  INV_X1 U6857 ( .A(n5366), .ZN(n5367) );
  NAND2_X1 U6858 ( .A1(n7817), .A2(n5639), .ZN(n5378) );
  NOR2_X1 U6859 ( .A1(n5369), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5370) );
  OR2_X1 U6860 ( .A1(n5398), .A2(n5370), .ZN(n9128) );
  OR2_X1 U6861 ( .A1(n4319), .A2(n9128), .ZN(n5376) );
  INV_X1 U6862 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7812) );
  OR2_X1 U6863 ( .A1(n5075), .A2(n7812), .ZN(n5375) );
  INV_X1 U6864 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6865 ( .A1(n5738), .A2(n5371), .ZN(n5374) );
  INV_X1 U6866 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5372) );
  OR2_X1 U6867 ( .A1(n7862), .A2(n5372), .ZN(n5373) );
  NAND4_X1 U6868 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n9702)
         );
  NAND2_X1 U6869 ( .A1(n9702), .A2(n5697), .ZN(n5377) );
  NAND2_X1 U6870 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  XNOR2_X1 U6871 ( .A(n5379), .B(n6482), .ZN(n5383) );
  NAND2_X1 U6872 ( .A1(n7817), .A2(n5697), .ZN(n5382) );
  NAND2_X1 U6873 ( .A1(n5206), .A2(n9702), .ZN(n5381) );
  NAND2_X1 U6874 ( .A1(n5382), .A2(n5381), .ZN(n9120) );
  NAND2_X1 U6875 ( .A1(n9121), .A2(n9120), .ZN(n9031) );
  INV_X1 U6876 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6877 ( .A1(n5387), .A2(n5386), .ZN(n5390) );
  NAND2_X1 U6878 ( .A1(n5388), .A2(SI_15_), .ZN(n5389) );
  NAND2_X1 U6879 ( .A1(n5390), .A2(n5389), .ZN(n5418) );
  MUX2_X1 U6880 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n9136), .Z(n5419) );
  XNOR2_X1 U6881 ( .A(n5419), .B(SI_16_), .ZN(n5416) );
  XNOR2_X1 U6882 ( .A(n5418), .B(n5416), .ZN(n6967) );
  NAND2_X1 U6883 ( .A1(n6967), .A2(n9137), .ZN(n5397) );
  INV_X1 U6884 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U6885 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5393) );
  XNOR2_X1 U6886 ( .A(n5393), .B(n5392), .ZN(n9449) );
  OAI22_X1 U6887 ( .A1(n5394), .A2(n6968), .B1(n6631), .B2(n9449), .ZN(n5395)
         );
  INV_X1 U6888 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U6889 ( .A1(n9719), .A2(n5682), .ZN(n5407) );
  OR2_X1 U6890 ( .A1(n5398), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6891 ( .A1(n5399), .A2(n5429), .ZN(n9711) );
  OR2_X1 U6892 ( .A1(n9711), .A2(n4320), .ZN(n5405) );
  NAND2_X1 U6893 ( .A1(n7859), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5404) );
  INV_X1 U6894 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5400) );
  OR2_X1 U6895 ( .A1(n5738), .A2(n5400), .ZN(n5403) );
  INV_X1 U6896 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5401) );
  OR2_X1 U6897 ( .A1(n7862), .A2(n5401), .ZN(n5402) );
  NAND4_X1 U6898 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n9690)
         );
  NAND2_X1 U6899 ( .A1(n9690), .A2(n5697), .ZN(n5406) );
  NAND2_X1 U6900 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  XNOR2_X1 U6901 ( .A(n5408), .B(n5694), .ZN(n5410) );
  AND2_X1 U6902 ( .A1(n5206), .A2(n9690), .ZN(n5409) );
  AOI21_X1 U6903 ( .B1(n9719), .B2(n5697), .A(n5409), .ZN(n5411) );
  NAND2_X1 U6904 ( .A1(n5410), .A2(n5411), .ZN(n5415) );
  INV_X1 U6905 ( .A(n5410), .ZN(n5413) );
  INV_X1 U6906 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6907 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  AND2_X1 U6908 ( .A1(n5415), .A2(n5414), .ZN(n9033) );
  NAND2_X1 U6909 ( .A1(n9030), .A2(n5415), .ZN(n9042) );
  INV_X1 U6910 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U6911 ( .A1(n5418), .A2(n5417), .ZN(n5421) );
  NAND2_X1 U6912 ( .A1(n5419), .A2(SI_16_), .ZN(n5420) );
  INV_X1 U6913 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7035) );
  INV_X1 U6914 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7033) );
  MUX2_X1 U6915 ( .A(n7035), .B(n7033), .S(n9136), .Z(n5423) );
  INV_X1 U6916 ( .A(SI_17_), .ZN(n5422) );
  NAND2_X1 U6917 ( .A1(n5423), .A2(n5422), .ZN(n5444) );
  INV_X1 U6918 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U6919 ( .A1(n5424), .A2(SI_17_), .ZN(n5425) );
  NAND2_X1 U6920 ( .A1(n5444), .A2(n5425), .ZN(n5443) );
  XNOR2_X1 U6921 ( .A(n5442), .B(n5443), .ZN(n7032) );
  NAND2_X1 U6922 ( .A1(n7032), .A2(n9137), .ZN(n5428) );
  XNOR2_X1 U6923 ( .A(n5426), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U6924 ( .A1(n5060), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5061), .B2(
        n9463), .ZN(n5427) );
  NAND2_X1 U6925 ( .A1(n6271), .A2(n5682), .ZN(n5435) );
  NAND2_X1 U6926 ( .A1(n5104), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5433) );
  INV_X1 U6927 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9469) );
  OR2_X1 U6928 ( .A1(n5075), .A2(n9469), .ZN(n5432) );
  INV_X1 U6929 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9450) );
  OR2_X1 U6930 ( .A1(n5738), .A2(n9450), .ZN(n5431) );
  INV_X1 U6931 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9045) );
  AOI21_X1 U6932 ( .B1(n5429), .B2(n9045), .A(n5449), .ZN(n9694) );
  INV_X1 U6933 ( .A(n9694), .ZN(n9047) );
  OR2_X1 U6934 ( .A1(n4319), .A2(n9047), .ZN(n5430) );
  NAND4_X1 U6935 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n9703)
         );
  NAND2_X1 U6936 ( .A1(n9703), .A2(n5697), .ZN(n5434) );
  NAND2_X1 U6937 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  XNOR2_X1 U6938 ( .A(n5436), .B(n6482), .ZN(n5438) );
  AND2_X1 U6939 ( .A1(n5206), .A2(n9703), .ZN(n5437) );
  AOI21_X1 U6940 ( .B1(n6271), .B2(n5697), .A(n5437), .ZN(n5439) );
  XNOR2_X1 U6941 ( .A(n5438), .B(n5439), .ZN(n9043) );
  NAND2_X1 U6942 ( .A1(n9042), .A2(n9043), .ZN(n9041) );
  INV_X1 U6943 ( .A(n5438), .ZN(n5440) );
  NAND2_X1 U6944 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  NAND2_X1 U6945 ( .A1(n9041), .A2(n5441), .ZN(n5460) );
  INV_X1 U6946 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7140) );
  INV_X1 U6947 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7105) );
  MUX2_X1 U6948 ( .A(n7140), .B(n7105), .S(n9136), .Z(n5462) );
  XNOR2_X1 U6949 ( .A(n5462), .B(SI_18_), .ZN(n5461) );
  XNOR2_X1 U6950 ( .A(n5465), .B(n5461), .ZN(n7104) );
  NAND2_X1 U6951 ( .A1(n7104), .A2(n9137), .ZN(n5448) );
  NAND2_X1 U6952 ( .A1(n5445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U6953 ( .A(n5446), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9486) );
  AOI22_X1 U6954 ( .A1(n9486), .A2(n5061), .B1(n5060), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6955 ( .A1(n9781), .A2(n5682), .ZN(n5455) );
  NAND2_X1 U6956 ( .A1(n5104), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5453) );
  INV_X1 U6957 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9473) );
  OR2_X1 U6958 ( .A1(n5075), .A2(n9473), .ZN(n5452) );
  INV_X1 U6959 ( .A(n5472), .ZN(n5474) );
  OAI21_X1 U6960 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(n5449), .A(n5474), .ZN(
        n9671) );
  OR2_X1 U6961 ( .A1(n4320), .A2(n9671), .ZN(n5451) );
  INV_X1 U6962 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6402) );
  OR2_X1 U6963 ( .A1(n5738), .A2(n6402), .ZN(n5450) );
  NAND4_X1 U6964 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n9689)
         );
  NAND2_X1 U6965 ( .A1(n9689), .A2(n5697), .ZN(n5454) );
  NAND2_X1 U6966 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  XNOR2_X1 U6967 ( .A(n5456), .B(n5694), .ZN(n5459) );
  NAND2_X1 U6968 ( .A1(n9781), .A2(n5697), .ZN(n5458) );
  NAND2_X1 U6969 ( .A1(n5206), .A2(n9689), .ZN(n5457) );
  NAND2_X1 U6970 ( .A1(n5458), .A2(n5457), .ZN(n9098) );
  INV_X1 U6971 ( .A(n5461), .ZN(n5464) );
  INV_X1 U6972 ( .A(n5462), .ZN(n5463) );
  INV_X1 U6973 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7276) );
  INV_X1 U6974 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7278) );
  MUX2_X1 U6975 ( .A(n7276), .B(n7278), .S(n9136), .Z(n5467) );
  INV_X1 U6976 ( .A(SI_19_), .ZN(n5466) );
  NAND2_X1 U6977 ( .A1(n5467), .A2(n5466), .ZN(n5491) );
  INV_X1 U6978 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U6979 ( .A1(n5468), .A2(SI_19_), .ZN(n5469) );
  NAND2_X1 U6980 ( .A1(n5491), .A2(n5469), .ZN(n5492) );
  XNOR2_X1 U6981 ( .A(n5493), .B(n5492), .ZN(n7275) );
  NAND2_X1 U6982 ( .A1(n7275), .A2(n9137), .ZN(n5471) );
  AOI22_X1 U6983 ( .A1(n9496), .A2(n5061), .B1(n5060), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6984 ( .A1(n9777), .A2(n5682), .ZN(n5482) );
  NAND2_X1 U6985 ( .A1(n5104), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5480) );
  INV_X1 U6986 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9657) );
  OR2_X1 U6987 ( .A1(n5075), .A2(n9657), .ZN(n5479) );
  INV_X1 U6988 ( .A(n5501), .ZN(n5503) );
  INV_X1 U6989 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6990 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  NAND2_X1 U6991 ( .A1(n5503), .A2(n5475), .ZN(n9656) );
  OR2_X1 U6992 ( .A1(n4320), .A2(n9656), .ZN(n5478) );
  INV_X1 U6993 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5476) );
  OR2_X1 U6994 ( .A1(n5738), .A2(n5476), .ZN(n5477) );
  NAND4_X1 U6995 ( .A1(n5480), .A2(n5479), .A3(n5478), .A4(n5477), .ZN(n9678)
         );
  NAND2_X1 U6996 ( .A1(n9678), .A2(n5697), .ZN(n5481) );
  NAND2_X1 U6997 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  XNOR2_X1 U6998 ( .A(n5483), .B(n5694), .ZN(n5485) );
  AND2_X1 U6999 ( .A1(n5206), .A2(n9678), .ZN(n5484) );
  AOI21_X1 U7000 ( .B1(n9777), .B2(n5697), .A(n5484), .ZN(n5486) );
  NAND2_X1 U7001 ( .A1(n5485), .A2(n5486), .ZN(n5490) );
  INV_X1 U7002 ( .A(n5485), .ZN(n5488) );
  INV_X1 U7003 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U7004 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  NAND2_X1 U7005 ( .A1(n8995), .A2(n5490), .ZN(n9058) );
  INV_X1 U7006 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7353) );
  INV_X1 U7007 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7394) );
  MUX2_X1 U7008 ( .A(n7353), .B(n7394), .S(n9136), .Z(n5495) );
  INV_X1 U7009 ( .A(SI_20_), .ZN(n5494) );
  NAND2_X1 U7010 ( .A1(n5495), .A2(n5494), .ZN(n5515) );
  INV_X1 U7011 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U7012 ( .A1(n5496), .A2(SI_20_), .ZN(n5497) );
  XNOR2_X1 U7013 ( .A(n5514), .B(n5513), .ZN(n7352) );
  NAND2_X1 U7014 ( .A1(n7352), .A2(n9137), .ZN(n5499) );
  NAND2_X1 U7015 ( .A1(n5060), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7016 ( .A1(n7859), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5509) );
  INV_X1 U7017 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5500) );
  OR2_X1 U7018 ( .A1(n5738), .A2(n5500), .ZN(n5508) );
  INV_X1 U7019 ( .A(n5520), .ZN(n5522) );
  INV_X1 U7020 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7021 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  NAND2_X1 U7022 ( .A1(n5522), .A2(n5504), .ZN(n9645) );
  OR2_X1 U7023 ( .A1(n4319), .A2(n9645), .ZN(n5507) );
  INV_X1 U7024 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5505) );
  OR2_X1 U7025 ( .A1(n7862), .A2(n5505), .ZN(n5506) );
  NAND4_X1 U7026 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n9401)
         );
  AOI22_X1 U7027 ( .A1(n9772), .A2(n5697), .B1(n5206), .B2(n9401), .ZN(n5533)
         );
  NAND2_X1 U7028 ( .A1(n9772), .A2(n5682), .ZN(n5511) );
  NAND2_X1 U7029 ( .A1(n9401), .A2(n5697), .ZN(n5510) );
  NAND2_X1 U7030 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  XNOR2_X1 U7031 ( .A(n5512), .B(n5694), .ZN(n5534) );
  XOR2_X1 U7032 ( .A(n5533), .B(n5534), .Z(n9059) );
  INV_X1 U7033 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7411) );
  INV_X1 U7034 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7437) );
  MUX2_X1 U7035 ( .A(n7411), .B(n7437), .S(n9136), .Z(n5540) );
  XNOR2_X1 U7036 ( .A(n5540), .B(SI_21_), .ZN(n5539) );
  XNOR2_X1 U7037 ( .A(n5544), .B(n5539), .ZN(n7410) );
  NAND2_X1 U7038 ( .A1(n7410), .A2(n9137), .ZN(n5518) );
  NAND2_X1 U7039 ( .A1(n5060), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7040 ( .A1(n9767), .A2(n5682), .ZN(n5530) );
  NAND2_X1 U7041 ( .A1(n7859), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5528) );
  INV_X1 U7042 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5519) );
  OR2_X1 U7043 ( .A1(n5738), .A2(n5519), .ZN(n5527) );
  INV_X1 U7044 ( .A(n5551), .ZN(n5552) );
  INV_X1 U7045 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7046 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  NAND2_X1 U7047 ( .A1(n5552), .A2(n5523), .ZN(n9629) );
  OR2_X1 U7048 ( .A1(n4319), .A2(n9629), .ZN(n5526) );
  INV_X1 U7049 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5524) );
  OR2_X1 U7050 ( .A1(n7862), .A2(n5524), .ZN(n5525) );
  NAND4_X1 U7051 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n9614)
         );
  NAND2_X1 U7052 ( .A1(n9614), .A2(n5697), .ZN(n5529) );
  NAND2_X1 U7053 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  XNOR2_X1 U7054 ( .A(n5531), .B(n6482), .ZN(n5538) );
  AND2_X1 U7055 ( .A1(n5206), .A2(n9614), .ZN(n5532) );
  AOI21_X1 U7056 ( .B1(n9767), .B2(n5697), .A(n5532), .ZN(n5536) );
  XNOR2_X1 U7057 ( .A(n5538), .B(n5536), .ZN(n9003) );
  NAND2_X1 U7058 ( .A1(n5534), .A2(n5533), .ZN(n9004) );
  INV_X1 U7059 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7060 ( .A1(n5538), .A2(n5537), .ZN(n8974) );
  INV_X1 U7061 ( .A(n5539), .ZN(n5543) );
  INV_X1 U7062 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7063 ( .A1(n5541), .A2(SI_21_), .ZN(n5542) );
  INV_X1 U7064 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7603) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U7066 ( .A(n7603), .B(n7600), .S(n9136), .Z(n5546) );
  INV_X1 U7067 ( .A(SI_22_), .ZN(n5545) );
  NAND2_X1 U7068 ( .A1(n5546), .A2(n5545), .ZN(n5565) );
  INV_X1 U7069 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7070 ( .A1(n5547), .A2(SI_22_), .ZN(n5548) );
  NAND2_X1 U7071 ( .A1(n5565), .A2(n5548), .ZN(n5566) );
  NAND2_X1 U7072 ( .A1(n7599), .A2(n9137), .ZN(n5550) );
  NAND2_X1 U7073 ( .A1(n5060), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7074 ( .A1(n9762), .A2(n5697), .ZN(n5561) );
  NAND2_X1 U7075 ( .A1(n5104), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5559) );
  INV_X1 U7076 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9608) );
  OR2_X1 U7077 ( .A1(n5075), .A2(n9608), .ZN(n5558) );
  INV_X1 U7078 ( .A(n5575), .ZN(n5554) );
  INV_X1 U7079 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U7080 ( .A1(n5552), .A2(n9078), .ZN(n5553) );
  NAND2_X1 U7081 ( .A1(n5554), .A2(n5553), .ZN(n9607) );
  OR2_X1 U7082 ( .A1(n4320), .A2(n9607), .ZN(n5557) );
  INV_X1 U7083 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5555) );
  OR2_X1 U7084 ( .A1(n5738), .A2(n5555), .ZN(n5556) );
  NAND4_X1 U7085 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n9400)
         );
  NAND2_X1 U7086 ( .A1(n5206), .A2(n9400), .ZN(n5560) );
  NAND2_X1 U7087 ( .A1(n8974), .A2(n9076), .ZN(n5585) );
  NAND2_X1 U7088 ( .A1(n9762), .A2(n5682), .ZN(n5563) );
  NAND2_X1 U7089 ( .A1(n9400), .A2(n5697), .ZN(n5562) );
  NAND2_X1 U7090 ( .A1(n5563), .A2(n5562), .ZN(n5564) );
  XNOR2_X1 U7091 ( .A(n5564), .B(n5694), .ZN(n5586) );
  NAND2_X1 U7092 ( .A1(n5586), .A2(n8974), .ZN(n8973) );
  INV_X1 U7093 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7610) );
  INV_X1 U7094 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7606) );
  MUX2_X1 U7095 ( .A(n7610), .B(n7606), .S(n9136), .Z(n5569) );
  INV_X1 U7096 ( .A(SI_23_), .ZN(n5568) );
  NAND2_X1 U7097 ( .A1(n5569), .A2(n5568), .ZN(n5596) );
  INV_X1 U7098 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7099 ( .A1(n5570), .A2(SI_23_), .ZN(n5571) );
  AND2_X1 U7100 ( .A1(n5596), .A2(n5571), .ZN(n5594) );
  XNOR2_X1 U7101 ( .A(n5595), .B(n5594), .ZN(n7608) );
  NAND2_X1 U7102 ( .A1(n7608), .A2(n9137), .ZN(n5573) );
  NAND2_X1 U7103 ( .A1(n5060), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7104 ( .A1(n9757), .A2(n5682), .ZN(n5582) );
  NAND2_X1 U7105 ( .A1(n7859), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5580) );
  INV_X1 U7106 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5574) );
  OR2_X1 U7107 ( .A1(n5738), .A2(n5574), .ZN(n5579) );
  NAND2_X1 U7108 ( .A1(n5575), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5604) );
  OAI21_X1 U7109 ( .B1(n5575), .B2(P1_REG3_REG_23__SCAN_IN), .A(n5604), .ZN(
        n9596) );
  OR2_X1 U7110 ( .A1(n4319), .A2(n9596), .ZN(n5578) );
  INV_X1 U7111 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5576) );
  OR2_X1 U7112 ( .A1(n7862), .A2(n5576), .ZN(n5577) );
  NAND4_X1 U7113 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n9615)
         );
  NAND2_X1 U7114 ( .A1(n9615), .A2(n5697), .ZN(n5581) );
  NAND2_X1 U7115 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  XNOR2_X1 U7116 ( .A(n5583), .B(n5694), .ZN(n5588) );
  AND2_X1 U7117 ( .A1(n5206), .A2(n9615), .ZN(n5584) );
  AOI21_X1 U7118 ( .B1(n9757), .B2(n5697), .A(n5584), .ZN(n5589) );
  NOR2_X1 U7119 ( .A1(n5588), .A2(n5589), .ZN(n8971) );
  AOI21_X1 U7120 ( .B1(n5585), .B2(n8973), .A(n8971), .ZN(n5593) );
  INV_X1 U7121 ( .A(n5586), .ZN(n8975) );
  INV_X1 U7122 ( .A(n9076), .ZN(n5587) );
  NOR3_X1 U7123 ( .A1(n8971), .A2(n8975), .A3(n5587), .ZN(n5592) );
  INV_X1 U7124 ( .A(n5588), .ZN(n5591) );
  INV_X1 U7125 ( .A(n5589), .ZN(n5590) );
  INV_X1 U7126 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7839) );
  INV_X1 U7127 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7752) );
  MUX2_X1 U7128 ( .A(n7839), .B(n7752), .S(n9136), .Z(n5598) );
  INV_X1 U7129 ( .A(SI_24_), .ZN(n5597) );
  NAND2_X1 U7130 ( .A1(n5598), .A2(n5597), .ZN(n5622) );
  INV_X1 U7131 ( .A(n5598), .ZN(n5599) );
  NAND2_X1 U7132 ( .A1(n5599), .A2(SI_24_), .ZN(n5600) );
  AND2_X1 U7133 ( .A1(n5622), .A2(n5600), .ZN(n5620) );
  XNOR2_X1 U7134 ( .A(n5621), .B(n5620), .ZN(n7751) );
  NAND2_X1 U7135 ( .A1(n7751), .A2(n9137), .ZN(n5602) );
  NAND2_X1 U7136 ( .A1(n5060), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7137 ( .A1(n9752), .A2(n5682), .ZN(n5611) );
  NAND2_X1 U7138 ( .A1(n7859), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5609) );
  INV_X1 U7139 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5603) );
  OR2_X1 U7140 ( .A1(n5738), .A2(n5603), .ZN(n5608) );
  INV_X1 U7141 ( .A(n5604), .ZN(n5605) );
  NAND2_X1 U7142 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5605), .ZN(n5631) );
  OAI21_X1 U7143 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n5605), .A(n5631), .ZN(
        n9579) );
  OR2_X1 U7144 ( .A1(n4320), .A2(n9579), .ZN(n5607) );
  INV_X1 U7145 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6310) );
  OR2_X1 U7146 ( .A1(n7862), .A2(n6310), .ZN(n5606) );
  NAND4_X1 U7147 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n9399)
         );
  NAND2_X1 U7148 ( .A1(n9399), .A2(n5697), .ZN(n5610) );
  NAND2_X1 U7149 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  XNOR2_X1 U7150 ( .A(n5612), .B(n5694), .ZN(n5614) );
  AND2_X1 U7151 ( .A1(n5206), .A2(n9399), .ZN(n5613) );
  AOI21_X1 U7152 ( .B1(n9752), .B2(n5697), .A(n5613), .ZN(n5615) );
  NAND2_X1 U7153 ( .A1(n5614), .A2(n5615), .ZN(n5619) );
  INV_X1 U7154 ( .A(n5614), .ZN(n5617) );
  INV_X1 U7155 ( .A(n5615), .ZN(n5616) );
  NAND2_X1 U7156 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  NAND2_X1 U7157 ( .A1(n5619), .A2(n5618), .ZN(n9051) );
  INV_X1 U7158 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7797) );
  INV_X1 U7159 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7799) );
  MUX2_X1 U7160 ( .A(n7797), .B(n7799), .S(n9136), .Z(n5624) );
  INV_X1 U7161 ( .A(SI_25_), .ZN(n5623) );
  NAND2_X1 U7162 ( .A1(n5624), .A2(n5623), .ZN(n5646) );
  INV_X1 U7163 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7164 ( .A1(n5625), .A2(SI_25_), .ZN(n5626) );
  AND2_X1 U7165 ( .A1(n5646), .A2(n5626), .ZN(n5644) );
  NAND2_X1 U7166 ( .A1(n5060), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7167 ( .A1(n7859), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5637) );
  INV_X1 U7168 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5629) );
  OR2_X1 U7169 ( .A1(n7862), .A2(n5629), .ZN(n5636) );
  INV_X1 U7170 ( .A(n5631), .ZN(n5630) );
  NAND2_X1 U7171 ( .A1(n5630), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5656) );
  INV_X1 U7172 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U7173 ( .A1(n9025), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U7174 ( .A1(n5656), .A2(n5632), .ZN(n9557) );
  OR2_X1 U7175 ( .A1(n4319), .A2(n9557), .ZN(n5635) );
  INV_X1 U7176 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5633) );
  OR2_X1 U7177 ( .A1(n5738), .A2(n5633), .ZN(n5634) );
  NAND4_X1 U7178 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n9574)
         );
  AND2_X1 U7179 ( .A1(n5206), .A2(n9574), .ZN(n5638) );
  AOI21_X1 U7180 ( .B1(n9746), .B2(n5697), .A(n5638), .ZN(n5641) );
  AOI22_X1 U7181 ( .A1(n9746), .A2(n5639), .B1(n5697), .B2(n9574), .ZN(n5640)
         );
  XNOR2_X1 U7182 ( .A(n5640), .B(n5694), .ZN(n5643) );
  XOR2_X1 U7183 ( .A(n5641), .B(n5643), .Z(n9024) );
  INV_X1 U7184 ( .A(n5641), .ZN(n5642) );
  INV_X1 U7185 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7803) );
  INV_X1 U7186 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7805) );
  MUX2_X1 U7187 ( .A(n7803), .B(n7805), .S(n9136), .Z(n5648) );
  INV_X1 U7188 ( .A(SI_26_), .ZN(n6407) );
  NAND2_X1 U7189 ( .A1(n5648), .A2(n6407), .ZN(n5672) );
  INV_X1 U7190 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U7191 ( .A1(n5649), .A2(SI_26_), .ZN(n5650) );
  AND2_X1 U7192 ( .A1(n5672), .A2(n5650), .ZN(n5670) );
  NAND2_X1 U7193 ( .A1(n5060), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7194 ( .A1(n9742), .A2(n5682), .ZN(n5663) );
  NAND2_X1 U7195 ( .A1(n7859), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5661) );
  INV_X1 U7196 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5653) );
  OR2_X1 U7197 ( .A1(n7862), .A2(n5653), .ZN(n5660) );
  INV_X1 U7198 ( .A(n5656), .ZN(n5654) );
  NAND2_X1 U7199 ( .A1(n5654), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5686) );
  INV_X1 U7200 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7201 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  NAND2_X1 U7202 ( .A1(n5686), .A2(n5657), .ZN(n9547) );
  OR2_X1 U7203 ( .A1(n4320), .A2(n9547), .ZN(n5659) );
  INV_X1 U7204 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6420) );
  OR2_X1 U7205 ( .A1(n5738), .A2(n6420), .ZN(n5658) );
  NAND4_X1 U7206 ( .A1(n5661), .A2(n5660), .A3(n5659), .A4(n5658), .ZN(n9398)
         );
  NAND2_X1 U7207 ( .A1(n9398), .A2(n5697), .ZN(n5662) );
  NAND2_X1 U7208 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  XNOR2_X1 U7209 ( .A(n5664), .B(n5694), .ZN(n5666) );
  AND2_X1 U7210 ( .A1(n5206), .A2(n9398), .ZN(n5665) );
  AOI21_X1 U7211 ( .B1(n9742), .B2(n5697), .A(n5665), .ZN(n5667) );
  XNOR2_X1 U7212 ( .A(n5666), .B(n5667), .ZN(n9109) );
  INV_X1 U7213 ( .A(n5666), .ZN(n5669) );
  INV_X1 U7214 ( .A(n5667), .ZN(n5668) );
  INV_X1 U7215 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6099) );
  INV_X1 U7216 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7826) );
  MUX2_X1 U7217 ( .A(n6099), .B(n7826), .S(n9136), .Z(n5674) );
  INV_X1 U7218 ( .A(SI_27_), .ZN(n5673) );
  NAND2_X1 U7219 ( .A1(n5674), .A2(n5673), .ZN(n6111) );
  INV_X1 U7220 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U7221 ( .A1(n5675), .A2(SI_27_), .ZN(n5676) );
  AND2_X1 U7222 ( .A1(n6111), .A2(n5676), .ZN(n5677) );
  NAND2_X1 U7223 ( .A1(n5060), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7224 ( .A1(n6298), .A2(n5682), .ZN(n5693) );
  NAND2_X1 U7225 ( .A1(n7859), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5691) );
  INV_X1 U7226 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5683) );
  OR2_X1 U7227 ( .A1(n5738), .A2(n5683), .ZN(n5690) );
  INV_X1 U7228 ( .A(n5686), .ZN(n5684) );
  NAND2_X1 U7229 ( .A1(n5684), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5736) );
  INV_X1 U7230 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7231 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  NAND2_X1 U7232 ( .A1(n5736), .A2(n5687), .ZN(n7954) );
  OR2_X1 U7233 ( .A1(n4319), .A2(n7954), .ZN(n5689) );
  OR2_X1 U7234 ( .A1(n7862), .A2(n6305), .ZN(n5688) );
  NAND4_X1 U7235 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n9397)
         );
  NAND2_X1 U7236 ( .A1(n9397), .A2(n5697), .ZN(n5692) );
  NAND2_X1 U7237 ( .A1(n5693), .A2(n5692), .ZN(n5695) );
  XNOR2_X1 U7238 ( .A(n5695), .B(n5694), .ZN(n5699) );
  AND2_X1 U7239 ( .A1(n5206), .A2(n9397), .ZN(n5696) );
  AOI21_X1 U7240 ( .B1(n6298), .B2(n5697), .A(n5696), .ZN(n5698) );
  NAND2_X1 U7241 ( .A1(n5699), .A2(n5698), .ZN(n6494) );
  OAI21_X1 U7242 ( .B1(n5699), .B2(n5698), .A(n6494), .ZN(n5702) );
  OAI21_X1 U7243 ( .B1(n9108), .B2(n5701), .A(n5702), .ZN(n5700) );
  INV_X1 U7244 ( .A(n5700), .ZN(n5725) );
  INV_X1 U7245 ( .A(n6267), .ZN(n9242) );
  AND2_X1 U7246 ( .A1(n9376), .A2(n9204), .ZN(n7246) );
  NAND2_X1 U7247 ( .A1(n9242), .A2(n7246), .ZN(n9996) );
  NAND2_X1 U7248 ( .A1(n9388), .A2(n9375), .ZN(n5730) );
  AND2_X1 U7249 ( .A1(n9996), .A2(n5730), .ZN(n5743) );
  NAND2_X1 U7250 ( .A1(n5704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U7251 ( .A(n5706), .B(n5705), .ZN(n6632) );
  AND2_X1 U7252 ( .A1(n6632), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6626) );
  INV_X1 U7253 ( .A(n5707), .ZN(n7801) );
  NAND2_X1 U7254 ( .A1(n7801), .A2(P1_B_REG_SCAN_IN), .ZN(n5709) );
  INV_X1 U7255 ( .A(n5708), .ZN(n7753) );
  MUX2_X1 U7256 ( .A(P1_B_REG_SCAN_IN), .B(n5709), .S(n7753), .Z(n5710) );
  NAND2_X1 U7257 ( .A1(n5710), .A2(n5711), .ZN(n6670) );
  INV_X1 U7258 ( .A(n6670), .ZN(n5722) );
  INV_X1 U7259 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5712) );
  INV_X1 U7260 ( .A(n5711), .ZN(n7807) );
  AND2_X1 U7261 ( .A1(n7807), .A2(n7753), .ZN(n6672) );
  AOI21_X1 U7262 ( .B1(n5722), .B2(n5712), .A(n6672), .ZN(n6904) );
  INV_X1 U7263 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5713) );
  AND2_X1 U7264 ( .A1(n7807), .A2(n7801), .ZN(n6674) );
  AOI21_X1 U7265 ( .B1(n5722), .B2(n5713), .A(n6674), .ZN(n7221) );
  NOR4_X1 U7266 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5717) );
  NOR4_X1 U7267 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5716) );
  NOR4_X1 U7268 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5715) );
  NOR4_X1 U7269 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5714) );
  NAND4_X1 U7270 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n5724)
         );
  NOR2_X1 U7271 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .ZN(
        n5721) );
  NOR4_X1 U7272 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5720) );
  NOR4_X1 U7273 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5719) );
  NOR4_X1 U7274 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5718) );
  NAND4_X1 U7275 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n5723)
         );
  OAI21_X1 U7276 ( .B1(n5724), .B2(n5723), .A(n5722), .ZN(n6301) );
  AND3_X1 U7277 ( .A1(n6904), .A2(n7221), .A3(n6301), .ZN(n5731) );
  INV_X1 U7278 ( .A(n5731), .ZN(n5746) );
  INV_X1 U7279 ( .A(n7246), .ZN(n6266) );
  OR2_X1 U7280 ( .A1(n6266), .A2(n9197), .ZN(n7228) );
  INV_X1 U7281 ( .A(n7228), .ZN(n5726) );
  NAND2_X1 U7282 ( .A1(n9380), .A2(n5726), .ZN(n5727) );
  NOR2_X1 U7283 ( .A1(n5746), .A2(n5727), .ZN(n5729) );
  NAND2_X1 U7284 ( .A1(n9197), .A2(n7246), .ZN(n9670) );
  NOR2_X1 U7285 ( .A1(n9384), .A2(n9670), .ZN(n6303) );
  OR2_X1 U7286 ( .A1(n5729), .A2(n9897), .ZN(n9082) );
  INV_X1 U7287 ( .A(n5730), .ZN(n9194) );
  AND2_X1 U7288 ( .A1(n6267), .A2(n9194), .ZN(n9381) );
  NAND2_X1 U7289 ( .A1(n9381), .A2(n9380), .ZN(n5745) );
  INV_X1 U7290 ( .A(n5745), .ZN(n5732) );
  NAND2_X1 U7291 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  OR2_X1 U7292 ( .A1(n5733), .A2(n6679), .ZN(n9126) );
  NOR2_X1 U7293 ( .A1(n9126), .A2(n9564), .ZN(n5750) );
  INV_X1 U7294 ( .A(n6679), .ZN(n7828) );
  NAND2_X1 U7295 ( .A1(n7859), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5742) );
  INV_X1 U7296 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5734) );
  OR2_X1 U7297 ( .A1(n7862), .A2(n5734), .ZN(n5741) );
  INV_X1 U7298 ( .A(n5736), .ZN(n5735) );
  NAND2_X1 U7299 ( .A1(n5735), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7848) );
  INV_X1 U7300 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U7301 ( .A1(n5736), .A2(n6497), .ZN(n5737) );
  NAND2_X1 U7302 ( .A1(n7848), .A2(n5737), .ZN(n9523) );
  OR2_X1 U7303 ( .A1(n4320), .A2(n9523), .ZN(n5740) );
  INV_X1 U7304 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6344) );
  OR2_X1 U7305 ( .A1(n5738), .A2(n6344), .ZN(n5739) );
  INV_X1 U7306 ( .A(n5743), .ZN(n5744) );
  NAND3_X1 U7307 ( .A1(n5745), .A2(n7228), .A3(n5744), .ZN(n5747) );
  NAND2_X1 U7308 ( .A1(n5747), .A2(n5746), .ZN(n6789) );
  NAND2_X1 U7309 ( .A1(n9242), .A2(n9194), .ZN(n6300) );
  NAND4_X1 U7310 ( .A1(n6789), .A2(n6300), .A3(n6628), .A4(n6632), .ZN(n5748)
         );
  OAI22_X1 U7311 ( .A1(n9115), .A2(n7866), .B1(n9129), .B2(n7954), .ZN(n5749)
         );
  AOI211_X1 U7312 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n5750), 
        .B(n5749), .ZN(n5751) );
  NAND3_X1 U7313 ( .A1(n5752), .A2(n4903), .A3(n5751), .ZN(P1_U3214) );
  INV_X1 U7314 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5994) );
  INV_X1 U7315 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5755) );
  INV_X1 U7316 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5756) );
  NOR2_X1 U7317 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5757) );
  INV_X1 U7318 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5758) );
  INV_X1 U7319 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5759) );
  INV_X1 U7320 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5763) );
  NOR2_X1 U7321 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5764) );
  INV_X1 U7322 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5783) );
  AND2_X2 U7323 ( .A1(n8202), .A2(n5769), .ZN(n5857) );
  NAND2_X1 U7324 ( .A1(n7985), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5782) );
  AND2_X2 U7325 ( .A1(n8202), .A2(n5777), .ZN(n5858) );
  INV_X2 U7326 ( .A(n5790), .ZN(n7986) );
  NAND2_X1 U7327 ( .A1(n7986), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5781) );
  INV_X1 U7328 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5773) );
  INV_X1 U7329 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5775) );
  INV_X1 U7330 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7743) );
  NAND2_X1 U7331 ( .A1(n5792), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7332 ( .A1(n5933), .A2(n5776), .ZN(n8749) );
  NAND2_X1 U7333 ( .A1(n6132), .A2(n8749), .ZN(n5780) );
  AND2_X4 U7334 ( .A1(n5778), .A2(n5777), .ZN(n6118) );
  NAND2_X1 U7335 ( .A1(n6118), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5779) );
  NAND4_X1 U7336 ( .A1(n5782), .A2(n5781), .A3(n5780), .A4(n5779), .ZN(n8759)
         );
  NAND2_X2 U7337 ( .A1(n5821), .A2(n6650), .ZN(n7984) );
  NAND2_X1 U7338 ( .A1(n6783), .A2(n7975), .ZN(n5789) );
  NAND2_X1 U7339 ( .A1(n5968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7340 ( .A1(n5928), .A2(n4598), .ZN(n5798) );
  NAND2_X1 U7341 ( .A1(n5798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U7342 ( .A(n5787), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6616) );
  AOI22_X1 U7343 ( .A1(n6013), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6012), .B2(
        n6616), .ZN(n5788) );
  INV_X1 U7344 ( .A(n8941), .ZN(n5926) );
  NAND2_X1 U7345 ( .A1(n7986), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7346 ( .A1(n6118), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7347 ( .A1(n5916), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7348 ( .A1(n5792), .A2(n5791), .ZN(n8765) );
  NAND2_X1 U7349 ( .A1(n6132), .A2(n8765), .ZN(n5794) );
  NAND2_X1 U7350 ( .A1(n7985), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7351 ( .A1(n6705), .A2(n7975), .ZN(n5801) );
  INV_X1 U7352 ( .A(n5928), .ZN(n5797) );
  NAND2_X1 U7353 ( .A1(n5797), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5799) );
  AND2_X1 U7354 ( .A1(n5799), .A2(n5798), .ZN(n6614) );
  AOI22_X1 U7355 ( .A1(n6013), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6012), .B2(
        n6614), .ZN(n5800) );
  NAND2_X1 U7356 ( .A1(n5801), .A2(n5800), .ZN(n8769) );
  INV_X1 U7357 ( .A(n8769), .ZN(n10073) );
  OR2_X1 U7358 ( .A1(n7984), .A2(n6677), .ZN(n5806) );
  OR2_X1 U7359 ( .A1(n7983), .A2(n6676), .ZN(n5805) );
  NAND2_X1 U7360 ( .A1(n5896), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  XNOR2_X1 U7361 ( .A(n5803), .B(n5802), .ZN(n6675) );
  OR2_X1 U7362 ( .A1(n5821), .A2(n6675), .ZN(n5804) );
  NAND2_X1 U7363 ( .A1(n7986), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7364 ( .A1(n7985), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7365 ( .A1(n5890), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7366 ( .A1(n5902), .A2(n5807), .ZN(n7717) );
  NAND2_X1 U7367 ( .A1(n6132), .A2(n7717), .ZN(n5809) );
  NAND2_X1 U7368 ( .A1(n6118), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7369 ( .A1(n5824), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7370 ( .A1(n6118), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7371 ( .A1(n5857), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5812) );
  OR2_X1 U7372 ( .A1(n5821), .A2(n7010), .ZN(n5815) );
  NAND2_X1 U7373 ( .A1(n6118), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7374 ( .A1(n5858), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7375 ( .A1(n5824), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7376 ( .A1(n5857), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7377 ( .A1(n6650), .A2(SI_0_), .ZN(n5820) );
  XNOR2_X1 U7378 ( .A(n5820), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8956) );
  MUX2_X1 U7379 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8956), .S(n5821), .Z(n7029) );
  NAND2_X1 U7380 ( .A1(n8392), .A2(n7029), .ZN(n7096) );
  NAND2_X1 U7381 ( .A1(n7097), .A2(n7096), .ZN(n5823) );
  INV_X1 U7382 ( .A(n6976), .ZN(n6977) );
  OR2_X1 U7383 ( .A1(n8390), .A2(n6977), .ZN(n5822) );
  NAND2_X1 U7384 ( .A1(n5823), .A2(n5822), .ZN(n7385) );
  NAND2_X1 U7385 ( .A1(n5824), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U7386 ( .A1(n5858), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7387 ( .A1(n6118), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7388 ( .A1(n5857), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5825) );
  INV_X1 U7389 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6656) );
  OR2_X1 U7390 ( .A1(n7983), .A2(n6656), .ZN(n5833) );
  OR2_X1 U7391 ( .A1(n7984), .A2(n6655), .ZN(n5832) );
  OR2_X1 U7392 ( .A1(n5821), .A2(n7038), .ZN(n5831) );
  OR2_X1 U7393 ( .A1(n8389), .A2(n7088), .ZN(n8045) );
  NAND2_X1 U7394 ( .A1(n8389), .A2(n7088), .ZN(n6147) );
  NAND2_X1 U7395 ( .A1(n8045), .A2(n6147), .ZN(n8041) );
  NAND2_X1 U7396 ( .A1(n7385), .A2(n8041), .ZN(n5835) );
  INV_X1 U7397 ( .A(n7088), .ZN(n7383) );
  OR2_X1 U7398 ( .A1(n8389), .A2(n7383), .ZN(n5834) );
  NAND2_X1 U7399 ( .A1(n5824), .A2(n6928), .ZN(n5839) );
  NAND2_X1 U7400 ( .A1(n5858), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7401 ( .A1(n6118), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7402 ( .A1(n5857), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5836) );
  OR2_X1 U7403 ( .A1(n7983), .A2(n6658), .ZN(n5844) );
  OR2_X1 U7404 ( .A1(n7984), .A2(n6657), .ZN(n5843) );
  NAND2_X1 U7405 ( .A1(n5840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7406 ( .A(n5841), .B(n5753), .ZN(n6939) );
  OR2_X1 U7407 ( .A1(n5821), .A2(n6939), .ZN(n5842) );
  OR2_X1 U7408 ( .A1(n8388), .A2(n7346), .ZN(n8052) );
  NAND2_X1 U7409 ( .A1(n8388), .A2(n7346), .ZN(n6148) );
  NAND2_X1 U7410 ( .A1(n8052), .A2(n6148), .ZN(n7204) );
  OR2_X1 U7411 ( .A1(n8388), .A2(n7212), .ZN(n7338) );
  NAND2_X1 U7412 ( .A1(n5858), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7413 ( .A1(n5857), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7414 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5845) );
  NAND2_X1 U7415 ( .A1(n5859), .A2(n5845), .ZN(n10034) );
  NAND2_X1 U7416 ( .A1(n5824), .A2(n10034), .ZN(n5847) );
  NAND2_X1 U7417 ( .A1(n6118), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5846) );
  NAND4_X1 U7418 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .ZN(n8387)
         );
  OR2_X1 U7419 ( .A1(n7984), .A2(n6651), .ZN(n5855) );
  OR2_X1 U7420 ( .A1(n7983), .A2(n6652), .ZN(n5854) );
  NAND2_X1 U7421 ( .A1(n5850), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  INV_X1 U7422 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U7423 ( .A(n5852), .B(n5851), .ZN(n7118) );
  OR2_X1 U7424 ( .A1(n5821), .A2(n7118), .ZN(n5853) );
  INV_X1 U7425 ( .A(n7875), .ZN(n10032) );
  OR2_X1 U7426 ( .A1(n8387), .A2(n10032), .ZN(n5856) );
  AND2_X1 U7427 ( .A1(n7338), .A2(n5856), .ZN(n7415) );
  NAND2_X1 U7428 ( .A1(n5857), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7429 ( .A1(n5858), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7430 ( .A1(n5859), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7431 ( .A1(n5876), .A2(n5860), .ZN(n7448) );
  NAND2_X1 U7432 ( .A1(n6132), .A2(n7448), .ZN(n5862) );
  NAND2_X1 U7433 ( .A1(n6118), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5861) );
  NAND4_X2 U7434 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(n8386)
         );
  OR2_X1 U7435 ( .A1(n5866), .A2(n5865), .ZN(n5868) );
  XNOR2_X1 U7436 ( .A(n5868), .B(n5867), .ZN(n6659) );
  OR2_X1 U7437 ( .A1(n7984), .A2(n6661), .ZN(n5870) );
  INV_X1 U7438 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6660) );
  OR2_X1 U7439 ( .A1(n7983), .A2(n6660), .ZN(n5869) );
  OAI211_X1 U7440 ( .C1(n5821), .C2(n6659), .A(n5870), .B(n5869), .ZN(n7421)
         );
  NOR2_X1 U7441 ( .A1(n8386), .A2(n7421), .ZN(n5872) );
  INV_X1 U7442 ( .A(n5872), .ZN(n5871) );
  AND2_X1 U7443 ( .A1(n7415), .A2(n5871), .ZN(n5873) );
  NAND2_X1 U7444 ( .A1(n7412), .A2(n10032), .ZN(n7417) );
  AOI21_X2 U7445 ( .B1(n7416), .B2(n5873), .A(n4375), .ZN(n5875) );
  NAND2_X1 U7446 ( .A1(n8386), .A2(n7421), .ZN(n5874) );
  NAND2_X1 U7447 ( .A1(n7985), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7448 ( .A1(n7986), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U7449 ( .A1(n5876), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7450 ( .A1(n5888), .A2(n5877), .ZN(n7645) );
  NAND2_X1 U7451 ( .A1(n6132), .A2(n7645), .ZN(n5879) );
  NAND2_X1 U7452 ( .A1(n6118), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7453 ( .A1(n5882), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  MUX2_X1 U7454 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5883), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5884) );
  NAND2_X1 U7455 ( .A1(n5884), .A2(n4363), .ZN(n6664) );
  OR2_X1 U7456 ( .A1(n7984), .A2(n6665), .ZN(n5886) );
  OR2_X1 U7457 ( .A1(n7983), .A2(n6666), .ZN(n5885) );
  OAI211_X1 U7458 ( .C1(n5821), .C2(n6664), .A(n5886), .B(n5885), .ZN(n7635)
         );
  INV_X1 U7459 ( .A(n8385), .ZN(n7443) );
  NAND2_X1 U7460 ( .A1(n5888), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7461 ( .A1(n5890), .A2(n5889), .ZN(n10023) );
  NAND2_X1 U7462 ( .A1(n6132), .A2(n10023), .ZN(n5894) );
  NAND2_X1 U7463 ( .A1(n7986), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7464 ( .A1(n6118), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7465 ( .A1(n7985), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5891) );
  OR2_X1 U7466 ( .A1(n7984), .A2(n6668), .ZN(n5900) );
  OR2_X1 U7467 ( .A1(n7983), .A2(n6667), .ZN(n5899) );
  NAND2_X1 U7468 ( .A1(n4363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5895) );
  MUX2_X1 U7469 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5895), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5897) );
  NAND2_X1 U7470 ( .A1(n5897), .A2(n5896), .ZN(n7329) );
  OR2_X1 U7471 ( .A1(n5821), .A2(n7329), .ZN(n5898) );
  NAND2_X1 U7472 ( .A1(n8383), .A2(n10056), .ZN(n8079) );
  NAND2_X1 U7473 ( .A1(n8072), .A2(n8079), .ZN(n7613) );
  NAND2_X1 U7474 ( .A1(n7985), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7475 ( .A1(n7986), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7476 ( .A1(n5902), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7477 ( .A1(n5914), .A2(n5903), .ZN(n7770) );
  NAND2_X1 U7478 ( .A1(n6132), .A2(n7770), .ZN(n5905) );
  NAND2_X1 U7479 ( .A1(n6118), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5904) );
  OR2_X1 U7480 ( .A1(n5908), .A2(n5865), .ZN(n5910) );
  XNOR2_X1 U7481 ( .A(n5910), .B(n5909), .ZN(n7474) );
  INV_X1 U7482 ( .A(n7474), .ZN(n6538) );
  AOI22_X1 U7483 ( .A1(n6013), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6012), .B2(
        n6538), .ZN(n5912) );
  NAND2_X1 U7484 ( .A1(n6687), .A2(n7975), .ZN(n5911) );
  NAND2_X1 U7485 ( .A1(n8777), .A2(n10061), .ZN(n5913) );
  NAND2_X1 U7486 ( .A1(n7986), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7487 ( .A1(n7985), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7488 ( .A1(n5914), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7489 ( .A1(n5916), .A2(n5915), .ZN(n8781) );
  NAND2_X1 U7490 ( .A1(n6132), .A2(n8781), .ZN(n5918) );
  NAND2_X1 U7491 ( .A1(n6118), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7492 ( .A1(n6691), .A2(n7975), .ZN(n5924) );
  NAND2_X1 U7493 ( .A1(n5921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7494 ( .A(n5922), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6543) );
  AOI22_X1 U7495 ( .A1(n6013), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6012), .B2(
        n6543), .ZN(n5923) );
  NAND2_X1 U7496 ( .A1(n5924), .A2(n5923), .ZN(n8786) );
  NAND2_X1 U7497 ( .A1(n8762), .A2(n8786), .ZN(n5925) );
  NAND2_X1 U7498 ( .A1(n8769), .A2(n8779), .ZN(n8091) );
  NAND2_X1 U7499 ( .A1(n6796), .A2(n7975), .ZN(n5930) );
  OR2_X1 U7500 ( .A1(n5966), .A2(n5865), .ZN(n5927) );
  NAND2_X1 U7501 ( .A1(n5928), .A2(n5927), .ZN(n5940) );
  XNOR2_X1 U7502 ( .A(n5940), .B(n5965), .ZN(n6618) );
  AOI22_X1 U7503 ( .A1(n6013), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6012), .B2(
        n6618), .ZN(n5929) );
  NAND2_X1 U7504 ( .A1(n7985), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7505 ( .A1(n7986), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5937) );
  INV_X1 U7506 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7507 ( .A1(n5933), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7508 ( .A1(n5943), .A2(n5934), .ZN(n8738) );
  NAND2_X1 U7509 ( .A1(n6132), .A2(n8738), .ZN(n5936) );
  NAND2_X1 U7510 ( .A1(n6118), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5935) );
  NAND4_X1 U7511 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n8746)
         );
  NAND2_X1 U7512 ( .A1(n8841), .A2(n8746), .ZN(n8099) );
  NAND2_X1 U7513 ( .A1(n5939), .A2(n8099), .ZN(n8732) );
  NAND2_X1 U7514 ( .A1(n6861), .A2(n7975), .ZN(n5942) );
  OAI21_X1 U7515 ( .B1(n5940), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7516 ( .A(n5950), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6619) );
  AOI22_X1 U7517 ( .A1(n6013), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6012), .B2(
        n6619), .ZN(n5941) );
  NAND2_X1 U7518 ( .A1(n7985), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7519 ( .A1(n7986), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7520 ( .A1(n5943), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7521 ( .A1(n5957), .A2(n5944), .ZN(n8720) );
  NAND2_X1 U7522 ( .A1(n6132), .A2(n8720), .ZN(n5946) );
  NAND2_X1 U7523 ( .A1(n6118), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5945) );
  NOR2_X1 U7524 ( .A1(n8222), .A2(n8734), .ZN(n5949) );
  NAND2_X1 U7525 ( .A1(n6874), .A2(n7975), .ZN(n5954) );
  NAND2_X1 U7526 ( .A1(n5950), .A2(n5964), .ZN(n5951) );
  NAND2_X1 U7527 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7528 ( .A(n5952), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8426) );
  AOI22_X1 U7529 ( .A1(n6013), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6012), .B2(
        n8426), .ZN(n5953) );
  NAND2_X1 U7530 ( .A1(n5954), .A2(n5953), .ZN(n7901) );
  NAND2_X1 U7531 ( .A1(n7986), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7532 ( .A1(n7985), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5961) );
  INV_X1 U7533 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7534 ( .A1(n5957), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7535 ( .A1(n5972), .A2(n5958), .ZN(n8713) );
  NAND2_X1 U7536 ( .A1(n6132), .A2(n8713), .ZN(n5960) );
  NAND2_X1 U7537 ( .A1(n6118), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7538 ( .A1(n7901), .A2(n8699), .ZN(n8109) );
  NAND2_X1 U7539 ( .A1(n7901), .A2(n8699), .ZN(n8125) );
  NAND2_X1 U7540 ( .A1(n8109), .A2(n8125), .ZN(n8711) );
  AOI22_X1 U7541 ( .A1(n8708), .A2(n8711), .B1(n8699), .B2(n8932), .ZN(n8694)
         );
  NAND2_X1 U7542 ( .A1(n6967), .A2(n7975), .ZN(n5971) );
  NAND4_X1 U7543 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n5967)
         );
  OR2_X1 U7544 ( .A1(n5980), .A2(n5865), .ZN(n5969) );
  XNOR2_X1 U7545 ( .A(n5969), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8433) );
  AOI22_X1 U7546 ( .A1(n6013), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6012), .B2(
        n8433), .ZN(n5970) );
  NAND2_X1 U7547 ( .A1(n7985), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7548 ( .A1(n7986), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7549 ( .A1(n5972), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7550 ( .A1(n5985), .A2(n5973), .ZN(n8704) );
  NAND2_X1 U7551 ( .A1(n6132), .A2(n8704), .ZN(n5975) );
  NAND2_X1 U7552 ( .A1(n6118), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7553 ( .A1(n8925), .A2(n8710), .ZN(n8653) );
  NAND2_X1 U7554 ( .A1(n8654), .A2(n8653), .ZN(n8695) );
  NAND2_X1 U7555 ( .A1(n8694), .A2(n8695), .ZN(n8701) );
  INV_X1 U7556 ( .A(n8710), .ZN(n8687) );
  NAND2_X1 U7557 ( .A1(n8925), .A2(n8687), .ZN(n5978) );
  NAND2_X1 U7558 ( .A1(n8701), .A2(n5978), .ZN(n8685) );
  NAND2_X1 U7559 ( .A1(n7032), .A2(n7975), .ZN(n5983) );
  INV_X1 U7560 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7561 ( .A1(n5992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7562 ( .A(n5981), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8468) );
  AOI22_X1 U7563 ( .A1(n6013), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6012), .B2(
        n8468), .ZN(n5982) );
  NAND2_X1 U7564 ( .A1(n7985), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7565 ( .A1(n7986), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5989) );
  INV_X1 U7566 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7567 ( .A1(n5985), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7568 ( .A1(n5999), .A2(n5986), .ZN(n8690) );
  NAND2_X1 U7569 ( .A1(n6132), .A2(n8690), .ZN(n5988) );
  NAND2_X1 U7570 ( .A1(n6118), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7571 ( .A1(n8919), .A2(n8698), .ZN(n8669) );
  NAND2_X1 U7572 ( .A1(n8670), .A2(n8669), .ZN(n8684) );
  INV_X1 U7573 ( .A(n8698), .ZN(n8675) );
  NAND2_X1 U7574 ( .A1(n8919), .A2(n8675), .ZN(n5991) );
  NAND2_X1 U7575 ( .A1(n7104), .A2(n7975), .ZN(n5998) );
  INV_X1 U7576 ( .A(n5995), .ZN(n5993) );
  NAND2_X1 U7577 ( .A1(n5993), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7578 ( .A1(n5995), .A2(n5994), .ZN(n6009) );
  AND2_X1 U7579 ( .A1(n5996), .A2(n6009), .ZN(n8496) );
  AOI22_X1 U7580 ( .A1(n6013), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6012), .B2(
        n8496), .ZN(n5997) );
  NAND2_X1 U7581 ( .A1(n7986), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7582 ( .A1(n6118), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7583 ( .A1(n5999), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7584 ( .A1(n6018), .A2(n6000), .ZN(n8679) );
  NAND2_X1 U7585 ( .A1(n6132), .A2(n8679), .ZN(n6002) );
  NAND2_X1 U7586 ( .A1(n7985), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6001) );
  NAND4_X1 U7587 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n8686)
         );
  NAND2_X1 U7588 ( .A1(n8352), .A2(n6005), .ZN(n6006) );
  NAND2_X1 U7589 ( .A1(n8913), .A2(n8686), .ZN(n6007) );
  NAND2_X1 U7590 ( .A1(n6008), .A2(n6007), .ZN(n8662) );
  NAND2_X1 U7591 ( .A1(n7275), .A2(n7975), .ZN(n6015) );
  NAND2_X1 U7592 ( .A1(n6009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6011) );
  INV_X1 U7593 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7594 ( .A(n6011), .B(n6010), .ZN(n6174) );
  AOI22_X1 U7595 ( .A1(n6013), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8194), .B2(
        n6012), .ZN(n6014) );
  NAND2_X1 U7596 ( .A1(n7986), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7597 ( .A1(n6118), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6022) );
  INV_X1 U7598 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7599 ( .A1(n6018), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7600 ( .A1(n6027), .A2(n6019), .ZN(n8666) );
  NAND2_X1 U7601 ( .A1(n6132), .A2(n8666), .ZN(n6021) );
  NAND2_X1 U7602 ( .A1(n7985), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7603 ( .A1(n8907), .A2(n8645), .ZN(n8113) );
  NAND2_X1 U7604 ( .A1(n8130), .A2(n8113), .ZN(n8659) );
  NAND2_X1 U7605 ( .A1(n8907), .A2(n8676), .ZN(n6024) );
  NAND2_X1 U7606 ( .A1(n7352), .A2(n7975), .ZN(n6026) );
  OR2_X1 U7607 ( .A1(n7983), .A2(n7353), .ZN(n6025) );
  NAND2_X1 U7608 ( .A1(n7985), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7609 ( .A1(n7986), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7610 ( .A1(n6027), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7611 ( .A1(n6036), .A2(n6028), .ZN(n8649) );
  NAND2_X1 U7612 ( .A1(n6132), .A2(n8649), .ZN(n6030) );
  NAND2_X1 U7613 ( .A1(n6118), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7614 ( .A1(n8650), .A2(n8251), .ZN(n8133) );
  NAND2_X1 U7615 ( .A1(n7410), .A2(n7975), .ZN(n6034) );
  OR2_X1 U7616 ( .A1(n7983), .A2(n7411), .ZN(n6033) );
  NAND2_X1 U7617 ( .A1(n7985), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7618 ( .A1(n7986), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6040) );
  INV_X1 U7619 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7620 ( .A1(n6036), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7621 ( .A1(n6044), .A2(n6037), .ZN(n8637) );
  NAND2_X1 U7622 ( .A1(n6132), .A2(n8637), .ZN(n6039) );
  NAND2_X1 U7623 ( .A1(n6118), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7624 ( .A1(n8896), .A2(n8646), .ZN(n8137) );
  NAND2_X1 U7625 ( .A1(n8138), .A2(n8137), .ZN(n8628) );
  NAND2_X1 U7626 ( .A1(n7599), .A2(n7975), .ZN(n6043) );
  OR2_X1 U7627 ( .A1(n7983), .A2(n7603), .ZN(n6042) );
  NAND2_X1 U7628 ( .A1(n6044), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7629 ( .A1(n6050), .A2(n6045), .ZN(n8625) );
  AOI22_X1 U7630 ( .A1(n8625), .A2(n6132), .B1(n6118), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6047) );
  AOI22_X1 U7631 ( .A1(n7985), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n7986), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7632 ( .A1(n8890), .A2(n7927), .ZN(n8141) );
  NAND2_X1 U7633 ( .A1(n8143), .A2(n8141), .ZN(n8136) );
  INV_X1 U7634 ( .A(n8136), .ZN(n6077) );
  NAND2_X1 U7635 ( .A1(n7608), .A2(n7975), .ZN(n6049) );
  OR2_X1 U7636 ( .A1(n7983), .A2(n7610), .ZN(n6048) );
  INV_X1 U7637 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U7638 ( .A1(n6050), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7639 ( .A1(n6057), .A2(n6051), .ZN(n8609) );
  NAND2_X1 U7640 ( .A1(n8609), .A2(n6132), .ZN(n6053) );
  AOI22_X1 U7641 ( .A1(n6118), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n7986), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7642 ( .A1(n8884), .A2(n8622), .ZN(n8590) );
  INV_X1 U7643 ( .A(n8590), .ZN(n6079) );
  OR2_X1 U7644 ( .A1(n8588), .A2(n6079), .ZN(n8567) );
  NAND2_X1 U7645 ( .A1(n7751), .A2(n7975), .ZN(n6056) );
  OR2_X1 U7646 ( .A1(n7983), .A2(n7839), .ZN(n6055) );
  INV_X1 U7647 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6061) );
  INV_X1 U7648 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U7649 ( .A1(n6057), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7650 ( .A1(n6066), .A2(n6058), .ZN(n8599) );
  NAND2_X1 U7651 ( .A1(n8599), .A2(n6132), .ZN(n6060) );
  AOI22_X1 U7652 ( .A1(n7985), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n7986), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7653 ( .A1(n8878), .A2(n8606), .ZN(n8570) );
  NAND2_X1 U7654 ( .A1(n7796), .A2(n7975), .ZN(n6063) );
  OR2_X1 U7655 ( .A1(n7983), .A2(n7797), .ZN(n6062) );
  INV_X1 U7656 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7657 ( .A1(n6066), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7658 ( .A1(n6088), .A2(n6067), .ZN(n8579) );
  NAND2_X1 U7659 ( .A1(n8579), .A2(n6132), .ZN(n6073) );
  INV_X1 U7660 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7661 ( .A1(n7985), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7662 ( .A1(n7986), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6068) );
  OAI211_X1 U7663 ( .C1(n6070), .C2(n6181), .A(n6069), .B(n6068), .ZN(n6071)
         );
  INV_X1 U7664 ( .A(n6071), .ZN(n6072) );
  NAND2_X1 U7665 ( .A1(n8268), .A2(n8358), .ZN(n8154) );
  INV_X1 U7666 ( .A(n8580), .ZN(n6074) );
  NAND2_X1 U7667 ( .A1(n8570), .A2(n6074), .ZN(n6083) );
  NAND2_X1 U7668 ( .A1(n8872), .A2(n8358), .ZN(n6084) );
  INV_X1 U7669 ( .A(n8890), .ZN(n8331) );
  NAND2_X1 U7670 ( .A1(n8331), .A2(n7927), .ZN(n6078) );
  NAND2_X1 U7671 ( .A1(n7919), .A2(n8646), .ZN(n8618) );
  INV_X1 U7672 ( .A(n8650), .ZN(n8901) );
  NAND2_X1 U7673 ( .A1(n8901), .A2(n8251), .ZN(n8630) );
  OR2_X1 U7674 ( .A1(n6079), .A2(n8589), .ZN(n6082) );
  OR2_X1 U7675 ( .A1(n8878), .A2(n8606), .ZN(n6080) );
  INV_X1 U7676 ( .A(n8884), .ZN(n6170) );
  NAND2_X1 U7677 ( .A1(n6170), .A2(n8327), .ZN(n8591) );
  AND2_X1 U7678 ( .A1(n6080), .A2(n8591), .ZN(n6081) );
  NAND2_X1 U7679 ( .A1(n7802), .A2(n7975), .ZN(n6087) );
  OR2_X1 U7680 ( .A1(n7983), .A2(n7803), .ZN(n6086) );
  NAND2_X1 U7681 ( .A1(n6088), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7682 ( .A1(n6104), .A2(n6089), .ZN(n8563) );
  NAND2_X1 U7683 ( .A1(n8563), .A2(n6132), .ZN(n6094) );
  INV_X1 U7684 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U7685 ( .A1(n7985), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7686 ( .A1(n7986), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6090) );
  OAI211_X1 U7687 ( .C1(n8562), .C2(n6181), .A(n6091), .B(n6090), .ZN(n6092)
         );
  INV_X1 U7688 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7689 ( .A1(n8867), .A2(n8550), .ZN(n6095) );
  NAND2_X1 U7690 ( .A1(n8559), .A2(n6095), .ZN(n6098) );
  INV_X1 U7691 ( .A(n8867), .ZN(n6096) );
  NAND2_X1 U7692 ( .A1(n6096), .A2(n8576), .ZN(n6097) );
  NAND2_X1 U7693 ( .A1(n7820), .A2(n7975), .ZN(n6101) );
  OR2_X1 U7694 ( .A1(n7983), .A2(n6099), .ZN(n6100) );
  INV_X1 U7695 ( .A(n6104), .ZN(n6103) );
  INV_X1 U7696 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7697 ( .A1(n6103), .A2(n6102), .ZN(n6116) );
  NAND2_X1 U7698 ( .A1(n6104), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7699 ( .A1(n6116), .A2(n6105), .ZN(n8554) );
  NAND2_X1 U7700 ( .A1(n8554), .A2(n6132), .ZN(n6110) );
  INV_X1 U7701 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U7702 ( .A1(n7986), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7703 ( .A1(n7985), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U7704 ( .C1(n8553), .C2(n6181), .A(n6107), .B(n6106), .ZN(n6108)
         );
  INV_X1 U7705 ( .A(n6108), .ZN(n6109) );
  INV_X1 U7706 ( .A(n8537), .ZN(n8560) );
  INV_X1 U7707 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6415) );
  INV_X1 U7708 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n6113) );
  MUX2_X1 U7709 ( .A(n6415), .B(n6113), .S(n7969), .Z(n6127) );
  XNOR2_X1 U7710 ( .A(n6127), .B(SI_28_), .ZN(n6124) );
  NAND2_X1 U7711 ( .A1(n7827), .A2(n7975), .ZN(n6115) );
  OR2_X1 U7712 ( .A1(n7983), .A2(n6415), .ZN(n6114) );
  NAND2_X1 U7713 ( .A1(n6116), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7714 ( .A1(n8521), .A2(n6117), .ZN(n8542) );
  NAND2_X1 U7715 ( .A1(n8542), .A2(n6132), .ZN(n6123) );
  INV_X1 U7716 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U7717 ( .A1(n7985), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7718 ( .A1(n6118), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6119) );
  OAI211_X1 U7719 ( .C1(n5790), .C2(n6457), .A(n6120), .B(n6119), .ZN(n6121)
         );
  INV_X1 U7720 ( .A(n6121), .ZN(n6122) );
  INV_X1 U7721 ( .A(SI_28_), .ZN(n6126) );
  NAND2_X1 U7722 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  INV_X1 U7723 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8954) );
  INV_X1 U7724 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6129) );
  MUX2_X1 U7725 ( .A(n8954), .B(n6129), .S(n7969), .Z(n7965) );
  NAND2_X1 U7726 ( .A1(n7844), .A2(n7975), .ZN(n6131) );
  OR2_X1 U7727 ( .A1(n7983), .A2(n8954), .ZN(n6130) );
  INV_X1 U7728 ( .A(n8521), .ZN(n6133) );
  NAND2_X1 U7729 ( .A1(n6133), .A2(n6132), .ZN(n7991) );
  INV_X1 U7730 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U7731 ( .A1(n7986), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7732 ( .A1(n7985), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6134) );
  OAI211_X1 U7733 ( .C1(n6181), .C2(n8527), .A(n6135), .B(n6134), .ZN(n6136)
         );
  INV_X1 U7734 ( .A(n6136), .ZN(n6137) );
  NAND2_X1 U7735 ( .A1(n8530), .A2(n8538), .ZN(n7994) );
  INV_X1 U7736 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7737 ( .A1(n6139), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6140) );
  XNOR2_X1 U7738 ( .A(n6140), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U7739 ( .A1(n8194), .A2(n8197), .ZN(n6234) );
  NAND2_X1 U7740 ( .A1(n6141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6142) );
  XNOR2_X1 U7741 ( .A(n6142), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U7742 ( .A1(n4376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6143) );
  MUX2_X1 U7743 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6143), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6144) );
  NAND2_X1 U7744 ( .A1(n6144), .A2(n6141), .ZN(n8190) );
  INV_X1 U7745 ( .A(n8190), .ZN(n6209) );
  NAND2_X1 U7746 ( .A1(n8033), .A2(n6209), .ZN(n6145) );
  NAND2_X1 U7747 ( .A1(n6234), .A2(n6145), .ZN(n8755) );
  NAND2_X1 U7748 ( .A1(n6146), .A2(n8755), .ZN(n6187) );
  INV_X1 U7749 ( .A(n7029), .ZN(n7054) );
  NAND2_X1 U7750 ( .A1(n8006), .A2(n8037), .ZN(n7095) );
  NAND2_X1 U7751 ( .A1(n7095), .A2(n8039), .ZN(n7378) );
  AND2_X1 U7752 ( .A1(n6148), .A2(n6147), .ZN(n8046) );
  NAND2_X1 U7753 ( .A1(n7378), .A2(n8046), .ZN(n6151) );
  INV_X1 U7754 ( .A(n6148), .ZN(n8060) );
  OAI21_X1 U7755 ( .B1(n8060), .B2(n8045), .A(n8052), .ZN(n6149) );
  INV_X1 U7756 ( .A(n6149), .ZN(n6150) );
  NAND2_X1 U7757 ( .A1(n6151), .A2(n6150), .ZN(n7336) );
  NAND2_X1 U7758 ( .A1(n8387), .A2(n7875), .ZN(n8053) );
  NAND2_X1 U7759 ( .A1(n7412), .A2(n8053), .ZN(n7334) );
  INV_X1 U7760 ( .A(n7421), .ZN(n10046) );
  NAND2_X1 U7761 ( .A1(n8386), .A2(n10046), .ZN(n8062) );
  INV_X1 U7762 ( .A(n8062), .ZN(n6152) );
  OR2_X1 U7763 ( .A1(n8386), .A2(n10046), .ZN(n8055) );
  OR2_X1 U7764 ( .A1(n8385), .A2(n10051), .ZN(n8063) );
  NAND2_X1 U7765 ( .A1(n8385), .A2(n10051), .ZN(n8064) );
  NAND2_X1 U7766 ( .A1(n8063), .A2(n8064), .ZN(n7480) );
  NAND2_X1 U7767 ( .A1(n8384), .A2(n8073), .ZN(n8078) );
  INV_X1 U7768 ( .A(n8079), .ZN(n6153) );
  OR2_X1 U7769 ( .A1(n8382), .A2(n10061), .ZN(n8075) );
  NAND2_X1 U7770 ( .A1(n8382), .A2(n10061), .ZN(n8080) );
  NAND2_X1 U7771 ( .A1(n8075), .A2(n8080), .ZN(n8013) );
  INV_X1 U7772 ( .A(n8013), .ZN(n6154) );
  NAND2_X1 U7773 ( .A1(n10067), .A2(n8762), .ZN(n8089) );
  OR2_X1 U7774 ( .A1(n8762), .A2(n10067), .ZN(n8752) );
  AND2_X1 U7775 ( .A1(n8091), .A2(n8752), .ZN(n8088) );
  NAND2_X1 U7776 ( .A1(n8753), .A2(n8088), .ZN(n6155) );
  NAND2_X1 U7777 ( .A1(n6155), .A2(n8093), .ZN(n8742) );
  OR2_X1 U7778 ( .A1(n8941), .A2(n8735), .ZN(n8095) );
  NAND2_X1 U7779 ( .A1(n8941), .A2(n8735), .ZN(n8096) );
  NAND2_X1 U7780 ( .A1(n8742), .A2(n8743), .ZN(n6156) );
  INV_X1 U7781 ( .A(n8746), .ZN(n8218) );
  NAND2_X1 U7782 ( .A1(n8841), .A2(n8218), .ZN(n6157) );
  OR2_X1 U7783 ( .A1(n8722), .A2(n8734), .ZN(n7876) );
  AND2_X1 U7784 ( .A1(n8722), .A2(n8734), .ZN(n8106) );
  NAND2_X1 U7785 ( .A1(n6158), .A2(n8109), .ZN(n8693) );
  INV_X1 U7786 ( .A(n8130), .ZN(n6161) );
  NAND2_X1 U7787 ( .A1(n8913), .A2(n6005), .ZN(n8122) );
  INV_X1 U7788 ( .A(n8122), .ZN(n8003) );
  AND2_X1 U7789 ( .A1(n8120), .A2(n8670), .ZN(n6159) );
  AND2_X1 U7790 ( .A1(n8669), .A2(n8122), .ZN(n8656) );
  AND2_X1 U7791 ( .A1(n8656), .A2(n8113), .ZN(n6160) );
  AND2_X1 U7792 ( .A1(n8653), .A2(n6165), .ZN(n6162) );
  NAND2_X1 U7793 ( .A1(n8693), .A2(n6162), .ZN(n6167) );
  AND2_X1 U7794 ( .A1(n8654), .A2(n6163), .ZN(n6164) );
  NAND2_X1 U7795 ( .A1(n6167), .A2(n6166), .ZN(n8640) );
  INV_X1 U7796 ( .A(n8132), .ZN(n6168) );
  INV_X1 U7797 ( .A(n8137), .ZN(n6169) );
  NAND2_X1 U7798 ( .A1(n8878), .A2(n8577), .ZN(n8001) );
  NAND2_X1 U7799 ( .A1(n8884), .A2(n8327), .ZN(n8585) );
  AND2_X1 U7800 ( .A1(n8001), .A2(n8585), .ZN(n8149) );
  INV_X1 U7801 ( .A(n8878), .ZN(n8597) );
  NAND2_X1 U7802 ( .A1(n6174), .A2(n8190), .ZN(n6974) );
  OR2_X1 U7803 ( .A1(n6974), .A2(n8171), .ZN(n6979) );
  INV_X1 U7804 ( .A(n8197), .ZN(n7601) );
  INV_X1 U7805 ( .A(n8033), .ZN(n8036) );
  INV_X1 U7806 ( .A(n7382), .ZN(n10072) );
  OAI21_X1 U7807 ( .B1(n8197), .B2(n8190), .A(n10072), .ZN(n6175) );
  NOR2_X1 U7808 ( .A1(n8194), .A2(n6175), .ZN(n6176) );
  AND2_X1 U7809 ( .A1(n6979), .A2(n6176), .ZN(n7757) );
  INV_X1 U7810 ( .A(n6177), .ZN(n6567) );
  NAND2_X1 U7811 ( .A1(n6567), .A2(n8493), .ZN(n6178) );
  NAND2_X1 U7812 ( .A1(n5821), .A2(n6178), .ZN(n6978) );
  INV_X1 U7813 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U7814 ( .A1(n7985), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7815 ( .A1(n7986), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6179) );
  OAI211_X1 U7816 ( .C1(n8525), .C2(n6181), .A(n6180), .B(n6179), .ZN(n6182)
         );
  INV_X1 U7817 ( .A(n6182), .ZN(n6183) );
  AND2_X1 U7818 ( .A1(n7991), .A2(n6183), .ZN(n7993) );
  NAND2_X1 U7819 ( .A1(n6978), .A2(n8185), .ZN(n8780) );
  AND2_X1 U7820 ( .A1(n5821), .A2(P2_B_REG_SCAN_IN), .ZN(n6184) );
  OR2_X1 U7821 ( .A1(n8780), .A2(n6184), .ZN(n8519) );
  OAI22_X1 U7822 ( .A1(n8208), .A2(n8778), .B1(n7993), .B2(n8519), .ZN(n6185)
         );
  INV_X1 U7823 ( .A(n7384), .ZN(n6189) );
  OR2_X1 U7824 ( .A1(n6189), .A2(n8197), .ZN(n10062) );
  NAND2_X1 U7825 ( .A1(n6190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7826 ( .A1(n6226), .A2(n5760), .ZN(n6191) );
  NAND2_X1 U7827 ( .A1(n6191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7828 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  NAND2_X1 U7829 ( .A1(n6197), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7830 ( .A(n6193), .B(n6192), .ZN(n7798) );
  OR2_X1 U7831 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  NAND2_X1 U7832 ( .A1(n6197), .A2(n6196), .ZN(n7840) );
  XNOR2_X1 U7833 ( .A(n7840), .B(P2_B_REG_SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7834 ( .A1(n7798), .A2(n6198), .ZN(n6202) );
  AND2_X1 U7835 ( .A1(n4393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7836 ( .A1(n6202), .A2(n6203), .ZN(n6703) );
  OR2_X1 U7837 ( .A1(n6703), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6205) );
  INV_X1 U7838 ( .A(n6203), .ZN(n7804) );
  NAND2_X1 U7839 ( .A1(n7798), .A2(n7804), .ZN(n6204) );
  NAND2_X1 U7840 ( .A1(n6205), .A2(n6204), .ZN(n7019) );
  INV_X1 U7841 ( .A(n7019), .ZN(n8948) );
  INV_X1 U7842 ( .A(n6703), .ZN(n6207) );
  INV_X1 U7843 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7844 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  NAND2_X1 U7845 ( .A1(n7804), .A2(n7840), .ZN(n6836) );
  AND2_X2 U7846 ( .A1(n6208), .A2(n6836), .ZN(n7017) );
  NAND2_X1 U7847 ( .A1(n8948), .A2(n7017), .ZN(n6237) );
  INV_X1 U7848 ( .A(n7017), .ZN(n7015) );
  AND2_X1 U7849 ( .A1(n7384), .A2(n7382), .ZN(n6887) );
  NAND3_X1 U7850 ( .A1(n6174), .A2(n8197), .A3(n6209), .ZN(n6210) );
  NAND2_X1 U7851 ( .A1(n6210), .A2(n8171), .ZN(n6227) );
  INV_X1 U7852 ( .A(n6227), .ZN(n7018) );
  OAI21_X1 U7853 ( .B1(n7015), .B2(n6887), .A(n7018), .ZN(n6211) );
  AND2_X1 U7854 ( .A1(n6237), .A2(n6211), .ZN(n6230) );
  NAND2_X1 U7855 ( .A1(n6974), .A2(n8185), .ZN(n6214) );
  INV_X1 U7856 ( .A(n7798), .ZN(n6213) );
  NOR2_X1 U7857 ( .A1(n7840), .A2(n7804), .ZN(n6212) );
  NAND2_X1 U7858 ( .A1(n6213), .A2(n6212), .ZN(n6570) );
  NAND2_X1 U7859 ( .A1(n6214), .A2(n6570), .ZN(n6889) );
  NOR2_X1 U7860 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n6218) );
  NOR4_X1 U7861 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6217) );
  NOR4_X1 U7862 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6216) );
  NOR4_X1 U7863 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6215) );
  NAND4_X1 U7864 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n6224)
         );
  NOR4_X1 U7865 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6222) );
  NOR4_X1 U7866 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6221) );
  NOR4_X1 U7867 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6220) );
  NOR4_X1 U7868 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6219) );
  NAND4_X1 U7869 ( .A1(n6222), .A2(n6221), .A3(n6220), .A4(n6219), .ZN(n6223)
         );
  NOR2_X1 U7870 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NOR2_X1 U7871 ( .A1(n6703), .A2(n6225), .ZN(n6236) );
  XNOR2_X1 U7872 ( .A(n6226), .B(n5760), .ZN(n7112) );
  NAND2_X1 U7873 ( .A1(n7112), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6512) );
  OR3_X1 U7874 ( .A1(n6889), .A2(n6236), .A3(n6512), .ZN(n7016) );
  AND2_X1 U7875 ( .A1(n7019), .A2(n6227), .ZN(n6228) );
  NOR2_X1 U7876 ( .A1(n7016), .A2(n6228), .ZN(n6229) );
  AND2_X2 U7877 ( .A1(n6230), .A2(n6229), .ZN(n10092) );
  INV_X1 U7878 ( .A(n6231), .ZN(n6232) );
  NAND2_X1 U7879 ( .A1(n10092), .A2(n7382), .ZN(n8838) );
  NAND2_X1 U7880 ( .A1(n6232), .A2(n4901), .ZN(P2_U3488) );
  NOR2_X1 U7881 ( .A1(n7017), .A2(n6236), .ZN(n6233) );
  AND2_X1 U7882 ( .A1(n6233), .A2(n7019), .ZN(n6896) );
  INV_X1 U7883 ( .A(n6512), .ZN(n6899) );
  OR2_X1 U7884 ( .A1(n8033), .A2(n8190), .ZN(n6971) );
  OR2_X1 U7885 ( .A1(n6234), .A2(n6971), .ZN(n6894) );
  NOR2_X1 U7886 ( .A1(n8185), .A2(n7382), .ZN(n6235) );
  NAND2_X1 U7887 ( .A1(n6894), .A2(n6235), .ZN(n6880) );
  OR2_X1 U7888 ( .A1(n7384), .A2(n10072), .ZN(n8736) );
  NAND2_X1 U7889 ( .A1(n6880), .A2(n8736), .ZN(n6890) );
  NAND2_X1 U7890 ( .A1(n6981), .A2(n6890), .ZN(n6241) );
  OR2_X1 U7891 ( .A1(n6237), .A2(n6236), .ZN(n6891) );
  INV_X1 U7892 ( .A(n8947), .ZN(n6238) );
  NOR2_X1 U7893 ( .A1(n6891), .A2(n6238), .ZN(n6886) );
  NAND2_X1 U7894 ( .A1(n6979), .A2(n6894), .ZN(n6239) );
  NAND2_X1 U7895 ( .A1(n6886), .A2(n6239), .ZN(n6240) );
  INV_X2 U7896 ( .A(n10080), .ZN(n10078) );
  NAND2_X1 U7897 ( .A1(n4340), .A2(n4905), .ZN(P2_U3456) );
  INV_X1 U7898 ( .A(n9400), .ZN(n9626) );
  XNOR2_X2 U7899 ( .A(n9413), .B(n9205), .ZN(n6941) );
  NAND2_X1 U7900 ( .A1(n6272), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U7901 ( .A1(n6941), .A2(n6942), .ZN(n6244) );
  OR2_X1 U7902 ( .A1(n9413), .A2(n9900), .ZN(n6243) );
  NAND2_X1 U7903 ( .A1(n6244), .A2(n6243), .ZN(n7215) );
  NAND2_X1 U7904 ( .A1(n7215), .A2(n9147), .ZN(n6246) );
  OR2_X1 U7905 ( .A1(n9411), .A2(n9201), .ZN(n6245) );
  NAND2_X1 U7906 ( .A1(n6246), .A2(n6245), .ZN(n7236) );
  NAND2_X1 U7907 ( .A1(n9878), .A2(n9921), .ZN(n9207) );
  NAND2_X1 U7908 ( .A1(n6278), .A2(n9207), .ZN(n7235) );
  NAND2_X1 U7909 ( .A1(n7236), .A2(n7235), .ZN(n6248) );
  OR2_X1 U7910 ( .A1(n9878), .A2(n7240), .ZN(n6247) );
  NAND2_X1 U7911 ( .A1(n6248), .A2(n6247), .ZN(n9886) );
  INV_X1 U7912 ( .A(n7079), .ZN(n9927) );
  XNOR2_X1 U7913 ( .A(n9410), .B(n9927), .ZN(n9887) );
  OR2_X1 U7914 ( .A1(n9410), .A2(n7079), .ZN(n6249) );
  NAND2_X1 U7915 ( .A1(n9880), .A2(n9933), .ZN(n9251) );
  NAND2_X1 U7916 ( .A1(n9253), .A2(n9251), .ZN(n9151) );
  INV_X1 U7917 ( .A(n9409), .ZN(n7254) );
  NAND2_X1 U7918 ( .A1(n7254), .A2(n6270), .ZN(n9254) );
  INV_X1 U7919 ( .A(n6270), .ZN(n9939) );
  NAND2_X1 U7920 ( .A1(n9939), .A2(n9409), .ZN(n9257) );
  NAND2_X1 U7921 ( .A1(n9254), .A2(n9257), .ZN(n9867) );
  NAND2_X1 U7922 ( .A1(n9866), .A2(n9867), .ZN(n6251) );
  NAND2_X1 U7923 ( .A1(n7254), .A2(n9939), .ZN(n6250) );
  INV_X1 U7924 ( .A(n9861), .ZN(n9834) );
  OR2_X1 U7925 ( .A1(n9945), .A2(n9834), .ZN(n9260) );
  NAND2_X1 U7926 ( .A1(n9834), .A2(n9945), .ZN(n9839) );
  NAND2_X1 U7927 ( .A1(n9260), .A2(n9839), .ZN(n7303) );
  OR2_X1 U7928 ( .A1(n9945), .A2(n9861), .ZN(n6252) );
  INV_X1 U7929 ( .A(n9408), .ZN(n7295) );
  NAND2_X1 U7930 ( .A1(n7590), .A2(n7295), .ZN(n9264) );
  NAND2_X1 U7931 ( .A1(n9843), .A2(n9264), .ZN(n9838) );
  INV_X1 U7932 ( .A(n9407), .ZN(n9836) );
  OR2_X1 U7933 ( .A1(n9960), .A2(n9836), .ZN(n9274) );
  NAND2_X1 U7934 ( .A1(n9960), .A2(n9836), .ZN(n9270) );
  OR2_X1 U7935 ( .A1(n7459), .A2(n7701), .ZN(n9279) );
  NAND2_X1 U7936 ( .A1(n7459), .A2(n7701), .ZN(n9276) );
  NAND2_X1 U7937 ( .A1(n9279), .A2(n9276), .ZN(n9145) );
  INV_X1 U7938 ( .A(n7459), .ZN(n9970) );
  INV_X1 U7939 ( .A(n9405), .ZN(n8989) );
  NAND2_X1 U7940 ( .A1(n7586), .A2(n8989), .ZN(n9281) );
  NAND2_X1 U7941 ( .A1(n7631), .A2(n9091), .ZN(n9282) );
  NAND2_X1 U7942 ( .A1(n9283), .A2(n9282), .ZN(n7624) );
  INV_X1 U7943 ( .A(n9403), .ZN(n9018) );
  OR2_X1 U7944 ( .A1(n7694), .A2(n9018), .ZN(n9289) );
  NAND2_X1 U7945 ( .A1(n7694), .A2(n9018), .ZN(n9288) );
  INV_X1 U7946 ( .A(n9402), .ZN(n9127) );
  NAND2_X1 U7947 ( .A1(n8968), .A2(n9127), .ZN(n9223) );
  INV_X1 U7948 ( .A(n8968), .ZN(n9997) );
  INV_X1 U7949 ( .A(n9702), .ZN(n9037) );
  NAND2_X1 U7950 ( .A1(n7817), .A2(n9037), .ZN(n9301) );
  INV_X1 U7951 ( .A(n9690), .ZN(n9046) );
  NAND2_X1 U7952 ( .A1(n9719), .A2(n9046), .ZN(n9306) );
  NAND2_X1 U7953 ( .A1(n9719), .A2(n9690), .ZN(n6255) );
  INV_X1 U7954 ( .A(n9703), .ZN(n6256) );
  NAND2_X1 U7955 ( .A1(n6271), .A2(n6256), .ZN(n9308) );
  OR2_X1 U7956 ( .A1(n9781), .A2(n9664), .ZN(n9229) );
  NAND2_X1 U7957 ( .A1(n9781), .A2(n9664), .ZN(n9312) );
  NAND2_X1 U7958 ( .A1(n9229), .A2(n9312), .ZN(n9165) );
  INV_X1 U7959 ( .A(n9777), .ZN(n9655) );
  INV_X1 U7960 ( .A(n9678), .ZN(n9643) );
  NAND2_X1 U7961 ( .A1(n9655), .A2(n9643), .ZN(n6257) );
  INV_X1 U7962 ( .A(n9401), .ZN(n9663) );
  NAND2_X1 U7963 ( .A1(n9767), .A2(n9614), .ZN(n6259) );
  NAND2_X1 U7964 ( .A1(n9633), .A2(n6260), .ZN(n6261) );
  NAND2_X1 U7965 ( .A1(n9752), .A2(n9592), .ZN(n9341) );
  NAND2_X1 U7966 ( .A1(n9746), .A2(n9544), .ZN(n9347) );
  XOR2_X1 U7967 ( .A(n9356), .B(n7842), .Z(n7962) );
  INV_X1 U7968 ( .A(n6265), .ZN(n6268) );
  OAI21_X1 U7969 ( .B1(n6268), .B2(n6267), .A(n6266), .ZN(n6269) );
  OR2_X1 U7970 ( .A1(n9381), .A2(n6269), .ZN(n7579) );
  OR2_X1 U7971 ( .A1(n9384), .A2(n9388), .ZN(n9383) );
  NAND2_X1 U7972 ( .A1(n9369), .A2(n9197), .ZN(n6940) );
  INV_X1 U7973 ( .A(n9996), .ZN(n9959) );
  NOR2_X1 U7974 ( .A1(n6943), .A2(n9900), .ZN(n7227) );
  INV_X1 U7975 ( .A(n9960), .ZN(n7707) );
  NAND2_X1 U7976 ( .A1(n9853), .A2(n7707), .ZN(n7455) );
  INV_X1 U7977 ( .A(n7694), .ZN(n9991) );
  INV_X1 U7978 ( .A(n9719), .ZN(n9819) );
  INV_X1 U7979 ( .A(n6271), .ZN(n9812) );
  AOI211_X1 U7980 ( .C1(n6298), .C2(n9545), .A(n9670), .B(n9519), .ZN(n7953)
         );
  INV_X1 U7981 ( .A(n6941), .ZN(n6273) );
  NAND2_X1 U7982 ( .A1(n6273), .A2(n6946), .ZN(n6275) );
  INV_X1 U7983 ( .A(n9413), .ZN(n6902) );
  NAND2_X1 U7984 ( .A1(n6902), .A2(n9900), .ZN(n6274) );
  NAND2_X1 U7985 ( .A1(n6275), .A2(n6274), .ZN(n7216) );
  INV_X1 U7986 ( .A(n9147), .ZN(n7217) );
  INV_X1 U7987 ( .A(n9411), .ZN(n9202) );
  NAND2_X1 U7988 ( .A1(n9202), .A2(n9201), .ZN(n6276) );
  AND2_X1 U7989 ( .A1(n9410), .A2(n9927), .ZN(n9206) );
  INV_X1 U7990 ( .A(n9151), .ZN(n6279) );
  NAND2_X1 U7991 ( .A1(n6280), .A2(n9253), .ZN(n9859) );
  NAND2_X1 U7992 ( .A1(n9274), .A2(n9843), .ZN(n9265) );
  AND2_X1 U7993 ( .A1(n9264), .A2(n9839), .ZN(n9262) );
  AND2_X1 U7994 ( .A1(n6281), .A2(n9270), .ZN(n6283) );
  NAND2_X1 U7995 ( .A1(n6283), .A2(n9254), .ZN(n9214) );
  NAND2_X1 U7996 ( .A1(n9260), .A2(n9257), .ZN(n6282) );
  OR2_X1 U7997 ( .A1(n9265), .A2(n6282), .ZN(n9146) );
  NAND2_X1 U7998 ( .A1(n6283), .A2(n9146), .ZN(n9213) );
  INV_X1 U7999 ( .A(n9158), .ZN(n7572) );
  INV_X1 U8000 ( .A(n9276), .ZN(n7573) );
  NAND2_X1 U8001 ( .A1(n7575), .A2(n9278), .ZN(n7622) );
  INV_X1 U8002 ( .A(n7624), .ZN(n9159) );
  INV_X1 U8003 ( .A(n9160), .ZN(n9291) );
  INV_X1 U8004 ( .A(n6286), .ZN(n7809) );
  NAND2_X1 U8005 ( .A1(n7808), .A2(n9301), .ZN(n9700) );
  INV_X1 U8006 ( .A(n9306), .ZN(n9228) );
  INV_X1 U8007 ( .A(n9684), .ZN(n9687) );
  INV_X1 U8008 ( .A(n9165), .ZN(n9676) );
  XNOR2_X1 U8009 ( .A(n9777), .B(n9678), .ZN(n9144) );
  AND2_X1 U8010 ( .A1(n9777), .A2(n9643), .ZN(n9311) );
  NOR2_X1 U8011 ( .A1(n9767), .A2(n6260), .ZN(n6288) );
  INV_X1 U8012 ( .A(n9321), .ZN(n6287) );
  NAND2_X1 U8013 ( .A1(n9767), .A2(n6260), .ZN(n9329) );
  NAND2_X1 U8014 ( .A1(n9329), .A2(n9621), .ZN(n6289) );
  INV_X1 U8015 ( .A(n6288), .ZN(n9319) );
  OR2_X1 U8016 ( .A1(n9762), .A2(n9626), .ZN(n9142) );
  NAND2_X1 U8017 ( .A1(n9762), .A2(n9626), .ZN(n9143) );
  INV_X1 U8018 ( .A(n9586), .ZN(n9590) );
  INV_X1 U8019 ( .A(n9335), .ZN(n9572) );
  INV_X1 U8020 ( .A(n9340), .ZN(n6290) );
  INV_X1 U8021 ( .A(n9541), .ZN(n6291) );
  INV_X1 U8022 ( .A(n9180), .ZN(n9350) );
  XNOR2_X1 U8023 ( .A(n7853), .B(n9356), .ZN(n6294) );
  OR2_X1 U8024 ( .A1(n9384), .A2(n9376), .ZN(n6293) );
  NAND2_X1 U8025 ( .A1(n6293), .A2(n9386), .ZN(n9876) );
  INV_X1 U8026 ( .A(n9876), .ZN(n9842) );
  NAND2_X1 U8027 ( .A1(n6294), .A2(n9876), .ZN(n6297) );
  NAND2_X1 U8028 ( .A1(n6679), .A2(n9194), .ZN(n9835) );
  NAND2_X1 U8029 ( .A1(n7828), .A2(n9194), .ZN(n9833) );
  INV_X1 U8030 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U8031 ( .A1(n6297), .A2(n6296), .ZN(n7960) );
  OAI21_X1 U8032 ( .B1(n7962), .B2(n9963), .A(n6299), .ZN(n9739) );
  NAND2_X1 U8033 ( .A1(n6300), .A2(n9380), .ZN(n6790) );
  INV_X1 U8034 ( .A(n6301), .ZN(n6302) );
  NOR2_X1 U8035 ( .A1(n7220), .A2(n6904), .ZN(n6304) );
  NOR2_X1 U8036 ( .A1(n6303), .A2(n7221), .ZN(n6905) );
  AND2_X2 U8037 ( .A1(n6304), .A2(n6905), .ZN(n10004) );
  INV_X1 U8038 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8816) );
  AOI22_X1 U8039 ( .A1(n8816), .A2(keyinput124), .B1(n7803), .B2(keyinput115), 
        .ZN(n6307) );
  OAI221_X1 U8040 ( .B1(n8816), .B2(keyinput124), .C1(n7803), .C2(keyinput115), 
        .A(n6307), .ZN(n6315) );
  INV_X1 U8041 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8357) );
  AOI22_X1 U8042 ( .A1(n6497), .A2(keyinput64), .B1(keyinput105), .B2(n8357), 
        .ZN(n6308) );
  OAI221_X1 U8043 ( .B1(n6497), .B2(keyinput64), .C1(n8357), .C2(keyinput105), 
        .A(n6308), .ZN(n6314) );
  AOI22_X1 U8044 ( .A1(n6310), .A2(keyinput91), .B1(n6415), .B2(keyinput71), 
        .ZN(n6309) );
  OAI221_X1 U8045 ( .B1(n6310), .B2(keyinput91), .C1(n6415), .C2(keyinput71), 
        .A(n6309), .ZN(n6313) );
  INV_X1 U8046 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7496) );
  AOI22_X1 U8047 ( .A1(n6728), .A2(keyinput77), .B1(keyinput107), .B2(n7496), 
        .ZN(n6311) );
  OAI221_X1 U8048 ( .B1(n6728), .B2(keyinput77), .C1(n7496), .C2(keyinput107), 
        .A(n6311), .ZN(n6312) );
  NOR4_X1 U8049 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(n6475)
         );
  OAI22_X1 U8050 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput92), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(keyinput113), .ZN(n6316) );
  AOI221_X1 U8051 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput92), .C1(
        keyinput113), .C2(P2_DATAO_REG_4__SCAN_IN), .A(n6316), .ZN(n6323) );
  OAI22_X1 U8052 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput78), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(keyinput119), .ZN(n6317) );
  AOI221_X1 U8053 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput78), .C1(
        keyinput119), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n6317), .ZN(n6322) );
  OAI22_X1 U8054 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput87), .B1(
        keyinput75), .B2(P2_STATE_REG_SCAN_IN), .ZN(n6318) );
  AOI221_X1 U8055 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput87), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput75), .A(n6318), .ZN(n6321) );
  OAI22_X1 U8056 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput81), .B1(
        P2_REG2_REG_13__SCAN_IN), .B2(keyinput84), .ZN(n6319) );
  AOI221_X1 U8057 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput81), .C1(
        keyinput84), .C2(P2_REG2_REG_13__SCAN_IN), .A(n6319), .ZN(n6320) );
  NAND4_X1 U8058 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(n6342)
         );
  OAI22_X1 U8059 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput102), .B1(
        keyinput88), .B2(P2_REG0_REG_28__SCAN_IN), .ZN(n6324) );
  AOI221_X1 U8060 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput102), .C1(
        P2_REG0_REG_28__SCAN_IN), .C2(keyinput88), .A(n6324), .ZN(n6331) );
  OAI22_X1 U8061 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput109), .B1(
        keyinput125), .B2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6325) );
  AOI221_X1 U8062 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput109), .C1(
        P2_ADDR_REG_9__SCAN_IN), .C2(keyinput125), .A(n6325), .ZN(n6330) );
  OAI22_X1 U8063 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput110), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput70), .ZN(n6326) );
  AOI221_X1 U8064 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput110), .C1(
        keyinput70), .C2(P1_REG1_REG_18__SCAN_IN), .A(n6326), .ZN(n6329) );
  OAI22_X1 U8065 ( .A1(SI_5_), .A2(keyinput76), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(keyinput104), .ZN(n6327) );
  AOI221_X1 U8066 ( .B1(SI_5_), .B2(keyinput76), .C1(keyinput104), .C2(
        P2_REG2_REG_14__SCAN_IN), .A(n6327), .ZN(n6328) );
  NAND4_X1 U8067 ( .A1(n6331), .A2(n6330), .A3(n6329), .A4(n6328), .ZN(n6341)
         );
  OAI22_X1 U8068 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput90), .B1(
        keyinput118), .B2(P1_ADDR_REG_16__SCAN_IN), .ZN(n6332) );
  AOI221_X1 U8069 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput90), .C1(
        P1_ADDR_REG_16__SCAN_IN), .C2(keyinput118), .A(n6332), .ZN(n6339) );
  OAI22_X1 U8070 ( .A1(SI_15_), .A2(keyinput121), .B1(keyinput79), .B2(
        P2_REG3_REG_24__SCAN_IN), .ZN(n6333) );
  AOI221_X1 U8071 ( .B1(SI_15_), .B2(keyinput121), .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput79), .A(n6333), .ZN(n6338) );
  OAI22_X1 U8072 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput82), .B1(
        P2_REG0_REG_7__SCAN_IN), .B2(keyinput72), .ZN(n6334) );
  AOI221_X1 U8073 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput82), .C1(
        keyinput72), .C2(P2_REG0_REG_7__SCAN_IN), .A(n6334), .ZN(n6337) );
  OAI22_X1 U8074 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(keyinput74), .B1(
        P1_REG1_REG_30__SCAN_IN), .B2(keyinput117), .ZN(n6335) );
  AOI221_X1 U8075 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(keyinput74), .C1(
        keyinput117), .C2(P1_REG1_REG_30__SCAN_IN), .A(n6335), .ZN(n6336) );
  NAND4_X1 U8076 ( .A1(n6339), .A2(n6338), .A3(n6337), .A4(n6336), .ZN(n6340)
         );
  NOR3_X1 U8077 ( .A1(n6342), .A2(n6341), .A3(n6340), .ZN(n6384) );
  AOI22_X1 U8078 ( .A1(n4921), .A2(keyinput103), .B1(keyinput126), .B2(n6344), 
        .ZN(n6343) );
  OAI221_X1 U8079 ( .B1(n4921), .B2(keyinput103), .C1(n6344), .C2(keyinput126), 
        .A(n6343), .ZN(n6351) );
  INV_X1 U8080 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6500) );
  INV_X1 U8081 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U8082 ( .A1(n6500), .A2(keyinput99), .B1(n9910), .B2(keyinput120), 
        .ZN(n6345) );
  OAI221_X1 U8083 ( .B1(n6500), .B2(keyinput99), .C1(n9910), .C2(keyinput120), 
        .A(n6345), .ZN(n6350) );
  INV_X1 U8084 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9828) );
  INV_X1 U8085 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8906) );
  AOI22_X1 U8086 ( .A1(n9828), .A2(keyinput80), .B1(keyinput86), .B2(n8906), 
        .ZN(n6346) );
  OAI221_X1 U8087 ( .B1(n9828), .B2(keyinput80), .C1(n8906), .C2(keyinput86), 
        .A(n6346), .ZN(n6349) );
  INV_X1 U8088 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6695) );
  AOI22_X1 U8089 ( .A1(n6206), .A2(keyinput89), .B1(keyinput85), .B2(n6695), 
        .ZN(n6347) );
  OAI221_X1 U8090 ( .B1(n6206), .B2(keyinput89), .C1(n6695), .C2(keyinput85), 
        .A(n6347), .ZN(n6348) );
  NOR4_X1 U8091 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n6383)
         );
  INV_X1 U8092 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8636) );
  INV_X1 U8093 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U8094 ( .A1(n8636), .A2(keyinput101), .B1(n6704), .B2(keyinput66), 
        .ZN(n6352) );
  OAI221_X1 U8095 ( .B1(n8636), .B2(keyinput101), .C1(n6704), .C2(keyinput66), 
        .A(n6352), .ZN(n6360) );
  INV_X1 U8096 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9911) );
  INV_X1 U8097 ( .A(SI_16_), .ZN(n6354) );
  AOI22_X1 U8098 ( .A1(n9911), .A2(keyinput65), .B1(keyinput108), .B2(n6354), 
        .ZN(n6353) );
  OAI221_X1 U8099 ( .B1(n9911), .B2(keyinput65), .C1(n6354), .C2(keyinput108), 
        .A(n6353), .ZN(n6359) );
  INV_X1 U8100 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8448) );
  INV_X1 U8101 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8203) );
  AOI22_X1 U8102 ( .A1(n8448), .A2(keyinput68), .B1(n8203), .B2(keyinput122), 
        .ZN(n6355) );
  OAI221_X1 U8103 ( .B1(n8448), .B2(keyinput68), .C1(n8203), .C2(keyinput122), 
        .A(n6355), .ZN(n6358) );
  AOI22_X1 U8104 ( .A1(n6431), .A2(keyinput100), .B1(n7437), .B2(keyinput83), 
        .ZN(n6356) );
  OAI221_X1 U8105 ( .B1(n6431), .B2(keyinput100), .C1(n7437), .C2(keyinput83), 
        .A(n6356), .ZN(n6357) );
  NOR4_X1 U8106 ( .A1(n6360), .A2(n6359), .A3(n6358), .A4(n6357), .ZN(n6382)
         );
  AOI22_X1 U8107 ( .A1(n9608), .A2(keyinput95), .B1(n6845), .B2(keyinput123), 
        .ZN(n6361) );
  OAI221_X1 U8108 ( .B1(n9608), .B2(keyinput95), .C1(n6845), .C2(keyinput123), 
        .A(n6361), .ZN(n6362) );
  INV_X1 U8109 ( .A(n6362), .ZN(n6370) );
  XNOR2_X1 U8110 ( .A(keyinput93), .B(P1_ADDR_REG_6__SCAN_IN), .ZN(n6369) );
  XNOR2_X1 U8111 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput111), .ZN(n6366) );
  XNOR2_X1 U8112 ( .A(SI_4_), .B(keyinput98), .ZN(n6365) );
  XNOR2_X1 U8113 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput96), .ZN(n6364) );
  XNOR2_X1 U8114 ( .A(keyinput127), .B(P1_REG0_REG_10__SCAN_IN), .ZN(n6363) );
  AND4_X1 U8115 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n6368)
         );
  XNOR2_X1 U8116 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput114), .ZN(n6367) );
  NAND4_X1 U8117 ( .A1(n6370), .A2(n6369), .A3(n6368), .A4(n6367), .ZN(n6380)
         );
  OAI22_X1 U8118 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(keyinput69), .B1(
        keyinput112), .B2(P2_ADDR_REG_4__SCAN_IN), .ZN(n6371) );
  AOI221_X1 U8119 ( .B1(P1_REG3_REG_7__SCAN_IN), .B2(keyinput69), .C1(
        P2_ADDR_REG_4__SCAN_IN), .C2(keyinput112), .A(n6371), .ZN(n6378) );
  OAI22_X1 U8120 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput97), .B1(
        P1_REG2_REG_11__SCAN_IN), .B2(keyinput73), .ZN(n6372) );
  AOI221_X1 U8121 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput97), .C1(
        keyinput73), .C2(P1_REG2_REG_11__SCAN_IN), .A(n6372), .ZN(n6377) );
  OAI22_X1 U8122 ( .A1(SI_26_), .A2(keyinput94), .B1(P1_REG1_REG_1__SCAN_IN), 
        .B2(keyinput106), .ZN(n6373) );
  AOI221_X1 U8123 ( .B1(SI_26_), .B2(keyinput94), .C1(keyinput106), .C2(
        P1_REG1_REG_1__SCAN_IN), .A(n6373), .ZN(n6376) );
  OAI22_X1 U8124 ( .A1(SI_2_), .A2(keyinput67), .B1(keyinput116), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6374) );
  AOI221_X1 U8125 ( .B1(SI_2_), .B2(keyinput67), .C1(P2_REG0_REG_22__SCAN_IN), 
        .C2(keyinput116), .A(n6374), .ZN(n6375) );
  NAND4_X1 U8126 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n6379)
         );
  NOR2_X1 U8127 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  AND4_X1 U8128 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(n6474)
         );
  AOI22_X1 U8129 ( .A1(P2_D_REG_0__SCAN_IN), .A2(keyinput25), .B1(
        P1_REG1_REG_28__SCAN_IN), .B2(keyinput62), .ZN(n6385) );
  OAI221_X1 U8130 ( .B1(P2_D_REG_0__SCAN_IN), .B2(keyinput25), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput62), .A(n6385), .ZN(n6392) );
  AOI22_X1 U8131 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(keyinput54), .B1(
        P1_REG2_REG_11__SCAN_IN), .B2(keyinput9), .ZN(n6386) );
  OAI221_X1 U8132 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(keyinput54), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(keyinput9), .A(n6386), .ZN(n6391) );
  AOI22_X1 U8133 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput38), .B1(
        P1_REG3_REG_28__SCAN_IN), .B2(keyinput0), .ZN(n6387) );
  OAI221_X1 U8134 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput38), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput0), .A(n6387), .ZN(n6390) );
  AOI22_X1 U8135 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput55), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput17), .ZN(n6388) );
  OAI221_X1 U8136 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput55), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput17), .A(n6388), .ZN(n6389) );
  NOR4_X1 U8137 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .ZN(n6452)
         );
  AOI22_X1 U8138 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(keyinput61), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput11), .ZN(n6393) );
  OAI221_X1 U8139 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(keyinput61), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput11), .A(n6393), .ZN(n6400) );
  AOI22_X1 U8140 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput29), .B1(
        P2_ADDR_REG_17__SCAN_IN), .B2(keyinput4), .ZN(n6394) );
  OAI221_X1 U8141 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput29), .C1(
        P2_ADDR_REG_17__SCAN_IN), .C2(keyinput4), .A(n6394), .ZN(n6399) );
  AOI22_X1 U8142 ( .A1(P1_D_REG_27__SCAN_IN), .A2(keyinput56), .B1(
        P1_D_REG_25__SCAN_IN), .B2(keyinput1), .ZN(n6395) );
  OAI221_X1 U8143 ( .B1(P1_D_REG_27__SCAN_IN), .B2(keyinput56), .C1(
        P1_D_REG_25__SCAN_IN), .C2(keyinput1), .A(n6395), .ZN(n6398) );
  AOI22_X1 U8144 ( .A1(P1_REG0_REG_31__SCAN_IN), .A2(keyinput21), .B1(SI_5_), 
        .B2(keyinput12), .ZN(n6396) );
  OAI221_X1 U8145 ( .B1(P1_REG0_REG_31__SCAN_IN), .B2(keyinput21), .C1(SI_5_), 
        .C2(keyinput12), .A(n6396), .ZN(n6397) );
  NOR4_X1 U8146 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6451)
         );
  AOI22_X1 U8147 ( .A1(n7803), .A2(keyinput51), .B1(keyinput6), .B2(n6402), 
        .ZN(n6401) );
  OAI221_X1 U8148 ( .B1(n7803), .B2(keyinput51), .C1(n6402), .C2(keyinput6), 
        .A(n6401), .ZN(n6411) );
  AOI22_X1 U8149 ( .A1(n7496), .A2(keyinput43), .B1(n6704), .B2(keyinput2), 
        .ZN(n6403) );
  OAI221_X1 U8150 ( .B1(n7496), .B2(keyinput43), .C1(n6704), .C2(keyinput2), 
        .A(n6403), .ZN(n6410) );
  INV_X1 U8151 ( .A(SI_15_), .ZN(n6405) );
  AOI22_X1 U8152 ( .A1(n6405), .A2(keyinput57), .B1(n7606), .B2(keyinput28), 
        .ZN(n6404) );
  OAI221_X1 U8153 ( .B1(n6405), .B2(keyinput57), .C1(n7606), .C2(keyinput28), 
        .A(n6404), .ZN(n6409) );
  AOI22_X1 U8154 ( .A1(n7437), .A2(keyinput19), .B1(n6407), .B2(keyinput30), 
        .ZN(n6406) );
  OAI221_X1 U8155 ( .B1(n7437), .B2(keyinput19), .C1(n6407), .C2(keyinput30), 
        .A(n6406), .ZN(n6408) );
  NOR4_X1 U8156 ( .A1(n6411), .A2(n6410), .A3(n6409), .A4(n6408), .ZN(n6450)
         );
  AOI22_X1 U8157 ( .A1(n8357), .A2(keyinput41), .B1(n6845), .B2(keyinput59), 
        .ZN(n6412) );
  OAI221_X1 U8158 ( .B1(n8357), .B2(keyinput41), .C1(n6845), .C2(keyinput59), 
        .A(n6412), .ZN(n6413) );
  INV_X1 U8159 ( .A(n6413), .ZN(n6429) );
  INV_X1 U8160 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U8161 ( .A1(n6415), .A2(keyinput7), .B1(n6799), .B2(keyinput26), 
        .ZN(n6414) );
  OAI221_X1 U8162 ( .B1(n6415), .B2(keyinput7), .C1(n6799), .C2(keyinput26), 
        .A(n6414), .ZN(n6418) );
  AOI22_X1 U8163 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(keyinput53), .B1(
        P1_REG3_REG_7__SCAN_IN), .B2(keyinput5), .ZN(n6416) );
  OAI221_X1 U8164 ( .B1(P1_REG1_REG_30__SCAN_IN), .B2(keyinput53), .C1(
        P1_REG3_REG_7__SCAN_IN), .C2(keyinput5), .A(n6416), .ZN(n6417) );
  NOR2_X1 U8165 ( .A1(n6418), .A2(n6417), .ZN(n6428) );
  INV_X1 U8166 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8725) );
  AOI22_X1 U8167 ( .A1(n8725), .A2(keyinput40), .B1(n6420), .B2(keyinput47), 
        .ZN(n6419) );
  OAI221_X1 U8168 ( .B1(n8725), .B2(keyinput40), .C1(n6420), .C2(keyinput47), 
        .A(n6419), .ZN(n6423) );
  AOI22_X1 U8169 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput52), .B1(
        P1_REG3_REG_24__SCAN_IN), .B2(keyinput10), .ZN(n6421) );
  OAI221_X1 U8170 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput52), .C1(
        P1_REG3_REG_24__SCAN_IN), .C2(keyinput10), .A(n6421), .ZN(n6422) );
  NOR2_X1 U8171 ( .A1(n6423), .A2(n6422), .ZN(n6427) );
  AOI22_X1 U8172 ( .A1(n8301), .A2(keyinput15), .B1(n9608), .B2(keyinput31), 
        .ZN(n6424) );
  OAI221_X1 U8173 ( .B1(n8301), .B2(keyinput15), .C1(n9608), .C2(keyinput31), 
        .A(n6424), .ZN(n6425) );
  INV_X1 U8174 ( .A(n6425), .ZN(n6426) );
  NAND4_X1 U8175 ( .A1(n6429), .A2(n6428), .A3(n6427), .A4(n6426), .ZN(n6448)
         );
  INV_X1 U8176 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U8177 ( .A1(n9974), .A2(keyinput63), .B1(n6678), .B2(keyinput33), 
        .ZN(n6430) );
  OAI221_X1 U8178 ( .B1(n9974), .B2(keyinput63), .C1(n6678), .C2(keyinput33), 
        .A(n6430), .ZN(n6437) );
  XNOR2_X1 U8179 ( .A(n6431), .B(keyinput36), .ZN(n6435) );
  XNOR2_X1 U8180 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput27), .ZN(n6434) );
  XNOR2_X1 U8181 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput23), .ZN(n6433) );
  XNOR2_X1 U8182 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput32), .ZN(n6432) );
  NAND4_X1 U8183 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n6436)
         );
  NOR2_X1 U8184 ( .A1(n6437), .A2(n6436), .ZN(n6446) );
  AOI22_X1 U8185 ( .A1(n6968), .A2(keyinput18), .B1(keyinput60), .B2(n8816), 
        .ZN(n6438) );
  OAI221_X1 U8186 ( .B1(n6968), .B2(keyinput18), .C1(n8816), .C2(keyinput60), 
        .A(n6438), .ZN(n6444) );
  XNOR2_X1 U8187 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput14), .ZN(n6442) );
  XNOR2_X1 U8188 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput50), .ZN(n6441) );
  XNOR2_X1 U8189 ( .A(SI_4_), .B(keyinput34), .ZN(n6440) );
  XNOR2_X1 U8190 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput42), .ZN(n6439) );
  NAND4_X1 U8191 ( .A1(n6442), .A2(n6441), .A3(n6440), .A4(n6439), .ZN(n6443)
         );
  NOR2_X1 U8192 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  NAND2_X1 U8193 ( .A1(n6446), .A2(n6445), .ZN(n6447) );
  NOR2_X1 U8194 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND4_X1 U8195 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n6473)
         );
  AOI22_X1 U8196 ( .A1(n8203), .A2(keyinput58), .B1(n4921), .B2(keyinput39), 
        .ZN(n6453) );
  AOI22_X1 U8197 ( .A1(n6728), .A2(keyinput13), .B1(keyinput22), .B2(n8906), 
        .ZN(n6454) );
  OAI221_X1 U8198 ( .B1(n6728), .B2(keyinput13), .C1(n8906), .C2(keyinput22), 
        .A(n6454), .ZN(n6460) );
  AOI22_X1 U8199 ( .A1(n8636), .A2(keyinput37), .B1(n9828), .B2(keyinput16), 
        .ZN(n6455) );
  OAI221_X1 U8200 ( .B1(n8636), .B2(keyinput37), .C1(n9828), .C2(keyinput16), 
        .A(n6455), .ZN(n6459) );
  INV_X1 U8201 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10066) );
  AOI22_X1 U8202 ( .A1(n10066), .A2(keyinput45), .B1(n6457), .B2(keyinput24), 
        .ZN(n6456) );
  OAI221_X1 U8203 ( .B1(n10066), .B2(keyinput45), .C1(n6457), .C2(keyinput24), 
        .A(n6456), .ZN(n6458) );
  NOR4_X1 U8204 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n6471)
         );
  AOI22_X1 U8205 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput48), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(keyinput49), .ZN(n6462) );
  OAI221_X1 U8206 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput48), .C1(
        P2_DATAO_REG_4__SCAN_IN), .C2(keyinput49), .A(n6462), .ZN(n6469) );
  AOI22_X1 U8207 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput46), .B1(SI_16_), 
        .B2(keyinput44), .ZN(n6463) );
  OAI221_X1 U8208 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput46), .C1(SI_16_), 
        .C2(keyinput44), .A(n6463), .ZN(n6468) );
  AOI22_X1 U8209 ( .A1(P2_REG0_REG_7__SCAN_IN), .A2(keyinput8), .B1(SI_2_), 
        .B2(keyinput3), .ZN(n6464) );
  OAI221_X1 U8210 ( .B1(P2_REG0_REG_7__SCAN_IN), .B2(keyinput8), .C1(SI_2_), 
        .C2(keyinput3), .A(n6464), .ZN(n6467) );
  AOI22_X1 U8211 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput20), .B1(
        P1_REG1_REG_29__SCAN_IN), .B2(keyinput35), .ZN(n6465) );
  OAI221_X1 U8212 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput20), .C1(
        P1_REG1_REG_29__SCAN_IN), .C2(keyinput35), .A(n6465), .ZN(n6466) );
  NOR4_X1 U8213 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n6470)
         );
  NAND2_X1 U8214 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  AOI211_X1 U8215 ( .C1(n6475), .C2(n6474), .A(n6473), .B(n6472), .ZN(n6476)
         );
  XNOR2_X1 U8216 ( .A(n6477), .B(n6476), .ZN(P1_U3517) );
  INV_X1 U8217 ( .A(n6493), .ZN(n6491) );
  NAND2_X1 U8218 ( .A1(n7827), .A2(n9137), .ZN(n6479) );
  NAND2_X1 U8219 ( .A1(n5060), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8220 ( .A1(n9735), .A2(n5639), .ZN(n6481) );
  OR2_X1 U8221 ( .A1(n7866), .A2(n5014), .ZN(n6480) );
  NAND2_X1 U8222 ( .A1(n6481), .A2(n6480), .ZN(n6483) );
  XNOR2_X1 U8223 ( .A(n6483), .B(n6482), .ZN(n6488) );
  NAND2_X1 U8224 ( .A1(n9735), .A2(n5697), .ZN(n6485) );
  OAI21_X1 U8225 ( .B1(n7866), .B2(n6486), .A(n6485), .ZN(n6487) );
  XNOR2_X1 U8226 ( .A(n6488), .B(n6487), .ZN(n6492) );
  NOR2_X1 U8227 ( .A1(n6495), .A2(n9122), .ZN(n6489) );
  AND2_X1 U8228 ( .A1(n6492), .A2(n6489), .ZN(n6490) );
  NAND2_X1 U8229 ( .A1(n6491), .A2(n6490), .ZN(n6511) );
  INV_X1 U8230 ( .A(n6492), .ZN(n6496) );
  NAND3_X1 U8231 ( .A1(n6493), .A2(n9113), .A3(n6496), .ZN(n6510) );
  INV_X1 U8232 ( .A(n6494), .ZN(n6495) );
  NAND3_X1 U8233 ( .A1(n6496), .A2(n6495), .A3(n9113), .ZN(n6508) );
  OAI22_X1 U8234 ( .A1(n9126), .A2(n9543), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6497), .ZN(n6506) );
  NAND2_X1 U8235 ( .A1(n7859), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6504) );
  INV_X1 U8236 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6498) );
  OR2_X1 U8237 ( .A1(n7862), .A2(n6498), .ZN(n6503) );
  OR2_X1 U8238 ( .A1(n4319), .A2(n7848), .ZN(n6502) );
  OR2_X1 U8239 ( .A1(n5738), .A2(n6500), .ZN(n6501) );
  OAI22_X1 U8240 ( .A1(n9129), .A2(n9523), .B1(n9530), .B2(n9115), .ZN(n6505)
         );
  AOI211_X1 U8241 ( .C1(n9735), .C2(n9082), .A(n6506), .B(n6505), .ZN(n6507)
         );
  NAND3_X1 U8242 ( .A1(n6511), .A2(n6510), .A3(n6509), .ZN(P1_U3220) );
  NAND2_X1 U8243 ( .A1(n6570), .A2(n8171), .ZN(n6513) );
  NAND2_X1 U8244 ( .A1(n6513), .A2(n7112), .ZN(n6596) );
  NAND2_X1 U8245 ( .A1(n6596), .A2(n5821), .ZN(n6514) );
  NAND2_X1 U8246 ( .A1(n6514), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  MUX2_X1 U8247 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4462), .Z(n6521) );
  XNOR2_X1 U8248 ( .A(n6516), .B(n7010), .ZN(n6996) );
  INV_X1 U8249 ( .A(n6987), .ZN(n6515) );
  AND2_X1 U8250 ( .A1(n6515), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6995) );
  INV_X1 U8251 ( .A(n7010), .ZN(n6518) );
  INV_X1 U8252 ( .A(n6516), .ZN(n6517) );
  OAI22_X1 U8253 ( .A1(n6996), .A2(n6995), .B1(n6518), .B2(n6517), .ZN(n7037)
         );
  MUX2_X1 U8254 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4462), .Z(n6519) );
  XOR2_X1 U8255 ( .A(n6939), .B(n6520), .Z(n6934) );
  NAND2_X1 U8256 ( .A1(n6935), .A2(n6934), .ZN(n6933) );
  OAI21_X1 U8257 ( .B1(n6520), .B2(n6939), .A(n6933), .ZN(n7133) );
  XNOR2_X1 U8258 ( .A(n6521), .B(n7118), .ZN(n7134) );
  NOR2_X1 U8259 ( .A1(n7133), .A2(n7134), .ZN(n7132) );
  XNOR2_X1 U8260 ( .A(n6522), .B(n6659), .ZN(n7061) );
  INV_X1 U8261 ( .A(n6522), .ZN(n6523) );
  OAI22_X1 U8262 ( .A1(n7062), .A2(n7061), .B1(n4831), .B2(n6523), .ZN(n7183)
         );
  INV_X1 U8263 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6525) );
  INV_X1 U8264 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6524) );
  MUX2_X1 U8265 ( .A(n6525), .B(n6524), .S(n4462), .Z(n6526) );
  INV_X1 U8266 ( .A(n6664), .ZN(n7200) );
  NAND2_X1 U8267 ( .A1(n6526), .A2(n7200), .ZN(n6527) );
  OAI21_X1 U8268 ( .B1(n6526), .B2(n7200), .A(n6527), .ZN(n7182) );
  NOR2_X1 U8269 ( .A1(n7183), .A2(n7182), .ZN(n7321) );
  INV_X1 U8270 ( .A(n6527), .ZN(n7320) );
  INV_X1 U8271 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6529) );
  INV_X1 U8272 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U8273 ( .A(n6529), .B(n6528), .S(n4462), .Z(n6530) );
  NAND2_X1 U8274 ( .A1(n6530), .A2(n4753), .ZN(n7362) );
  INV_X1 U8275 ( .A(n6530), .ZN(n6531) );
  NAND2_X1 U8276 ( .A1(n6531), .A2(n7329), .ZN(n6532) );
  AND2_X1 U8277 ( .A1(n7362), .A2(n6532), .ZN(n7319) );
  OAI21_X1 U8278 ( .B1(n7321), .B2(n7320), .A(n7319), .ZN(n7363) );
  INV_X1 U8279 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7618) );
  INV_X1 U8280 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6582) );
  MUX2_X1 U8281 ( .A(n7618), .B(n6582), .S(n4462), .Z(n6533) );
  INV_X1 U8282 ( .A(n6675), .ZN(n7374) );
  NAND2_X1 U8283 ( .A1(n6533), .A2(n7374), .ZN(n6536) );
  INV_X1 U8284 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U8285 ( .A1(n6534), .A2(n6675), .ZN(n6535) );
  NAND2_X1 U8286 ( .A1(n6536), .A2(n6535), .ZN(n7361) );
  INV_X1 U8287 ( .A(n6536), .ZN(n7467) );
  INV_X1 U8288 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7762) );
  INV_X1 U8289 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U8290 ( .A(n7762), .B(n6537), .S(n4462), .Z(n6539) );
  NAND2_X1 U8291 ( .A1(n6539), .A2(n6538), .ZN(n7540) );
  INV_X1 U8292 ( .A(n6539), .ZN(n6540) );
  NAND2_X1 U8293 ( .A1(n6540), .A2(n7474), .ZN(n6541) );
  AND2_X1 U8294 ( .A1(n7540), .A2(n6541), .ZN(n7466) );
  OAI21_X1 U8295 ( .B1(n7468), .B2(n7467), .A(n7466), .ZN(n7541) );
  INV_X1 U8296 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8784) );
  INV_X1 U8297 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10088) );
  MUX2_X1 U8298 ( .A(n8784), .B(n10088), .S(n4462), .Z(n6542) );
  NAND2_X1 U8299 ( .A1(n6542), .A2(n6543), .ZN(n6546) );
  INV_X1 U8300 ( .A(n6542), .ZN(n6544) );
  INV_X1 U8301 ( .A(n6543), .ZN(n7557) );
  NAND2_X1 U8302 ( .A1(n6544), .A2(n7557), .ZN(n6545) );
  NAND2_X1 U8303 ( .A1(n6546), .A2(n6545), .ZN(n7539) );
  AOI21_X1 U8304 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7651) );
  INV_X1 U8305 ( .A(n6546), .ZN(n7650) );
  INV_X1 U8306 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8767) );
  INV_X1 U8307 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8308 ( .A1(n6548), .A2(n6614), .ZN(n7736) );
  INV_X1 U8309 ( .A(n6548), .ZN(n6549) );
  INV_X1 U8310 ( .A(n6614), .ZN(n7658) );
  NAND2_X1 U8311 ( .A1(n6549), .A2(n7658), .ZN(n6550) );
  AND2_X1 U8312 ( .A1(n7736), .A2(n6550), .ZN(n7649) );
  OAI21_X1 U8313 ( .B1(n7651), .B2(n7650), .A(n7649), .ZN(n7737) );
  INV_X1 U8314 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8748) );
  INV_X1 U8315 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8844) );
  MUX2_X1 U8316 ( .A(n8748), .B(n8844), .S(n4462), .Z(n6551) );
  NAND2_X1 U8317 ( .A1(n6551), .A2(n6616), .ZN(n6554) );
  INV_X1 U8318 ( .A(n6551), .ZN(n6552) );
  INV_X1 U8319 ( .A(n6616), .ZN(n7745) );
  NAND2_X1 U8320 ( .A1(n6552), .A2(n7745), .ZN(n6553) );
  NAND2_X1 U8321 ( .A1(n6554), .A2(n6553), .ZN(n7735) );
  INV_X1 U8322 ( .A(n6554), .ZN(n7782) );
  INV_X1 U8323 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6555) );
  INV_X1 U8324 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8840) );
  MUX2_X1 U8325 ( .A(n6555), .B(n8840), .S(n4462), .Z(n6556) );
  NAND2_X1 U8326 ( .A1(n6556), .A2(n6618), .ZN(n6563) );
  INV_X1 U8327 ( .A(n6556), .ZN(n6557) );
  INV_X1 U8328 ( .A(n6618), .ZN(n7790) );
  NAND2_X1 U8329 ( .A1(n6557), .A2(n7790), .ZN(n6558) );
  AND2_X1 U8330 ( .A1(n6563), .A2(n6558), .ZN(n7781) );
  OAI21_X1 U8331 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7780) );
  INV_X1 U8332 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7883) );
  MUX2_X1 U8333 ( .A(n8725), .B(n7883), .S(n4462), .Z(n6559) );
  NAND2_X1 U8334 ( .A1(n6559), .A2(n6619), .ZN(n8395) );
  INV_X1 U8335 ( .A(n6559), .ZN(n6560) );
  INV_X1 U8336 ( .A(n6619), .ZN(n8402) );
  NAND2_X1 U8337 ( .A1(n6560), .A2(n8402), .ZN(n6561) );
  NAND2_X1 U8338 ( .A1(n8395), .A2(n6561), .ZN(n6562) );
  AOI21_X1 U8339 ( .B1(n7780), .B2(n6563), .A(n6562), .ZN(n8397) );
  INV_X1 U8340 ( .A(n8397), .ZN(n6565) );
  NAND3_X1 U8341 ( .A1(n7780), .A2(n6563), .A3(n6562), .ZN(n6564) );
  NAND2_X1 U8342 ( .A1(P2_U3893), .A2(n6177), .ZN(n8517) );
  AOI21_X1 U8343 ( .B1(n6565), .B2(n6564), .A(n8517), .ZN(n6625) );
  INV_X1 U8344 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6566) );
  NOR2_X1 U8345 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6566), .ZN(n8216) );
  NOR2_X1 U8346 ( .A1(n4462), .A2(P2_U3151), .ZN(n7821) );
  NAND2_X1 U8347 ( .A1(n6596), .A2(n7821), .ZN(n6568) );
  MUX2_X1 U8348 ( .A(n6568), .B(n8391), .S(n6567), .Z(n8506) );
  INV_X1 U8349 ( .A(n7112), .ZN(n6569) );
  NOR2_X1 U8350 ( .A1(n6570), .A2(n6569), .ZN(n6571) );
  INV_X1 U8351 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7526) );
  OAI22_X1 U8352 ( .A1(n8506), .A2(n8402), .B1(n8505), .B2(n7526), .ZN(n6624)
         );
  NAND2_X1 U8353 ( .A1(n7557), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6588) );
  OAI21_X1 U8354 ( .B1(n7557), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6588), .ZN(
        n7544) );
  INV_X1 U8355 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U8356 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10081), .S(n7038), .Z(n7045)
         );
  AND2_X1 U8357 ( .A1(n6993), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6572) );
  OAI21_X1 U8358 ( .B1(n7010), .B2(n6572), .A(n6573), .ZN(n7003) );
  INV_X1 U8359 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7002) );
  OR2_X1 U8360 ( .A1(n7003), .A2(n7002), .ZN(n7005) );
  NAND2_X1 U8361 ( .A1(n7005), .A2(n6573), .ZN(n7044) );
  NAND2_X1 U8362 ( .A1(n7045), .A2(n7044), .ZN(n7043) );
  NAND2_X1 U8363 ( .A1(n7038), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8364 ( .A1(n7043), .A2(n6574), .ZN(n6575) );
  INV_X1 U8365 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7873) );
  XNOR2_X1 U8366 ( .A(n7118), .B(n7873), .ZN(n7122) );
  NAND2_X1 U8367 ( .A1(n6576), .A2(n7122), .ZN(n7127) );
  NAND2_X1 U8368 ( .A1(n7118), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U8369 ( .A1(n7127), .A2(n6577), .ZN(n6578) );
  INV_X1 U8370 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10083) );
  MUX2_X1 U8371 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6524), .S(n6664), .Z(n7184)
         );
  NAND2_X1 U8372 ( .A1(n6579), .A2(n7184), .ZN(n7189) );
  NAND2_X1 U8373 ( .A1(n6664), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8374 ( .A1(n7189), .A2(n6580), .ZN(n6581) );
  XNOR2_X1 U8375 ( .A(n6675), .B(n6582), .ZN(n7366) );
  NAND2_X1 U8376 ( .A1(n6583), .A2(n7366), .ZN(n7371) );
  NAND2_X1 U8377 ( .A1(n6675), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8378 ( .A1(n7371), .A2(n6584), .ZN(n6585) );
  INV_X1 U8379 ( .A(n6588), .ZN(n6589) );
  NOR2_X1 U8380 ( .A1(n6614), .A2(n6590), .ZN(n6591) );
  XOR2_X1 U8381 ( .A(n6590), .B(n7658), .Z(n7648) );
  NOR2_X1 U8382 ( .A1(n6547), .A2(n7648), .ZN(n7647) );
  AOI22_X1 U8383 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6616), .B1(n7745), .B2(
        n8844), .ZN(n7733) );
  NOR2_X1 U8384 ( .A1(n7734), .A2(n7733), .ZN(n7732) );
  NOR2_X1 U8385 ( .A1(n6618), .A2(n6592), .ZN(n6593) );
  XNOR2_X1 U8386 ( .A(n6618), .B(n6592), .ZN(n7779) );
  NOR2_X1 U8387 ( .A1(n8840), .A2(n7779), .ZN(n7778) );
  AOI22_X1 U8388 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6619), .B1(n8402), .B2(
        n7883), .ZN(n6594) );
  NOR2_X1 U8389 ( .A1(n6595), .A2(n6594), .ZN(n8393) );
  AOI21_X1 U8390 ( .B1(n6595), .B2(n6594), .A(n8393), .ZN(n6622) );
  NOR2_X1 U8391 ( .A1(n6177), .A2(P2_U3151), .ZN(n7830) );
  AND2_X1 U8392 ( .A1(n6596), .A2(n7830), .ZN(n6986) );
  NAND2_X1 U8393 ( .A1(n7557), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6612) );
  OAI21_X1 U8394 ( .B1(n7557), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6612), .ZN(
        n7547) );
  INV_X1 U8395 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6597) );
  AND2_X1 U8396 ( .A1(n6993), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6598) );
  OAI21_X1 U8397 ( .B1(n7010), .B2(n6598), .A(n6599), .ZN(n6998) );
  INV_X1 U8398 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6997) );
  OR2_X1 U8399 ( .A1(n6998), .A2(n6997), .ZN(n7000) );
  NAND2_X1 U8400 ( .A1(n7000), .A2(n6599), .ZN(n7040) );
  NAND2_X1 U8401 ( .A1(n7038), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8402 ( .A1(n6601), .A2(n6939), .ZN(n6602) );
  OAI21_X1 U8403 ( .B1(n6601), .B2(n6939), .A(n6602), .ZN(n6926) );
  INV_X1 U8404 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8405 ( .A1(n6924), .A2(n6602), .ZN(n7120) );
  OR2_X1 U8406 ( .A1(n7118), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8407 ( .A1(n7118), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6604) );
  AND2_X1 U8408 ( .A1(n6603), .A2(n6604), .ZN(n7121) );
  INV_X1 U8409 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U8410 ( .A1(n7192), .A2(n4828), .ZN(n6605) );
  MUX2_X1 U8411 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6525), .S(n6664), .Z(n7190)
         );
  NAND2_X1 U8412 ( .A1(n6605), .A2(n7190), .ZN(n7194) );
  NAND2_X1 U8413 ( .A1(n6664), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8414 ( .A1(n7194), .A2(n6606), .ZN(n6607) );
  XNOR2_X1 U8415 ( .A(n6675), .B(n7618), .ZN(n7355) );
  NAND2_X1 U8416 ( .A1(n6608), .A2(n7355), .ZN(n7357) );
  NAND2_X1 U8417 ( .A1(n6675), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U8418 ( .A1(n7357), .A2(n6609), .ZN(n6610) );
  INV_X1 U8419 ( .A(n6612), .ZN(n6613) );
  AOI22_X1 U8420 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6616), .B1(n7745), .B2(
        n8748), .ZN(n7740) );
  XNOR2_X1 U8421 ( .A(n6618), .B(n6617), .ZN(n7787) );
  AOI22_X1 U8422 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6619), .B1(n8402), .B2(
        n8725), .ZN(n6620) );
  AOI21_X1 U8423 ( .B1(n4408), .B2(n6620), .A(n8401), .ZN(n6621) );
  AND2_X1 U8424 ( .A1(n6986), .A2(n8493), .ZN(n8509) );
  OAI22_X1 U8425 ( .A1(n6622), .A2(n8491), .B1(n6621), .B2(n8484), .ZN(n6623)
         );
  OR4_X1 U8426 ( .A1(n6625), .A2(n8216), .A3(n6624), .A4(n6623), .ZN(P2_U3196)
         );
  INV_X1 U8427 ( .A(n6626), .ZN(n6627) );
  OR2_X2 U8428 ( .A1(n6628), .A2(n6627), .ZN(n9412) );
  INV_X1 U8429 ( .A(n9412), .ZN(P1_U3973) );
  XNOR2_X1 U8430 ( .A(n6723), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6636) );
  OR2_X1 U8431 ( .A1(n6681), .A2(n6629), .ZN(n6635) );
  NOR3_X1 U8432 ( .A1(n6636), .A2(n6681), .A3(n6629), .ZN(n6722) );
  NAND2_X1 U8433 ( .A1(n9194), .A2(n6632), .ZN(n6630) );
  NAND2_X1 U8434 ( .A1(n6631), .A2(n6630), .ZN(n6638) );
  INV_X1 U8435 ( .A(n6638), .ZN(n6634) );
  OR2_X1 U8436 ( .A1(n6632), .A2(P1_U3086), .ZN(n9387) );
  INV_X1 U8437 ( .A(n9387), .ZN(n6633) );
  OR2_X1 U8438 ( .A1(n9380), .A2(n6633), .ZN(n6639) );
  AND2_X1 U8439 ( .A1(n6634), .A2(n6639), .ZN(n6683) );
  AND2_X1 U8440 ( .A1(n6683), .A2(n7858), .ZN(n9488) );
  INV_X1 U8441 ( .A(n9488), .ZN(n9491) );
  AOI211_X1 U8442 ( .C1(n6636), .C2(n6635), .A(n6722), .B(n9491), .ZN(n6644)
         );
  NAND2_X1 U8443 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6801) );
  XNOR2_X1 U8444 ( .A(n6723), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U8445 ( .A1(n6637), .A2(n6801), .ZN(n6709) );
  NOR2_X1 U8446 ( .A1(n6679), .A2(n7858), .ZN(n9379) );
  NAND2_X1 U8447 ( .A1(n6683), .A2(n9379), .ZN(n9484) );
  AOI211_X1 U8448 ( .C1(n6801), .C2(n6637), .A(n6709), .B(n9484), .ZN(n6643)
         );
  NAND2_X1 U8449 ( .A1(n6683), .A2(n6679), .ZN(n9490) );
  INV_X1 U8450 ( .A(n6723), .ZN(n6646) );
  NOR2_X1 U8451 ( .A1(n9490), .A2(n6646), .ZN(n6642) );
  NAND2_X1 U8452 ( .A1(n6639), .A2(n6638), .ZN(n9502) );
  INV_X1 U8453 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6640) );
  OAI22_X1 U8454 ( .A1(n9502), .A2(n6640), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6856), .ZN(n6641) );
  OR4_X1 U8455 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(P1_U3244)
         );
  AND2_X1 U8456 ( .A1(n9136), .A2(P1_U3086), .ZN(n7604) );
  INV_X2 U8457 ( .A(n7604), .ZN(n9807) );
  NOR2_X1 U8458 ( .A1(n9136), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9804) );
  AOI22_X1 U8459 ( .A1(n9804), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9417), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6645) );
  OAI21_X1 U8460 ( .B1(n6655), .B2(n9807), .A(n6645), .ZN(P1_U3353) );
  INV_X1 U8461 ( .A(n9804), .ZN(n7825) );
  OAI222_X1 U8462 ( .A1(n7825), .A2(n6647), .B1(n9807), .B2(n6653), .C1(
        P1_U3086), .C2(n6646), .ZN(P1_U3354) );
  INV_X1 U8463 ( .A(n6724), .ZN(n6782) );
  OAI222_X1 U8464 ( .A1(n7825), .A2(n6648), .B1(n9807), .B2(n6657), .C1(
        P1_U3086), .C2(n6782), .ZN(P1_U3352) );
  INV_X1 U8465 ( .A(n6725), .ZN(n6818) );
  OAI222_X1 U8466 ( .A1(n7825), .A2(n6649), .B1(n9807), .B2(n6651), .C1(
        P1_U3086), .C2(n6818), .ZN(P1_U3351) );
  AND2_X1 U8467 ( .A1(n7969), .A2(P2_U3151), .ZN(n8951) );
  INV_X2 U8468 ( .A(n8951), .ZN(n8953) );
  AND2_X1 U8469 ( .A1(n6650), .A2(P2_U3151), .ZN(n7607) );
  INV_X2 U8470 ( .A(n7607), .ZN(n8955) );
  OAI222_X1 U8471 ( .A1(n8953), .A2(n6652), .B1(n8955), .B2(n6651), .C1(
        P2_U3151), .C2(n7118), .ZN(P2_U3291) );
  OAI222_X1 U8472 ( .A1(n8953), .A2(n6654), .B1(n8955), .B2(n6653), .C1(
        P2_U3151), .C2(n7010), .ZN(P2_U3294) );
  OAI222_X1 U8473 ( .A1(n8953), .A2(n6656), .B1(n8955), .B2(n6655), .C1(
        P2_U3151), .C2(n7038), .ZN(P2_U3293) );
  OAI222_X1 U8474 ( .A1(n8953), .A2(n6658), .B1(n8955), .B2(n6657), .C1(
        P2_U3151), .C2(n6939), .ZN(P2_U3292) );
  OAI222_X1 U8475 ( .A1(n8953), .A2(n6660), .B1(n8955), .B2(n6661), .C1(
        P2_U3151), .C2(n6659), .ZN(P2_U3290) );
  INV_X1 U8476 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6662) );
  INV_X1 U8477 ( .A(n6720), .ZN(n6755) );
  OAI222_X1 U8478 ( .A1(n7825), .A2(n6662), .B1(n9807), .B2(n6661), .C1(
        P1_U3086), .C2(n6755), .ZN(P1_U3350) );
  OAI222_X1 U8479 ( .A1(n7825), .A2(n6663), .B1(n9807), .B2(n6665), .C1(
        P1_U3086), .C2(n6743), .ZN(P1_U3349) );
  OAI222_X1 U8480 ( .A1(n8953), .A2(n6666), .B1(n8955), .B2(n6665), .C1(
        P2_U3151), .C2(n6664), .ZN(P2_U3289) );
  OAI222_X1 U8481 ( .A1(n8953), .A2(n6667), .B1(n8955), .B2(n6668), .C1(
        P2_U3151), .C2(n7329), .ZN(P2_U3288) );
  INV_X1 U8482 ( .A(n6716), .ZN(n6767) );
  OAI222_X1 U8483 ( .A1(n7825), .A2(n6669), .B1(n9807), .B2(n6668), .C1(
        P1_U3086), .C2(n6767), .ZN(P1_U3348) );
  AND2_X1 U8484 ( .A1(n9380), .A2(n6670), .ZN(n9912) );
  NAND2_X1 U8485 ( .A1(n9913), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6671) );
  OAI21_X1 U8486 ( .B1(n9913), .B2(n6672), .A(n6671), .ZN(P1_U3439) );
  NAND2_X1 U8487 ( .A1(n9913), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6673) );
  OAI21_X1 U8488 ( .B1(n9913), .B2(n6674), .A(n6673), .ZN(P1_U3440) );
  INV_X1 U8489 ( .A(n9502), .ZN(n9478) );
  NOR2_X1 U8490 ( .A1(n9478), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8491 ( .A(n7858), .ZN(n6680) );
  AOI21_X1 U8492 ( .B1(n6680), .B2(n7250), .A(n6679), .ZN(n6805) );
  OAI21_X1 U8493 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n6680), .A(n6805), .ZN(
        n6682) );
  XNOR2_X1 U8494 ( .A(n6682), .B(n6681), .ZN(n6686) );
  INV_X1 U8495 ( .A(n6683), .ZN(n6685) );
  AOI22_X1 U8496 ( .A1(n9478), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6684) );
  OAI21_X1 U8497 ( .B1(n6686), .B2(n6685), .A(n6684), .ZN(P1_U3243) );
  INV_X1 U8498 ( .A(n6687), .ZN(n6690) );
  AOI22_X1 U8499 ( .A1(n6842), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9804), .ZN(n6688) );
  OAI21_X1 U8500 ( .B1(n6690), .B2(n9807), .A(n6688), .ZN(P1_U3346) );
  OAI222_X1 U8501 ( .A1(n8955), .A2(n6690), .B1(n7474), .B2(P2_U3151), .C1(
        n6689), .C2(n8953), .ZN(P2_U3286) );
  INV_X1 U8502 ( .A(n6691), .ZN(n6693) );
  OAI222_X1 U8503 ( .A1(n8955), .A2(n6693), .B1(n7557), .B2(P2_U3151), .C1(
        n6692), .C2(n8953), .ZN(P2_U3285) );
  INV_X1 U8504 ( .A(n6909), .ZN(n6914) );
  OAI222_X1 U8505 ( .A1(n7825), .A2(n6694), .B1(n9807), .B2(n6693), .C1(n6914), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8506 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6700) );
  INV_X1 U8507 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8508 ( .A1(n7859), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6697) );
  OR2_X1 U8509 ( .A1(n7862), .A2(n6695), .ZN(n6696) );
  OAI211_X1 U8510 ( .C1(n5738), .C2(n6698), .A(n6697), .B(n6696), .ZN(n9507)
         );
  NAND2_X1 U8511 ( .A1(n9507), .A2(P1_U3973), .ZN(n6699) );
  OAI21_X1 U8512 ( .B1(P1_U3973), .B2(n6700), .A(n6699), .ZN(P1_U3585) );
  INV_X1 U8513 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U8514 ( .A1(n6272), .A2(P1_U3973), .ZN(n6701) );
  OAI21_X1 U8515 ( .B1(P1_U3973), .B2(n6702), .A(n6701), .ZN(P1_U3554) );
  AND2_X1 U8516 ( .A1(n8947), .A2(n6703), .ZN(n6835) );
  NOR2_X1 U8517 ( .A1(n6835), .A2(n6704), .ZN(P2_U3247) );
  INV_X1 U8518 ( .A(n6705), .ZN(n6707) );
  INV_X1 U8519 ( .A(n7149), .ZN(n7142) );
  OAI222_X1 U8520 ( .A1(n7825), .A2(n6706), .B1(n9807), .B2(n6707), .C1(
        P1_U3086), .C2(n7142), .ZN(P1_U3344) );
  OAI222_X1 U8521 ( .A1(n8953), .A2(n6708), .B1(n8955), .B2(n6707), .C1(
        P2_U3151), .C2(n7658), .ZN(P2_U3284) );
  AOI21_X1 U8522 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6723), .A(n6709), .ZN(
        n9424) );
  XNOR2_X1 U8523 ( .A(n9417), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9423) );
  NOR2_X1 U8524 ( .A1(n9424), .A2(n9423), .ZN(n9422) );
  AOI21_X1 U8525 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n9417), .A(n9422), .ZN(
        n6772) );
  XNOR2_X1 U8526 ( .A(n6724), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6771) );
  NOR2_X1 U8527 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  AOI21_X1 U8528 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6724), .A(n6770), .ZN(
        n6808) );
  NAND2_X1 U8529 ( .A1(n6725), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6710) );
  OAI21_X1 U8530 ( .B1(n6725), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6710), .ZN(
        n6807) );
  NOR2_X1 U8531 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  INV_X1 U8532 ( .A(n6710), .ZN(n6711) );
  NOR2_X1 U8533 ( .A1(n6806), .A2(n6711), .ZN(n6748) );
  AOI22_X1 U8534 ( .A1(n6720), .A2(n7259), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n6755), .ZN(n6747) );
  AOI22_X1 U8535 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6743), .B1(n6718), .B2(
        n5131), .ZN(n6736) );
  NAND2_X1 U8536 ( .A1(n6716), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6712) );
  OAI21_X1 U8537 ( .B1(n6716), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6712), .ZN(
        n6759) );
  NOR2_X1 U8538 ( .A1(n6760), .A2(n6759), .ZN(n6758) );
  NAND2_X1 U8539 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6828), .ZN(n6713) );
  OAI21_X1 U8540 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6828), .A(n6713), .ZN(
        n6714) );
  AOI211_X1 U8541 ( .C1(n6715), .C2(n6714), .A(n6827), .B(n9484), .ZN(n6734)
         );
  NAND2_X1 U8542 ( .A1(n6716), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6727) );
  MUX2_X1 U8543 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6717), .S(n6716), .Z(n6762)
         );
  MUX2_X1 U8544 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6719), .S(n6718), .Z(n6739)
         );
  MUX2_X1 U8545 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6721), .S(n6720), .Z(n6750)
         );
  INV_X1 U8546 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6726) );
  AOI21_X1 U8547 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n6723), .A(n6722), .ZN(
        n9421) );
  MUX2_X1 U8548 ( .A(n5022), .B(P1_REG1_REG_2__SCAN_IN), .S(n9417), .Z(n9420)
         );
  NOR2_X1 U8549 ( .A1(n9421), .A2(n9420), .ZN(n9419) );
  INV_X1 U8550 ( .A(n9419), .ZN(n6775) );
  NAND2_X1 U8551 ( .A1(n9417), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6774) );
  MUX2_X1 U8552 ( .A(n5048), .B(P1_REG1_REG_3__SCAN_IN), .S(n6724), .Z(n6773)
         );
  AOI21_X1 U8553 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n6777) );
  AOI21_X1 U8554 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6724), .A(n6777), .ZN(
        n6811) );
  MUX2_X1 U8555 ( .A(n6726), .B(P1_REG1_REG_4__SCAN_IN), .S(n6725), .Z(n6810)
         );
  OR2_X1 U8556 ( .A1(n6811), .A2(n6810), .ZN(n6813) );
  OAI21_X1 U8557 ( .B1(n6726), .B2(n6818), .A(n6813), .ZN(n6751) );
  NAND2_X1 U8558 ( .A1(n6750), .A2(n6751), .ZN(n6749) );
  OAI21_X1 U8559 ( .B1(n6755), .B2(n6721), .A(n6749), .ZN(n6740) );
  NAND2_X1 U8560 ( .A1(n6739), .A2(n6740), .ZN(n6738) );
  OAI21_X1 U8561 ( .B1(n6743), .B2(n6719), .A(n6738), .ZN(n6763) );
  NAND2_X1 U8562 ( .A1(n6762), .A2(n6763), .ZN(n6761) );
  NAND2_X1 U8563 ( .A1(n6727), .A2(n6761), .ZN(n6730) );
  MUX2_X1 U8564 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6728), .S(n6828), .Z(n6729)
         );
  NAND2_X1 U8565 ( .A1(n6729), .A2(n6730), .ZN(n6819) );
  OAI211_X1 U8566 ( .C1(n6730), .C2(n6729), .A(n6819), .B(n9488), .ZN(n6732)
         );
  AND2_X1 U8567 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7596) );
  AOI21_X1 U8568 ( .B1(n9478), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7596), .ZN(
        n6731) );
  OAI211_X1 U8569 ( .C1(n9490), .C2(n6820), .A(n6732), .B(n6731), .ZN(n6733)
         );
  OR2_X1 U8570 ( .A1(n6734), .A2(n6733), .ZN(P1_U3251) );
  AOI211_X1 U8571 ( .C1(n6737), .C2(n6736), .A(n6735), .B(n9484), .ZN(n6745)
         );
  OAI211_X1 U8572 ( .C1(n6740), .C2(n6739), .A(n9488), .B(n6738), .ZN(n6742)
         );
  AND2_X1 U8573 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7272) );
  AOI21_X1 U8574 ( .B1(n9478), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7272), .ZN(
        n6741) );
  OAI211_X1 U8575 ( .C1(n9490), .C2(n6743), .A(n6742), .B(n6741), .ZN(n6744)
         );
  OR2_X1 U8576 ( .A1(n6745), .A2(n6744), .ZN(P1_U3249) );
  AOI211_X1 U8577 ( .C1(n6748), .C2(n6747), .A(n6746), .B(n9484), .ZN(n6757)
         );
  OAI211_X1 U8578 ( .C1(n6751), .C2(n6750), .A(n9488), .B(n6749), .ZN(n6754)
         );
  NAND2_X1 U8579 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7160) );
  INV_X1 U8580 ( .A(n7160), .ZN(n6752) );
  AOI21_X1 U8581 ( .B1(n9478), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6752), .ZN(
        n6753) );
  OAI211_X1 U8582 ( .C1(n9490), .C2(n6755), .A(n6754), .B(n6753), .ZN(n6756)
         );
  OR2_X1 U8583 ( .A1(n6757), .A2(n6756), .ZN(P1_U3248) );
  AOI211_X1 U8584 ( .C1(n6760), .C2(n6759), .A(n6758), .B(n9484), .ZN(n6769)
         );
  OAI211_X1 U8585 ( .C1(n6763), .C2(n6762), .A(n9488), .B(n6761), .ZN(n6766)
         );
  INV_X1 U8586 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6764) );
  NOR2_X1 U8587 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6764), .ZN(n7297) );
  AOI21_X1 U8588 ( .B1(n9478), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7297), .ZN(
        n6765) );
  OAI211_X1 U8589 ( .C1(n9490), .C2(n6767), .A(n6766), .B(n6765), .ZN(n6768)
         );
  OR2_X1 U8590 ( .A1(n6769), .A2(n6768), .ZN(P1_U3250) );
  AOI211_X1 U8591 ( .C1(n6772), .C2(n6771), .A(n6770), .B(n9484), .ZN(n6779)
         );
  AND3_X1 U8592 ( .A1(n6775), .A2(n6774), .A3(n6773), .ZN(n6776) );
  NOR3_X1 U8593 ( .A1(n9491), .A2(n6777), .A3(n6776), .ZN(n6778) );
  NOR2_X1 U8594 ( .A1(n6779), .A2(n6778), .ZN(n6781) );
  AND2_X1 U8595 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6957) );
  AOI21_X1 U8596 ( .B1(n9478), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6957), .ZN(
        n6780) );
  OAI211_X1 U8597 ( .C1(n6782), .C2(n9490), .A(n6781), .B(n6780), .ZN(P1_U3246) );
  INV_X1 U8598 ( .A(n6783), .ZN(n6785) );
  INV_X1 U8599 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6784) );
  OAI222_X1 U8600 ( .A1(n8955), .A2(n6785), .B1(n7745), .B2(P2_U3151), .C1(
        n6784), .C2(n8953), .ZN(P2_U3283) );
  INV_X1 U8601 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6786) );
  INV_X1 U8602 ( .A(n7170), .ZN(n7174) );
  OAI222_X1 U8603 ( .A1(n7825), .A2(n6786), .B1(P1_U3086), .B2(n7174), .C1(
        n6785), .C2(n9807), .ZN(P1_U3343) );
  INV_X1 U8604 ( .A(n9113), .ZN(n9122) );
  XNOR2_X1 U8605 ( .A(n6788), .B(n6787), .ZN(n6800) );
  INV_X1 U8606 ( .A(n9115), .ZN(n9132) );
  INV_X1 U8607 ( .A(n6789), .ZN(n6791) );
  NOR2_X1 U8608 ( .A1(n6791), .A2(n6790), .ZN(n6869) );
  OAI22_X1 U8609 ( .A1(n6869), .A2(n6792), .B1(n9135), .B2(n7252), .ZN(n6793)
         );
  AOI21_X1 U8610 ( .B1(n9132), .B2(n9413), .A(n6793), .ZN(n6794) );
  OAI21_X1 U8611 ( .B1(n9122), .B2(n6800), .A(n6794), .ZN(P1_U3232) );
  INV_X1 U8612 ( .A(n6835), .ZN(n6795) );
  AND2_X1 U8613 ( .A1(n6795), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8614 ( .A1(n6795), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8615 ( .A1(n6795), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8616 ( .A1(n6795), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8617 ( .A1(n6795), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8618 ( .A1(n6795), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8619 ( .A1(n6795), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8620 ( .A1(n6795), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8621 ( .A1(n6795), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8622 ( .A1(n6795), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8623 ( .A1(n6795), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8624 ( .A1(n6795), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8625 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6797) );
  INV_X1 U8626 ( .A(n6796), .ZN(n6798) );
  INV_X1 U8627 ( .A(n7403), .ZN(n7396) );
  OAI222_X1 U8628 ( .A1(n7825), .A2(n6797), .B1(n9807), .B2(n6798), .C1(
        P1_U3086), .C2(n7396), .ZN(P1_U3342) );
  OAI222_X1 U8629 ( .A1(n8953), .A2(n6799), .B1(n8955), .B2(n6798), .C1(
        P2_U3151), .C2(n7790), .ZN(P2_U3282) );
  NAND3_X1 U8630 ( .A1(n6800), .A2(n7858), .A3(n7828), .ZN(n6804) );
  INV_X1 U8631 ( .A(n6801), .ZN(n6802) );
  AOI21_X1 U8632 ( .B1(n9379), .B2(n6802), .A(n9412), .ZN(n6803) );
  OAI211_X1 U8633 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6805), .A(n6804), .B(n6803), .ZN(n9429) );
  AND2_X1 U8634 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7078) );
  AOI21_X1 U8635 ( .B1(n6808), .B2(n6807), .A(n6806), .ZN(n6809) );
  INV_X1 U8636 ( .A(n6809), .ZN(n6815) );
  NAND2_X1 U8637 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  NAND3_X1 U8638 ( .A1(n9488), .A2(n6813), .A3(n6812), .ZN(n6814) );
  OAI21_X1 U8639 ( .B1(n9484), .B2(n6815), .A(n6814), .ZN(n6816) );
  AOI211_X1 U8640 ( .C1(n9478), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n7078), .B(
        n6816), .ZN(n6817) );
  OAI211_X1 U8641 ( .C1(n9490), .C2(n6818), .A(n9429), .B(n6817), .ZN(P1_U3247) );
  INV_X1 U8642 ( .A(n9490), .ZN(n9418) );
  OAI21_X1 U8643 ( .B1(n6820), .B2(n6728), .A(n6819), .ZN(n6823) );
  MUX2_X1 U8644 ( .A(n6821), .B(P1_REG1_REG_9__SCAN_IN), .S(n6842), .Z(n6822)
         );
  NOR2_X1 U8645 ( .A1(n6822), .A2(n6823), .ZN(n6843) );
  AOI21_X1 U8646 ( .B1(n6823), .B2(n6822), .A(n6843), .ZN(n6826) );
  NOR2_X1 U8647 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6824), .ZN(n7704) );
  AOI21_X1 U8648 ( .B1(n9478), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7704), .ZN(
        n6825) );
  OAI21_X1 U8649 ( .B1(n9491), .B2(n6826), .A(n6825), .ZN(n6833) );
  NOR2_X1 U8650 ( .A1(n6842), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6829) );
  AOI21_X1 U8651 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6842), .A(n6829), .ZN(
        n6830) );
  AOI221_X1 U8652 ( .B1(n6831), .B2(n6839), .C1(n6830), .C2(n6839), .A(n9484), 
        .ZN(n6832) );
  AOI211_X1 U8653 ( .C1(n9418), .C2(n6842), .A(n6833), .B(n6832), .ZN(n6834)
         );
  INV_X1 U8654 ( .A(n6834), .ZN(P1_U3252) );
  INV_X1 U8655 ( .A(n6836), .ZN(n6837) );
  AOI22_X1 U8656 ( .A1(n6795), .A2(n6206), .B1(n6899), .B2(n6837), .ZN(
        P2_U3376) );
  NAND2_X1 U8657 ( .A1(n6909), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8658 ( .B1(n6909), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6838), .ZN(
        n6841) );
  AOI211_X1 U8659 ( .C1(n6841), .C2(n6840), .A(n6908), .B(n9484), .ZN(n6851)
         );
  NOR2_X1 U8660 ( .A1(n6842), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U8661 ( .A1(n6844), .A2(n6843), .ZN(n6847) );
  MUX2_X1 U8662 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6845), .S(n6909), .Z(n6846)
         );
  NAND2_X1 U8663 ( .A1(n6846), .A2(n6847), .ZN(n6913) );
  OAI211_X1 U8664 ( .C1(n6847), .C2(n6846), .A(n6913), .B(n9488), .ZN(n6849)
         );
  AND2_X1 U8665 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8992) );
  AOI21_X1 U8666 ( .B1(n9478), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n8992), .ZN(
        n6848) );
  OAI211_X1 U8667 ( .C1(n9490), .C2(n6914), .A(n6849), .B(n6848), .ZN(n6850)
         );
  OR2_X1 U8668 ( .A1(n6851), .A2(n6850), .ZN(P1_U3253) );
  INV_X1 U8669 ( .A(n6853), .ZN(n6854) );
  AOI21_X1 U8670 ( .B1(n6855), .B2(n6852), .A(n6854), .ZN(n6860) );
  INV_X1 U8671 ( .A(n9126), .ZN(n9105) );
  NOR2_X1 U8672 ( .A1(n9115), .A2(n9202), .ZN(n6858) );
  OAI22_X1 U8673 ( .A1(n6869), .A2(n6856), .B1(n9205), .B2(n9135), .ZN(n6857)
         );
  AOI211_X1 U8674 ( .C1(n9105), .C2(n6272), .A(n6858), .B(n6857), .ZN(n6859)
         );
  OAI21_X1 U8675 ( .B1(n6860), .B2(n9122), .A(n6859), .ZN(P1_U3222) );
  AND2_X1 U8676 ( .A1(n6795), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8677 ( .A1(n6795), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8678 ( .A1(n6795), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8679 ( .A1(n6795), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8680 ( .A1(n6795), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8681 ( .A1(n6795), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8682 ( .A1(n6795), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8683 ( .A1(n6795), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8684 ( .A1(n6795), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8685 ( .A1(n6795), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8686 ( .A1(n6795), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8687 ( .A1(n6795), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8688 ( .A1(n6795), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8689 ( .A1(n6795), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8690 ( .A1(n6795), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8691 ( .A1(n6795), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8692 ( .A1(n6795), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  INV_X1 U8693 ( .A(n6861), .ZN(n6863) );
  OAI222_X1 U8694 ( .A1(n7825), .A2(n6862), .B1(n9807), .B2(n6863), .C1(
        P1_U3086), .C2(n7681), .ZN(P1_U3341) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6864) );
  OAI222_X1 U8696 ( .A1(n8953), .A2(n6864), .B1(n8955), .B2(n6863), .C1(
        P2_U3151), .C2(n8402), .ZN(P2_U3281) );
  INV_X1 U8697 ( .A(n6866), .ZN(n6867) );
  NAND3_X1 U8698 ( .A1(n6867), .A2(n6853), .A3(n5020), .ZN(n6868) );
  AOI21_X1 U8699 ( .B1(n6865), .B2(n6868), .A(n9122), .ZN(n6873) );
  OAI22_X1 U8700 ( .A1(n6869), .A2(n9414), .B1(n9917), .B2(n9135), .ZN(n6872)
         );
  INV_X1 U8701 ( .A(n9878), .ZN(n6870) );
  OAI22_X1 U8702 ( .A1(n6902), .A2(n9126), .B1(n9115), .B2(n6870), .ZN(n6871)
         );
  OR3_X1 U8703 ( .A1(n6873), .A2(n6872), .A3(n6871), .ZN(P1_U3237) );
  INV_X1 U8704 ( .A(n6874), .ZN(n6876) );
  OAI222_X1 U8705 ( .A1(n7825), .A2(n6875), .B1(n9807), .B2(n6876), .C1(
        P1_U3086), .C2(n9437), .ZN(P1_U3340) );
  INV_X1 U8706 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6877) );
  INV_X1 U8707 ( .A(n8426), .ZN(n8407) );
  OAI222_X1 U8708 ( .A1(n8953), .A2(n6877), .B1(n8955), .B2(n6876), .C1(
        P2_U3151), .C2(n8407), .ZN(P2_U3280) );
  NAND2_X1 U8709 ( .A1(n8392), .A2(n7054), .ZN(n8035) );
  INV_X1 U8710 ( .A(n8035), .ZN(n6878) );
  OR2_X1 U8711 ( .A1(n6878), .A2(n8037), .ZN(n8008) );
  INV_X1 U8712 ( .A(n8008), .ZN(n7025) );
  INV_X1 U8713 ( .A(n6894), .ZN(n6879) );
  NAND2_X1 U8714 ( .A1(n6981), .A2(n6879), .ZN(n6883) );
  INV_X1 U8715 ( .A(n6880), .ZN(n6881) );
  NAND2_X1 U8716 ( .A1(n6886), .A2(n6881), .ZN(n6882) );
  NAND2_X1 U8717 ( .A1(n6883), .A2(n6882), .ZN(n8344) );
  INV_X1 U8718 ( .A(n6978), .ZN(n6884) );
  NOR2_X1 U8719 ( .A1(n6884), .A2(n6979), .ZN(n6885) );
  NAND2_X1 U8720 ( .A1(n6981), .A2(n6885), .ZN(n8359) );
  INV_X1 U8721 ( .A(n8359), .ZN(n8371) );
  NAND2_X1 U8722 ( .A1(n6886), .A2(n7382), .ZN(n6888) );
  NAND2_X1 U8723 ( .A1(n6887), .A2(n8947), .ZN(n8782) );
  NAND2_X1 U8724 ( .A1(n6888), .A2(n8782), .ZN(n8362) );
  AOI22_X1 U8725 ( .A1(n8371), .A2(n8390), .B1(n8362), .B2(n7029), .ZN(n6901)
         );
  INV_X1 U8726 ( .A(n6889), .ZN(n6893) );
  NAND2_X1 U8727 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  OAI211_X1 U8728 ( .C1(n6896), .C2(n6894), .A(n6893), .B(n6892), .ZN(n6895)
         );
  NAND2_X1 U8729 ( .A1(n6895), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6898) );
  INV_X1 U8730 ( .A(n6979), .ZN(n7024) );
  NAND2_X1 U8731 ( .A1(n7024), .A2(n8947), .ZN(n8196) );
  OR2_X1 U8732 ( .A1(n6896), .A2(n8196), .ZN(n6897) );
  AND2_X1 U8733 ( .A1(n6898), .A2(n6897), .ZN(n7113) );
  NAND2_X1 U8734 ( .A1(n7113), .A2(n6899), .ZN(n7090) );
  NAND2_X1 U8735 ( .A1(n7090), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6900) );
  OAI211_X1 U8736 ( .C1(n7025), .C2(n8366), .A(n6901), .B(n6900), .ZN(P2_U3172) );
  NOR2_X1 U8737 ( .A1(n6902), .A2(n9835), .ZN(n7248) );
  AND2_X1 U8738 ( .A1(n6272), .A2(n7252), .ZN(n9199) );
  NOR2_X1 U8739 ( .A1(n6946), .A2(n9199), .ZN(n9149) );
  AOI21_X1 U8740 ( .B1(n9963), .B2(n9842), .A(n9149), .ZN(n6903) );
  AOI211_X1 U8741 ( .C1(n6943), .C2(n7246), .A(n7248), .B(n6903), .ZN(n6963)
         );
  INV_X1 U8742 ( .A(n6904), .ZN(n7222) );
  NOR2_X1 U8743 ( .A1(n7220), .A2(n7222), .ZN(n6906) );
  AND2_X2 U8744 ( .A1(n6906), .A2(n6905), .ZN(n10019) );
  NAND2_X1 U8745 ( .A1(n10017), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6907) );
  OAI21_X1 U8746 ( .B1(n6963), .B2(n10017), .A(n6907), .ZN(P1_U3522) );
  NAND2_X1 U8747 ( .A1(n7149), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6910) );
  OAI21_X1 U8748 ( .B1(n7149), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6910), .ZN(
        n6911) );
  AOI211_X1 U8749 ( .C1(n6912), .C2(n6911), .A(n7148), .B(n9484), .ZN(n6922)
         );
  OAI21_X1 U8750 ( .B1(n6914), .B2(n6845), .A(n6913), .ZN(n6917) );
  MUX2_X1 U8751 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6915), .S(n7149), .Z(n6916)
         );
  NAND2_X1 U8752 ( .A1(n6916), .A2(n6917), .ZN(n7141) );
  OAI211_X1 U8753 ( .C1(n6917), .C2(n6916), .A(n9488), .B(n7141), .ZN(n6920)
         );
  INV_X1 U8754 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U8755 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6918), .ZN(n9094) );
  AOI21_X1 U8756 ( .B1(n9478), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9094), .ZN(
        n6919) );
  OAI211_X1 U8757 ( .C1(n9490), .C2(n7142), .A(n6920), .B(n6919), .ZN(n6921)
         );
  OR2_X1 U8758 ( .A1(n6922), .A2(n6921), .ZN(P1_U3254) );
  OAI21_X1 U8759 ( .B1(n4419), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7125), .ZN(
        n6932) );
  INV_X1 U8760 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8761 ( .A1(n8505), .A2(n6923), .ZN(n6931) );
  INV_X1 U8762 ( .A(n6924), .ZN(n6925) );
  AOI21_X1 U8763 ( .B1(n6927), .B2(n6926), .A(n6925), .ZN(n6929) );
  OAI22_X1 U8764 ( .A1(n8484), .A2(n6929), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6928), .ZN(n6930) );
  AOI211_X1 U8765 ( .C1(n8514), .C2(n6932), .A(n6931), .B(n6930), .ZN(n6938)
         );
  OAI21_X1 U8766 ( .B1(n6935), .B2(n6934), .A(n6933), .ZN(n6936) );
  INV_X1 U8767 ( .A(n8517), .ZN(n8474) );
  NAND2_X1 U8768 ( .A1(n6936), .A2(n8474), .ZN(n6937) );
  OAI211_X1 U8769 ( .C1(n8506), .C2(n6939), .A(n6938), .B(n6937), .ZN(P2_U3185) );
  INV_X1 U8770 ( .A(n6940), .ZN(n9981) );
  XNOR2_X1 U8771 ( .A(n6941), .B(n6942), .ZN(n9898) );
  INV_X1 U8772 ( .A(n7227), .ZN(n6945) );
  AOI21_X1 U8773 ( .B1(n6943), .B2(n9900), .A(n9670), .ZN(n6944) );
  NAND2_X1 U8774 ( .A1(n6945), .A2(n6944), .ZN(n9905) );
  OAI21_X1 U8775 ( .B1(n9205), .B2(n9996), .A(n9905), .ZN(n6951) );
  INV_X1 U8776 ( .A(n7579), .ZN(n9847) );
  XNOR2_X1 U8777 ( .A(n6941), .B(n6946), .ZN(n6948) );
  AOI22_X1 U8778 ( .A1(n9879), .A2(n9411), .B1(n6272), .B2(n9877), .ZN(n6947)
         );
  OAI21_X1 U8779 ( .B1(n6948), .B2(n9842), .A(n6947), .ZN(n6949) );
  AOI21_X1 U8780 ( .B1(n9847), .B2(n9898), .A(n6949), .ZN(n9909) );
  INV_X1 U8781 ( .A(n9909), .ZN(n6950) );
  AOI211_X1 U8782 ( .C1(n9981), .C2(n9898), .A(n6951), .B(n6950), .ZN(n9914)
         );
  NAND2_X1 U8783 ( .A1(n10017), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6952) );
  OAI21_X1 U8784 ( .B1(n9914), .B2(n10017), .A(n6952), .ZN(P1_U3523) );
  OAI21_X1 U8785 ( .B1(n6956), .B2(n6953), .A(n6955), .ZN(n6961) );
  AOI22_X1 U8786 ( .A1(n9105), .A2(n9411), .B1(n9132), .B2(n9410), .ZN(n6959)
         );
  AOI21_X1 U8787 ( .B1(n9082), .B2(n7240), .A(n6957), .ZN(n6958) );
  OAI211_X1 U8788 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9129), .A(n6959), .B(
        n6958), .ZN(n6960) );
  AOI21_X1 U8789 ( .B1(n6961), .B2(n9113), .A(n6960), .ZN(n6962) );
  INV_X1 U8790 ( .A(n6962), .ZN(P1_U3218) );
  INV_X1 U8791 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6965) );
  OR2_X1 U8792 ( .A1(n6963), .A2(n10002), .ZN(n6964) );
  OAI21_X1 U8793 ( .B1(n10004), .B2(n6965), .A(n6964), .ZN(P1_U3453) );
  NAND2_X1 U8794 ( .A1(n9412), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6966) );
  OAI21_X1 U8795 ( .B1(n9530), .B2(n9412), .A(n6966), .ZN(P1_U3583) );
  INV_X1 U8796 ( .A(n6967), .ZN(n6969) );
  OAI222_X1 U8797 ( .A1(n7825), .A2(n6968), .B1(n9807), .B2(n6969), .C1(
        P1_U3086), .C2(n9449), .ZN(P1_U3339) );
  INV_X1 U8798 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6970) );
  INV_X1 U8799 ( .A(n8433), .ZN(n8449) );
  OAI222_X1 U8800 ( .A1(n8953), .A2(n6970), .B1(n8955), .B2(n6969), .C1(
        P2_U3151), .C2(n8449), .ZN(P2_U3279) );
  INV_X1 U8801 ( .A(n6971), .ZN(n6972) );
  NAND2_X1 U8802 ( .A1(n7017), .A2(n6972), .ZN(n6975) );
  NAND2_X1 U8803 ( .A1(n8033), .A2(n8190), .ZN(n6973) );
  AOI21_X1 U8804 ( .B1(n7936), .B2(n7054), .A(n8037), .ZN(n7086) );
  XOR2_X1 U8805 ( .A(n7085), .B(n7086), .Z(n6985) );
  INV_X1 U8806 ( .A(n6977), .ZN(n7165) );
  NOR2_X1 U8807 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  AOI22_X1 U8808 ( .A1(n8371), .A2(n8389), .B1(n8347), .B2(n8392), .ZN(n6982)
         );
  OAI21_X1 U8809 ( .B1(n7165), .B2(n8378), .A(n6982), .ZN(n6983) );
  AOI21_X1 U8810 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7090), .A(n6983), .ZN(
        n6984) );
  OAI21_X1 U8811 ( .B1(n6985), .B2(n8366), .A(n6984), .ZN(P2_U3162) );
  INV_X1 U8812 ( .A(n8505), .ZN(n8488) );
  NOR2_X1 U8813 ( .A1(n8474), .A2(n6986), .ZN(n6990) );
  AOI21_X1 U8814 ( .B1(n6993), .B2(n6987), .A(n6995), .ZN(n6989) );
  INV_X1 U8815 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6988) );
  OAI22_X1 U8816 ( .A1(n6990), .A2(n6989), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6988), .ZN(n6991) );
  AOI21_X1 U8817 ( .B1(n8488), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6991), .ZN(
        n6992) );
  OAI21_X1 U8818 ( .B1(n6993), .B2(n8506), .A(n6992), .ZN(P2_U3182) );
  NAND2_X1 U8819 ( .A1(n9412), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6994) );
  OAI21_X1 U8820 ( .B1(n7866), .B2(n9412), .A(n6994), .ZN(P1_U3582) );
  XNOR2_X1 U8821 ( .A(n6996), .B(n6995), .ZN(n7014) );
  INV_X1 U8822 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U8823 ( .A1(n6998), .A2(n6997), .ZN(n6999) );
  NAND2_X1 U8824 ( .A1(n7000), .A2(n6999), .ZN(n7001) );
  NAND2_X1 U8825 ( .A1(n8509), .A2(n7001), .ZN(n7008) );
  NAND2_X1 U8826 ( .A1(n7003), .A2(n7002), .ZN(n7004) );
  NAND2_X1 U8827 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  NAND2_X1 U8828 ( .A1(n8514), .A2(n7006), .ZN(n7007) );
  OAI211_X1 U8829 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7009), .A(n7008), .B(n7007), .ZN(n7012) );
  NOR2_X1 U8830 ( .A1(n8506), .A2(n7010), .ZN(n7011) );
  AOI211_X1 U8831 ( .C1(n8488), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7012), .B(
        n7011), .ZN(n7013) );
  OAI21_X1 U8832 ( .B1(n8517), .B2(n7014), .A(n7013), .ZN(P2_U3183) );
  NAND2_X1 U8833 ( .A1(n7015), .A2(n7019), .ZN(n7023) );
  INV_X1 U8834 ( .A(n7016), .ZN(n7022) );
  NAND2_X1 U8835 ( .A1(n7017), .A2(n7018), .ZN(n7021) );
  OR2_X1 U8836 ( .A1(n7019), .A2(n7018), .ZN(n7020) );
  NAND4_X1 U8837 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n7028)
         );
  INV_X2 U8838 ( .A(n8739), .ZN(n10038) );
  NOR3_X1 U8839 ( .A1(n7025), .A2(n7024), .A3(n7382), .ZN(n7027) );
  NAND2_X1 U8840 ( .A1(n8390), .A2(n8760), .ZN(n7053) );
  INV_X1 U8841 ( .A(n7053), .ZN(n7026) );
  OAI21_X1 U8842 ( .B1(n7027), .B2(n7026), .A(n10038), .ZN(n7031) );
  OR2_X1 U8843 ( .A1(n7028), .A2(n8736), .ZN(n8715) );
  AOI22_X1 U8844 ( .A1(n10031), .A2(n7029), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10033), .ZN(n7030) );
  OAI211_X1 U8845 ( .C1(n4439), .C2(n10038), .A(n7031), .B(n7030), .ZN(
        P2_U3233) );
  INV_X1 U8846 ( .A(n7032), .ZN(n7034) );
  INV_X1 U8847 ( .A(n9463), .ZN(n9470) );
  OAI222_X1 U8848 ( .A1(n7825), .A2(n7033), .B1(n9807), .B2(n7034), .C1(
        P1_U3086), .C2(n9470), .ZN(P1_U3338) );
  INV_X1 U8849 ( .A(n8468), .ZN(n8451) );
  OAI222_X1 U8850 ( .A1(n8953), .A2(n7035), .B1(n8955), .B2(n7034), .C1(
        P2_U3151), .C2(n8451), .ZN(P2_U3278) );
  XNOR2_X1 U8851 ( .A(n7037), .B(n7036), .ZN(n7052) );
  INV_X1 U8852 ( .A(n8506), .ZN(n8476) );
  OAI21_X1 U8853 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(n7042) );
  AOI22_X1 U8854 ( .A1(n8509), .A2(n7042), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7049) );
  NAND2_X1 U8855 ( .A1(n8488), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n7048) );
  OAI21_X1 U8856 ( .B1(n7045), .B2(n7044), .A(n7043), .ZN(n7046) );
  NAND2_X1 U8857 ( .A1(n8514), .A2(n7046), .ZN(n7047) );
  NAND3_X1 U8858 ( .A1(n7049), .A2(n7048), .A3(n7047), .ZN(n7050) );
  AOI21_X1 U8859 ( .B1(n4434), .B2(n8476), .A(n7050), .ZN(n7051) );
  OAI21_X1 U8860 ( .B1(n8517), .B2(n7052), .A(n7051), .ZN(P2_U3184) );
  INV_X1 U8861 ( .A(n10062), .ZN(n10043) );
  OR2_X1 U8862 ( .A1(n7757), .A2(n10043), .ZN(n8834) );
  INV_X1 U8863 ( .A(n8834), .ZN(n10074) );
  INV_X1 U8864 ( .A(n8755), .ZN(n8775) );
  NAND2_X1 U8865 ( .A1(n10074), .A2(n8775), .ZN(n7056) );
  OAI21_X1 U8866 ( .B1(n10072), .B2(n7054), .A(n7053), .ZN(n7055) );
  AOI21_X1 U8867 ( .B1(n8008), .B2(n7056), .A(n7055), .ZN(n7060) );
  MUX2_X1 U8868 ( .A(n7060), .B(n4438), .S(n10090), .Z(n7057) );
  INV_X1 U8869 ( .A(n7057), .ZN(P2_U3459) );
  INV_X1 U8870 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7058) );
  OR2_X1 U8871 ( .A1(n10078), .A2(n7058), .ZN(n7059) );
  OAI21_X1 U8872 ( .B1(n7060), .B2(n10080), .A(n7059), .ZN(P2_U3390) );
  XNOR2_X1 U8873 ( .A(n7062), .B(n7061), .ZN(n7073) );
  INV_X1 U8874 ( .A(n7192), .ZN(n7063) );
  AOI21_X1 U8875 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(n7066) );
  NAND2_X1 U8876 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7442) );
  OAI21_X1 U8877 ( .B1(n8484), .B2(n7066), .A(n7442), .ZN(n7070) );
  NAND2_X1 U8878 ( .A1(n7067), .A2(n10083), .ZN(n7068) );
  AOI21_X1 U8879 ( .B1(n7187), .B2(n7068), .A(n8491), .ZN(n7069) );
  AOI211_X1 U8880 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n8488), .A(n7070), .B(
        n7069), .ZN(n7072) );
  NAND2_X1 U8881 ( .A1(n8476), .A2(n4831), .ZN(n7071) );
  OAI211_X1 U8882 ( .C1(n7073), .C2(n8517), .A(n7072), .B(n7071), .ZN(P2_U3187) );
  INV_X1 U8883 ( .A(n7075), .ZN(n7076) );
  AOI211_X1 U8884 ( .C1(n7077), .C2(n7074), .A(n9122), .B(n7076), .ZN(n7083)
         );
  AOI22_X1 U8885 ( .A1(n9105), .A2(n9878), .B1(n9132), .B2(n9880), .ZN(n7081)
         );
  AOI21_X1 U8886 ( .B1(n9082), .B2(n7079), .A(n7078), .ZN(n7080) );
  OAI211_X1 U8887 ( .C1(n9881), .C2(n9129), .A(n7081), .B(n7080), .ZN(n7082)
         );
  OR2_X1 U8888 ( .A1(n7083), .A2(n7082), .ZN(P1_U3230) );
  XNOR2_X1 U8889 ( .A(n7383), .B(n7438), .ZN(n7106) );
  XNOR2_X1 U8890 ( .A(n7106), .B(n8389), .ZN(n7107) );
  OAI22_X1 U8891 ( .A1(n7086), .A2(n7085), .B1(n7084), .B2(n8390), .ZN(n7108)
         );
  XOR2_X1 U8892 ( .A(n7107), .B(n7108), .Z(n7092) );
  AOI22_X1 U8893 ( .A1(n8371), .A2(n8388), .B1(n8347), .B2(n8390), .ZN(n7087)
         );
  OAI21_X1 U8894 ( .B1(n7088), .B2(n8378), .A(n7087), .ZN(n7089) );
  AOI21_X1 U8895 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7090), .A(n7089), .ZN(
        n7091) );
  OAI21_X1 U8896 ( .B1(n7092), .B2(n8366), .A(n7091), .ZN(P2_U3177) );
  INV_X1 U8897 ( .A(n8037), .ZN(n7093) );
  NAND2_X1 U8898 ( .A1(n7093), .A2(n7097), .ZN(n7094) );
  NAND2_X1 U8899 ( .A1(n7095), .A2(n7094), .ZN(n7834) );
  XNOR2_X1 U8900 ( .A(n7097), .B(n7096), .ZN(n7098) );
  NAND2_X1 U8901 ( .A1(n7098), .A2(n8755), .ZN(n7100) );
  AOI22_X1 U8902 ( .A1(n8761), .A2(n8392), .B1(n8389), .B2(n8760), .ZN(n7099)
         );
  NAND2_X1 U8903 ( .A1(n7100), .A2(n7099), .ZN(n7833) );
  AOI21_X1 U8904 ( .B1(n8834), .B2(n7834), .A(n7833), .ZN(n7167) );
  INV_X1 U8905 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7101) );
  OAI22_X1 U8906 ( .A1(n7165), .A2(n8934), .B1(n10078), .B2(n7101), .ZN(n7102)
         );
  INV_X1 U8907 ( .A(n7102), .ZN(n7103) );
  OAI21_X1 U8908 ( .B1(n7167), .B2(n10080), .A(n7103), .ZN(P2_U3393) );
  INV_X1 U8909 ( .A(n9486), .ZN(n9481) );
  INV_X1 U8910 ( .A(n7104), .ZN(n7139) );
  OAI222_X1 U8911 ( .A1(P1_U3086), .A2(n9481), .B1(n9807), .B2(n7139), .C1(
        n7105), .C2(n7825), .ZN(P1_U3337) );
  INV_X1 U8912 ( .A(n8389), .ZN(n7111) );
  AOI22_X1 U8913 ( .A1(n7108), .A2(n7107), .B1(n7111), .B2(n7106), .ZN(n7110)
         );
  XNOR2_X1 U8914 ( .A(n7212), .B(n7438), .ZN(n7280) );
  XNOR2_X1 U8915 ( .A(n7280), .B(n8388), .ZN(n7109) );
  OAI211_X1 U8916 ( .C1(n7110), .C2(n7109), .A(n7279), .B(n8344), .ZN(n7117)
         );
  INV_X1 U8917 ( .A(n8347), .ZN(n8373) );
  INV_X1 U8918 ( .A(n8387), .ZN(n7441) );
  OAI22_X1 U8919 ( .A1(n8373), .A2(n7111), .B1(n7441), .B2(n8359), .ZN(n7115)
         );
  OR2_X1 U8920 ( .A1(n7112), .A2(P2_U3151), .ZN(n8200) );
  MUX2_X1 U8921 ( .A(n8375), .B(P2_U3151), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7114) );
  AOI211_X1 U8922 ( .C1(n7212), .C2(n8362), .A(n7115), .B(n7114), .ZN(n7116)
         );
  NAND2_X1 U8923 ( .A1(n7117), .A2(n7116), .ZN(P2_U3158) );
  INV_X1 U8924 ( .A(n7118), .ZN(n7137) );
  INV_X1 U8925 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7497) );
  OAI21_X1 U8926 ( .B1(n7121), .B2(n7120), .A(n7119), .ZN(n7130) );
  NAND2_X1 U8927 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7283) );
  INV_X1 U8928 ( .A(n7283), .ZN(n7129) );
  INV_X1 U8929 ( .A(n7122), .ZN(n7124) );
  NAND3_X1 U8930 ( .A1(n7125), .A2(n7124), .A3(n7123), .ZN(n7126) );
  AOI21_X1 U8931 ( .B1(n7127), .B2(n7126), .A(n8491), .ZN(n7128) );
  AOI211_X1 U8932 ( .C1(n8509), .C2(n7130), .A(n7129), .B(n7128), .ZN(n7131)
         );
  OAI21_X1 U8933 ( .B1(n7497), .B2(n8505), .A(n7131), .ZN(n7136) );
  AOI211_X1 U8934 ( .C1(n7134), .C2(n7133), .A(n8517), .B(n7132), .ZN(n7135)
         );
  AOI211_X1 U8935 ( .C1(n8476), .C2(n7137), .A(n7136), .B(n7135), .ZN(n7138)
         );
  INV_X1 U8936 ( .A(n7138), .ZN(P2_U3186) );
  INV_X1 U8937 ( .A(n8496), .ZN(n8464) );
  OAI222_X1 U8938 ( .A1(n8953), .A2(n7140), .B1(n8464), .B2(P2_U3151), .C1(
        n8955), .C2(n7139), .ZN(P2_U3277) );
  OAI21_X1 U8939 ( .B1(n7142), .B2(n6915), .A(n7141), .ZN(n7145) );
  MUX2_X1 U8940 ( .A(n7143), .B(P1_REG1_REG_12__SCAN_IN), .S(n7170), .Z(n7144)
         );
  NOR2_X1 U8941 ( .A1(n7145), .A2(n7144), .ZN(n7173) );
  AOI21_X1 U8942 ( .B1(n7145), .B2(n7144), .A(n7173), .ZN(n7147) );
  AND2_X1 U8943 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9021) );
  AOI21_X1 U8944 ( .B1(n9478), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9021), .ZN(
        n7146) );
  OAI21_X1 U8945 ( .B1(n9491), .B2(n7147), .A(n7146), .ZN(n7154) );
  NOR2_X1 U8946 ( .A1(n7170), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7150) );
  AOI21_X1 U8947 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7170), .A(n7150), .ZN(
        n7151) );
  AOI221_X1 U8948 ( .B1(n7152), .B2(n7169), .C1(n7151), .C2(n7169), .A(n9484), 
        .ZN(n7153) );
  AOI211_X1 U8949 ( .C1(n9418), .C2(n7170), .A(n7154), .B(n7153), .ZN(n7155)
         );
  INV_X1 U8950 ( .A(n7155), .ZN(P1_U3255) );
  NAND2_X1 U8951 ( .A1(n7157), .A2(n7156), .ZN(n7159) );
  XNOR2_X1 U8952 ( .A(n7159), .B(n7158), .ZN(n7164) );
  INV_X1 U8953 ( .A(n9410), .ZN(n7256) );
  OAI21_X1 U8954 ( .B1(n9126), .B2(n7256), .A(n7160), .ZN(n7162) );
  OAI22_X1 U8955 ( .A1(n9129), .A2(n7258), .B1(n7254), .B2(n9115), .ZN(n7161)
         );
  AOI211_X1 U8956 ( .C1(n7261), .C2(n9082), .A(n7162), .B(n7161), .ZN(n7163)
         );
  OAI21_X1 U8957 ( .B1(n7164), .B2(n9122), .A(n7163), .ZN(P1_U3227) );
  AOI22_X1 U8958 ( .A1(n8845), .A2(n6977), .B1(n10090), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7166) );
  OAI21_X1 U8959 ( .B1(n7167), .B2(n10090), .A(n7166), .ZN(P2_U3460) );
  NAND2_X1 U8960 ( .A1(n7403), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7168) );
  OAI21_X1 U8961 ( .B1(n7403), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7168), .ZN(
        n7172) );
  AOI211_X1 U8962 ( .C1(n7172), .C2(n7171), .A(n7402), .B(n9484), .ZN(n7181)
         );
  AOI21_X1 U8963 ( .B1(n7174), .B2(n7143), .A(n7173), .ZN(n7177) );
  MUX2_X1 U8964 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7175), .S(n7403), .Z(n7176)
         );
  NAND2_X1 U8965 ( .A1(n7176), .A2(n7177), .ZN(n7395) );
  OAI211_X1 U8966 ( .C1(n7177), .C2(n7176), .A(n9488), .B(n7395), .ZN(n7179)
         );
  AND2_X1 U8967 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9070) );
  AOI21_X1 U8968 ( .B1(n9478), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9070), .ZN(
        n7178) );
  OAI211_X1 U8969 ( .C1(n9490), .C2(n7396), .A(n7179), .B(n7178), .ZN(n7180)
         );
  OR2_X1 U8970 ( .A1(n7181), .A2(n7180), .ZN(P1_U3256) );
  AOI21_X1 U8971 ( .B1(n7183), .B2(n7182), .A(n7321), .ZN(n7202) );
  INV_X1 U8972 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7501) );
  INV_X1 U8973 ( .A(n7184), .ZN(n7186) );
  NAND3_X1 U8974 ( .A1(n7187), .A2(n7186), .A3(n7185), .ZN(n7188) );
  AOI21_X1 U8975 ( .B1(n7189), .B2(n7188), .A(n8491), .ZN(n7197) );
  INV_X1 U8976 ( .A(n7190), .ZN(n7191) );
  NAND3_X1 U8977 ( .A1(n7192), .A2(n7191), .A3(n4828), .ZN(n7193) );
  AOI21_X1 U8978 ( .B1(n7194), .B2(n7193), .A(n8484), .ZN(n7196) );
  INV_X1 U8979 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7195) );
  NOR2_X1 U8980 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7195), .ZN(n7634) );
  NOR3_X1 U8981 ( .A1(n7197), .A2(n7196), .A3(n7634), .ZN(n7198) );
  OAI21_X1 U8982 ( .B1(n7501), .B2(n8505), .A(n7198), .ZN(n7199) );
  AOI21_X1 U8983 ( .B1(n7200), .B2(n8476), .A(n7199), .ZN(n7201) );
  OAI21_X1 U8984 ( .B1(n7202), .B2(n8517), .A(n7201), .ZN(P2_U3188) );
  INV_X1 U8985 ( .A(n8041), .ZN(n8004) );
  NAND2_X1 U8986 ( .A1(n7378), .A2(n8004), .ZN(n7380) );
  NAND2_X1 U8987 ( .A1(n7380), .A2(n8045), .ZN(n7203) );
  INV_X1 U8988 ( .A(n7204), .ZN(n8005) );
  NAND2_X1 U8989 ( .A1(n7203), .A2(n8005), .ZN(n7335) );
  OAI21_X1 U8990 ( .B1(n7203), .B2(n8005), .A(n7335), .ZN(n7350) );
  XNOR2_X1 U8991 ( .A(n7205), .B(n7204), .ZN(n7206) );
  NAND2_X1 U8992 ( .A1(n7206), .A2(n8755), .ZN(n7208) );
  AOI22_X1 U8993 ( .A1(n8761), .A2(n8389), .B1(n8387), .B2(n8760), .ZN(n7207)
         );
  NAND2_X1 U8994 ( .A1(n7208), .A2(n7207), .ZN(n7347) );
  AOI21_X1 U8995 ( .B1(n8834), .B2(n7350), .A(n7347), .ZN(n7214) );
  INV_X1 U8996 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7209) );
  OAI22_X1 U8997 ( .A1(n7346), .A2(n8934), .B1(n10078), .B2(n7209), .ZN(n7210)
         );
  INV_X1 U8998 ( .A(n7210), .ZN(n7211) );
  OAI21_X1 U8999 ( .B1(n7214), .B2(n10080), .A(n7211), .ZN(P2_U3399) );
  AOI22_X1 U9000 ( .A1(n8845), .A2(n7212), .B1(n10090), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7213) );
  OAI21_X1 U9001 ( .B1(n7214), .B2(n10090), .A(n7213), .ZN(P2_U3462) );
  XNOR2_X1 U9002 ( .A(n7215), .B(n9147), .ZN(n9919) );
  XNOR2_X1 U9003 ( .A(n7216), .B(n7217), .ZN(n7218) );
  AOI222_X1 U9004 ( .A1(n9876), .A2(n7218), .B1(n9413), .B2(n9877), .C1(n9878), 
        .C2(n9879), .ZN(n9916) );
  OAI21_X1 U9005 ( .B1(n9414), .B2(n9710), .A(n9916), .ZN(n7219) );
  AOI21_X1 U9006 ( .B1(n9847), .B2(n9919), .A(n7219), .ZN(n7232) );
  INV_X1 U9007 ( .A(n7220), .ZN(n7224) );
  AND2_X1 U9008 ( .A1(n7222), .A2(n7221), .ZN(n7223) );
  NAND2_X1 U9009 ( .A1(n7224), .A2(n7223), .ZN(n7225) );
  NAND2_X2 U9010 ( .A1(n7225), .A2(n9710), .ZN(n9713) );
  OR2_X1 U9011 ( .A1(n4321), .A2(n7237), .ZN(n7589) );
  INV_X1 U9012 ( .A(n7589), .ZN(n9899) );
  INV_X1 U9013 ( .A(n7239), .ZN(n7226) );
  INV_X1 U9014 ( .A(n9670), .ZN(n9890) );
  OAI211_X1 U9015 ( .C1(n9917), .C2(n7227), .A(n7226), .B(n9890), .ZN(n9915)
         );
  AOI22_X1 U9016 ( .A1(n9901), .A2(n9201), .B1(n4321), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n7229) );
  OAI21_X1 U9017 ( .B1(n9904), .B2(n9915), .A(n7229), .ZN(n7230) );
  AOI21_X1 U9018 ( .B1(n9899), .B2(n9919), .A(n7230), .ZN(n7231) );
  OAI21_X1 U9019 ( .B1(n7232), .B2(n4321), .A(n7231), .ZN(P1_U3291) );
  INV_X1 U9020 ( .A(n7235), .ZN(n9148) );
  XNOR2_X1 U9021 ( .A(n7233), .B(n9148), .ZN(n7234) );
  AOI222_X1 U9022 ( .A1(n9410), .A2(n9879), .B1(n9411), .B2(n9877), .C1(n9876), 
        .C2(n7234), .ZN(n9922) );
  XNOR2_X1 U9023 ( .A(n7236), .B(n7235), .ZN(n9925) );
  AND2_X1 U9024 ( .A1(n7579), .A2(n7237), .ZN(n7238) );
  INV_X1 U9025 ( .A(n9709), .ZN(n9894) );
  OAI211_X1 U9026 ( .C1(n7239), .C2(n9921), .A(n9890), .B(n9888), .ZN(n9920)
         );
  NAND2_X1 U9027 ( .A1(n9901), .A2(n7240), .ZN(n7243) );
  AOI22_X1 U9028 ( .A1(n4321), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9897), .B2(
        n7241), .ZN(n7242) );
  OAI211_X1 U9029 ( .C1(n9920), .C2(n9904), .A(n7243), .B(n7242), .ZN(n7244)
         );
  AOI21_X1 U9030 ( .B1(n9925), .B2(n9894), .A(n7244), .ZN(n7245) );
  OAI21_X1 U9031 ( .B1(n9922), .B2(n4321), .A(n7245), .ZN(P1_U3290) );
  AOI21_X1 U9032 ( .B1(n9893), .B2(n9890), .A(n9901), .ZN(n7253) );
  NOR3_X1 U9033 ( .A1(n9149), .A2(n7246), .A3(n9381), .ZN(n7247) );
  AOI211_X1 U9034 ( .C1(n9897), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7248), .B(
        n7247), .ZN(n7249) );
  MUX2_X1 U9035 ( .A(n7250), .B(n7249), .S(n9713), .Z(n7251) );
  OAI21_X1 U9036 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(P1_U3293) );
  XNOR2_X1 U9037 ( .A(n9252), .B(n9151), .ZN(n7255) );
  OAI222_X1 U9038 ( .A1(n9833), .A2(n7256), .B1(n7255), .B2(n9842), .C1(n9835), 
        .C2(n7254), .ZN(n9934) );
  INV_X1 U9039 ( .A(n9934), .ZN(n7265) );
  XNOR2_X1 U9040 ( .A(n7257), .B(n9151), .ZN(n9936) );
  OAI211_X1 U9041 ( .C1(n9889), .C2(n9933), .A(n9868), .B(n9890), .ZN(n9932)
         );
  OAI22_X1 U9042 ( .A1(n9713), .A2(n7259), .B1(n7258), .B2(n9710), .ZN(n7260)
         );
  AOI21_X1 U9043 ( .B1(n9901), .B2(n7261), .A(n7260), .ZN(n7262) );
  OAI21_X1 U9044 ( .B1(n9932), .B2(n9904), .A(n7262), .ZN(n7263) );
  AOI21_X1 U9045 ( .B1(n9936), .B2(n9894), .A(n7263), .ZN(n7264) );
  OAI21_X1 U9046 ( .B1(n7265), .B2(n4321), .A(n7264), .ZN(P1_U3288) );
  NAND2_X1 U9047 ( .A1(n7268), .A2(n7267), .ZN(n7269) );
  XNOR2_X1 U9048 ( .A(n7266), .B(n7269), .ZN(n7270) );
  NAND2_X1 U9049 ( .A1(n7270), .A2(n9113), .ZN(n7274) );
  OAI22_X1 U9050 ( .A1(n9129), .A2(n9862), .B1(n9834), .B2(n9115), .ZN(n7271)
         );
  AOI211_X1 U9051 ( .C1(n9105), .C2(n9880), .A(n7272), .B(n7271), .ZN(n7273)
         );
  OAI211_X1 U9052 ( .C1(n9939), .C2(n9135), .A(n7274), .B(n7273), .ZN(P1_U3239) );
  INV_X1 U9053 ( .A(n7275), .ZN(n7277) );
  OAI222_X1 U9054 ( .A1(n8953), .A2(n7276), .B1(n8955), .B2(n7277), .C1(n6174), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9055 ( .A1(n7825), .A2(n7278), .B1(n9807), .B2(n7277), .C1(
        P1_U3086), .C2(n9384), .ZN(P1_U3336) );
  XNOR2_X1 U9056 ( .A(n7438), .B(n7875), .ZN(n7439) );
  XNOR2_X1 U9057 ( .A(n7439), .B(n8387), .ZN(n7282) );
  INV_X1 U9058 ( .A(n8388), .ZN(n7341) );
  AOI21_X1 U9059 ( .B1(n7282), .B2(n7281), .A(n4414), .ZN(n7288) );
  OAI21_X1 U9060 ( .B1(n8373), .B2(n7341), .A(n7283), .ZN(n7284) );
  AOI21_X1 U9061 ( .B1(n8371), .B2(n8386), .A(n7284), .ZN(n7285) );
  OAI21_X1 U9062 ( .B1(n7875), .B2(n8378), .A(n7285), .ZN(n7286) );
  AOI21_X1 U9063 ( .B1(n10034), .B2(n8375), .A(n7286), .ZN(n7287) );
  OAI21_X1 U9064 ( .B1(n7288), .B2(n8366), .A(n7287), .ZN(P2_U3170) );
  NAND2_X1 U9065 ( .A1(n8391), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7289) );
  OAI21_X1 U9066 ( .B1(n7993), .B2(n8391), .A(n7289), .ZN(P2_U3521) );
  NAND2_X1 U9067 ( .A1(n8391), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7290) );
  OAI21_X1 U9068 ( .B1(n8538), .B2(n8391), .A(n7290), .ZN(P2_U3520) );
  XOR2_X1 U9069 ( .A(n7293), .B(n7292), .Z(n7294) );
  XNOR2_X1 U9070 ( .A(n7291), .B(n7294), .ZN(n7300) );
  OAI22_X1 U9071 ( .A1(n9129), .A2(n7311), .B1(n7295), .B2(n9115), .ZN(n7296)
         );
  AOI211_X1 U9072 ( .C1(n9105), .C2(n9409), .A(n7297), .B(n7296), .ZN(n7299)
         );
  NAND2_X1 U9073 ( .A1(n9082), .A2(n9945), .ZN(n7298) );
  OAI211_X1 U9074 ( .C1(n7300), .C2(n9122), .A(n7299), .B(n7298), .ZN(P1_U3213) );
  XNOR2_X1 U9075 ( .A(n7301), .B(n7303), .ZN(n9946) );
  INV_X1 U9076 ( .A(n9946), .ZN(n7318) );
  NAND2_X1 U9077 ( .A1(n9859), .A2(n9257), .ZN(n7304) );
  NAND2_X1 U9078 ( .A1(n7304), .A2(n9254), .ZN(n7302) );
  NAND2_X1 U9079 ( .A1(n7302), .A2(n4682), .ZN(n9840) );
  NAND3_X1 U9080 ( .A1(n7304), .A2(n9254), .A3(n7303), .ZN(n7305) );
  AOI21_X1 U9081 ( .B1(n9840), .B2(n7305), .A(n9842), .ZN(n7310) );
  AND2_X1 U9082 ( .A1(n9946), .A2(n9847), .ZN(n7309) );
  NAND2_X1 U9083 ( .A1(n9408), .A2(n9879), .ZN(n7307) );
  NAND2_X1 U9084 ( .A1(n9409), .A2(n9877), .ZN(n7306) );
  NAND2_X1 U9085 ( .A1(n7307), .A2(n7306), .ZN(n7308) );
  OR3_X1 U9086 ( .A1(n7310), .A2(n7309), .A3(n7308), .ZN(n9951) );
  NAND2_X1 U9087 ( .A1(n9951), .A2(n9713), .ZN(n7317) );
  OAI22_X1 U9088 ( .A1(n9713), .A2(n7312), .B1(n7311), .B2(n9710), .ZN(n7315)
         );
  AOI21_X1 U9089 ( .B1(n9869), .B2(n9945), .A(n9670), .ZN(n7313) );
  NAND2_X1 U9090 ( .A1(n7313), .A2(n9852), .ZN(n9947) );
  NOR2_X1 U9091 ( .A1(n9947), .A2(n9904), .ZN(n7314) );
  AOI211_X1 U9092 ( .C1(n9901), .C2(n9945), .A(n7315), .B(n7314), .ZN(n7316)
         );
  OAI211_X1 U9093 ( .C1(n7318), .C2(n7589), .A(n7317), .B(n7316), .ZN(P1_U3286) );
  OR3_X1 U9094 ( .A1(n7321), .A2(n7320), .A3(n7319), .ZN(n7322) );
  AOI21_X1 U9095 ( .B1(n7363), .B2(n7322), .A(n8517), .ZN(n7333) );
  INV_X1 U9096 ( .A(n7369), .ZN(n7323) );
  AOI21_X1 U9097 ( .B1(n6528), .B2(n7324), .A(n7323), .ZN(n7326) );
  NAND2_X1 U9098 ( .A1(n8488), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U9099 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7669) );
  OAI211_X1 U9100 ( .C1(n8491), .C2(n7326), .A(n7325), .B(n7669), .ZN(n7332)
         );
  INV_X1 U9101 ( .A(n7359), .ZN(n7327) );
  AOI21_X1 U9102 ( .B1(n6529), .B2(n7328), .A(n7327), .ZN(n7330) );
  OAI22_X1 U9103 ( .A1(n7330), .A2(n8484), .B1(n8506), .B2(n7329), .ZN(n7331)
         );
  OR3_X1 U9104 ( .A1(n7333), .A2(n7332), .A3(n7331), .ZN(P2_U3189) );
  NAND3_X1 U9105 ( .A1(n7335), .A2(n7334), .A3(n8052), .ZN(n7337) );
  NAND2_X1 U9106 ( .A1(n7336), .A2(n8050), .ZN(n7413) );
  NAND2_X1 U9107 ( .A1(n7337), .A2(n7413), .ZN(n10028) );
  INV_X1 U9108 ( .A(n8386), .ZN(n7342) );
  NAND2_X1 U9109 ( .A1(n7416), .A2(n7338), .ZN(n7339) );
  XNOR2_X1 U9110 ( .A(n7339), .B(n8050), .ZN(n7340) );
  OAI222_X1 U9111 ( .A1(n8780), .A2(n7342), .B1(n8778), .B2(n7341), .C1(n8775), 
        .C2(n7340), .ZN(n10027) );
  AOI21_X1 U9112 ( .B1(n8834), .B2(n10028), .A(n10027), .ZN(n7872) );
  INV_X1 U9113 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7343) );
  OAI22_X1 U9114 ( .A1(n7875), .A2(n8934), .B1(n10078), .B2(n7343), .ZN(n7344)
         );
  INV_X1 U9115 ( .A(n7344), .ZN(n7345) );
  OAI21_X1 U9116 ( .B1(n7872), .B2(n10080), .A(n7345), .ZN(P2_U3402) );
  AND2_X1 U9117 ( .A1(n7384), .A2(n8033), .ZN(n7381) );
  OR2_X1 U9118 ( .A1(n7757), .A2(n7381), .ZN(n10029) );
  OAI22_X1 U9119 ( .A1(n8715), .A2(n7346), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8782), .ZN(n7349) );
  MUX2_X1 U9120 ( .A(n7347), .B(P2_REG2_REG_3__SCAN_IN), .S(n8739), .Z(n7348)
         );
  AOI211_X1 U9121 ( .C1(n8717), .C2(n7350), .A(n7349), .B(n7348), .ZN(n7351)
         );
  INV_X1 U9122 ( .A(n7351), .ZN(P2_U3230) );
  INV_X1 U9123 ( .A(n7352), .ZN(n7393) );
  OAI222_X1 U9124 ( .A1(n8955), .A2(n7393), .B1(P2_U3151), .B2(n8190), .C1(
        n7353), .C2(n8953), .ZN(P2_U3275) );
  INV_X1 U9125 ( .A(n7354), .ZN(n7356) );
  NOR2_X1 U9126 ( .A1(n7356), .A2(n7355), .ZN(n7360) );
  INV_X1 U9127 ( .A(n7357), .ZN(n7358) );
  AOI21_X1 U9128 ( .B1(n7360), .B2(n7359), .A(n7358), .ZN(n7377) );
  AND3_X1 U9129 ( .A1(n7363), .A2(n7362), .A3(n7361), .ZN(n7364) );
  OAI21_X1 U9130 ( .B1(n7468), .B2(n7364), .A(n8474), .ZN(n7376) );
  INV_X1 U9131 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7506) );
  NOR2_X1 U9132 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4429), .ZN(n7713) );
  INV_X1 U9133 ( .A(n7713), .ZN(n7365) );
  OAI21_X1 U9134 ( .B1(n8505), .B2(n7506), .A(n7365), .ZN(n7373) );
  INV_X1 U9135 ( .A(n7366), .ZN(n7368) );
  NAND3_X1 U9136 ( .A1(n7369), .A2(n7368), .A3(n7367), .ZN(n7370) );
  AOI21_X1 U9137 ( .B1(n7371), .B2(n7370), .A(n8491), .ZN(n7372) );
  AOI211_X1 U9138 ( .C1(n8476), .C2(n7374), .A(n7373), .B(n7372), .ZN(n7375)
         );
  OAI211_X1 U9139 ( .C1(n7377), .C2(n8484), .A(n7376), .B(n7375), .ZN(P2_U3190) );
  OR2_X1 U9140 ( .A1(n7378), .A2(n8004), .ZN(n7379) );
  NAND2_X1 U9141 ( .A1(n7380), .A2(n7379), .ZN(n10042) );
  INV_X1 U9142 ( .A(n10042), .ZN(n7392) );
  NAND2_X1 U9143 ( .A1(n10038), .A2(n7381), .ZN(n8533) );
  NAND2_X1 U9144 ( .A1(n7383), .A2(n7382), .ZN(n10039) );
  NOR2_X1 U9145 ( .A1(n10039), .A2(n7384), .ZN(n7389) );
  XNOR2_X1 U9146 ( .A(n7385), .B(n8004), .ZN(n7388) );
  NAND2_X1 U9147 ( .A1(n10042), .A2(n7757), .ZN(n7387) );
  AOI22_X1 U9148 ( .A1(n8761), .A2(n8390), .B1(n8388), .B2(n8760), .ZN(n7386)
         );
  OAI211_X1 U9149 ( .C1(n8775), .C2(n7388), .A(n7387), .B(n7386), .ZN(n10040)
         );
  AOI211_X1 U9150 ( .C1(n10033), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7389), .B(
        n10040), .ZN(n7390) );
  MUX2_X1 U9151 ( .A(n6597), .B(n7390), .S(n10038), .Z(n7391) );
  OAI21_X1 U9152 ( .B1(n7392), .B2(n8533), .A(n7391), .ZN(P2_U3231) );
  OAI222_X1 U9153 ( .A1(n7825), .A2(n7394), .B1(n9807), .B2(n7393), .C1(n9197), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U9154 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7401) );
  OAI21_X1 U9155 ( .B1(n7396), .B2(n7175), .A(n7395), .ZN(n7399) );
  MUX2_X1 U9156 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7397), .S(n7678), .Z(n7398)
         );
  NAND2_X1 U9157 ( .A1(n7398), .A2(n7399), .ZN(n7680) );
  OAI211_X1 U9158 ( .C1(n7399), .C2(n7398), .A(n9488), .B(n7680), .ZN(n7400)
         );
  NAND2_X1 U9159 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8964) );
  OAI211_X1 U9160 ( .C1(n9502), .C2(n7401), .A(n7400), .B(n8964), .ZN(n7408)
         );
  NAND2_X1 U9161 ( .A1(n7678), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7404) );
  OAI21_X1 U9162 ( .B1(n7678), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7404), .ZN(
        n7405) );
  AOI211_X1 U9163 ( .C1(n7406), .C2(n7405), .A(n7677), .B(n9484), .ZN(n7407)
         );
  AOI211_X1 U9164 ( .C1(n9418), .C2(n7678), .A(n7408), .B(n7407), .ZN(n7409)
         );
  INV_X1 U9165 ( .A(n7409), .ZN(P1_U3257) );
  INV_X1 U9166 ( .A(n7410), .ZN(n7436) );
  OAI222_X1 U9167 ( .A1(n8955), .A2(n7436), .B1(P2_U3151), .B2(n8036), .C1(
        n7411), .C2(n8953), .ZN(P2_U3274) );
  NAND2_X1 U9168 ( .A1(n7413), .A2(n7412), .ZN(n7414) );
  NAND2_X1 U9169 ( .A1(n8055), .A2(n8062), .ZN(n8007) );
  XNOR2_X1 U9170 ( .A(n7414), .B(n8007), .ZN(n10047) );
  NAND2_X1 U9171 ( .A1(n7416), .A2(n7415), .ZN(n7418) );
  AND2_X1 U9172 ( .A1(n7418), .A2(n7417), .ZN(n7419) );
  XNOR2_X1 U9173 ( .A(n7419), .B(n8007), .ZN(n7420) );
  AOI222_X1 U9174 ( .A1(n8755), .A2(n7420), .B1(n8385), .B2(n8760), .C1(n8387), 
        .C2(n8761), .ZN(n10045) );
  MUX2_X1 U9175 ( .A(n7065), .B(n10045), .S(n10038), .Z(n7423) );
  AOI22_X1 U9176 ( .A1(n10031), .A2(n7421), .B1(n10033), .B2(n7448), .ZN(n7422) );
  OAI211_X1 U9177 ( .C1(n8789), .C2(n10047), .A(n7423), .B(n7422), .ZN(
        P2_U3228) );
  XNOR2_X1 U9178 ( .A(n7424), .B(n4409), .ZN(n9964) );
  NAND2_X1 U9179 ( .A1(n9840), .A2(n9262), .ZN(n9837) );
  NAND2_X1 U9180 ( .A1(n9837), .A2(n9843), .ZN(n7425) );
  XNOR2_X1 U9181 ( .A(n7425), .B(n4409), .ZN(n7427) );
  AND2_X1 U9182 ( .A1(n9408), .A2(n9877), .ZN(n7426) );
  AOI21_X1 U9183 ( .B1(n7427), .B2(n9876), .A(n7426), .ZN(n9967) );
  OAI21_X1 U9184 ( .B1(n7702), .B2(n9710), .A(n9967), .ZN(n7428) );
  NAND2_X1 U9185 ( .A1(n7428), .A2(n9713), .ZN(n7435) );
  XNOR2_X1 U9186 ( .A(n9853), .B(n9960), .ZN(n7429) );
  NAND2_X1 U9187 ( .A1(n7429), .A2(n9890), .ZN(n7431) );
  NAND2_X1 U9188 ( .A1(n9406), .A2(n9879), .ZN(n7430) );
  NAND2_X1 U9189 ( .A1(n7431), .A2(n7430), .ZN(n9962) );
  OAI22_X1 U9190 ( .A1(n7707), .A2(n9884), .B1(n9713), .B2(n7432), .ZN(n7433)
         );
  AOI21_X1 U9191 ( .B1(n9962), .B2(n9893), .A(n7433), .ZN(n7434) );
  OAI211_X1 U9192 ( .C1(n9964), .C2(n9709), .A(n7435), .B(n7434), .ZN(P1_U3284) );
  OAI222_X1 U9193 ( .A1(n7825), .A2(n7437), .B1(n9807), .B2(n7436), .C1(n9204), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U9194 ( .A(n7940), .B(n10046), .ZN(n7638) );
  XNOR2_X1 U9195 ( .A(n7638), .B(n8386), .ZN(n7639) );
  INV_X1 U9196 ( .A(n7439), .ZN(n7440) );
  XOR2_X1 U9197 ( .A(n7639), .B(n7640), .Z(n7450) );
  INV_X1 U9198 ( .A(n7442), .ZN(n7445) );
  NOR2_X1 U9199 ( .A1(n8359), .A2(n7443), .ZN(n7444) );
  AOI211_X1 U9200 ( .C1(n8347), .C2(n8387), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OAI21_X1 U9201 ( .B1(n10046), .B2(n8378), .A(n7446), .ZN(n7447) );
  AOI21_X1 U9202 ( .B1(n7448), .B2(n8375), .A(n7447), .ZN(n7449) );
  OAI21_X1 U9203 ( .B1(n7450), .B2(n8366), .A(n7449), .ZN(P2_U3167) );
  XNOR2_X1 U9204 ( .A(n7451), .B(n9145), .ZN(n9973) );
  INV_X1 U9205 ( .A(n9973), .ZN(n7463) );
  INV_X1 U9206 ( .A(n7452), .ZN(n7574) );
  AOI21_X1 U9207 ( .B1(n9145), .B2(n7453), .A(n7574), .ZN(n7454) );
  OAI222_X1 U9208 ( .A1(n9833), .A2(n9836), .B1(n9835), .B2(n8989), .C1(n9842), 
        .C2(n7454), .ZN(n9971) );
  INV_X1 U9209 ( .A(n7455), .ZN(n7456) );
  OAI211_X1 U9210 ( .C1(n7456), .C2(n9970), .A(n9890), .B(n7581), .ZN(n9969)
         );
  OAI22_X1 U9211 ( .A1(n9713), .A2(n7457), .B1(n8990), .B2(n9710), .ZN(n7458)
         );
  AOI21_X1 U9212 ( .B1(n9901), .B2(n7459), .A(n7458), .ZN(n7460) );
  OAI21_X1 U9213 ( .B1(n9969), .B2(n9904), .A(n7460), .ZN(n7461) );
  AOI21_X1 U9214 ( .B1(n9971), .B2(n9713), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9215 ( .B1(n7463), .B2(n9709), .A(n7462), .ZN(P1_U3283) );
  AOI21_X1 U9216 ( .B1(n7465), .B2(n7762), .A(n7464), .ZN(n7479) );
  INV_X1 U9217 ( .A(n7541), .ZN(n7470) );
  NOR3_X1 U9218 ( .A1(n7468), .A2(n7467), .A3(n7466), .ZN(n7469) );
  OAI21_X1 U9219 ( .B1(n7470), .B2(n7469), .A(n8474), .ZN(n7478) );
  AOI21_X1 U9220 ( .B1(n7472), .B2(n6537), .A(n7471), .ZN(n7473) );
  NOR2_X1 U9221 ( .A1(n7473), .A2(n8491), .ZN(n7476) );
  AND2_X1 U9222 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7771) );
  INV_X1 U9223 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7510) );
  OAI22_X1 U9224 ( .A1(n8506), .A2(n7474), .B1(n7510), .B2(n8505), .ZN(n7475)
         );
  NOR3_X1 U9225 ( .A1(n7476), .A2(n7771), .A3(n7475), .ZN(n7477) );
  OAI211_X1 U9226 ( .C1(n7479), .C2(n8484), .A(n7478), .B(n7477), .ZN(P2_U3191) );
  INV_X1 U9227 ( .A(n7480), .ZN(n8010) );
  XNOR2_X1 U9228 ( .A(n7481), .B(n8010), .ZN(n10052) );
  XNOR2_X1 U9229 ( .A(n7482), .B(n8010), .ZN(n7483) );
  NAND2_X1 U9230 ( .A1(n7483), .A2(n8755), .ZN(n7485) );
  AOI22_X1 U9231 ( .A1(n8761), .A2(n8386), .B1(n8384), .B2(n8760), .ZN(n7484)
         );
  NAND2_X1 U9232 ( .A1(n7485), .A2(n7484), .ZN(n10054) );
  MUX2_X1 U9233 ( .A(n10054), .B(P2_REG2_REG_6__SCAN_IN), .S(n8739), .Z(n7486)
         );
  INV_X1 U9234 ( .A(n7486), .ZN(n7488) );
  AOI22_X1 U9235 ( .A1(n10031), .A2(n7635), .B1(n10033), .B2(n7645), .ZN(n7487) );
  OAI211_X1 U9236 ( .C1(n10052), .C2(n8789), .A(n7488), .B(n7487), .ZN(
        P2_U3227) );
  NOR2_X1 U9237 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7535) );
  INV_X1 U9238 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7532) );
  INV_X1 U9239 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8436) );
  INV_X1 U9240 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7530) );
  INV_X1 U9241 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8406) );
  NOR2_X1 U9242 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7528) );
  NOR2_X1 U9243 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7525) );
  NOR2_X1 U9244 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7522) );
  NOR2_X1 U9245 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7519) );
  NOR2_X1 U9246 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7516) );
  NOR2_X1 U9247 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7513) );
  NOR2_X1 U9248 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7509) );
  NOR2_X1 U9249 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7505) );
  NOR2_X1 U9250 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7503) );
  NOR2_X1 U9251 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7499) );
  NAND2_X1 U9252 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7494) );
  XOR2_X1 U9253 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10129) );
  NAND2_X1 U9254 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7492) );
  AOI21_X1 U9255 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10094) );
  NAND2_X1 U9256 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7489) );
  NOR2_X1 U9257 ( .A1(n6640), .A2(n7489), .ZN(n10093) );
  NOR2_X1 U9258 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10093), .ZN(n7490) );
  NOR2_X1 U9259 ( .A1(n10094), .A2(n7490), .ZN(n10127) );
  XOR2_X1 U9260 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10126) );
  NAND2_X1 U9261 ( .A1(n10127), .A2(n10126), .ZN(n7491) );
  NAND2_X1 U9262 ( .A1(n7492), .A2(n7491), .ZN(n10128) );
  NAND2_X1 U9263 ( .A1(n10129), .A2(n10128), .ZN(n7493) );
  NAND2_X1 U9264 ( .A1(n7494), .A2(n7493), .ZN(n10131) );
  AOI22_X1 U9265 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n7496), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n7497), .ZN(n10130) );
  NOR2_X1 U9266 ( .A1(n10131), .A2(n10130), .ZN(n7495) );
  AOI21_X1 U9267 ( .B1(n7497), .B2(n7496), .A(n7495), .ZN(n10117) );
  XNOR2_X1 U9268 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10116) );
  NOR2_X1 U9269 ( .A1(n10117), .A2(n10116), .ZN(n7498) );
  NOR2_X1 U9270 ( .A1(n7499), .A2(n7498), .ZN(n10125) );
  INV_X1 U9271 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7500) );
  AOI22_X1 U9272 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7501), .B1(
        P2_ADDR_REG_6__SCAN_IN), .B2(n7500), .ZN(n10124) );
  NOR2_X1 U9273 ( .A1(n10125), .A2(n10124), .ZN(n7502) );
  NOR2_X1 U9274 ( .A1(n7503), .A2(n7502), .ZN(n10121) );
  XNOR2_X1 U9275 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10120) );
  NOR2_X1 U9276 ( .A1(n10121), .A2(n10120), .ZN(n7504) );
  NOR2_X1 U9277 ( .A1(n7505), .A2(n7504), .ZN(n10123) );
  INV_X1 U9278 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7507) );
  AOI22_X1 U9279 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n7507), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n7506), .ZN(n10122) );
  NOR2_X1 U9280 ( .A1(n10123), .A2(n10122), .ZN(n7508) );
  NOR2_X1 U9281 ( .A1(n7509), .A2(n7508), .ZN(n10119) );
  INV_X1 U9282 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7511) );
  AOI22_X1 U9283 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7511), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7510), .ZN(n10118) );
  NOR2_X1 U9284 ( .A1(n10119), .A2(n10118), .ZN(n7512) );
  NOR2_X1 U9285 ( .A1(n7513), .A2(n7512), .ZN(n10115) );
  INV_X1 U9286 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7514) );
  INV_X1 U9287 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7551) );
  AOI22_X1 U9288 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7514), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7551), .ZN(n10114) );
  NOR2_X1 U9289 ( .A1(n10115), .A2(n10114), .ZN(n7515) );
  NOR2_X1 U9290 ( .A1(n7516), .A2(n7515), .ZN(n10113) );
  INV_X1 U9291 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7517) );
  INV_X1 U9292 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7657) );
  AOI22_X1 U9293 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7517), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7657), .ZN(n10112) );
  NOR2_X1 U9294 ( .A1(n10113), .A2(n10112), .ZN(n7518) );
  NOR2_X1 U9295 ( .A1(n7519), .A2(n7518), .ZN(n10111) );
  INV_X1 U9296 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7520) );
  INV_X1 U9297 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7744) );
  AOI22_X1 U9298 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7520), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7744), .ZN(n10110) );
  NOR2_X1 U9299 ( .A1(n10111), .A2(n10110), .ZN(n7521) );
  NOR2_X1 U9300 ( .A1(n7522), .A2(n7521), .ZN(n10109) );
  INV_X1 U9301 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7523) );
  INV_X1 U9302 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7789) );
  AOI22_X1 U9303 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7523), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n7789), .ZN(n10108) );
  NOR2_X1 U9304 ( .A1(n10109), .A2(n10108), .ZN(n7524) );
  NOR2_X1 U9305 ( .A1(n7525), .A2(n7524), .ZN(n10107) );
  AOI22_X1 U9306 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7401), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n7526), .ZN(n10106) );
  NOR2_X1 U9307 ( .A1(n10107), .A2(n10106), .ZN(n7527) );
  NOR2_X1 U9308 ( .A1(n7528), .A2(n7527), .ZN(n10105) );
  AOI22_X1 U9309 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n8406), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(n7530), .ZN(n10104) );
  NOR2_X1 U9310 ( .A1(n10105), .A2(n10104), .ZN(n7529) );
  AOI21_X1 U9311 ( .B1(n7530), .B2(n8406), .A(n7529), .ZN(n10103) );
  AOI22_X1 U9312 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n8436), .B1(
        P2_ADDR_REG_16__SCAN_IN), .B2(n7532), .ZN(n10102) );
  NOR2_X1 U9313 ( .A1(n10103), .A2(n10102), .ZN(n7531) );
  AOI21_X1 U9314 ( .B1(n7532), .B2(n8436), .A(n7531), .ZN(n10101) );
  INV_X1 U9315 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7533) );
  AOI22_X1 U9316 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7533), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8448), .ZN(n10100) );
  NOR2_X1 U9317 ( .A1(n10101), .A2(n10100), .ZN(n7534) );
  NOR2_X1 U9318 ( .A1(n7535), .A2(n7534), .ZN(n10097) );
  NAND2_X1 U9319 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10097), .ZN(n7536) );
  INV_X1 U9320 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10098) );
  NOR2_X1 U9321 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10097), .ZN(n10096) );
  AOI21_X1 U9322 ( .B1(n7536), .B2(n10098), .A(n10096), .ZN(n7538) );
  XNOR2_X1 U9323 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7537) );
  XNOR2_X1 U9324 ( .A(n7538), .B(n7537), .ZN(ADD_1068_U4) );
  AND3_X1 U9325 ( .A1(n7541), .A2(n7540), .A3(n7539), .ZN(n7542) );
  OAI21_X1 U9326 ( .B1(n7651), .B2(n7542), .A(n8474), .ZN(n7556) );
  AOI21_X1 U9327 ( .B1(n4415), .B2(n7544), .A(n7543), .ZN(n7545) );
  NOR2_X1 U9328 ( .A1(n8491), .A2(n7545), .ZN(n7554) );
  AOI21_X1 U9329 ( .B1(n7548), .B2(n7547), .A(n7546), .ZN(n7549) );
  NOR2_X1 U9330 ( .A1(n8484), .A2(n7549), .ZN(n7553) );
  INV_X1 U9331 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7550) );
  NOR2_X1 U9332 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7550), .ZN(n8233) );
  NOR2_X1 U9333 ( .A1(n8505), .A2(n7551), .ZN(n7552) );
  NOR4_X1 U9334 ( .A1(n7554), .A2(n7553), .A3(n8233), .A4(n7552), .ZN(n7555)
         );
  OAI211_X1 U9335 ( .C1(n8506), .C2(n7557), .A(n7556), .B(n7555), .ZN(P2_U3192) );
  INV_X1 U9336 ( .A(n7558), .ZN(n7560) );
  OAI21_X1 U9337 ( .B1(n7560), .B2(n4580), .A(n7559), .ZN(n10021) );
  OAI211_X1 U9338 ( .C1(n7562), .C2(n8069), .A(n7561), .B(n8755), .ZN(n7564)
         );
  AOI22_X1 U9339 ( .A1(n8761), .A2(n8385), .B1(n8383), .B2(n8760), .ZN(n7563)
         );
  AND2_X1 U9340 ( .A1(n7564), .A2(n7563), .ZN(n10020) );
  OAI21_X1 U9341 ( .B1(n10074), .B2(n10021), .A(n10020), .ZN(n7569) );
  OAI22_X1 U9342 ( .A1(n8838), .A2(n8073), .B1(n10092), .B2(n6528), .ZN(n7565)
         );
  AOI21_X1 U9343 ( .B1(n7569), .B2(n10092), .A(n7565), .ZN(n7566) );
  INV_X1 U9344 ( .A(n7566), .ZN(P2_U3466) );
  INV_X1 U9345 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7567) );
  OAI22_X1 U9346 ( .A1(n8073), .A2(n8934), .B1(n10078), .B2(n7567), .ZN(n7568)
         );
  AOI21_X1 U9347 ( .B1(n7569), .B2(n10078), .A(n7568), .ZN(n7570) );
  INV_X1 U9348 ( .A(n7570), .ZN(P2_U3411) );
  XNOR2_X1 U9349 ( .A(n7571), .B(n7572), .ZN(n9975) );
  AOI22_X1 U9350 ( .A1(n9879), .A2(n9404), .B1(n9406), .B2(n9877), .ZN(n7578)
         );
  OAI21_X1 U9351 ( .B1(n7574), .B2(n7573), .A(n7572), .ZN(n7576) );
  NAND3_X1 U9352 ( .A1(n7576), .A2(n7575), .A3(n9876), .ZN(n7577) );
  OAI211_X1 U9353 ( .C1(n9975), .C2(n7579), .A(n7578), .B(n7577), .ZN(n9978)
         );
  NAND2_X1 U9354 ( .A1(n9978), .A2(n9713), .ZN(n7588) );
  OAI22_X1 U9355 ( .A1(n9713), .A2(n7580), .B1(n9092), .B2(n9710), .ZN(n7585)
         );
  INV_X1 U9356 ( .A(n7586), .ZN(n9977) );
  INV_X1 U9357 ( .A(n7581), .ZN(n7583) );
  INV_X1 U9358 ( .A(n7628), .ZN(n7582) );
  OAI211_X1 U9359 ( .C1(n9977), .C2(n7583), .A(n7582), .B(n9890), .ZN(n9976)
         );
  NOR2_X1 U9360 ( .A1(n9976), .A2(n9904), .ZN(n7584) );
  AOI211_X1 U9361 ( .C1(n9901), .C2(n7586), .A(n7585), .B(n7584), .ZN(n7587)
         );
  OAI211_X1 U9362 ( .C1(n9975), .C2(n7589), .A(n7588), .B(n7587), .ZN(P1_U3282) );
  INV_X1 U9363 ( .A(n7590), .ZN(n9954) );
  OAI21_X1 U9364 ( .B1(n7593), .B2(n7591), .A(n7592), .ZN(n7594) );
  NAND2_X1 U9365 ( .A1(n7594), .A2(n9113), .ZN(n7598) );
  OAI22_X1 U9366 ( .A1(n9129), .A2(n9848), .B1(n9836), .B2(n9115), .ZN(n7595)
         );
  AOI211_X1 U9367 ( .C1(n9105), .C2(n9861), .A(n7596), .B(n7595), .ZN(n7597)
         );
  OAI211_X1 U9368 ( .C1(n9954), .C2(n9135), .A(n7598), .B(n7597), .ZN(P1_U3221) );
  INV_X1 U9369 ( .A(n7599), .ZN(n7602) );
  OAI222_X1 U9370 ( .A1(n7825), .A2(n7600), .B1(n9807), .B2(n7602), .C1(
        P1_U3086), .C2(n9376), .ZN(P1_U3333) );
  OAI222_X1 U9371 ( .A1(n8953), .A2(n7603), .B1(n8955), .B2(n7602), .C1(n7601), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  NAND2_X1 U9372 ( .A1(n7608), .A2(n7604), .ZN(n7605) );
  OAI211_X1 U9373 ( .C1(n7606), .C2(n7825), .A(n7605), .B(n9387), .ZN(P1_U3332) );
  NAND2_X1 U9374 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  OAI211_X1 U9375 ( .C1(n7610), .C2(n8953), .A(n7609), .B(n8200), .ZN(P2_U3272) );
  INV_X1 U9376 ( .A(n7613), .ZN(n8011) );
  XNOR2_X1 U9377 ( .A(n7611), .B(n8011), .ZN(n10057) );
  OAI211_X1 U9378 ( .C1(n7614), .C2(n7613), .A(n7612), .B(n8755), .ZN(n7616)
         );
  AOI22_X1 U9379 ( .A1(n8382), .A2(n8760), .B1(n8761), .B2(n8384), .ZN(n7615)
         );
  NAND2_X1 U9380 ( .A1(n7616), .A2(n7615), .ZN(n10059) );
  NAND2_X1 U9381 ( .A1(n10059), .A2(n10038), .ZN(n7621) );
  INV_X1 U9382 ( .A(n7717), .ZN(n7617) );
  OAI22_X1 U9383 ( .A1(n10038), .A2(n7618), .B1(n7617), .B2(n8782), .ZN(n7619)
         );
  AOI21_X1 U9384 ( .B1(n10031), .B2(n4592), .A(n7619), .ZN(n7620) );
  OAI211_X1 U9385 ( .C1(n10057), .C2(n8789), .A(n7621), .B(n7620), .ZN(
        P2_U3225) );
  XNOR2_X1 U9386 ( .A(n4425), .B(n7624), .ZN(n7623) );
  AOI222_X1 U9387 ( .A1(n9876), .A2(n7623), .B1(n9405), .B2(n9877), .C1(n9403), 
        .C2(n9879), .ZN(n9984) );
  XNOR2_X1 U9388 ( .A(n7625), .B(n7624), .ZN(n9987) );
  NAND2_X1 U9389 ( .A1(n9987), .A2(n9894), .ZN(n7633) );
  OAI22_X1 U9390 ( .A1(n9713), .A2(n7626), .B1(n9019), .B2(n9710), .ZN(n7630)
         );
  INV_X1 U9391 ( .A(n7691), .ZN(n7627) );
  OAI211_X1 U9392 ( .C1(n9985), .C2(n7628), .A(n7627), .B(n9890), .ZN(n9983)
         );
  NOR2_X1 U9393 ( .A1(n9983), .A2(n9904), .ZN(n7629) );
  AOI211_X1 U9394 ( .C1(n9901), .C2(n7631), .A(n7630), .B(n7629), .ZN(n7632)
         );
  OAI211_X1 U9395 ( .C1(n4321), .C2(n9984), .A(n7633), .B(n7632), .ZN(P1_U3281) );
  AOI21_X1 U9396 ( .B1(n8347), .B2(n8386), .A(n7634), .ZN(n7637) );
  NAND2_X1 U9397 ( .A1(n8362), .A2(n7635), .ZN(n7636) );
  OAI211_X1 U9398 ( .C1(n7666), .C2(n8359), .A(n7637), .B(n7636), .ZN(n7644)
         );
  XNOR2_X1 U9399 ( .A(n7940), .B(n10051), .ZN(n7664) );
  XNOR2_X1 U9400 ( .A(n7664), .B(n8385), .ZN(n7642) );
  NOR2_X2 U9401 ( .A1(n7641), .A2(n7642), .ZN(n7665) );
  AOI211_X1 U9402 ( .C1(n7642), .C2(n7641), .A(n8366), .B(n7665), .ZN(n7643)
         );
  AOI211_X1 U9403 ( .C1(n7645), .C2(n8375), .A(n7644), .B(n7643), .ZN(n7646)
         );
  INV_X1 U9404 ( .A(n7646), .ZN(P2_U3179) );
  AOI21_X1 U9405 ( .B1(n6547), .B2(n7648), .A(n7647), .ZN(n7663) );
  INV_X1 U9406 ( .A(n7737), .ZN(n7653) );
  NOR3_X1 U9407 ( .A1(n7651), .A2(n7650), .A3(n7649), .ZN(n7652) );
  OAI21_X1 U9408 ( .B1(n7653), .B2(n7652), .A(n8474), .ZN(n7662) );
  AOI21_X1 U9409 ( .B1(n8767), .B2(n7655), .A(n7654), .ZN(n7656) );
  NOR2_X1 U9410 ( .A1(n7656), .A2(n8484), .ZN(n7660) );
  AND2_X1 U9411 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8336) );
  OAI22_X1 U9412 ( .A1(n8506), .A2(n7658), .B1(n8505), .B2(n7657), .ZN(n7659)
         );
  NOR3_X1 U9413 ( .A1(n7660), .A2(n8336), .A3(n7659), .ZN(n7661) );
  OAI211_X1 U9414 ( .C1(n7663), .C2(n8491), .A(n7662), .B(n7661), .ZN(P2_U3193) );
  INV_X1 U9415 ( .A(n10023), .ZN(n7676) );
  INV_X1 U9416 ( .A(n8375), .ZN(n7675) );
  XNOR2_X1 U9417 ( .A(n7940), .B(n8073), .ZN(n7708) );
  XNOR2_X1 U9418 ( .A(n7708), .B(n7666), .ZN(n7667) );
  OAI21_X1 U9419 ( .B1(n4413), .B2(n7667), .A(n7711), .ZN(n7668) );
  NAND2_X1 U9420 ( .A1(n7668), .A2(n8344), .ZN(n7674) );
  INV_X1 U9421 ( .A(n8073), .ZN(n10024) );
  INV_X1 U9422 ( .A(n7669), .ZN(n7670) );
  AOI21_X1 U9423 ( .B1(n8347), .B2(n8385), .A(n7670), .ZN(n7671) );
  OAI21_X1 U9424 ( .B1(n7768), .B2(n8359), .A(n7671), .ZN(n7672) );
  AOI21_X1 U9425 ( .B1(n10024), .B2(n8362), .A(n7672), .ZN(n7673) );
  OAI211_X1 U9426 ( .C1(n7676), .C2(n7675), .A(n7674), .B(n7673), .ZN(P2_U3153) );
  NOR2_X1 U9427 ( .A1(n7812), .A2(n7679), .ZN(n9439) );
  AOI211_X1 U9428 ( .C1(n7812), .C2(n7679), .A(n9439), .B(n9484), .ZN(n7686)
         );
  OAI21_X1 U9429 ( .B1(n7397), .B2(n7681), .A(n7680), .ZN(n9430) );
  XNOR2_X1 U9430 ( .A(n9437), .B(n9430), .ZN(n7682) );
  NAND2_X1 U9431 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7682), .ZN(n9432) );
  OAI211_X1 U9432 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7682), .A(n9488), .B(
        n9432), .ZN(n7684) );
  AND2_X1 U9433 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9131) );
  AOI21_X1 U9434 ( .B1(n9478), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9131), .ZN(
        n7683) );
  OAI211_X1 U9435 ( .C1(n9490), .C2(n9437), .A(n7684), .B(n7683), .ZN(n7685)
         );
  OR2_X1 U9436 ( .A1(n7686), .A2(n7685), .ZN(P1_U3258) );
  OAI21_X1 U9437 ( .B1(n4407), .B2(n9160), .A(n7687), .ZN(n7688) );
  AOI222_X1 U9438 ( .A1(n9876), .A2(n7688), .B1(n9404), .B2(n9877), .C1(n9402), 
        .C2(n9879), .ZN(n9990) );
  XNOR2_X1 U9439 ( .A(n7689), .B(n9160), .ZN(n9993) );
  NAND2_X1 U9440 ( .A1(n9993), .A2(n9894), .ZN(n7696) );
  OAI22_X1 U9441 ( .A1(n9713), .A2(n7690), .B1(n9068), .B2(n9710), .ZN(n7693)
         );
  OAI211_X1 U9442 ( .C1(n7691), .C2(n9991), .A(n9890), .B(n7725), .ZN(n9989)
         );
  NOR2_X1 U9443 ( .A1(n9989), .A2(n9904), .ZN(n7692) );
  AOI211_X1 U9444 ( .C1(n9901), .C2(n7694), .A(n7693), .B(n7692), .ZN(n7695)
         );
  OAI211_X1 U9445 ( .C1(n4321), .C2(n9990), .A(n7696), .B(n7695), .ZN(P1_U3280) );
  OAI21_X1 U9446 ( .B1(n7699), .B2(n7697), .A(n7698), .ZN(n7700) );
  NAND2_X1 U9447 ( .A1(n7700), .A2(n9113), .ZN(n7706) );
  OAI22_X1 U9448 ( .A1(n9129), .A2(n7702), .B1(n7701), .B2(n9115), .ZN(n7703)
         );
  AOI211_X1 U9449 ( .C1(n9105), .C2(n9408), .A(n7704), .B(n7703), .ZN(n7705)
         );
  OAI211_X1 U9450 ( .C1(n7707), .C2(n9135), .A(n7706), .B(n7705), .ZN(P1_U3231) );
  INV_X1 U9451 ( .A(n7708), .ZN(n7709) );
  XNOR2_X1 U9452 ( .A(n7940), .B(n10056), .ZN(n7766) );
  XNOR2_X1 U9453 ( .A(n7766), .B(n8383), .ZN(n7712) );
  XNOR2_X1 U9454 ( .A(n7769), .B(n7712), .ZN(n7719) );
  NOR2_X1 U9455 ( .A1(n8378), .A2(n10056), .ZN(n7716) );
  AOI21_X1 U9456 ( .B1(n8347), .B2(n8384), .A(n7713), .ZN(n7714) );
  OAI21_X1 U9457 ( .B1(n8777), .B2(n8359), .A(n7714), .ZN(n7715) );
  AOI211_X1 U9458 ( .C1(n7717), .C2(n8375), .A(n7716), .B(n7715), .ZN(n7718)
         );
  OAI21_X1 U9459 ( .B1(n7719), .B2(n8366), .A(n7718), .ZN(P2_U3161) );
  XNOR2_X1 U9460 ( .A(n7720), .B(n9162), .ZN(n10001) );
  INV_X1 U9461 ( .A(n10001), .ZN(n7731) );
  XNOR2_X1 U9462 ( .A(n7721), .B(n4663), .ZN(n7722) );
  NAND2_X1 U9463 ( .A1(n7722), .A2(n9876), .ZN(n7724) );
  AOI22_X1 U9464 ( .A1(n9879), .A2(n9702), .B1(n9403), .B2(n9877), .ZN(n7723)
         );
  NAND2_X1 U9465 ( .A1(n7724), .A2(n7723), .ZN(n9999) );
  OAI211_X1 U9466 ( .C1(n4774), .C2(n9997), .A(n9890), .B(n7813), .ZN(n9995)
         );
  OAI22_X1 U9467 ( .A1(n9713), .A2(n7726), .B1(n8965), .B2(n9710), .ZN(n7727)
         );
  AOI21_X1 U9468 ( .B1(n8968), .B2(n9901), .A(n7727), .ZN(n7728) );
  OAI21_X1 U9469 ( .B1(n9995), .B2(n9904), .A(n7728), .ZN(n7729) );
  AOI21_X1 U9470 ( .B1(n9999), .B2(n9713), .A(n7729), .ZN(n7730) );
  OAI21_X1 U9471 ( .B1(n7731), .B2(n9709), .A(n7730), .ZN(P1_U3279) );
  AOI21_X1 U9472 ( .B1(n7734), .B2(n7733), .A(n7732), .ZN(n7750) );
  AND3_X1 U9473 ( .A1(n7737), .A2(n7736), .A3(n7735), .ZN(n7738) );
  OAI21_X1 U9474 ( .B1(n7783), .B2(n7738), .A(n8474), .ZN(n7749) );
  AOI21_X1 U9475 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7742) );
  NOR2_X1 U9476 ( .A1(n7742), .A2(n8484), .ZN(n7747) );
  NOR2_X1 U9477 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7743), .ZN(n8257) );
  OAI22_X1 U9478 ( .A1(n8506), .A2(n7745), .B1(n8505), .B2(n7744), .ZN(n7746)
         );
  NOR3_X1 U9479 ( .A1(n7747), .A2(n8257), .A3(n7746), .ZN(n7748) );
  OAI211_X1 U9480 ( .C1(n7750), .C2(n8491), .A(n7749), .B(n7748), .ZN(P2_U3194) );
  INV_X1 U9481 ( .A(n7751), .ZN(n7841) );
  OAI222_X1 U9482 ( .A1(P1_U3086), .A2(n7753), .B1(n9807), .B2(n7841), .C1(
        n7752), .C2(n7825), .ZN(P1_U3331) );
  XOR2_X1 U9483 ( .A(n7754), .B(n8013), .Z(n7758) );
  INV_X1 U9484 ( .A(n7758), .ZN(n10063) );
  XNOR2_X1 U9485 ( .A(n7755), .B(n8013), .ZN(n7760) );
  OAI22_X1 U9486 ( .A1(n7768), .A2(n8778), .B1(n7889), .B2(n8780), .ZN(n7756)
         );
  AOI21_X1 U9487 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7759) );
  OAI21_X1 U9488 ( .B1(n7760), .B2(n8775), .A(n7759), .ZN(n10065) );
  NAND2_X1 U9489 ( .A1(n10065), .A2(n10038), .ZN(n7765) );
  INV_X1 U9490 ( .A(n7770), .ZN(n7761) );
  OAI22_X1 U9491 ( .A1(n10038), .A2(n7762), .B1(n7761), .B2(n8782), .ZN(n7763)
         );
  AOI21_X1 U9492 ( .B1(n10031), .B2(n7775), .A(n7763), .ZN(n7764) );
  OAI211_X1 U9493 ( .C1(n10063), .C2(n8533), .A(n7765), .B(n7764), .ZN(
        P2_U3224) );
  INV_X1 U9494 ( .A(n7766), .ZN(n7767) );
  XNOR2_X1 U9495 ( .A(n10061), .B(n7940), .ZN(n7886) );
  XNOR2_X1 U9496 ( .A(n7886), .B(n8777), .ZN(n7887) );
  XNOR2_X1 U9497 ( .A(n7888), .B(n7887), .ZN(n7777) );
  NAND2_X1 U9498 ( .A1(n8375), .A2(n7770), .ZN(n7773) );
  AOI21_X1 U9499 ( .B1(n8347), .B2(n8383), .A(n7771), .ZN(n7772) );
  OAI211_X1 U9500 ( .C1(n7889), .C2(n8359), .A(n7773), .B(n7772), .ZN(n7774)
         );
  AOI21_X1 U9501 ( .B1(n7775), .B2(n8362), .A(n7774), .ZN(n7776) );
  OAI21_X1 U9502 ( .B1(n7777), .B2(n8366), .A(n7776), .ZN(P2_U3171) );
  AOI21_X1 U9503 ( .B1(n8840), .B2(n7779), .A(n7778), .ZN(n7795) );
  INV_X1 U9504 ( .A(n7780), .ZN(n7785) );
  NOR3_X1 U9505 ( .A1(n7783), .A2(n7782), .A3(n7781), .ZN(n7784) );
  OAI21_X1 U9506 ( .B1(n7785), .B2(n7784), .A(n8474), .ZN(n7794) );
  AOI21_X1 U9507 ( .B1(n6555), .B2(n7787), .A(n7786), .ZN(n7788) );
  NOR2_X1 U9508 ( .A1(n7788), .A2(n8484), .ZN(n7792) );
  AND2_X1 U9509 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8316) );
  OAI22_X1 U9510 ( .A1(n8506), .A2(n7790), .B1(n8505), .B2(n7789), .ZN(n7791)
         );
  NOR3_X1 U9511 ( .A1(n7792), .A2(n8316), .A3(n7791), .ZN(n7793) );
  OAI211_X1 U9512 ( .C1(n7795), .C2(n8491), .A(n7794), .B(n7793), .ZN(P2_U3195) );
  INV_X1 U9513 ( .A(n7796), .ZN(n7800) );
  OAI222_X1 U9514 ( .A1(n8955), .A2(n7800), .B1(P2_U3151), .B2(n7798), .C1(
        n7797), .C2(n8953), .ZN(P2_U3270) );
  OAI222_X1 U9515 ( .A1(P1_U3086), .A2(n7801), .B1(n9807), .B2(n7800), .C1(
        n7799), .C2(n7825), .ZN(P1_U3330) );
  INV_X1 U9516 ( .A(n7802), .ZN(n7806) );
  OAI222_X1 U9517 ( .A1(n8955), .A2(n7806), .B1(P2_U3151), .B2(n7804), .C1(
        n7803), .C2(n8953), .ZN(P2_U3269) );
  OAI222_X1 U9518 ( .A1(P1_U3086), .A2(n7807), .B1(n9807), .B2(n7806), .C1(
        n7805), .C2(n7825), .ZN(P1_U3329) );
  OAI21_X1 U9519 ( .B1(n7809), .B2(n9298), .A(n7808), .ZN(n7810) );
  AOI222_X1 U9520 ( .A1(n9876), .A2(n7810), .B1(n9402), .B2(n9877), .C1(n9690), 
        .C2(n9879), .ZN(n9824) );
  XNOR2_X1 U9521 ( .A(n7811), .B(n9298), .ZN(n9827) );
  NAND2_X1 U9522 ( .A1(n9827), .A2(n9894), .ZN(n7819) );
  OAI22_X1 U9523 ( .A1(n9713), .A2(n7812), .B1(n9128), .B2(n9710), .ZN(n7816)
         );
  INV_X1 U9524 ( .A(n7817), .ZN(n9825) );
  INV_X1 U9525 ( .A(n9716), .ZN(n7814) );
  OAI211_X1 U9526 ( .C1(n9825), .C2(n4777), .A(n7814), .B(n9890), .ZN(n9823)
         );
  NOR2_X1 U9527 ( .A1(n9823), .A2(n9904), .ZN(n7815) );
  AOI211_X1 U9528 ( .C1(n9901), .C2(n7817), .A(n7816), .B(n7815), .ZN(n7818)
         );
  OAI211_X1 U9529 ( .C1(n4321), .C2(n9824), .A(n7819), .B(n7818), .ZN(P1_U3278) );
  INV_X1 U9530 ( .A(n7820), .ZN(n7823) );
  AOI21_X1 U9531 ( .B1(n8951), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7821), .ZN(
        n7822) );
  OAI21_X1 U9532 ( .B1(n7823), .B2(n8955), .A(n7822), .ZN(P2_U3268) );
  INV_X1 U9533 ( .A(n7827), .ZN(n7832) );
  AOI22_X1 U9534 ( .A1(n7828), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9804), .ZN(n7829) );
  OAI21_X1 U9535 ( .B1(n7832), .B2(n9807), .A(n7829), .ZN(P1_U3327) );
  AOI21_X1 U9536 ( .B1(n8951), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7830), .ZN(
        n7831) );
  OAI21_X1 U9537 ( .B1(n7832), .B2(n8955), .A(n7831), .ZN(P2_U3267) );
  MUX2_X1 U9538 ( .A(n7833), .B(P2_REG2_REG_1__SCAN_IN), .S(n8739), .Z(n7838)
         );
  NAND2_X1 U9539 ( .A1(n7834), .A2(n8717), .ZN(n7836) );
  AOI22_X1 U9540 ( .A1(n10031), .A2(n6977), .B1(n10033), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U9541 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  OR2_X1 U9542 ( .A1(n7838), .A2(n7837), .ZN(P2_U3232) );
  OAI222_X1 U9543 ( .A1(n8955), .A2(n7841), .B1(P2_U3151), .B2(n7840), .C1(
        n7839), .C2(n8953), .ZN(P2_U3271) );
  NAND2_X1 U9544 ( .A1(n9735), .A2(n7866), .ZN(n9359) );
  INV_X1 U9545 ( .A(n7866), .ZN(n7843) );
  NAND2_X1 U9546 ( .A1(n7844), .A2(n9137), .ZN(n7846) );
  NAND2_X1 U9547 ( .A1(n5060), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U9548 ( .A1(n9728), .A2(n9530), .ZN(n9364) );
  AOI211_X1 U9549 ( .C1(n9728), .C2(n9520), .A(n9670), .B(n9512), .ZN(n9730)
         );
  INV_X1 U9550 ( .A(n9728), .ZN(n7851) );
  INV_X1 U9551 ( .A(n7848), .ZN(n7849) );
  AOI22_X1 U9552 ( .A1(n4321), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n7849), .B2(
        n9897), .ZN(n7850) );
  OAI21_X1 U9553 ( .B1(n7851), .B2(n9884), .A(n7850), .ZN(n7852) );
  AOI21_X1 U9554 ( .B1(n9730), .B2(n9893), .A(n7852), .ZN(n7871) );
  INV_X1 U9555 ( .A(n9358), .ZN(n7854) );
  XNOR2_X1 U9556 ( .A(n7855), .B(n4501), .ZN(n7856) );
  INV_X1 U9557 ( .A(P1_B_REG_SCAN_IN), .ZN(n7857) );
  OAI21_X1 U9558 ( .B1(n7858), .B2(n7857), .A(n9879), .ZN(n9505) );
  NAND2_X1 U9559 ( .A1(n7859), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7865) );
  INV_X1 U9560 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7860) );
  OR2_X1 U9561 ( .A1(n5738), .A2(n7860), .ZN(n7864) );
  INV_X1 U9562 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n7861) );
  OR2_X1 U9563 ( .A1(n7862), .A2(n7861), .ZN(n7863) );
  AND3_X1 U9564 ( .A1(n7865), .A2(n7864), .A3(n7863), .ZN(n9243) );
  OAI22_X1 U9565 ( .A1(n7866), .A2(n9833), .B1(n9505), .B2(n9243), .ZN(n7867)
         );
  NAND2_X1 U9566 ( .A1(n9731), .A2(n9713), .ZN(n7870) );
  OAI211_X1 U9567 ( .C1(n9733), .C2(n9709), .A(n7871), .B(n7870), .ZN(P1_U3356) );
  MUX2_X1 U9568 ( .A(n7873), .B(n7872), .S(n10092), .Z(n7874) );
  OAI21_X1 U9569 ( .B1(n7875), .B2(n8838), .A(n7874), .ZN(P2_U3463) );
  INV_X1 U9570 ( .A(n7876), .ZN(n8107) );
  OR2_X1 U9571 ( .A1(n8107), .A2(n8106), .ZN(n8104) );
  XNOR2_X1 U9572 ( .A(n7877), .B(n8104), .ZN(n8726) );
  INV_X1 U9573 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7880) );
  XOR2_X1 U9574 ( .A(n8104), .B(n7878), .Z(n7879) );
  INV_X1 U9575 ( .A(n8699), .ZN(n8380) );
  AOI222_X1 U9576 ( .A1(n8755), .A2(n7879), .B1(n8380), .B2(n8760), .C1(n8746), 
        .C2(n8761), .ZN(n8724) );
  MUX2_X1 U9577 ( .A(n7880), .B(n8724), .S(n10078), .Z(n7882) );
  NAND2_X1 U9578 ( .A1(n8722), .A2(n8942), .ZN(n7881) );
  OAI211_X1 U9579 ( .C1(n8726), .C2(n8945), .A(n7882), .B(n7881), .ZN(P2_U3432) );
  NAND2_X1 U9580 ( .A1(n10092), .A2(n8834), .ZN(n8848) );
  MUX2_X1 U9581 ( .A(n7883), .B(n8724), .S(n10092), .Z(n7885) );
  NAND2_X1 U9582 ( .A1(n8722), .A2(n8845), .ZN(n7884) );
  OAI211_X1 U9583 ( .C1(n8848), .C2(n8726), .A(n7885), .B(n7884), .ZN(P2_U3473) );
  XNOR2_X1 U9584 ( .A(n8786), .B(n7940), .ZN(n8230) );
  NAND2_X1 U9585 ( .A1(n7890), .A2(n7889), .ZN(n8332) );
  XNOR2_X1 U9586 ( .A(n8757), .B(n7936), .ZN(n8334) );
  OR2_X1 U9587 ( .A1(n8334), .A2(n8779), .ZN(n7892) );
  XNOR2_X1 U9588 ( .A(n8941), .B(n7940), .ZN(n7893) );
  XNOR2_X1 U9589 ( .A(n7893), .B(n8759), .ZN(n8255) );
  NAND2_X1 U9590 ( .A1(n8256), .A2(n8255), .ZN(n7895) );
  OR2_X1 U9591 ( .A1(n7893), .A2(n8735), .ZN(n7894) );
  NAND2_X1 U9592 ( .A1(n7895), .A2(n7894), .ZN(n8315) );
  XNOR2_X1 U9593 ( .A(n8841), .B(n7940), .ZN(n7896) );
  XNOR2_X1 U9594 ( .A(n7896), .B(n8746), .ZN(n8314) );
  INV_X1 U9595 ( .A(n7896), .ZN(n7897) );
  AOI21_X2 U9596 ( .B1(n8315), .B2(n8314), .A(n4904), .ZN(n8214) );
  XNOR2_X1 U9597 ( .A(n8222), .B(n7940), .ZN(n7898) );
  XNOR2_X1 U9598 ( .A(n7898), .B(n8734), .ZN(n8213) );
  NAND2_X1 U9599 ( .A1(n8214), .A2(n8213), .ZN(n8212) );
  INV_X1 U9600 ( .A(n7898), .ZN(n7899) );
  NAND2_X2 U9601 ( .A1(n8212), .A2(n7900), .ZN(n8271) );
  XNOR2_X1 U9602 ( .A(n7901), .B(n7940), .ZN(n7908) );
  XNOR2_X1 U9603 ( .A(n7908), .B(n8699), .ZN(n8367) );
  XNOR2_X1 U9604 ( .A(n8919), .B(n7940), .ZN(n7902) );
  NAND2_X1 U9605 ( .A1(n7902), .A2(n8698), .ZN(n7906) );
  INV_X1 U9606 ( .A(n7902), .ZN(n7903) );
  NAND2_X1 U9607 ( .A1(n7903), .A2(n8675), .ZN(n7904) );
  INV_X1 U9608 ( .A(n8284), .ZN(n7905) );
  XNOR2_X1 U9609 ( .A(n8925), .B(n7940), .ZN(n7907) );
  NAND2_X1 U9610 ( .A1(n7907), .A2(n8710), .ZN(n8283) );
  NOR2_X1 U9611 ( .A1(n7905), .A2(n8283), .ZN(n7911) );
  OR2_X1 U9612 ( .A1(n8367), .A2(n7911), .ZN(n8287) );
  INV_X1 U9613 ( .A(n7906), .ZN(n8342) );
  OAI21_X1 U9614 ( .B1(n7907), .B2(n8710), .A(n8283), .ZN(n8274) );
  INV_X1 U9615 ( .A(n7908), .ZN(n7909) );
  AND2_X1 U9616 ( .A1(n7909), .A2(n8380), .ZN(n8273) );
  NOR2_X1 U9617 ( .A1(n8274), .A2(n8273), .ZN(n8272) );
  AND2_X1 U9618 ( .A1(n8272), .A2(n8284), .ZN(n7910) );
  OR2_X1 U9619 ( .A1(n7911), .A2(n7910), .ZN(n8288) );
  XNOR2_X1 U9620 ( .A(n8913), .B(n7438), .ZN(n7914) );
  XNOR2_X1 U9621 ( .A(n7914), .B(n8686), .ZN(n8341) );
  INV_X1 U9622 ( .A(n7914), .ZN(n7915) );
  XNOR2_X1 U9623 ( .A(n8907), .B(n7936), .ZN(n7916) );
  NAND2_X1 U9624 ( .A1(n7916), .A2(n8676), .ZN(n8238) );
  XNOR2_X1 U9625 ( .A(n8650), .B(n7438), .ZN(n7917) );
  XNOR2_X1 U9626 ( .A(n7917), .B(n8251), .ZN(n8308) );
  INV_X1 U9627 ( .A(n7917), .ZN(n7918) );
  INV_X1 U9628 ( .A(n8251), .ZN(n8663) );
  XNOR2_X1 U9629 ( .A(n7919), .B(n7940), .ZN(n7920) );
  XNOR2_X1 U9630 ( .A(n7920), .B(n8646), .ZN(n8248) );
  NAND2_X1 U9631 ( .A1(n8247), .A2(n8248), .ZN(n7923) );
  INV_X1 U9632 ( .A(n7920), .ZN(n7921) );
  NAND2_X1 U9633 ( .A1(n7921), .A2(n8646), .ZN(n7922) );
  NAND2_X1 U9634 ( .A1(n7923), .A2(n7922), .ZN(n8323) );
  INV_X1 U9635 ( .A(n8323), .ZN(n7925) );
  XNOR2_X1 U9636 ( .A(n8890), .B(n7438), .ZN(n7926) );
  XNOR2_X1 U9637 ( .A(n7926), .B(n7927), .ZN(n8322) );
  INV_X1 U9638 ( .A(n7926), .ZN(n7928) );
  INV_X1 U9639 ( .A(n7927), .ZN(n8634) );
  NAND2_X1 U9640 ( .A1(n7928), .A2(n8634), .ZN(n7929) );
  XNOR2_X1 U9642 ( .A(n8878), .B(n7940), .ZN(n8298) );
  XNOR2_X1 U9643 ( .A(n8884), .B(n7940), .ZN(n7930) );
  OAI22_X1 U9644 ( .A1(n8298), .A2(n8577), .B1(n8327), .B2(n7930), .ZN(n7934)
         );
  INV_X1 U9645 ( .A(n7930), .ZN(n8296) );
  OAI21_X1 U9646 ( .B1(n8296), .B2(n8622), .A(n8606), .ZN(n7932) );
  NOR2_X1 U9647 ( .A1(n8606), .A2(n8622), .ZN(n7931) );
  AOI22_X1 U9648 ( .A1(n7932), .A2(n8298), .B1(n7931), .B2(n7930), .ZN(n7933)
         );
  XNOR2_X1 U9649 ( .A(n7935), .B(n8358), .ZN(n8264) );
  XNOR2_X1 U9650 ( .A(n8867), .B(n7936), .ZN(n7937) );
  NAND2_X1 U9651 ( .A1(n7937), .A2(n8550), .ZN(n8353) );
  INV_X1 U9652 ( .A(n7937), .ZN(n7938) );
  NAND2_X1 U9653 ( .A1(n7938), .A2(n8576), .ZN(n8354) );
  NAND2_X1 U9654 ( .A1(n7939), .A2(n8354), .ZN(n8204) );
  XNOR2_X1 U9655 ( .A(n8861), .B(n7940), .ZN(n7941) );
  XNOR2_X1 U9656 ( .A(n7941), .B(n8537), .ZN(n8205) );
  OAI22_X1 U9657 ( .A1(n8204), .A2(n8205), .B1(n8537), .B2(n7941), .ZN(n7946)
         );
  INV_X1 U9658 ( .A(n7942), .ZN(n7944) );
  XNOR2_X1 U9659 ( .A(n8541), .B(n7438), .ZN(n7945) );
  XNOR2_X1 U9660 ( .A(n7946), .B(n7945), .ZN(n7947) );
  NAND2_X1 U9661 ( .A1(n7947), .A2(n8344), .ZN(n7952) );
  AOI22_X1 U9662 ( .A1(n8560), .A2(n8347), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7949) );
  NAND2_X1 U9663 ( .A1(n8542), .A2(n8375), .ZN(n7948) );
  OAI211_X1 U9664 ( .C1(n8538), .C2(n8359), .A(n7949), .B(n7948), .ZN(n7950)
         );
  AOI21_X1 U9665 ( .B1(n8178), .B2(n8362), .A(n7950), .ZN(n7951) );
  NAND2_X1 U9666 ( .A1(n7952), .A2(n7951), .ZN(P2_U3160) );
  NAND2_X1 U9667 ( .A1(n7953), .A2(n9893), .ZN(n7957) );
  INV_X1 U9668 ( .A(n7954), .ZN(n7955) );
  AOI22_X1 U9669 ( .A1(n4321), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n7955), .B2(
        n9897), .ZN(n7956) );
  OAI211_X1 U9670 ( .C1(n7958), .C2(n9884), .A(n7957), .B(n7956), .ZN(n7959)
         );
  AOI21_X1 U9671 ( .B1(n7960), .B2(n9713), .A(n7959), .ZN(n7961) );
  OAI21_X1 U9672 ( .B1(n7962), .B2(n9709), .A(n7961), .ZN(P1_U3266) );
  INV_X1 U9673 ( .A(SI_29_), .ZN(n7963) );
  INV_X1 U9674 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7970) );
  MUX2_X1 U9675 ( .A(n8203), .B(n7970), .S(n7969), .Z(n7972) );
  INV_X1 U9676 ( .A(SI_30_), .ZN(n7971) );
  NAND2_X1 U9677 ( .A1(n7972), .A2(n7971), .ZN(n7978) );
  INV_X1 U9678 ( .A(n7972), .ZN(n7973) );
  NAND2_X1 U9679 ( .A1(n7973), .A2(SI_30_), .ZN(n7974) );
  NAND2_X1 U9680 ( .A1(n7978), .A2(n7974), .ZN(n7979) );
  NAND2_X1 U9681 ( .A1(n9138), .A2(n7975), .ZN(n7977) );
  OR2_X1 U9682 ( .A1(n7983), .A2(n8203), .ZN(n7976) );
  INV_X1 U9683 ( .A(n8176), .ZN(n8181) );
  MUX2_X1 U9684 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n9136), .Z(n7981) );
  XNOR2_X1 U9685 ( .A(n7981), .B(SI_31_), .ZN(n7982) );
  NAND2_X1 U9686 ( .A1(n6118), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U9687 ( .A1(n7985), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U9688 ( .A1(n7986), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7987) );
  AND3_X1 U9689 ( .A1(n7989), .A2(n7988), .A3(n7987), .ZN(n7990) );
  AND2_X1 U9690 ( .A1(n7991), .A2(n7990), .ZN(n8520) );
  NAND2_X1 U9691 ( .A1(n7999), .A2(n8520), .ZN(n8183) );
  INV_X1 U9692 ( .A(n8183), .ZN(n8028) );
  INV_X1 U9693 ( .A(n7992), .ZN(n7997) );
  NAND2_X1 U9694 ( .A1(n8791), .A2(n7993), .ZN(n8182) );
  AND2_X1 U9695 ( .A1(n8182), .A2(n7994), .ZN(n8174) );
  INV_X1 U9696 ( .A(n8174), .ZN(n7996) );
  INV_X1 U9697 ( .A(n8791), .ZN(n8854) );
  INV_X1 U9698 ( .A(n8520), .ZN(n8379) );
  NAND2_X1 U9699 ( .A1(n8851), .A2(n8379), .ZN(n8187) );
  OAI21_X1 U9700 ( .B1(n8854), .B2(n7999), .A(n8187), .ZN(n7995) );
  INV_X1 U9701 ( .A(n8187), .ZN(n8027) );
  NAND2_X1 U9702 ( .A1(n8176), .A2(n8182), .ZN(n8025) );
  INV_X1 U9703 ( .A(n8000), .ZN(n8159) );
  INV_X1 U9704 ( .A(n8585), .ZN(n8002) );
  OR2_X1 U9705 ( .A1(n8145), .A2(n8002), .ZN(n8604) );
  INV_X1 U9706 ( .A(n8604), .ZN(n8602) );
  INV_X1 U9707 ( .A(n8659), .ZN(n8661) );
  OR2_X1 U9708 ( .A1(n8124), .A2(n8003), .ZN(n8674) );
  AND4_X1 U9709 ( .A1(n8050), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(n8012)
         );
  NOR2_X1 U9710 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  NAND4_X1 U9711 ( .A1(n8012), .A2(n8011), .A3(n8010), .A4(n8009), .ZN(n8014)
         );
  NAND2_X1 U9712 ( .A1(n8752), .A2(n8089), .ZN(n8774) );
  NOR4_X1 U9713 ( .A1(n8014), .A2(n8069), .A3(n8774), .A4(n8013), .ZN(n8016)
         );
  INV_X1 U9714 ( .A(n8757), .ZN(n8015) );
  NAND4_X1 U9715 ( .A1(n8016), .A2(n8743), .A3(n8015), .A4(n8732), .ZN(n8017)
         );
  OR4_X1 U9716 ( .A1(n8104), .A2(n8695), .A3(n8017), .A4(n8711), .ZN(n8018) );
  NOR3_X1 U9717 ( .A1(n8674), .A2(n8684), .A3(n8018), .ZN(n8019) );
  NAND4_X1 U9718 ( .A1(n8631), .A2(n8643), .A3(n8661), .A4(n8019), .ZN(n8020)
         );
  NOR2_X1 U9719 ( .A1(n8020), .A2(n8136), .ZN(n8021) );
  NAND4_X1 U9720 ( .A1(n8580), .A2(n8594), .A3(n8602), .A4(n8021), .ZN(n8022)
         );
  NOR3_X1 U9721 ( .A1(n8028), .A2(n8027), .A3(n8026), .ZN(n8029) );
  NAND2_X1 U9722 ( .A1(n8035), .A2(n8033), .ZN(n8034) );
  NAND2_X1 U9723 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  NOR2_X1 U9724 ( .A1(n8040), .A2(n8185), .ZN(n8042) );
  NOR2_X1 U9725 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  NAND2_X1 U9726 ( .A1(n8044), .A2(n8043), .ZN(n8049) );
  AND2_X1 U9727 ( .A1(n8052), .A2(n8045), .ZN(n8047) );
  MUX2_X1 U9728 ( .A(n8047), .B(n8046), .S(n8185), .Z(n8048) );
  NAND2_X1 U9729 ( .A1(n8049), .A2(n8048), .ZN(n8051) );
  INV_X1 U9730 ( .A(n8052), .ZN(n8054) );
  OAI211_X1 U9731 ( .C1(n8061), .C2(n8054), .A(n8062), .B(n8053), .ZN(n8058)
         );
  AND2_X1 U9732 ( .A1(n8063), .A2(n8055), .ZN(n8057) );
  INV_X1 U9733 ( .A(n8064), .ZN(n8056) );
  AOI21_X1 U9734 ( .B1(n8058), .B2(n8057), .A(n8056), .ZN(n8067) );
  NAND2_X1 U9735 ( .A1(n8065), .A2(n8064), .ZN(n8066) );
  MUX2_X1 U9736 ( .A(n8067), .B(n8066), .S(n8171), .Z(n8071) );
  NAND2_X1 U9737 ( .A1(n8072), .A2(n8075), .ZN(n8081) );
  NAND2_X1 U9738 ( .A1(n8080), .A2(n8079), .ZN(n8068) );
  MUX2_X1 U9739 ( .A(n8081), .B(n8068), .S(n8185), .Z(n8077) );
  NOR2_X1 U9740 ( .A1(n8077), .A2(n8069), .ZN(n8070) );
  NAND2_X1 U9741 ( .A1(n8071), .A2(n8070), .ZN(n8087) );
  OAI21_X1 U9742 ( .B1(n8073), .B2(n8384), .A(n8072), .ZN(n8074) );
  INV_X1 U9743 ( .A(n8074), .ZN(n8076) );
  OAI211_X1 U9744 ( .C1(n8077), .C2(n8076), .A(n8752), .B(n8075), .ZN(n8084)
         );
  AND2_X1 U9745 ( .A1(n8079), .A2(n8078), .ZN(n8082) );
  OAI211_X1 U9746 ( .C1(n8082), .C2(n8081), .A(n8089), .B(n8080), .ZN(n8083)
         );
  MUX2_X1 U9747 ( .A(n8084), .B(n8083), .S(n8171), .Z(n8085) );
  INV_X1 U9748 ( .A(n8085), .ZN(n8086) );
  NAND2_X1 U9749 ( .A1(n8087), .A2(n8086), .ZN(n8090) );
  AOI21_X1 U9750 ( .B1(n8090), .B2(n8088), .A(n4861), .ZN(n8094) );
  NAND2_X1 U9751 ( .A1(n8090), .A2(n8089), .ZN(n8092) );
  MUX2_X1 U9752 ( .A(n8096), .B(n8095), .S(n8185), .Z(n8097) );
  INV_X1 U9753 ( .A(n8099), .ZN(n8101) );
  INV_X1 U9754 ( .A(n8841), .ZN(n8935) );
  MUX2_X1 U9755 ( .A(n8218), .B(n8935), .S(n8185), .Z(n8100) );
  AOI21_X1 U9756 ( .B1(n8102), .B2(n8101), .A(n8100), .ZN(n8103) );
  MUX2_X1 U9757 ( .A(n8107), .B(n8106), .S(n8171), .Z(n8108) );
  INV_X1 U9758 ( .A(n8711), .ZN(n8707) );
  INV_X1 U9759 ( .A(n8109), .ZN(n8110) );
  XNOR2_X1 U9760 ( .A(n8653), .B(n8171), .ZN(n8111) );
  NOR2_X1 U9761 ( .A1(n8112), .A2(n8111), .ZN(n8118) );
  NAND3_X1 U9762 ( .A1(n8133), .A2(n8185), .A3(n8113), .ZN(n8116) );
  NAND3_X1 U9763 ( .A1(n8120), .A2(n8171), .A3(n8670), .ZN(n8115) );
  AOI21_X1 U9764 ( .B1(n8122), .B2(n8669), .A(n8171), .ZN(n8114) );
  AOI21_X1 U9765 ( .B1(n8116), .B2(n8115), .A(n8114), .ZN(n8117) );
  INV_X1 U9766 ( .A(n8907), .ZN(n8242) );
  AOI21_X1 U9767 ( .B1(n8124), .B2(n8676), .A(n8242), .ZN(n8119) );
  AOI211_X1 U9768 ( .C1(n8645), .C2(n8120), .A(n8171), .B(n8119), .ZN(n8129)
         );
  NAND3_X1 U9769 ( .A1(n8907), .A2(n8645), .A3(n8171), .ZN(n8121) );
  OAI21_X1 U9770 ( .B1(n8185), .B2(n8122), .A(n8121), .ZN(n8128) );
  NAND3_X1 U9771 ( .A1(n8670), .A2(n8171), .A3(n8654), .ZN(n8123) );
  AOI211_X1 U9772 ( .C1(n8126), .C2(n8125), .A(n8124), .B(n8123), .ZN(n8127)
         );
  AOI21_X1 U9773 ( .B1(n8643), .B2(n8130), .A(n8185), .ZN(n8131) );
  NAND2_X1 U9774 ( .A1(n8138), .A2(n8132), .ZN(n8135) );
  NAND2_X1 U9775 ( .A1(n8137), .A2(n8133), .ZN(n8134) );
  MUX2_X1 U9776 ( .A(n8135), .B(n8134), .S(n8171), .Z(n8140) );
  MUX2_X1 U9777 ( .A(n8138), .B(n8137), .S(n8185), .Z(n8139) );
  AND2_X1 U9778 ( .A1(n8585), .A2(n8141), .ZN(n8142) );
  MUX2_X1 U9779 ( .A(n8143), .B(n8142), .S(n8171), .Z(n8144) );
  NOR2_X1 U9780 ( .A1(n8148), .A2(n8145), .ZN(n8147) );
  AOI21_X1 U9781 ( .B1(n8150), .B2(n8147), .A(n8146), .ZN(n8152) );
  AOI21_X1 U9782 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8151) );
  MUX2_X1 U9783 ( .A(n8152), .B(n8151), .S(n8185), .Z(n8153) );
  INV_X1 U9784 ( .A(n8154), .ZN(n8157) );
  INV_X1 U9785 ( .A(n8155), .ZN(n8156) );
  MUX2_X1 U9786 ( .A(n8157), .B(n8156), .S(n8171), .Z(n8158) );
  NOR2_X1 U9787 ( .A1(n8558), .A2(n8158), .ZN(n8162) );
  MUX2_X1 U9788 ( .A(n8160), .B(n8159), .S(n8185), .Z(n8161) );
  NAND2_X1 U9789 ( .A1(n8538), .A2(n8185), .ZN(n8165) );
  INV_X1 U9790 ( .A(n8166), .ZN(n8168) );
  MUX2_X1 U9791 ( .A(n8168), .B(n8167), .S(n8171), .Z(n8169) );
  NOR3_X1 U9792 ( .A1(n8170), .A2(n8172), .A3(n8169), .ZN(n8180) );
  MUX2_X1 U9793 ( .A(n8551), .B(n8178), .S(n8171), .Z(n8179) );
  INV_X1 U9794 ( .A(n8172), .ZN(n8173) );
  AOI21_X1 U9795 ( .B1(n8185), .B2(n8182), .A(n8181), .ZN(n8184) );
  OAI21_X1 U9796 ( .B1(n8186), .B2(n8184), .A(n8183), .ZN(n8189) );
  AND2_X1 U9797 ( .A1(n8186), .A2(n8171), .ZN(n8188) );
  OAI21_X1 U9798 ( .B1(n8189), .B2(n8188), .A(n8187), .ZN(n8191) );
  NAND2_X1 U9799 ( .A1(n8191), .A2(n8190), .ZN(n8192) );
  NAND2_X1 U9800 ( .A1(n8193), .A2(n8192), .ZN(n8195) );
  XNOR2_X1 U9801 ( .A(n8195), .B(n8194), .ZN(n8201) );
  NOR3_X1 U9802 ( .A1(n8196), .A2(n8493), .A3(n6177), .ZN(n8199) );
  OAI21_X1 U9803 ( .B1(n8200), .B2(n8197), .A(P2_B_REG_SCAN_IN), .ZN(n8198) );
  OAI22_X1 U9804 ( .A1(n8201), .A2(n8200), .B1(n8199), .B2(n8198), .ZN(
        P2_U3296) );
  INV_X1 U9805 ( .A(n9138), .ZN(n9803) );
  OAI222_X1 U9806 ( .A1(n8953), .A2(n8203), .B1(n8955), .B2(n9803), .C1(
        P2_U3151), .C2(n8202), .ZN(P2_U3265) );
  XNOR2_X1 U9807 ( .A(n8204), .B(n8205), .ZN(n8211) );
  AOI22_X1 U9808 ( .A1(n8550), .A2(n8347), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8207) );
  NAND2_X1 U9809 ( .A1(n8554), .A2(n8375), .ZN(n8206) );
  OAI211_X1 U9810 ( .C1(n8208), .C2(n8359), .A(n8207), .B(n8206), .ZN(n8209)
         );
  AOI21_X1 U9811 ( .B1(n8861), .B2(n8362), .A(n8209), .ZN(n8210) );
  OAI21_X1 U9812 ( .B1(n8211), .B2(n8366), .A(n8210), .ZN(P2_U3154) );
  OAI21_X1 U9813 ( .B1(n8214), .B2(n8213), .A(n8212), .ZN(n8215) );
  NAND2_X1 U9814 ( .A1(n8215), .A2(n8344), .ZN(n8221) );
  AOI21_X1 U9815 ( .B1(n8371), .B2(n8380), .A(n8216), .ZN(n8217) );
  OAI21_X1 U9816 ( .B1(n8218), .B2(n8373), .A(n8217), .ZN(n8219) );
  AOI21_X1 U9817 ( .B1(n8720), .B2(n8375), .A(n8219), .ZN(n8220) );
  OAI211_X1 U9818 ( .C1(n8222), .C2(n8378), .A(n8221), .B(n8220), .ZN(P2_U3155) );
  XNOR2_X1 U9819 ( .A(n8223), .B(n8296), .ZN(n8297) );
  XNOR2_X1 U9820 ( .A(n8297), .B(n8327), .ZN(n8228) );
  NAND2_X1 U9821 ( .A1(n8375), .A2(n8609), .ZN(n8225) );
  AOI22_X1 U9822 ( .A1(n8347), .A2(n8634), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8224) );
  OAI211_X1 U9823 ( .C1(n8577), .C2(n8359), .A(n8225), .B(n8224), .ZN(n8226)
         );
  AOI21_X1 U9824 ( .B1(n8884), .B2(n8362), .A(n8226), .ZN(n8227) );
  OAI21_X1 U9825 ( .B1(n8228), .B2(n8366), .A(n8227), .ZN(P2_U3156) );
  OAI21_X1 U9826 ( .B1(n8231), .B2(n8230), .A(n8229), .ZN(n8232) );
  NAND2_X1 U9827 ( .A1(n8232), .A2(n8344), .ZN(n8237) );
  AOI21_X1 U9828 ( .B1(n8347), .B2(n8382), .A(n8233), .ZN(n8234) );
  OAI21_X1 U9829 ( .B1(n8779), .B2(n8359), .A(n8234), .ZN(n8235) );
  AOI21_X1 U9830 ( .B1(n8781), .B2(n8375), .A(n8235), .ZN(n8236) );
  OAI211_X1 U9831 ( .C1(n10067), .C2(n8378), .A(n8237), .B(n8236), .ZN(
        P2_U3157) );
  NAND2_X1 U9832 ( .A1(n4412), .A2(n8238), .ZN(n8239) );
  XNOR2_X1 U9833 ( .A(n8240), .B(n8239), .ZN(n8246) );
  NAND2_X1 U9834 ( .A1(n8347), .A2(n8686), .ZN(n8241) );
  NAND2_X1 U9835 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8503) );
  OAI211_X1 U9836 ( .C1(n8251), .C2(n8359), .A(n8241), .B(n8503), .ZN(n8244)
         );
  NOR2_X1 U9837 ( .A1(n8242), .A2(n8378), .ZN(n8243) );
  AOI211_X1 U9838 ( .C1(n8666), .C2(n8375), .A(n8244), .B(n8243), .ZN(n8245)
         );
  OAI21_X1 U9839 ( .B1(n8246), .B2(n8366), .A(n8245), .ZN(P2_U3159) );
  XOR2_X1 U9840 ( .A(n8248), .B(n8247), .Z(n8254) );
  NAND2_X1 U9841 ( .A1(n8375), .A2(n8637), .ZN(n8250) );
  AOI22_X1 U9842 ( .A1(n8371), .A2(n8634), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8249) );
  OAI211_X1 U9843 ( .C1(n8251), .C2(n8373), .A(n8250), .B(n8249), .ZN(n8252)
         );
  AOI21_X1 U9844 ( .B1(n8896), .B2(n8362), .A(n8252), .ZN(n8253) );
  OAI21_X1 U9845 ( .B1(n8254), .B2(n8366), .A(n8253), .ZN(P2_U3163) );
  XNOR2_X1 U9846 ( .A(n8256), .B(n8255), .ZN(n8262) );
  NAND2_X1 U9847 ( .A1(n8375), .A2(n8749), .ZN(n8259) );
  AOI21_X1 U9848 ( .B1(n8371), .B2(n8746), .A(n8257), .ZN(n8258) );
  OAI211_X1 U9849 ( .C1(n8779), .C2(n8373), .A(n8259), .B(n8258), .ZN(n8260)
         );
  AOI21_X1 U9850 ( .B1(n8941), .B2(n8362), .A(n8260), .ZN(n8261) );
  OAI21_X1 U9851 ( .B1(n8262), .B2(n8366), .A(n8261), .ZN(P2_U3164) );
  XOR2_X1 U9852 ( .A(n8264), .B(n8263), .Z(n8270) );
  AOI22_X1 U9853 ( .A1(n8550), .A2(n8371), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8266) );
  NAND2_X1 U9854 ( .A1(n8375), .A2(n8579), .ZN(n8265) );
  OAI211_X1 U9855 ( .C1(n8577), .C2(n8373), .A(n8266), .B(n8265), .ZN(n8267)
         );
  AOI21_X1 U9856 ( .B1(n8268), .B2(n8362), .A(n8267), .ZN(n8269) );
  OAI21_X1 U9857 ( .B1(n8270), .B2(n8366), .A(n8269), .ZN(P2_U3165) );
  INV_X1 U9858 ( .A(n8925), .ZN(n8282) );
  OR2_X1 U9859 ( .A1(n8271), .A2(n8367), .ZN(n8368) );
  AND2_X1 U9860 ( .A1(n8368), .A2(n8272), .ZN(n8286) );
  INV_X1 U9861 ( .A(n8273), .ZN(n8276) );
  INV_X1 U9862 ( .A(n8274), .ZN(n8275) );
  AOI21_X1 U9863 ( .B1(n8368), .B2(n8276), .A(n8275), .ZN(n8277) );
  OAI21_X1 U9864 ( .B1(n8286), .B2(n8277), .A(n8344), .ZN(n8281) );
  NAND2_X1 U9865 ( .A1(n8347), .A2(n8380), .ZN(n8278) );
  NAND2_X1 U9866 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8434) );
  OAI211_X1 U9867 ( .C1(n8698), .C2(n8359), .A(n8278), .B(n8434), .ZN(n8279)
         );
  AOI21_X1 U9868 ( .B1(n8704), .B2(n8375), .A(n8279), .ZN(n8280) );
  OAI211_X1 U9869 ( .C1(n8282), .C2(n8378), .A(n8281), .B(n8280), .ZN(P2_U3166) );
  INV_X1 U9870 ( .A(n8919), .ZN(n8295) );
  INV_X1 U9871 ( .A(n8283), .ZN(n8285) );
  NOR3_X1 U9872 ( .A1(n8286), .A2(n8285), .A3(n8284), .ZN(n8290) );
  OR2_X1 U9873 ( .A1(n8271), .A2(n8287), .ZN(n8289) );
  OAI21_X1 U9874 ( .B1(n8290), .B2(n4912), .A(n8344), .ZN(n8294) );
  NAND2_X1 U9875 ( .A1(n8347), .A2(n8687), .ZN(n8291) );
  NAND2_X1 U9876 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8454) );
  OAI211_X1 U9877 ( .C1(n6005), .C2(n8359), .A(n8291), .B(n8454), .ZN(n8292)
         );
  AOI21_X1 U9878 ( .B1(n8690), .B2(n8375), .A(n8292), .ZN(n8293) );
  OAI211_X1 U9879 ( .C1(n8295), .C2(n8378), .A(n8294), .B(n8293), .ZN(P2_U3168) );
  OAI22_X1 U9880 ( .A1(n8297), .A2(n8622), .B1(n8296), .B2(n8223), .ZN(n8300)
         );
  XNOR2_X1 U9881 ( .A(n8298), .B(n8577), .ZN(n8299) );
  XNOR2_X1 U9882 ( .A(n8300), .B(n8299), .ZN(n8306) );
  NOR2_X1 U9883 ( .A1(n8373), .A2(n8327), .ZN(n8303) );
  OAI22_X1 U9884 ( .A1(n8358), .A2(n8359), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8301), .ZN(n8302) );
  AOI211_X1 U9885 ( .C1(n8599), .C2(n8375), .A(n8303), .B(n8302), .ZN(n8305)
         );
  NAND2_X1 U9886 ( .A1(n8878), .A2(n8362), .ZN(n8304) );
  OAI211_X1 U9887 ( .C1(n8306), .C2(n8366), .A(n8305), .B(n8304), .ZN(P2_U3169) );
  XOR2_X1 U9888 ( .A(n8308), .B(n8307), .Z(n8313) );
  NAND2_X1 U9889 ( .A1(n8375), .A2(n8649), .ZN(n8310) );
  INV_X1 U9890 ( .A(n8646), .ZN(n8621) );
  AOI22_X1 U9891 ( .A1(n8371), .A2(n8621), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8309) );
  OAI211_X1 U9892 ( .C1(n8645), .C2(n8373), .A(n8310), .B(n8309), .ZN(n8311)
         );
  AOI21_X1 U9893 ( .B1(n8650), .B2(n8362), .A(n8311), .ZN(n8312) );
  OAI21_X1 U9894 ( .B1(n8313), .B2(n8366), .A(n8312), .ZN(P2_U3173) );
  XNOR2_X1 U9895 ( .A(n8315), .B(n8314), .ZN(n8321) );
  NAND2_X1 U9896 ( .A1(n8375), .A2(n8738), .ZN(n8318) );
  AOI21_X1 U9897 ( .B1(n8347), .B2(n8759), .A(n8316), .ZN(n8317) );
  OAI211_X1 U9898 ( .C1(n8734), .C2(n8359), .A(n8318), .B(n8317), .ZN(n8319)
         );
  AOI21_X1 U9899 ( .B1(n8841), .B2(n8362), .A(n8319), .ZN(n8320) );
  OAI21_X1 U9900 ( .B1(n8321), .B2(n8366), .A(n8320), .ZN(P2_U3174) );
  AOI21_X1 U9901 ( .B1(n8323), .B2(n8322), .A(n8366), .ZN(n8325) );
  NAND2_X1 U9902 ( .A1(n8325), .A2(n8324), .ZN(n8330) );
  AOI22_X1 U9903 ( .A1(n8347), .A2(n8621), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8326) );
  OAI21_X1 U9904 ( .B1(n8327), .B2(n8359), .A(n8326), .ZN(n8328) );
  AOI21_X1 U9905 ( .B1(n8625), .B2(n8375), .A(n8328), .ZN(n8329) );
  OAI211_X1 U9906 ( .C1(n8331), .C2(n8378), .A(n8330), .B(n8329), .ZN(P2_U3175) );
  AND2_X1 U9907 ( .A1(n8229), .A2(n8332), .ZN(n8335) );
  OAI211_X1 U9908 ( .C1(n8335), .C2(n8334), .A(n8344), .B(n8333), .ZN(n8340)
         );
  AOI21_X1 U9909 ( .B1(n8347), .B2(n8762), .A(n8336), .ZN(n8337) );
  OAI21_X1 U9910 ( .B1(n8735), .B2(n8359), .A(n8337), .ZN(n8338) );
  AOI21_X1 U9911 ( .B1(n8765), .B2(n8375), .A(n8338), .ZN(n8339) );
  OAI211_X1 U9912 ( .C1(n10073), .C2(n8378), .A(n8340), .B(n8339), .ZN(
        P2_U3176) );
  NOR3_X1 U9913 ( .A1(n4912), .A2(n8342), .A3(n8341), .ZN(n8346) );
  INV_X1 U9914 ( .A(n8343), .ZN(n8345) );
  OAI21_X1 U9915 ( .B1(n8346), .B2(n8345), .A(n8344), .ZN(n8351) );
  AND2_X1 U9916 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8487) );
  AOI21_X1 U9917 ( .B1(n8347), .B2(n8675), .A(n8487), .ZN(n8348) );
  OAI21_X1 U9918 ( .B1(n8645), .B2(n8359), .A(n8348), .ZN(n8349) );
  AOI21_X1 U9919 ( .B1(n8679), .B2(n8375), .A(n8349), .ZN(n8350) );
  OAI211_X1 U9920 ( .C1(n8352), .C2(n8378), .A(n8351), .B(n8350), .ZN(P2_U3178) );
  NAND2_X1 U9921 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  XNOR2_X1 U9922 ( .A(n8356), .B(n8355), .ZN(n8365) );
  OAI22_X1 U9923 ( .A1(n8358), .A2(n8373), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8357), .ZN(n8361) );
  NOR2_X1 U9924 ( .A1(n8537), .A2(n8359), .ZN(n8360) );
  AOI211_X1 U9925 ( .C1(n8563), .C2(n8375), .A(n8361), .B(n8360), .ZN(n8364)
         );
  NAND2_X1 U9926 ( .A1(n8867), .A2(n8362), .ZN(n8363) );
  OAI211_X1 U9927 ( .C1(n8365), .C2(n8366), .A(n8364), .B(n8363), .ZN(P2_U3180) );
  AOI21_X1 U9928 ( .B1(n8271), .B2(n8367), .A(n8366), .ZN(n8369) );
  NAND2_X1 U9929 ( .A1(n8369), .A2(n8368), .ZN(n8377) );
  AND2_X1 U9930 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8410) );
  AOI21_X1 U9931 ( .B1(n8371), .B2(n8687), .A(n8410), .ZN(n8372) );
  OAI21_X1 U9932 ( .B1(n8734), .B2(n8373), .A(n8372), .ZN(n8374) );
  AOI21_X1 U9933 ( .B1(n8713), .B2(n8375), .A(n8374), .ZN(n8376) );
  OAI211_X1 U9934 ( .C1(n8932), .C2(n8378), .A(n8377), .B(n8376), .ZN(P2_U3181) );
  MUX2_X1 U9935 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8379), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8551), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9937 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8560), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9938 ( .A(n8550), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8391), .Z(
        P2_U3517) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8595), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8606), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9941 ( .A(n8622), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8391), .Z(
        P2_U3514) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8634), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8621), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8663), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8676), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9946 ( .A(n8686), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8391), .Z(
        P2_U3509) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8675), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8687), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8380), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8381), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9951 ( .A(n8746), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8391), .Z(
        P2_U3504) );
  MUX2_X1 U9952 ( .A(n8759), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8391), .Z(
        P2_U3503) );
  INV_X1 U9953 ( .A(n8779), .ZN(n8745) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8745), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8762), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8382), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9957 ( .A(n8383), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8391), .Z(
        P2_U3499) );
  MUX2_X1 U9958 ( .A(n8384), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8391), .Z(
        P2_U3498) );
  MUX2_X1 U9959 ( .A(n8385), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8391), .Z(
        P2_U3497) );
  MUX2_X1 U9960 ( .A(n8386), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8391), .Z(
        P2_U3496) );
  MUX2_X1 U9961 ( .A(n8387), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8391), .Z(
        P2_U3495) );
  MUX2_X1 U9962 ( .A(n8388), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8391), .Z(
        P2_U3494) );
  MUX2_X1 U9963 ( .A(n8389), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8391), .Z(
        P2_U3493) );
  MUX2_X1 U9964 ( .A(n8390), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8391), .Z(
        P2_U3492) );
  MUX2_X1 U9965 ( .A(n8392), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8391), .Z(
        P2_U3491) );
  INV_X1 U9966 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8836) );
  XOR2_X1 U9967 ( .A(n8414), .B(n8407), .Z(n8394) );
  NOR2_X1 U9968 ( .A1(n8836), .A2(n8394), .ZN(n8415) );
  AOI21_X1 U9969 ( .B1(n8836), .B2(n8394), .A(n8415), .ZN(n8413) );
  INV_X1 U9970 ( .A(n8395), .ZN(n8396) );
  NOR2_X1 U9971 ( .A1(n8397), .A2(n8396), .ZN(n8399) );
  MUX2_X1 U9972 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4462), .Z(n8419) );
  XNOR2_X1 U9973 ( .A(n8419), .B(n8407), .ZN(n8398) );
  AOI21_X1 U9974 ( .B1(n8399), .B2(n8398), .A(n8420), .ZN(n8400) );
  NOR2_X1 U9975 ( .A1(n8400), .A2(n8517), .ZN(n8411) );
  INV_X1 U9976 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8404) );
  AOI21_X1 U9977 ( .B1(n8404), .B2(n8403), .A(n8427), .ZN(n8405) );
  NOR2_X1 U9978 ( .A1(n8405), .A2(n8484), .ZN(n8409) );
  OAI22_X1 U9979 ( .A1(n8506), .A2(n8407), .B1(n8505), .B2(n8406), .ZN(n8408)
         );
  NOR4_X1 U9980 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n8412)
         );
  OAI21_X1 U9981 ( .B1(n8413), .B2(n8491), .A(n8412), .ZN(P2_U3197) );
  NOR2_X1 U9982 ( .A1(n8426), .A2(n8414), .ZN(n8416) );
  INV_X1 U9983 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8830) );
  AOI22_X1 U9984 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8433), .B1(n8449), .B2(
        n8830), .ZN(n8417) );
  NOR2_X1 U9985 ( .A1(n8418), .A2(n8417), .ZN(n8442) );
  AOI21_X1 U9986 ( .B1(n8418), .B2(n8417), .A(n8442), .ZN(n8441) );
  INV_X1 U9987 ( .A(n8419), .ZN(n8421) );
  AOI21_X1 U9988 ( .B1(n8426), .B2(n8421), .A(n8420), .ZN(n8446) );
  INV_X1 U9989 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8703) );
  MUX2_X1 U9990 ( .A(n8703), .B(n8830), .S(n4462), .Z(n8422) );
  NOR2_X1 U9991 ( .A1(n8422), .A2(n8433), .ZN(n8445) );
  INV_X1 U9992 ( .A(n8445), .ZN(n8423) );
  NAND2_X1 U9993 ( .A1(n8422), .A2(n8433), .ZN(n8444) );
  NAND2_X1 U9994 ( .A1(n8423), .A2(n8444), .ZN(n8424) );
  XNOR2_X1 U9995 ( .A(n8446), .B(n8424), .ZN(n8439) );
  NOR2_X1 U9996 ( .A1(n8426), .A2(n8425), .ZN(n8428) );
  MUX2_X1 U9997 ( .A(n8703), .B(P2_REG2_REG_16__SCAN_IN), .S(n8433), .Z(n8429)
         );
  INV_X1 U9998 ( .A(n8429), .ZN(n8430) );
  AOI21_X1 U9999 ( .B1(n8431), .B2(n8430), .A(n4392), .ZN(n8432) );
  NOR2_X1 U10000 ( .A1(n8432), .A2(n8484), .ZN(n8438) );
  NAND2_X1 U10001 ( .A1(n8476), .A2(n8433), .ZN(n8435) );
  OAI211_X1 U10002 ( .C1(n8436), .C2(n8505), .A(n8435), .B(n8434), .ZN(n8437)
         );
  AOI211_X1 U10003 ( .C1(n8439), .C2(n8474), .A(n8438), .B(n8437), .ZN(n8440)
         );
  OAI21_X1 U10004 ( .B1(n8441), .B2(n8491), .A(n8440), .ZN(P2_U3198) );
  INV_X1 U10005 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8827) );
  XNOR2_X1 U10006 ( .A(n8468), .B(n8461), .ZN(n8443) );
  AOI21_X1 U10007 ( .B1(n8827), .B2(n8443), .A(n8462), .ZN(n8460) );
  MUX2_X1 U10008 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4462), .Z(n8466) );
  XNOR2_X1 U10009 ( .A(n8466), .B(n8468), .ZN(n8469) );
  XNOR2_X1 U10010 ( .A(n8470), .B(n8469), .ZN(n8447) );
  NAND2_X1 U10011 ( .A1(n8447), .A2(n8474), .ZN(n8459) );
  NOR2_X1 U10012 ( .A1(n8505), .A2(n8448), .ZN(n8457) );
  INV_X1 U10013 ( .A(n8481), .ZN(n8450) );
  OAI21_X1 U10014 ( .B1(n4366), .B2(n8451), .A(n8450), .ZN(n8453) );
  INV_X1 U10015 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8452) );
  NOR2_X1 U10016 ( .A1(n8452), .A2(n8453), .ZN(n8482) );
  AOI21_X1 U10017 ( .B1(n8453), .B2(n8452), .A(n8482), .ZN(n8455) );
  OAI21_X1 U10018 ( .B1(n8484), .B2(n8455), .A(n8454), .ZN(n8456) );
  AOI211_X1 U10019 ( .C1(n8476), .C2(n8468), .A(n8457), .B(n8456), .ZN(n8458)
         );
  OAI211_X1 U10020 ( .C1(n8460), .C2(n8491), .A(n8459), .B(n8458), .ZN(
        P2_U3199) );
  NOR2_X1 U10021 ( .A1(n8468), .A2(n8461), .ZN(n8463) );
  NAND2_X1 U10022 ( .A1(n8464), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8510) );
  OAI21_X1 U10023 ( .B1(n8464), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8510), .ZN(
        n8465) );
  AOI21_X1 U10024 ( .B1(n4368), .B2(n8465), .A(n8511), .ZN(n8492) );
  INV_X1 U10025 ( .A(n8466), .ZN(n8467) );
  AOI22_X1 U10026 ( .A1(n8470), .A2(n8469), .B1(n8468), .B2(n8467), .ZN(n8472)
         );
  MUX2_X1 U10027 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4462), .Z(n8471) );
  NOR2_X1 U10028 ( .A1(n8472), .A2(n8471), .ZN(n8494) );
  NAND2_X1 U10029 ( .A1(n8472), .A2(n8471), .ZN(n8495) );
  INV_X1 U10030 ( .A(n8495), .ZN(n8473) );
  NOR2_X1 U10031 ( .A1(n8494), .A2(n8473), .ZN(n8477) );
  INV_X1 U10032 ( .A(n8477), .ZN(n8475) );
  NAND2_X1 U10033 ( .A1(n8475), .A2(n8474), .ZN(n8479) );
  AOI21_X1 U10034 ( .B1(n8477), .B2(P2_U3893), .A(n8476), .ZN(n8478) );
  MUX2_X1 U10035 ( .A(n8479), .B(n8478), .S(n8496), .Z(n8490) );
  INV_X1 U10036 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8678) );
  OR2_X1 U10037 ( .A1(n8496), .A2(n8678), .ZN(n8499) );
  NAND2_X1 U10038 ( .A1(n8496), .A2(n8678), .ZN(n8480) );
  AND2_X1 U10039 ( .A1(n8499), .A2(n8480), .ZN(n8483) );
  OAI21_X1 U10040 ( .B1(n8482), .B2(n8481), .A(n8483), .ZN(n8500) );
  OR3_X1 U10041 ( .A1(n8483), .A2(n8482), .A3(n8481), .ZN(n8485) );
  AOI21_X1 U10042 ( .B1(n8500), .B2(n8485), .A(n8484), .ZN(n8486) );
  XNOR2_X1 U10043 ( .A(n6174), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8512) );
  XNOR2_X1 U10044 ( .A(n6174), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8501) );
  MUX2_X1 U10045 ( .A(n8512), .B(n8501), .S(n8493), .Z(n8498) );
  AOI21_X1 U10046 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8497) );
  XOR2_X1 U10047 ( .A(n8498), .B(n8497), .Z(n8518) );
  INV_X1 U10048 ( .A(n8501), .ZN(n8502) );
  OAI21_X1 U10049 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8508) );
  NOR2_X1 U10050 ( .A1(n8506), .A2(n6174), .ZN(n8507) );
  XNOR2_X1 U10051 ( .A(n8513), .B(n8512), .ZN(n8515) );
  NAND2_X1 U10052 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  NOR2_X1 U10053 ( .A1(n8520), .A2(n8519), .ZN(n8849) );
  NOR2_X1 U10054 ( .A1(n8521), .A2(n8782), .ZN(n8528) );
  AOI21_X1 U10055 ( .B1(n8849), .B2(n10038), .A(n8528), .ZN(n8523) );
  NAND2_X1 U10056 ( .A1(n8739), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8522) );
  OAI211_X1 U10057 ( .C1(n8851), .C2(n8715), .A(n8523), .B(n8522), .ZN(
        P2_U3202) );
  NAND2_X1 U10058 ( .A1(n8791), .A2(n10031), .ZN(n8524) );
  OAI211_X1 U10059 ( .C1(n10038), .C2(n8525), .A(n8524), .B(n8523), .ZN(
        P2_U3203) );
  NAND2_X1 U10060 ( .A1(n8526), .A2(n10038), .ZN(n8532) );
  NOR2_X1 U10061 ( .A1(n10038), .A2(n8527), .ZN(n8529) );
  AOI211_X1 U10062 ( .C1(n8530), .C2(n10031), .A(n8529), .B(n8528), .ZN(n8531)
         );
  OAI211_X1 U10063 ( .C1(n8534), .C2(n8533), .A(n8532), .B(n8531), .ZN(
        P2_U3204) );
  XNOR2_X1 U10064 ( .A(n8536), .B(n8535), .ZN(n8540) );
  OAI22_X1 U10065 ( .A1(n8538), .A2(n8780), .B1(n8537), .B2(n8778), .ZN(n8539)
         );
  XNOR2_X1 U10066 ( .A(n4389), .B(n8541), .ZN(n8856) );
  INV_X1 U10067 ( .A(n8856), .ZN(n8545) );
  AOI22_X1 U10068 ( .A1(n8542), .A2(n10033), .B1(n8739), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8543) );
  OAI21_X1 U10069 ( .B1(n8796), .B2(n8715), .A(n8543), .ZN(n8544) );
  AOI21_X1 U10070 ( .B1(n8545), .B2(n8717), .A(n8544), .ZN(n8546) );
  OAI21_X1 U10071 ( .B1(n8795), .B2(n8739), .A(n8546), .ZN(P2_U3205) );
  XOR2_X1 U10072 ( .A(n8548), .B(n8547), .Z(n8864) );
  XNOR2_X1 U10073 ( .A(n8549), .B(n8548), .ZN(n8552) );
  AOI222_X1 U10074 ( .A1(n8755), .A2(n8552), .B1(n8551), .B2(n8760), .C1(n8550), .C2(n8761), .ZN(n8859) );
  MUX2_X1 U10075 ( .A(n8553), .B(n8859), .S(n10038), .Z(n8556) );
  AOI22_X1 U10076 ( .A1(n8861), .A2(n10031), .B1(n10033), .B2(n8554), .ZN(
        n8555) );
  OAI211_X1 U10077 ( .C1(n8864), .C2(n8789), .A(n8556), .B(n8555), .ZN(
        P2_U3206) );
  XNOR2_X1 U10078 ( .A(n8557), .B(n8558), .ZN(n8870) );
  XNOR2_X1 U10079 ( .A(n8559), .B(n8558), .ZN(n8561) );
  AOI222_X1 U10080 ( .A1(n8755), .A2(n8561), .B1(n8560), .B2(n8760), .C1(n8595), .C2(n8761), .ZN(n8865) );
  MUX2_X1 U10081 ( .A(n8562), .B(n8865), .S(n10038), .Z(n8565) );
  AOI22_X1 U10082 ( .A1(n8867), .A2(n10031), .B1(n10033), .B2(n8563), .ZN(
        n8564) );
  OAI211_X1 U10083 ( .C1(n8870), .C2(n8789), .A(n8565), .B(n8564), .ZN(
        P2_U3207) );
  NOR2_X1 U10084 ( .A1(n8872), .A2(n8736), .ZN(n8578) );
  OR2_X1 U10085 ( .A1(n8566), .A2(n8567), .ZN(n8569) );
  NAND2_X1 U10086 ( .A1(n8569), .A2(n8568), .ZN(n8571) );
  NAND2_X1 U10087 ( .A1(n8571), .A2(n8570), .ZN(n8574) );
  AOI21_X1 U10088 ( .B1(n8580), .B2(n8574), .A(n4913), .ZN(n8575) );
  OAI222_X1 U10089 ( .A1(n8778), .A2(n8577), .B1(n8780), .B2(n8576), .C1(n8775), .C2(n8575), .ZN(n8871) );
  AOI211_X1 U10090 ( .C1(n10033), .C2(n8579), .A(n8578), .B(n8871), .ZN(n8584)
         );
  XOR2_X1 U10091 ( .A(n8581), .B(n8580), .Z(n8873) );
  INV_X1 U10092 ( .A(n8873), .ZN(n8582) );
  AOI22_X1 U10093 ( .A1(n8582), .A2(n8717), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8739), .ZN(n8583) );
  OAI21_X1 U10094 ( .B1(n8584), .B2(n8739), .A(n8583), .ZN(P2_U3208) );
  NAND2_X1 U10095 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  NAND2_X1 U10097 ( .A1(n8605), .A2(n8590), .ZN(n8592) );
  NAND2_X1 U10098 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  XOR2_X1 U10099 ( .A(n8594), .B(n8593), .Z(n8596) );
  AOI222_X1 U10100 ( .A1(n8755), .A2(n8596), .B1(n8595), .B2(n8760), .C1(n8622), .C2(n8761), .ZN(n8876) );
  OAI21_X1 U10101 ( .B1(n8597), .B2(n8736), .A(n8876), .ZN(n8598) );
  NAND2_X1 U10102 ( .A1(n8598), .A2(n10038), .ZN(n8601) );
  AOI22_X1 U10103 ( .A1(n8739), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n10033), 
        .B2(n8599), .ZN(n8600) );
  OAI211_X1 U10104 ( .C1(n8881), .C2(n8789), .A(n8601), .B(n8600), .ZN(
        P2_U3209) );
  XNOR2_X1 U10105 ( .A(n8603), .B(n8602), .ZN(n8887) );
  INV_X1 U10106 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8608) );
  XNOR2_X1 U10107 ( .A(n8605), .B(n8604), .ZN(n8607) );
  AOI222_X1 U10108 ( .A1(n8755), .A2(n8607), .B1(n8606), .B2(n8760), .C1(n8634), .C2(n8761), .ZN(n8882) );
  MUX2_X1 U10109 ( .A(n8608), .B(n8882), .S(n10038), .Z(n8611) );
  AOI22_X1 U10110 ( .A1(n8884), .A2(n10031), .B1(n10033), .B2(n8609), .ZN(
        n8610) );
  OAI211_X1 U10111 ( .C1(n8887), .C2(n8789), .A(n8611), .B(n8610), .ZN(
        P2_U3210) );
  XNOR2_X1 U10112 ( .A(n8612), .B(n6077), .ZN(n8893) );
  INV_X1 U10113 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8624) );
  AND2_X1 U10114 ( .A1(n8614), .A2(n8613), .ZN(n8620) );
  OR2_X1 U10115 ( .A1(n8566), .A2(n8615), .ZN(n8617) );
  NAND3_X1 U10116 ( .A1(n8633), .A2(n6077), .A3(n8618), .ZN(n8619) );
  NAND2_X1 U10117 ( .A1(n8620), .A2(n8619), .ZN(n8623) );
  AOI222_X1 U10118 ( .A1(n8755), .A2(n8623), .B1(n8622), .B2(n8760), .C1(n8621), .C2(n8761), .ZN(n8888) );
  MUX2_X1 U10119 ( .A(n8624), .B(n8888), .S(n10038), .Z(n8627) );
  AOI22_X1 U10120 ( .A1(n8890), .A2(n10031), .B1(n10033), .B2(n8625), .ZN(
        n8626) );
  OAI211_X1 U10121 ( .C1(n8893), .C2(n8789), .A(n8627), .B(n8626), .ZN(
        P2_U3211) );
  XNOR2_X1 U10122 ( .A(n8629), .B(n8628), .ZN(n8899) );
  OR2_X1 U10123 ( .A1(n8566), .A2(n8643), .ZN(n8641) );
  NAND3_X1 U10124 ( .A1(n8641), .A2(n8631), .A3(n8630), .ZN(n8632) );
  NAND2_X1 U10125 ( .A1(n8633), .A2(n8632), .ZN(n8635) );
  AOI222_X1 U10126 ( .A1(n8755), .A2(n8635), .B1(n8634), .B2(n8760), .C1(n8663), .C2(n8761), .ZN(n8894) );
  MUX2_X1 U10127 ( .A(n8636), .B(n8894), .S(n10038), .Z(n8639) );
  AOI22_X1 U10128 ( .A1(n8896), .A2(n10031), .B1(n10033), .B2(n8637), .ZN(
        n8638) );
  OAI211_X1 U10129 ( .C1(n8899), .C2(n8789), .A(n8639), .B(n8638), .ZN(
        P2_U3212) );
  XNOR2_X1 U10130 ( .A(n8640), .B(n8643), .ZN(n8902) );
  INV_X1 U10131 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8648) );
  INV_X1 U10132 ( .A(n8641), .ZN(n8642) );
  AOI21_X1 U10133 ( .B1(n8643), .B2(n8566), .A(n8642), .ZN(n8644) );
  OAI222_X1 U10134 ( .A1(n8780), .A2(n8646), .B1(n8778), .B2(n8645), .C1(n8775), .C2(n8644), .ZN(n8900) );
  INV_X1 U10135 ( .A(n8900), .ZN(n8647) );
  MUX2_X1 U10136 ( .A(n8648), .B(n8647), .S(n10038), .Z(n8652) );
  AOI22_X1 U10137 ( .A1(n8650), .A2(n10031), .B1(n10033), .B2(n8649), .ZN(
        n8651) );
  OAI211_X1 U10138 ( .C1(n8902), .C2(n8789), .A(n8652), .B(n8651), .ZN(
        P2_U3213) );
  NAND2_X1 U10139 ( .A1(n8693), .A2(n8653), .ZN(n8655) );
  NAND2_X1 U10140 ( .A1(n8655), .A2(n8654), .ZN(n8682) );
  NAND2_X1 U10141 ( .A1(n8682), .A2(n8656), .ZN(n8657) );
  AND2_X1 U10142 ( .A1(n8658), .A2(n8657), .ZN(n8660) );
  XNOR2_X1 U10143 ( .A(n8660), .B(n8659), .ZN(n8910) );
  INV_X1 U10144 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8665) );
  XNOR2_X1 U10145 ( .A(n8662), .B(n8661), .ZN(n8664) );
  AOI222_X1 U10146 ( .A1(n8755), .A2(n8664), .B1(n8663), .B2(n8760), .C1(n8686), .C2(n8761), .ZN(n8905) );
  MUX2_X1 U10147 ( .A(n8665), .B(n8905), .S(n10038), .Z(n8668) );
  AOI22_X1 U10148 ( .A1(n8907), .A2(n10031), .B1(n10033), .B2(n8666), .ZN(
        n8667) );
  OAI211_X1 U10149 ( .C1(n8910), .C2(n8789), .A(n8668), .B(n8667), .ZN(
        P2_U3214) );
  NAND2_X1 U10150 ( .A1(n8682), .A2(n8669), .ZN(n8671) );
  NAND2_X1 U10151 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  XOR2_X1 U10152 ( .A(n8674), .B(n8672), .Z(n8916) );
  XOR2_X1 U10153 ( .A(n8674), .B(n8673), .Z(n8677) );
  AOI222_X1 U10154 ( .A1(n8755), .A2(n8677), .B1(n8676), .B2(n8760), .C1(n8675), .C2(n8761), .ZN(n8911) );
  MUX2_X1 U10155 ( .A(n8678), .B(n8911), .S(n10038), .Z(n8681) );
  AOI22_X1 U10156 ( .A1(n8913), .A2(n10031), .B1(n10033), .B2(n8679), .ZN(
        n8680) );
  OAI211_X1 U10157 ( .C1(n8916), .C2(n8789), .A(n8681), .B(n8680), .ZN(
        P2_U3215) );
  XOR2_X1 U10158 ( .A(n8684), .B(n8682), .Z(n8922) );
  OAI211_X1 U10159 ( .C1(n8685), .C2(n8684), .A(n8683), .B(n8755), .ZN(n8689)
         );
  AOI22_X1 U10160 ( .A1(n8687), .A2(n8761), .B1(n8760), .B2(n8686), .ZN(n8688)
         );
  MUX2_X1 U10161 ( .A(n8452), .B(n8917), .S(n10038), .Z(n8692) );
  AOI22_X1 U10162 ( .A1(n8919), .A2(n10031), .B1(n10033), .B2(n8690), .ZN(
        n8691) );
  OAI211_X1 U10163 ( .C1(n8922), .C2(n8789), .A(n8692), .B(n8691), .ZN(
        P2_U3216) );
  XOR2_X1 U10164 ( .A(n8693), .B(n8695), .Z(n8928) );
  INV_X1 U10165 ( .A(n8694), .ZN(n8697) );
  INV_X1 U10166 ( .A(n8695), .ZN(n8696) );
  AOI21_X1 U10167 ( .B1(n8697), .B2(n8696), .A(n8775), .ZN(n8702) );
  OAI22_X1 U10168 ( .A1(n8699), .A2(n8778), .B1(n8698), .B2(n8780), .ZN(n8700)
         );
  AOI21_X1 U10169 ( .B1(n8702), .B2(n8701), .A(n8700), .ZN(n8923) );
  MUX2_X1 U10170 ( .A(n8703), .B(n8923), .S(n10038), .Z(n8706) );
  AOI22_X1 U10171 ( .A1(n8925), .A2(n10031), .B1(n10033), .B2(n8704), .ZN(
        n8705) );
  OAI211_X1 U10172 ( .C1(n8928), .C2(n8789), .A(n8706), .B(n8705), .ZN(
        P2_U3217) );
  XNOR2_X1 U10173 ( .A(n8708), .B(n8707), .ZN(n8709) );
  OAI222_X1 U10174 ( .A1(n8780), .A2(n8710), .B1(n8778), .B2(n8734), .C1(n8775), .C2(n8709), .ZN(n8833) );
  INV_X1 U10175 ( .A(n8833), .ZN(n8719) );
  XNOR2_X1 U10176 ( .A(n8712), .B(n8711), .ZN(n8835) );
  AOI22_X1 U10177 ( .A1(n8739), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n10033), 
        .B2(n8713), .ZN(n8714) );
  OAI21_X1 U10178 ( .B1(n8932), .B2(n8715), .A(n8714), .ZN(n8716) );
  AOI21_X1 U10179 ( .B1(n8835), .B2(n8717), .A(n8716), .ZN(n8718) );
  OAI21_X1 U10180 ( .B1(n8719), .B2(n8739), .A(n8718), .ZN(P2_U3218) );
  INV_X1 U10181 ( .A(n8736), .ZN(n8721) );
  AOI22_X1 U10182 ( .A1(n8722), .A2(n8721), .B1(n10033), .B2(n8720), .ZN(n8723) );
  AOI21_X1 U10183 ( .B1(n8724), .B2(n8723), .A(n8739), .ZN(n8728) );
  OAI22_X1 U10184 ( .A1(n8726), .A2(n8789), .B1(n8725), .B2(n10038), .ZN(n8727) );
  OR2_X1 U10185 ( .A1(n8728), .A2(n8727), .ZN(P2_U3219) );
  XNOR2_X1 U10186 ( .A(n8729), .B(n8732), .ZN(n8936) );
  AOI21_X1 U10187 ( .B1(n8732), .B2(n8731), .A(n8730), .ZN(n8733) );
  OAI222_X1 U10188 ( .A1(n8778), .A2(n8735), .B1(n8780), .B2(n8734), .C1(n8775), .C2(n8733), .ZN(n8933) );
  INV_X1 U10189 ( .A(n8933), .ZN(n8839) );
  OAI21_X1 U10190 ( .B1(n8935), .B2(n8736), .A(n8839), .ZN(n8737) );
  NAND2_X1 U10191 ( .A1(n8737), .A2(n10038), .ZN(n8741) );
  AOI22_X1 U10192 ( .A1(n8739), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10033), 
        .B2(n8738), .ZN(n8740) );
  OAI211_X1 U10193 ( .C1(n8936), .C2(n8789), .A(n8741), .B(n8740), .ZN(
        P2_U3220) );
  XNOR2_X1 U10194 ( .A(n8742), .B(n8743), .ZN(n8946) );
  XNOR2_X1 U10195 ( .A(n8744), .B(n8743), .ZN(n8747) );
  AOI222_X1 U10196 ( .A1(n8755), .A2(n8747), .B1(n8746), .B2(n8760), .C1(n8745), .C2(n8761), .ZN(n8939) );
  MUX2_X1 U10197 ( .A(n8748), .B(n8939), .S(n10038), .Z(n8751) );
  AOI22_X1 U10198 ( .A1(n8941), .A2(n10031), .B1(n10033), .B2(n8749), .ZN(
        n8750) );
  OAI211_X1 U10199 ( .C1(n8946), .C2(n8789), .A(n8751), .B(n8750), .ZN(
        P2_U3221) );
  NAND2_X1 U10200 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  XNOR2_X1 U10201 ( .A(n8754), .B(n8757), .ZN(n10075) );
  OAI211_X1 U10202 ( .C1(n8758), .C2(n8757), .A(n8756), .B(n8755), .ZN(n8764)
         );
  AOI22_X1 U10203 ( .A1(n8762), .A2(n8761), .B1(n8760), .B2(n8759), .ZN(n8763)
         );
  NAND2_X1 U10204 ( .A1(n8764), .A2(n8763), .ZN(n10077) );
  NAND2_X1 U10205 ( .A1(n10077), .A2(n10038), .ZN(n8771) );
  INV_X1 U10206 ( .A(n8765), .ZN(n8766) );
  OAI22_X1 U10207 ( .A1(n10038), .A2(n8767), .B1(n8766), .B2(n8782), .ZN(n8768) );
  AOI21_X1 U10208 ( .B1(n10031), .B2(n8769), .A(n8768), .ZN(n8770) );
  OAI211_X1 U10209 ( .C1(n8789), .C2(n10075), .A(n8771), .B(n8770), .ZN(
        P2_U3222) );
  XNOR2_X1 U10210 ( .A(n8772), .B(n8774), .ZN(n10068) );
  XOR2_X1 U10211 ( .A(n8774), .B(n8773), .Z(n8776) );
  OAI222_X1 U10212 ( .A1(n8780), .A2(n8779), .B1(n8778), .B2(n8777), .C1(n8776), .C2(n8775), .ZN(n10070) );
  NAND2_X1 U10213 ( .A1(n10070), .A2(n10038), .ZN(n8788) );
  INV_X1 U10214 ( .A(n8781), .ZN(n8783) );
  OAI22_X1 U10215 ( .A1(n10038), .A2(n8784), .B1(n8783), .B2(n8782), .ZN(n8785) );
  AOI21_X1 U10216 ( .B1(n10031), .B2(n8786), .A(n8785), .ZN(n8787) );
  OAI211_X1 U10217 ( .C1(n8789), .C2(n10068), .A(n8788), .B(n8787), .ZN(
        P2_U3223) );
  NAND2_X1 U10218 ( .A1(n8849), .A2(n10092), .ZN(n8792) );
  NAND2_X1 U10219 ( .A1(n10090), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8790) );
  OAI211_X1 U10220 ( .C1(n8851), .C2(n8838), .A(n8792), .B(n8790), .ZN(
        P2_U3490) );
  INV_X1 U10221 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U10222 ( .A1(n8791), .A2(n8845), .ZN(n8793) );
  OAI211_X1 U10223 ( .C1(n10092), .C2(n8794), .A(n8793), .B(n8792), .ZN(
        P2_U3489) );
  OAI21_X1 U10224 ( .B1(n8796), .B2(n10072), .A(n8795), .ZN(n8855) );
  MUX2_X1 U10225 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8855), .S(n10092), .Z(
        n8798) );
  NOR2_X1 U10226 ( .A1(n8856), .A2(n8848), .ZN(n8797) );
  OR2_X1 U10227 ( .A1(n8798), .A2(n8797), .ZN(P2_U3487) );
  INV_X1 U10228 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8799) );
  MUX2_X1 U10229 ( .A(n8799), .B(n8859), .S(n10092), .Z(n8801) );
  NAND2_X1 U10230 ( .A1(n8861), .A2(n8845), .ZN(n8800) );
  OAI211_X1 U10231 ( .C1(n8864), .C2(n8848), .A(n8801), .B(n8800), .ZN(
        P2_U3486) );
  INV_X1 U10232 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10233 ( .A(n8802), .B(n8865), .S(n10092), .Z(n8804) );
  NAND2_X1 U10234 ( .A1(n8867), .A2(n8845), .ZN(n8803) );
  OAI211_X1 U10235 ( .C1(n8848), .C2(n8870), .A(n8804), .B(n8803), .ZN(
        P2_U3485) );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8871), .S(n10092), .Z(
        n8806) );
  OAI22_X1 U10237 ( .A1(n8873), .A2(n8848), .B1(n8872), .B2(n8838), .ZN(n8805)
         );
  OR2_X1 U10238 ( .A1(n8806), .A2(n8805), .ZN(P2_U3484) );
  INV_X1 U10239 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8807) );
  MUX2_X1 U10240 ( .A(n8807), .B(n8876), .S(n10092), .Z(n8809) );
  NAND2_X1 U10241 ( .A1(n8878), .A2(n8845), .ZN(n8808) );
  OAI211_X1 U10242 ( .C1(n8848), .C2(n8881), .A(n8809), .B(n8808), .ZN(
        P2_U3483) );
  MUX2_X1 U10243 ( .A(n8810), .B(n8882), .S(n10092), .Z(n8812) );
  NAND2_X1 U10244 ( .A1(n8884), .A2(n8845), .ZN(n8811) );
  OAI211_X1 U10245 ( .C1(n8887), .C2(n8848), .A(n8812), .B(n8811), .ZN(
        P2_U3482) );
  INV_X1 U10246 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8813) );
  MUX2_X1 U10247 ( .A(n8813), .B(n8888), .S(n10092), .Z(n8815) );
  NAND2_X1 U10248 ( .A1(n8890), .A2(n8845), .ZN(n8814) );
  OAI211_X1 U10249 ( .C1(n8893), .C2(n8848), .A(n8815), .B(n8814), .ZN(
        P2_U3481) );
  MUX2_X1 U10250 ( .A(n8816), .B(n8894), .S(n10092), .Z(n8818) );
  NAND2_X1 U10251 ( .A1(n8896), .A2(n8845), .ZN(n8817) );
  OAI211_X1 U10252 ( .C1(n8848), .C2(n8899), .A(n8818), .B(n8817), .ZN(
        P2_U3480) );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8900), .S(n10092), .Z(
        n8820) );
  OAI22_X1 U10254 ( .A1(n8902), .A2(n8848), .B1(n8901), .B2(n8838), .ZN(n8819)
         );
  OR2_X1 U10255 ( .A1(n8820), .A2(n8819), .ZN(P2_U3479) );
  INV_X1 U10256 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8821) );
  MUX2_X1 U10257 ( .A(n8821), .B(n8905), .S(n10092), .Z(n8823) );
  NAND2_X1 U10258 ( .A1(n8907), .A2(n8845), .ZN(n8822) );
  OAI211_X1 U10259 ( .C1(n8848), .C2(n8910), .A(n8823), .B(n8822), .ZN(
        P2_U3478) );
  INV_X1 U10260 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8824) );
  MUX2_X1 U10261 ( .A(n8824), .B(n8911), .S(n10092), .Z(n8826) );
  NAND2_X1 U10262 ( .A1(n8913), .A2(n8845), .ZN(n8825) );
  OAI211_X1 U10263 ( .C1(n8916), .C2(n8848), .A(n8826), .B(n8825), .ZN(
        P2_U3477) );
  MUX2_X1 U10264 ( .A(n8827), .B(n8917), .S(n10092), .Z(n8829) );
  NAND2_X1 U10265 ( .A1(n8919), .A2(n8845), .ZN(n8828) );
  OAI211_X1 U10266 ( .C1(n8922), .C2(n8848), .A(n8829), .B(n8828), .ZN(
        P2_U3476) );
  MUX2_X1 U10267 ( .A(n8830), .B(n8923), .S(n10092), .Z(n8832) );
  NAND2_X1 U10268 ( .A1(n8925), .A2(n8845), .ZN(n8831) );
  OAI211_X1 U10269 ( .C1(n8928), .C2(n8848), .A(n8832), .B(n8831), .ZN(
        P2_U3475) );
  AOI21_X1 U10270 ( .B1(n8835), .B2(n8834), .A(n8833), .ZN(n8929) );
  MUX2_X1 U10271 ( .A(n8836), .B(n8929), .S(n10092), .Z(n8837) );
  OAI21_X1 U10272 ( .B1(n8932), .B2(n8838), .A(n8837), .ZN(P2_U3474) );
  MUX2_X1 U10273 ( .A(n8840), .B(n8839), .S(n10092), .Z(n8843) );
  NAND2_X1 U10274 ( .A1(n8841), .A2(n8845), .ZN(n8842) );
  OAI211_X1 U10275 ( .C1(n8848), .C2(n8936), .A(n8843), .B(n8842), .ZN(
        P2_U3472) );
  MUX2_X1 U10276 ( .A(n8844), .B(n8939), .S(n10092), .Z(n8847) );
  NAND2_X1 U10277 ( .A1(n8941), .A2(n8845), .ZN(n8846) );
  OAI211_X1 U10278 ( .C1(n8946), .C2(n8848), .A(n8847), .B(n8846), .ZN(
        P2_U3471) );
  NAND2_X1 U10279 ( .A1(n8849), .A2(n10078), .ZN(n8852) );
  NAND2_X1 U10280 ( .A1(n10080), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8850) );
  OAI211_X1 U10281 ( .C1(n8851), .C2(n8934), .A(n8852), .B(n8850), .ZN(
        P2_U3458) );
  NAND2_X1 U10282 ( .A1(n10080), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8853) );
  OAI211_X1 U10283 ( .C1(n8854), .C2(n8934), .A(n8853), .B(n8852), .ZN(
        P2_U3457) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8855), .S(n10078), .Z(
        n8858) );
  NOR2_X1 U10285 ( .A1(n8856), .A2(n8945), .ZN(n8857) );
  OR2_X1 U10286 ( .A1(n8858), .A2(n8857), .ZN(P2_U3455) );
  INV_X1 U10287 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8860) );
  MUX2_X1 U10288 ( .A(n8860), .B(n8859), .S(n10078), .Z(n8863) );
  NAND2_X1 U10289 ( .A1(n8861), .A2(n8942), .ZN(n8862) );
  OAI211_X1 U10290 ( .C1(n8864), .C2(n8945), .A(n8863), .B(n8862), .ZN(
        P2_U3454) );
  INV_X1 U10291 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U10292 ( .A(n8866), .B(n8865), .S(n10078), .Z(n8869) );
  NAND2_X1 U10293 ( .A1(n8867), .A2(n8942), .ZN(n8868) );
  OAI211_X1 U10294 ( .C1(n8870), .C2(n8945), .A(n8869), .B(n8868), .ZN(
        P2_U3453) );
  MUX2_X1 U10295 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8871), .S(n10078), .Z(
        n8875) );
  OAI22_X1 U10296 ( .A1(n8873), .A2(n8945), .B1(n8872), .B2(n8934), .ZN(n8874)
         );
  OR2_X1 U10297 ( .A1(n8875), .A2(n8874), .ZN(P2_U3452) );
  INV_X1 U10298 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8877) );
  MUX2_X1 U10299 ( .A(n8877), .B(n8876), .S(n10078), .Z(n8880) );
  NAND2_X1 U10300 ( .A1(n8878), .A2(n8942), .ZN(n8879) );
  OAI211_X1 U10301 ( .C1(n8881), .C2(n8945), .A(n8880), .B(n8879), .ZN(
        P2_U3451) );
  INV_X1 U10302 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8883) );
  MUX2_X1 U10303 ( .A(n8883), .B(n8882), .S(n10078), .Z(n8886) );
  NAND2_X1 U10304 ( .A1(n8884), .A2(n8942), .ZN(n8885) );
  OAI211_X1 U10305 ( .C1(n8887), .C2(n8945), .A(n8886), .B(n8885), .ZN(
        P2_U3450) );
  INV_X1 U10306 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U10307 ( .A(n8889), .B(n8888), .S(n10078), .Z(n8892) );
  NAND2_X1 U10308 ( .A1(n8890), .A2(n8942), .ZN(n8891) );
  OAI211_X1 U10309 ( .C1(n8893), .C2(n8945), .A(n8892), .B(n8891), .ZN(
        P2_U3449) );
  INV_X1 U10310 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10311 ( .A(n8895), .B(n8894), .S(n10078), .Z(n8898) );
  NAND2_X1 U10312 ( .A1(n8896), .A2(n8942), .ZN(n8897) );
  OAI211_X1 U10313 ( .C1(n8899), .C2(n8945), .A(n8898), .B(n8897), .ZN(
        P2_U3448) );
  MUX2_X1 U10314 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8900), .S(n10078), .Z(
        n8904) );
  OAI22_X1 U10315 ( .A1(n8902), .A2(n8945), .B1(n8901), .B2(n8934), .ZN(n8903)
         );
  OR2_X1 U10316 ( .A1(n8904), .A2(n8903), .ZN(P2_U3447) );
  MUX2_X1 U10317 ( .A(n8906), .B(n8905), .S(n10078), .Z(n8909) );
  NAND2_X1 U10318 ( .A1(n8907), .A2(n8942), .ZN(n8908) );
  OAI211_X1 U10319 ( .C1(n8910), .C2(n8945), .A(n8909), .B(n8908), .ZN(
        P2_U3446) );
  INV_X1 U10320 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8912) );
  MUX2_X1 U10321 ( .A(n8912), .B(n8911), .S(n10078), .Z(n8915) );
  NAND2_X1 U10322 ( .A1(n8913), .A2(n8942), .ZN(n8914) );
  OAI211_X1 U10323 ( .C1(n8916), .C2(n8945), .A(n8915), .B(n8914), .ZN(
        P2_U3444) );
  INV_X1 U10324 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8918) );
  MUX2_X1 U10325 ( .A(n8918), .B(n8917), .S(n10078), .Z(n8921) );
  NAND2_X1 U10326 ( .A1(n8919), .A2(n8942), .ZN(n8920) );
  OAI211_X1 U10327 ( .C1(n8922), .C2(n8945), .A(n8921), .B(n8920), .ZN(
        P2_U3441) );
  INV_X1 U10328 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8924) );
  MUX2_X1 U10329 ( .A(n8924), .B(n8923), .S(n10078), .Z(n8927) );
  NAND2_X1 U10330 ( .A1(n8925), .A2(n8942), .ZN(n8926) );
  OAI211_X1 U10331 ( .C1(n8928), .C2(n8945), .A(n8927), .B(n8926), .ZN(
        P2_U3438) );
  INV_X1 U10332 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8930) );
  MUX2_X1 U10333 ( .A(n8930), .B(n8929), .S(n10078), .Z(n8931) );
  OAI21_X1 U10334 ( .B1(n8932), .B2(n8934), .A(n8931), .ZN(P2_U3435) );
  MUX2_X1 U10335 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8933), .S(n10078), .Z(
        n8938) );
  OAI22_X1 U10336 ( .A1(n8936), .A2(n8945), .B1(n8935), .B2(n8934), .ZN(n8937)
         );
  OR2_X1 U10337 ( .A1(n8938), .A2(n8937), .ZN(P2_U3429) );
  INV_X1 U10338 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8940) );
  MUX2_X1 U10339 ( .A(n8940), .B(n8939), .S(n10078), .Z(n8944) );
  NAND2_X1 U10340 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  OAI211_X1 U10341 ( .C1(n8946), .C2(n8945), .A(n8944), .B(n8943), .ZN(
        P2_U3426) );
  MUX2_X1 U10342 ( .A(P2_D_REG_1__SCAN_IN), .B(n8948), .S(n8947), .Z(P2_U3377)
         );
  NOR4_X1 U10343 ( .A1(n8949), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5865), .ZN(n8950) );
  AOI21_X1 U10344 ( .B1(n8951), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8950), .ZN(
        n8952) );
  OAI21_X1 U10345 ( .B1(n9801), .B2(n8955), .A(n8952), .ZN(P2_U3264) );
  INV_X1 U10346 ( .A(n7844), .ZN(n9808) );
  OAI222_X1 U10347 ( .A1(n8955), .A2(n9808), .B1(n5777), .B2(P2_U3151), .C1(
        n8954), .C2(n8953), .ZN(P2_U3266) );
  MUX2_X1 U10348 ( .A(n8956), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10349 ( .A(n8957), .ZN(n8959) );
  NOR2_X1 U10350 ( .A1(n8959), .A2(n8958), .ZN(n8963) );
  XNOR2_X1 U10351 ( .A(n8961), .B(n8960), .ZN(n8962) );
  XNOR2_X1 U10352 ( .A(n8963), .B(n8962), .ZN(n8970) );
  OAI21_X1 U10353 ( .B1(n9115), .B2(n9037), .A(n8964), .ZN(n8967) );
  OAI22_X1 U10354 ( .A1(n9129), .A2(n8965), .B1(n9018), .B2(n9126), .ZN(n8966)
         );
  AOI211_X1 U10355 ( .C1(n8968), .C2(n9082), .A(n8967), .B(n8966), .ZN(n8969)
         );
  OAI21_X1 U10356 ( .B1(n8970), .B2(n9122), .A(n8969), .ZN(P1_U3215) );
  OR2_X1 U10357 ( .A1(n8971), .A2(n9052), .ZN(n8978) );
  INV_X1 U10358 ( .A(n8974), .ZN(n8976) );
  OAI21_X2 U10359 ( .B1(n9006), .B2(n8976), .A(n8975), .ZN(n9074) );
  INV_X1 U10360 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8979) );
  OAI22_X1 U10361 ( .A1(n9115), .A2(n9592), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8979), .ZN(n8981) );
  OAI22_X1 U10362 ( .A1(n9126), .A2(n9626), .B1(n9596), .B2(n9129), .ZN(n8980)
         );
  AOI211_X1 U10363 ( .C1(n9757), .C2(n9082), .A(n8981), .B(n8980), .ZN(n8982)
         );
  OAI21_X1 U10364 ( .B1(n8983), .B2(n9122), .A(n8982), .ZN(P1_U3216) );
  AND2_X1 U10365 ( .A1(n8984), .A2(n9085), .ZN(n8986) );
  OAI21_X1 U10366 ( .B1(n8987), .B2(n8986), .A(n8985), .ZN(n8988) );
  NAND2_X1 U10367 ( .A1(n8988), .A2(n9113), .ZN(n8994) );
  OAI22_X1 U10368 ( .A1(n9129), .A2(n8990), .B1(n8989), .B2(n9115), .ZN(n8991)
         );
  AOI211_X1 U10369 ( .C1(n9105), .C2(n9407), .A(n8992), .B(n8991), .ZN(n8993)
         );
  OAI211_X1 U10370 ( .C1(n9970), .C2(n9135), .A(n8994), .B(n8993), .ZN(
        P1_U3217) );
  INV_X1 U10371 ( .A(n8995), .ZN(n8998) );
  NOR3_X1 U10372 ( .A1(n9097), .A2(n9101), .A3(n8996), .ZN(n8997) );
  OAI21_X1 U10373 ( .B1(n8998), .B2(n8997), .A(n9113), .ZN(n9001) );
  AND2_X1 U10374 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9499) );
  OAI22_X1 U10375 ( .A1(n9129), .A2(n9656), .B1(n9664), .B2(n9126), .ZN(n8999)
         );
  AOI211_X1 U10376 ( .C1(n9132), .C2(n9401), .A(n9499), .B(n8999), .ZN(n9000)
         );
  OAI211_X1 U10377 ( .C1(n9655), .C2(n9135), .A(n9001), .B(n9000), .ZN(
        P1_U3219) );
  AOI21_X1 U10378 ( .B1(n9002), .B2(n9004), .A(n9003), .ZN(n9005) );
  OR3_X1 U10379 ( .A1(n9006), .A2(n9005), .A3(n9122), .ZN(n9010) );
  NOR2_X1 U10380 ( .A1(n9126), .A2(n9663), .ZN(n9008) );
  OAI22_X1 U10381 ( .A1(n9129), .A2(n9629), .B1(n9626), .B2(n9115), .ZN(n9007)
         );
  AOI211_X1 U10382 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n9008), 
        .B(n9007), .ZN(n9009) );
  OAI211_X1 U10383 ( .C1(n9633), .C2(n9135), .A(n9010), .B(n9009), .ZN(
        P1_U3223) );
  INV_X1 U10384 ( .A(n9011), .ZN(n9089) );
  INV_X1 U10385 ( .A(n9012), .ZN(n9014) );
  NOR3_X1 U10386 ( .A1(n9089), .A2(n9014), .A3(n9013), .ZN(n9017) );
  INV_X1 U10387 ( .A(n9015), .ZN(n9016) );
  OAI21_X1 U10388 ( .B1(n9017), .B2(n9016), .A(n9113), .ZN(n9023) );
  OAI22_X1 U10389 ( .A1(n9129), .A2(n9019), .B1(n9018), .B2(n9115), .ZN(n9020)
         );
  AOI211_X1 U10390 ( .C1(n9105), .C2(n9405), .A(n9021), .B(n9020), .ZN(n9022)
         );
  OAI211_X1 U10391 ( .C1(n9985), .C2(n9135), .A(n9023), .B(n9022), .ZN(
        P1_U3224) );
  AOI21_X1 U10392 ( .B1(n9024), .B2(n4394), .A(n9111), .ZN(n9029) );
  OAI22_X1 U10393 ( .A1(n9115), .A2(n9564), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9025), .ZN(n9027) );
  OAI22_X1 U10394 ( .A1(n9129), .A2(n9557), .B1(n9592), .B2(n9126), .ZN(n9026)
         );
  AOI211_X1 U10395 ( .C1(n9746), .C2(n9082), .A(n9027), .B(n9026), .ZN(n9028)
         );
  OAI21_X1 U10396 ( .B1(n9029), .B2(n9122), .A(n9028), .ZN(P1_U3225) );
  INV_X1 U10397 ( .A(n9030), .ZN(n9035) );
  AOI21_X1 U10398 ( .B1(n9031), .B2(n9032), .A(n9033), .ZN(n9034) );
  OAI21_X1 U10399 ( .B1(n9035), .B2(n9034), .A(n9113), .ZN(n9040) );
  INV_X1 U10400 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9036) );
  NOR2_X1 U10401 ( .A1(n9036), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9446) );
  OAI22_X1 U10402 ( .A1(n9129), .A2(n9711), .B1(n9037), .B2(n9126), .ZN(n9038)
         );
  AOI211_X1 U10403 ( .C1(n9132), .C2(n9703), .A(n9446), .B(n9038), .ZN(n9039)
         );
  OAI211_X1 U10404 ( .C1(n9819), .C2(n9135), .A(n9040), .B(n9039), .ZN(
        P1_U3226) );
  OAI21_X1 U10405 ( .B1(n9043), .B2(n9042), .A(n9041), .ZN(n9044) );
  NAND2_X1 U10406 ( .A1(n9044), .A2(n9113), .ZN(n9050) );
  NOR2_X1 U10407 ( .A1(n9045), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9460) );
  OAI22_X1 U10408 ( .A1(n9129), .A2(n9047), .B1(n9046), .B2(n9126), .ZN(n9048)
         );
  AOI211_X1 U10409 ( .C1(n9132), .C2(n9689), .A(n9460), .B(n9048), .ZN(n9049)
         );
  OAI211_X1 U10410 ( .C1(n9812), .C2(n9135), .A(n9050), .B(n9049), .ZN(
        P1_U3228) );
  INV_X1 U10411 ( .A(n9752), .ZN(n9583) );
  NOR2_X1 U10412 ( .A1(n9115), .A2(n9544), .ZN(n9055) );
  OAI22_X1 U10413 ( .A1(n9126), .A2(n9079), .B1(n9129), .B2(n9579), .ZN(n9054)
         );
  AOI211_X1 U10414 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n9055), 
        .B(n9054), .ZN(n9056) );
  OAI211_X1 U10415 ( .C1(n9583), .C2(n9135), .A(n9057), .B(n9056), .ZN(
        P1_U3229) );
  INV_X1 U10416 ( .A(n9772), .ZN(n9649) );
  OAI21_X1 U10417 ( .B1(n9059), .B2(n9058), .A(n9002), .ZN(n9060) );
  NAND2_X1 U10418 ( .A1(n9060), .A2(n9113), .ZN(n9064) );
  NOR2_X1 U10419 ( .A1(n9115), .A2(n6260), .ZN(n9062) );
  OAI22_X1 U10420 ( .A1(n9129), .A2(n9645), .B1(n9643), .B2(n9126), .ZN(n9061)
         );
  AOI211_X1 U10421 ( .C1(P1_REG3_REG_20__SCAN_IN), .C2(P1_U3086), .A(n9062), 
        .B(n9061), .ZN(n9063) );
  OAI211_X1 U10422 ( .C1(n9649), .C2(n9135), .A(n9064), .B(n9063), .ZN(
        P1_U3233) );
  OAI21_X1 U10423 ( .B1(n9066), .B2(n9065), .A(n8957), .ZN(n9067) );
  NAND2_X1 U10424 ( .A1(n9067), .A2(n9113), .ZN(n9072) );
  OAI22_X1 U10425 ( .A1(n9129), .A2(n9068), .B1(n9091), .B2(n9126), .ZN(n9069)
         );
  AOI211_X1 U10426 ( .C1(n9132), .C2(n9402), .A(n9070), .B(n9069), .ZN(n9071)
         );
  OAI211_X1 U10427 ( .C1(n9991), .C2(n9135), .A(n9072), .B(n9071), .ZN(
        P1_U3234) );
  INV_X1 U10428 ( .A(n9073), .ZN(n9075) );
  NAND2_X1 U10429 ( .A1(n9075), .A2(n9074), .ZN(n9077) );
  XNOR2_X1 U10430 ( .A(n9077), .B(n9076), .ZN(n9084) );
  OAI22_X1 U10431 ( .A1(n9126), .A2(n6260), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9078), .ZN(n9081) );
  OAI22_X1 U10432 ( .A1(n9129), .A2(n9607), .B1(n9079), .B2(n9115), .ZN(n9080)
         );
  AOI211_X1 U10433 ( .C1(n9762), .C2(n9082), .A(n9081), .B(n9080), .ZN(n9083)
         );
  OAI21_X1 U10434 ( .B1(n9084), .B2(n9122), .A(n9083), .ZN(P1_U3235) );
  INV_X1 U10435 ( .A(n8985), .ZN(n9088) );
  INV_X1 U10436 ( .A(n9085), .ZN(n9087) );
  NOR3_X1 U10437 ( .A1(n9088), .A2(n9087), .A3(n9086), .ZN(n9090) );
  OAI21_X1 U10438 ( .B1(n9090), .B2(n9089), .A(n9113), .ZN(n9096) );
  OAI22_X1 U10439 ( .A1(n9129), .A2(n9092), .B1(n9091), .B2(n9115), .ZN(n9093)
         );
  AOI211_X1 U10440 ( .C1(n9105), .C2(n9406), .A(n9094), .B(n9093), .ZN(n9095)
         );
  OAI211_X1 U10441 ( .C1(n9977), .C2(n9135), .A(n9096), .B(n9095), .ZN(
        P1_U3236) );
  INV_X1 U10442 ( .A(n9097), .ZN(n9102) );
  OAI21_X1 U10443 ( .B1(n9099), .B2(n9101), .A(n9098), .ZN(n9100) );
  OAI21_X1 U10444 ( .B1(n9102), .B2(n9101), .A(n9100), .ZN(n9103) );
  NAND2_X1 U10445 ( .A1(n9103), .A2(n9113), .ZN(n9107) );
  AND2_X1 U10446 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9477) );
  OAI22_X1 U10447 ( .A1(n9129), .A2(n9671), .B1(n9643), .B2(n9115), .ZN(n9104)
         );
  AOI211_X1 U10448 ( .C1(n9105), .C2(n9703), .A(n9477), .B(n9104), .ZN(n9106)
         );
  OAI211_X1 U10449 ( .C1(n4786), .C2(n9135), .A(n9107), .B(n9106), .ZN(
        P1_U3238) );
  INV_X1 U10450 ( .A(n9108), .ZN(n9114) );
  OAI21_X1 U10451 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(n9112) );
  NAND3_X1 U10452 ( .A1(n9114), .A2(n9113), .A3(n9112), .ZN(n9119) );
  NOR2_X1 U10453 ( .A1(n9126), .A2(n9544), .ZN(n9117) );
  OAI22_X1 U10454 ( .A1(n9129), .A2(n9547), .B1(n9543), .B2(n9115), .ZN(n9116)
         );
  AOI211_X1 U10455 ( .C1(P1_REG3_REG_26__SCAN_IN), .C2(P1_U3086), .A(n9117), 
        .B(n9116), .ZN(n9118) );
  OAI211_X1 U10456 ( .C1(n4780), .C2(n9135), .A(n9119), .B(n9118), .ZN(
        P1_U3240) );
  INV_X1 U10457 ( .A(n9032), .ZN(n9125) );
  AOI21_X1 U10458 ( .B1(n9121), .B2(n9032), .A(n9120), .ZN(n9123) );
  NOR2_X1 U10459 ( .A1(n9123), .A2(n9122), .ZN(n9124) );
  OAI21_X1 U10460 ( .B1(n9125), .B2(n9031), .A(n9124), .ZN(n9134) );
  OAI22_X1 U10461 ( .A1(n9129), .A2(n9128), .B1(n9127), .B2(n9126), .ZN(n9130)
         );
  AOI211_X1 U10462 ( .C1(n9132), .C2(n9690), .A(n9131), .B(n9130), .ZN(n9133)
         );
  OAI211_X1 U10463 ( .C1(n9825), .C2(n9135), .A(n9134), .B(n9133), .ZN(
        P1_U3241) );
  OR2_X1 U10464 ( .A1(n9724), .A2(n9507), .ZN(n9141) );
  NAND2_X1 U10465 ( .A1(n9138), .A2(n9137), .ZN(n9140) );
  NAND2_X1 U10466 ( .A1(n5060), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9139) );
  OR2_X1 U10467 ( .A1(n9503), .A2(n9243), .ZN(n9368) );
  NAND2_X1 U10468 ( .A1(n9141), .A2(n9368), .ZN(n9238) );
  NAND2_X1 U10469 ( .A1(n9724), .A2(n9507), .ZN(n9385) );
  NAND2_X1 U10470 ( .A1(n9336), .A2(n9142), .ZN(n9245) );
  INV_X1 U10471 ( .A(n9245), .ZN(n9169) );
  NAND2_X1 U10472 ( .A1(n9335), .A2(n9143), .ZN(n9246) );
  INV_X1 U10473 ( .A(n9246), .ZN(n9168) );
  INV_X1 U10474 ( .A(n9144), .ZN(n9660) );
  INV_X1 U10475 ( .A(n9145), .ZN(n9155) );
  INV_X1 U10476 ( .A(n9146), .ZN(n9154) );
  NOR2_X1 U10477 ( .A1(n6941), .A2(n9147), .ZN(n9150) );
  NAND4_X1 U10478 ( .A1(n9150), .A2(n9149), .A3(n9148), .A4(n9204), .ZN(n9152)
         );
  NOR3_X1 U10479 ( .A1(n9152), .A2(n9887), .A3(n9151), .ZN(n9153) );
  NAND3_X1 U10480 ( .A1(n9155), .A2(n9154), .A3(n9153), .ZN(n9156) );
  NOR2_X1 U10481 ( .A1(n9156), .A2(n9214), .ZN(n9157) );
  NAND4_X1 U10482 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n9161)
         );
  NOR2_X1 U10483 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  NAND3_X1 U10484 ( .A1(n9707), .A2(n9298), .A3(n9163), .ZN(n9164) );
  OR3_X1 U10485 ( .A1(n9165), .A2(n9684), .A3(n9164), .ZN(n9166) );
  NOR3_X1 U10486 ( .A1(n9640), .A2(n9660), .A3(n9166), .ZN(n9167) );
  XNOR2_X1 U10487 ( .A(n9767), .B(n9614), .ZN(n9623) );
  NAND4_X1 U10488 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9623), .ZN(n9170)
         );
  NOR2_X1 U10489 ( .A1(n9571), .A2(n9170), .ZN(n9171) );
  NAND2_X1 U10490 ( .A1(n9553), .A2(n9171), .ZN(n9172) );
  OR4_X1 U10491 ( .A1(n9356), .A2(n9529), .A3(n9541), .A4(n9172), .ZN(n9173)
         );
  NOR2_X1 U10492 ( .A1(n9362), .A2(n9173), .ZN(n9174) );
  NAND2_X1 U10493 ( .A1(n9503), .A2(n9243), .ZN(n9184) );
  NAND3_X1 U10494 ( .A1(n9385), .A2(n9174), .A3(n9184), .ZN(n9175) );
  OR2_X1 U10495 ( .A1(n9238), .A2(n9175), .ZN(n9193) );
  INV_X1 U10496 ( .A(n9193), .ZN(n9196) );
  NOR2_X1 U10497 ( .A1(n9384), .A2(n9197), .ZN(n9374) );
  NAND2_X1 U10498 ( .A1(n9363), .A2(n9358), .ZN(n9187) );
  AND2_X1 U10499 ( .A1(n9354), .A2(n9349), .ZN(n9198) );
  INV_X1 U10500 ( .A(n9341), .ZN(n9176) );
  NOR3_X1 U10501 ( .A1(n9176), .A2(n9247), .A3(n9246), .ZN(n9181) );
  NAND2_X1 U10502 ( .A1(n9245), .A2(n9335), .ZN(n9177) );
  NAND2_X1 U10503 ( .A1(n9177), .A2(n9340), .ZN(n9178) );
  NAND2_X1 U10504 ( .A1(n9178), .A2(n9341), .ZN(n9179) );
  NAND2_X1 U10505 ( .A1(n9537), .A2(n9179), .ZN(n9186) );
  AND2_X1 U10506 ( .A1(n9180), .A2(n9347), .ZN(n9345) );
  OAI21_X1 U10507 ( .B1(n9181), .B2(n9186), .A(n9345), .ZN(n9183) );
  NAND2_X1 U10508 ( .A1(n9359), .A2(n9182), .ZN(n9352) );
  AOI21_X1 U10509 ( .B1(n9198), .B2(n9183), .A(n9352), .ZN(n9185) );
  OAI211_X1 U10510 ( .C1(n9187), .C2(n9185), .A(n9364), .B(n9184), .ZN(n9235)
         );
  NOR2_X1 U10511 ( .A1(n9187), .A2(n9186), .ZN(n9237) );
  AND3_X1 U10512 ( .A1(n9237), .A2(n9198), .A3(n9188), .ZN(n9189) );
  AOI211_X1 U10513 ( .C1(n9724), .C2(n9503), .A(n9235), .B(n9189), .ZN(n9191)
         );
  AOI21_X1 U10514 ( .B1(n9507), .B2(n9368), .A(n9724), .ZN(n9190) );
  OAI21_X1 U10515 ( .B1(n9191), .B2(n9190), .A(n9385), .ZN(n9195) );
  INV_X1 U10516 ( .A(n9197), .ZN(n9192) );
  NAND2_X1 U10517 ( .A1(n9496), .A2(n9197), .ZN(n9241) );
  INV_X1 U10518 ( .A(n9198), .ZN(n9234) );
  AND2_X1 U10519 ( .A1(n9312), .A2(n9308), .ZN(n9324) );
  INV_X1 U10520 ( .A(n9249), .ZN(n9212) );
  INV_X1 U10521 ( .A(n9199), .ZN(n9200) );
  OAI21_X1 U10522 ( .B1(n9202), .B2(n9201), .A(n9200), .ZN(n9203) );
  AOI211_X1 U10523 ( .C1(n9205), .C2(n9413), .A(n9204), .B(n9203), .ZN(n9209)
         );
  INV_X1 U10524 ( .A(n9206), .ZN(n9208) );
  NAND3_X1 U10525 ( .A1(n9209), .A2(n9208), .A3(n9207), .ZN(n9211) );
  INV_X1 U10526 ( .A(n9251), .ZN(n9210) );
  AOI21_X1 U10527 ( .B1(n9212), .B2(n9211), .A(n9210), .ZN(n9215) );
  OAI21_X1 U10528 ( .B1(n9215), .B2(n9214), .A(n9213), .ZN(n9221) );
  NAND2_X1 U10529 ( .A1(n9283), .A2(n9278), .ZN(n9218) );
  INV_X1 U10530 ( .A(n9279), .ZN(n9216) );
  NOR2_X1 U10531 ( .A1(n9218), .A2(n9216), .ZN(n9272) );
  INV_X1 U10532 ( .A(n9272), .ZN(n9220) );
  AND2_X1 U10533 ( .A1(n9281), .A2(n9276), .ZN(n9217) );
  OAI21_X1 U10534 ( .B1(n9218), .B2(n9217), .A(n9282), .ZN(n9271) );
  INV_X1 U10535 ( .A(n9271), .ZN(n9219) );
  OAI211_X1 U10536 ( .C1(n9221), .C2(n9220), .A(n9219), .B(n9288), .ZN(n9222)
         );
  NAND3_X1 U10537 ( .A1(n9222), .A2(n9289), .A3(n9299), .ZN(n9226) );
  NAND2_X1 U10538 ( .A1(n9301), .A2(n9223), .ZN(n9293) );
  INV_X1 U10539 ( .A(n9293), .ZN(n9225) );
  INV_X1 U10540 ( .A(n9300), .ZN(n9224) );
  AOI21_X1 U10541 ( .B1(n9226), .B2(n9225), .A(n9224), .ZN(n9227) );
  AND2_X1 U10542 ( .A1(n9229), .A2(n9674), .ZN(n9309) );
  OAI211_X1 U10543 ( .C1(n9228), .C2(n9227), .A(n9309), .B(n9304), .ZN(n9231)
         );
  OR2_X1 U10544 ( .A1(n9777), .A2(n9643), .ZN(n9315) );
  AND2_X1 U10545 ( .A1(n9315), .A2(n9229), .ZN(n9326) );
  INV_X1 U10546 ( .A(n9326), .ZN(n9230) );
  AOI21_X1 U10547 ( .B1(n9324), .B2(n9231), .A(n9230), .ZN(n9232) );
  OAI211_X1 U10548 ( .C1(n9311), .C2(n9232), .A(n9319), .B(n9321), .ZN(n9233)
         );
  NOR2_X1 U10549 ( .A1(n9234), .A2(n9233), .ZN(n9236) );
  AOI21_X1 U10550 ( .B1(n9237), .B2(n9236), .A(n9235), .ZN(n9239) );
  OAI21_X1 U10551 ( .B1(n9239), .B2(n9238), .A(n9385), .ZN(n9240) );
  MUX2_X1 U10552 ( .A(n9242), .B(n9241), .S(n9240), .Z(n9378) );
  INV_X1 U10553 ( .A(n9243), .ZN(n9396) );
  INV_X1 U10554 ( .A(n9385), .ZN(n9244) );
  AOI21_X1 U10555 ( .B1(n9507), .B2(n9396), .A(n9244), .ZN(n9373) );
  MUX2_X1 U10556 ( .A(n9246), .B(n9245), .S(n9369), .Z(n9339) );
  NAND2_X1 U10557 ( .A1(n9247), .A2(n9369), .ZN(n9248) );
  AND2_X1 U10558 ( .A1(n9612), .A2(n9248), .ZN(n9334) );
  AND2_X1 U10559 ( .A1(n9300), .A2(n9369), .ZN(n9297) );
  NAND3_X1 U10560 ( .A1(n9249), .A2(n9251), .A3(n9257), .ZN(n9250) );
  NAND2_X1 U10561 ( .A1(n9252), .A2(n9251), .ZN(n9255) );
  NAND3_X1 U10562 ( .A1(n9255), .A2(n9254), .A3(n9253), .ZN(n9258) );
  INV_X1 U10563 ( .A(n9839), .ZN(n9256) );
  AOI21_X1 U10564 ( .B1(n9258), .B2(n9257), .A(n9256), .ZN(n9259) );
  AND2_X1 U10565 ( .A1(n9843), .A2(n9260), .ZN(n9261) );
  MUX2_X1 U10566 ( .A(n9262), .B(n9261), .S(n9369), .Z(n9263) );
  NAND2_X1 U10567 ( .A1(n9270), .A2(n9264), .ZN(n9266) );
  MUX2_X1 U10568 ( .A(n9266), .B(n9265), .S(n9383), .Z(n9267) );
  INV_X1 U10569 ( .A(n9267), .ZN(n9268) );
  NAND2_X1 U10570 ( .A1(n9269), .A2(n9268), .ZN(n9275) );
  NAND2_X1 U10571 ( .A1(n9275), .A2(n9270), .ZN(n9273) );
  AOI21_X1 U10572 ( .B1(n9273), .B2(n9272), .A(n9271), .ZN(n9287) );
  NAND2_X1 U10573 ( .A1(n9275), .A2(n9274), .ZN(n9277) );
  NAND2_X1 U10574 ( .A1(n9277), .A2(n9276), .ZN(n9280) );
  NAND3_X1 U10575 ( .A1(n9280), .A2(n9279), .A3(n9278), .ZN(n9285) );
  AND2_X1 U10576 ( .A1(n9282), .A2(n9281), .ZN(n9284) );
  AOI21_X1 U10577 ( .B1(n9285), .B2(n9284), .A(n6285), .ZN(n9286) );
  MUX2_X1 U10578 ( .A(n9287), .B(n9286), .S(n9369), .Z(n9292) );
  MUX2_X1 U10579 ( .A(n9289), .B(n9288), .S(n9383), .Z(n9290) );
  OAI211_X1 U10580 ( .C1(n9292), .C2(n9291), .A(n4663), .B(n9290), .ZN(n9295)
         );
  NAND2_X1 U10581 ( .A1(n9293), .A2(n9369), .ZN(n9294) );
  NAND2_X1 U10582 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  OAI21_X1 U10583 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9303) );
  NAND2_X1 U10584 ( .A1(n9300), .A2(n9299), .ZN(n9302) );
  AND2_X1 U10585 ( .A1(n9674), .A2(n9304), .ZN(n9305) );
  MUX2_X1 U10586 ( .A(n9306), .B(n9305), .S(n9383), .Z(n9307) );
  INV_X1 U10587 ( .A(n9308), .ZN(n9310) );
  OAI21_X1 U10588 ( .B1(n9325), .B2(n9310), .A(n9309), .ZN(n9313) );
  NAND3_X1 U10589 ( .A1(n9313), .A2(n9312), .A3(n4676), .ZN(n9320) );
  NAND2_X1 U10590 ( .A1(n9621), .A2(n9655), .ZN(n9314) );
  NAND2_X1 U10591 ( .A1(n9314), .A2(n9383), .ZN(n9316) );
  NAND3_X1 U10592 ( .A1(n9316), .A2(n9321), .A3(n9315), .ZN(n9318) );
  NAND3_X1 U10593 ( .A1(n9621), .A2(n9383), .A3(n9678), .ZN(n9317) );
  NAND2_X1 U10594 ( .A1(n9318), .A2(n9317), .ZN(n9328) );
  NAND4_X1 U10595 ( .A1(n9320), .A2(n9369), .A3(n9328), .A4(n9319), .ZN(n9333)
         );
  OAI21_X1 U10596 ( .B1(n9321), .B2(n6260), .A(n9767), .ZN(n9323) );
  NAND2_X1 U10597 ( .A1(n9321), .A2(n6260), .ZN(n9322) );
  NAND3_X1 U10598 ( .A1(n9323), .A2(n9383), .A3(n9322), .ZN(n9332) );
  NAND2_X1 U10599 ( .A1(n9327), .A2(n9326), .ZN(n9330) );
  NAND4_X1 U10600 ( .A1(n9330), .A2(n9383), .A3(n9329), .A4(n9328), .ZN(n9331)
         );
  AND4_X1 U10601 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n9338)
         );
  MUX2_X1 U10602 ( .A(n9336), .B(n9335), .S(n9369), .Z(n9337) );
  OAI211_X1 U10603 ( .C1(n9339), .C2(n9338), .A(n4644), .B(n9337), .ZN(n9343)
         );
  MUX2_X1 U10604 ( .A(n9341), .B(n9340), .S(n9369), .Z(n9342) );
  NAND2_X1 U10605 ( .A1(n9348), .A2(n9537), .ZN(n9346) );
  INV_X1 U10606 ( .A(n9349), .ZN(n9344) );
  AOI21_X1 U10607 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9351) );
  INV_X1 U10608 ( .A(n9352), .ZN(n9353) );
  MUX2_X1 U10609 ( .A(n9354), .B(n9353), .S(n9369), .Z(n9355) );
  OAI211_X1 U10610 ( .C1(n9357), .C2(n9356), .A(n9355), .B(n9358), .ZN(n9361)
         );
  MUX2_X1 U10611 ( .A(n9359), .B(n9358), .S(n9369), .Z(n9360) );
  MUX2_X1 U10612 ( .A(n9364), .B(n9363), .S(n9383), .Z(n9365) );
  MUX2_X1 U10613 ( .A(n9366), .B(n9369), .S(n9503), .Z(n9372) );
  INV_X1 U10614 ( .A(n9724), .ZN(n9371) );
  OAI211_X1 U10615 ( .C1(n9369), .C2(n9368), .A(n9367), .B(n9507), .ZN(n9370)
         );
  AOI22_X1 U10616 ( .A1(n9373), .A2(n9372), .B1(n9371), .B2(n9370), .ZN(n9392)
         );
  OAI211_X1 U10617 ( .C1(n9392), .C2(n9376), .A(n9375), .B(n9374), .ZN(n9377)
         );
  NAND3_X1 U10618 ( .A1(n9381), .A2(n9380), .A3(n9379), .ZN(n9382) );
  OAI211_X1 U10619 ( .C1(n9388), .C2(n9387), .A(n9382), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9394) );
  NOR3_X1 U10620 ( .A1(n9724), .A2(n9507), .A3(n9383), .ZN(n9391) );
  NOR2_X1 U10621 ( .A1(n9385), .A2(n9384), .ZN(n9389) );
  NOR4_X1 U10622 ( .A1(n9389), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n9390)
         );
  OAI21_X1 U10623 ( .B1(n9392), .B2(n9391), .A(n9390), .ZN(n9393) );
  NAND3_X1 U10624 ( .A1(n9395), .A2(n9394), .A3(n9393), .ZN(P1_U3242) );
  MUX2_X1 U10625 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9396), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10626 ( .A(n9397), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9412), .Z(
        P1_U3581) );
  MUX2_X1 U10627 ( .A(n9398), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9412), .Z(
        P1_U3580) );
  MUX2_X1 U10628 ( .A(n9574), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9412), .Z(
        P1_U3579) );
  MUX2_X1 U10629 ( .A(n9399), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9412), .Z(
        P1_U3578) );
  MUX2_X1 U10630 ( .A(n9615), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9412), .Z(
        P1_U3577) );
  MUX2_X1 U10631 ( .A(n9400), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9412), .Z(
        P1_U3576) );
  MUX2_X1 U10632 ( .A(n9614), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9412), .Z(
        P1_U3575) );
  MUX2_X1 U10633 ( .A(n9401), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9412), .Z(
        P1_U3574) );
  MUX2_X1 U10634 ( .A(n9678), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9412), .Z(
        P1_U3573) );
  MUX2_X1 U10635 ( .A(n9689), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9412), .Z(
        P1_U3572) );
  MUX2_X1 U10636 ( .A(n9703), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9412), .Z(
        P1_U3571) );
  MUX2_X1 U10637 ( .A(n9690), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9412), .Z(
        P1_U3570) );
  MUX2_X1 U10638 ( .A(n9702), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9412), .Z(
        P1_U3569) );
  MUX2_X1 U10639 ( .A(n9402), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9412), .Z(
        P1_U3568) );
  MUX2_X1 U10640 ( .A(n9403), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9412), .Z(
        P1_U3567) );
  MUX2_X1 U10641 ( .A(n9404), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9412), .Z(
        P1_U3566) );
  MUX2_X1 U10642 ( .A(n9405), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9412), .Z(
        P1_U3565) );
  MUX2_X1 U10643 ( .A(n9406), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9412), .Z(
        P1_U3564) );
  MUX2_X1 U10644 ( .A(n9407), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9412), .Z(
        P1_U3563) );
  MUX2_X1 U10645 ( .A(n9408), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9412), .Z(
        P1_U3562) );
  MUX2_X1 U10646 ( .A(n9861), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9412), .Z(
        P1_U3561) );
  MUX2_X1 U10647 ( .A(n9409), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9412), .Z(
        P1_U3560) );
  MUX2_X1 U10648 ( .A(n9880), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9412), .Z(
        P1_U3559) );
  MUX2_X1 U10649 ( .A(n9410), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9412), .Z(
        P1_U3558) );
  MUX2_X1 U10650 ( .A(n9878), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9412), .Z(
        P1_U3557) );
  MUX2_X1 U10651 ( .A(n9411), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9412), .Z(
        P1_U3556) );
  MUX2_X1 U10652 ( .A(n9413), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9412), .Z(
        P1_U3555) );
  INV_X1 U10653 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9415) );
  OAI22_X1 U10654 ( .A1(n9502), .A2(n9415), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9414), .ZN(n9416) );
  AOI21_X1 U10655 ( .B1(n9418), .B2(n9417), .A(n9416), .ZN(n9428) );
  AOI211_X1 U10656 ( .C1(n9421), .C2(n9420), .A(n9419), .B(n9491), .ZN(n9426)
         );
  AOI211_X1 U10657 ( .C1(n9424), .C2(n9423), .A(n9422), .B(n9484), .ZN(n9425)
         );
  NOR2_X1 U10658 ( .A1(n9426), .A2(n9425), .ZN(n9427) );
  NAND3_X1 U10659 ( .A1(n9429), .A2(n9428), .A3(n9427), .ZN(P1_U3245) );
  MUX2_X1 U10660 ( .A(n5400), .B(P1_REG1_REG_16__SCAN_IN), .S(n9449), .Z(n9435) );
  NAND2_X1 U10661 ( .A1(n9431), .A2(n9430), .ZN(n9433) );
  NAND2_X1 U10662 ( .A1(n9434), .A2(n9435), .ZN(n9453) );
  OAI21_X1 U10663 ( .B1(n9435), .B2(n9434), .A(n9453), .ZN(n9436) );
  NAND2_X1 U10664 ( .A1(n9436), .A2(n9488), .ZN(n9448) );
  NOR2_X1 U10665 ( .A1(n9438), .A2(n9437), .ZN(n9440) );
  NOR2_X1 U10666 ( .A1(n9440), .A2(n9439), .ZN(n9444) );
  INV_X1 U10667 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9712) );
  OR2_X1 U10668 ( .A1(n9449), .A2(n9712), .ZN(n9455) );
  NAND2_X1 U10669 ( .A1(n9449), .A2(n9712), .ZN(n9441) );
  NAND2_X1 U10670 ( .A1(n9455), .A2(n9441), .ZN(n9443) );
  INV_X1 U10671 ( .A(n9456), .ZN(n9442) );
  AOI211_X1 U10672 ( .C1(n9444), .C2(n9443), .A(n9442), .B(n9484), .ZN(n9445)
         );
  AOI211_X1 U10673 ( .C1(n9478), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9446), .B(
        n9445), .ZN(n9447) );
  OAI211_X1 U10674 ( .C1(n9490), .C2(n9449), .A(n9448), .B(n9447), .ZN(
        P1_U3259) );
  NAND2_X1 U10675 ( .A1(n9449), .A2(n5400), .ZN(n9451) );
  MUX2_X1 U10676 ( .A(n9450), .B(P1_REG1_REG_17__SCAN_IN), .S(n9463), .Z(n9452) );
  AOI21_X1 U10677 ( .B1(n9453), .B2(n9451), .A(n9452), .ZN(n9466) );
  AND3_X1 U10678 ( .A1(n9453), .A2(n9452), .A3(n9451), .ZN(n9454) );
  OAI21_X1 U10679 ( .B1(n9466), .B2(n9454), .A(n9488), .ZN(n9462) );
  XNOR2_X1 U10680 ( .A(n9463), .B(n9469), .ZN(n9457) );
  AOI221_X1 U10681 ( .B1(n9458), .B2(n9472), .C1(n9457), .C2(n9472), .A(n9484), 
        .ZN(n9459) );
  AOI211_X1 U10682 ( .C1(n9478), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9460), .B(
        n9459), .ZN(n9461) );
  OAI211_X1 U10683 ( .C1(n9490), .C2(n9470), .A(n9462), .B(n9461), .ZN(
        P1_U3260) );
  NOR2_X1 U10684 ( .A1(n9463), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9465) );
  XNOR2_X1 U10685 ( .A(n9486), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9464) );
  NOR3_X1 U10686 ( .A1(n9466), .A2(n9465), .A3(n9464), .ZN(n9485) );
  INV_X1 U10687 ( .A(n9485), .ZN(n9468) );
  OAI21_X1 U10688 ( .B1(n9466), .B2(n9465), .A(n9464), .ZN(n9467) );
  NAND3_X1 U10689 ( .A1(n9468), .A2(n9488), .A3(n9467), .ZN(n9480) );
  NAND2_X1 U10690 ( .A1(n9470), .A2(n9469), .ZN(n9471) );
  MUX2_X1 U10691 ( .A(n9473), .B(P1_REG2_REG_18__SCAN_IN), .S(n9486), .Z(n9474) );
  AOI211_X1 U10692 ( .C1(n9475), .C2(n9474), .A(n9482), .B(n9484), .ZN(n9476)
         );
  AOI211_X1 U10693 ( .C1(n9478), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9477), .B(
        n9476), .ZN(n9479) );
  OAI211_X1 U10694 ( .C1(n9490), .C2(n9481), .A(n9480), .B(n9479), .ZN(
        P1_U3261) );
  XNOR2_X1 U10695 ( .A(n9483), .B(n9657), .ZN(n9489) );
  INV_X1 U10696 ( .A(n9484), .ZN(n9494) );
  AOI21_X1 U10697 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9486), .A(n9485), .ZN(
        n9487) );
  XNOR2_X1 U10698 ( .A(n9487), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9492) );
  AOI22_X1 U10699 ( .A1(n9489), .A2(n9494), .B1(n9488), .B2(n9492), .ZN(n9498)
         );
  INV_X1 U10700 ( .A(n9489), .ZN(n9495) );
  OAI21_X1 U10701 ( .B1(n9492), .B2(n9491), .A(n9490), .ZN(n9493) );
  AOI21_X1 U10702 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9497) );
  MUX2_X1 U10703 ( .A(n9498), .B(n9497), .S(n9496), .Z(n9501) );
  INV_X1 U10704 ( .A(n9499), .ZN(n9500) );
  OAI211_X1 U10705 ( .C1(n4819), .C2(n9502), .A(n9501), .B(n9500), .ZN(
        P1_U3262) );
  NAND2_X1 U10706 ( .A1(n9727), .A2(n9512), .ZN(n9511) );
  XNOR2_X1 U10707 ( .A(n9724), .B(n9511), .ZN(n9504) );
  NAND2_X1 U10708 ( .A1(n9504), .A2(n9890), .ZN(n9723) );
  INV_X1 U10709 ( .A(n9505), .ZN(n9506) );
  NAND2_X1 U10710 ( .A1(n9507), .A2(n9506), .ZN(n9725) );
  OR2_X1 U10711 ( .A1(n4321), .A2(n9725), .ZN(n9513) );
  NAND2_X1 U10712 ( .A1(n4321), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9508) );
  OAI211_X1 U10713 ( .C1(n9724), .C2(n9884), .A(n9513), .B(n9508), .ZN(n9509)
         );
  INV_X1 U10714 ( .A(n9509), .ZN(n9510) );
  OAI21_X1 U10715 ( .B1(n9723), .B2(n9904), .A(n9510), .ZN(P1_U3263) );
  OAI211_X1 U10716 ( .C1(n9727), .C2(n9512), .A(n9890), .B(n9511), .ZN(n9726)
         );
  INV_X1 U10717 ( .A(n9513), .ZN(n9515) );
  NOR2_X1 U10718 ( .A1(n9727), .A2(n9884), .ZN(n9514) );
  AOI211_X1 U10719 ( .C1(n4321), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9515), .B(
        n9514), .ZN(n9516) );
  OAI21_X1 U10720 ( .B1(n9904), .B2(n9726), .A(n9516), .ZN(P1_U3264) );
  OAI21_X1 U10721 ( .B1(n9518), .B2(n9529), .A(n9517), .ZN(n9738) );
  INV_X1 U10722 ( .A(n9519), .ZN(n9522) );
  INV_X1 U10723 ( .A(n9520), .ZN(n9521) );
  INV_X1 U10724 ( .A(n9523), .ZN(n9524) );
  AOI22_X1 U10725 ( .A1(n4321), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9524), .B2(
        n9897), .ZN(n9525) );
  OAI21_X1 U10726 ( .B1(n9526), .B2(n9884), .A(n9525), .ZN(n9534) );
  AOI211_X1 U10727 ( .C1(n9529), .C2(n9528), .A(n9842), .B(n9527), .ZN(n9532)
         );
  OAI22_X1 U10728 ( .A1(n9543), .A2(n9833), .B1(n9530), .B2(n9835), .ZN(n9531)
         );
  NOR2_X1 U10729 ( .A1(n9737), .A2(n4321), .ZN(n9533) );
  AOI211_X1 U10730 ( .C1(n9734), .C2(n9893), .A(n9534), .B(n9533), .ZN(n9535)
         );
  OAI21_X1 U10731 ( .B1(n9709), .B2(n9738), .A(n9535), .ZN(P1_U3265) );
  XNOR2_X1 U10732 ( .A(n9536), .B(n9541), .ZN(n9744) );
  INV_X1 U10733 ( .A(n9561), .ZN(n9538) );
  NAND2_X1 U10734 ( .A1(n9538), .A2(n9537), .ZN(n9540) );
  AOI21_X1 U10735 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9542) );
  OAI222_X1 U10736 ( .A1(n9833), .A2(n9544), .B1(n9835), .B2(n9543), .C1(n9842), .C2(n9542), .ZN(n9740) );
  INV_X1 U10737 ( .A(n9545), .ZN(n9546) );
  AOI211_X1 U10738 ( .C1(n9742), .C2(n9555), .A(n9670), .B(n9546), .ZN(n9741)
         );
  NAND2_X1 U10739 ( .A1(n9741), .A2(n9893), .ZN(n9550) );
  INV_X1 U10740 ( .A(n9547), .ZN(n9548) );
  AOI22_X1 U10741 ( .A1(n4321), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9548), .B2(
        n9897), .ZN(n9549) );
  OAI211_X1 U10742 ( .C1(n4780), .C2(n9884), .A(n9550), .B(n9549), .ZN(n9551)
         );
  AOI21_X1 U10743 ( .B1(n9740), .B2(n9713), .A(n9551), .ZN(n9552) );
  OAI21_X1 U10744 ( .B1(n9744), .B2(n9709), .A(n9552), .ZN(P1_U3267) );
  XNOR2_X1 U10745 ( .A(n9554), .B(n9553), .ZN(n9749) );
  INV_X1 U10746 ( .A(n9555), .ZN(n9556) );
  AOI211_X1 U10747 ( .C1(n9746), .C2(n4784), .A(n9670), .B(n9556), .ZN(n9745)
         );
  INV_X1 U10748 ( .A(n9557), .ZN(n9558) );
  AOI22_X1 U10749 ( .A1(n4321), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9558), .B2(
        n9897), .ZN(n9559) );
  OAI21_X1 U10750 ( .B1(n9560), .B2(n9884), .A(n9559), .ZN(n9568) );
  AOI211_X1 U10751 ( .C1(n9563), .C2(n9562), .A(n9842), .B(n9561), .ZN(n9566)
         );
  OAI22_X1 U10752 ( .A1(n9564), .A2(n9835), .B1(n9592), .B2(n9833), .ZN(n9565)
         );
  NOR2_X1 U10753 ( .A1(n9566), .A2(n9565), .ZN(n9748) );
  NOR2_X1 U10754 ( .A1(n9748), .A2(n4321), .ZN(n9567) );
  AOI211_X1 U10755 ( .C1(n9745), .C2(n9893), .A(n9568), .B(n9567), .ZN(n9569)
         );
  OAI21_X1 U10756 ( .B1(n9749), .B2(n9709), .A(n9569), .ZN(P1_U3268) );
  XNOR2_X1 U10757 ( .A(n9570), .B(n9571), .ZN(n9754) );
  OAI21_X1 U10758 ( .B1(n9588), .B2(n9572), .A(n9571), .ZN(n9573) );
  NAND2_X1 U10759 ( .A1(n9573), .A2(n9876), .ZN(n9576) );
  AOI22_X1 U10760 ( .A1(n9879), .A2(n9574), .B1(n9615), .B2(n9877), .ZN(n9575)
         );
  OAI21_X1 U10761 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9750) );
  AOI211_X1 U10762 ( .C1(n9752), .C2(n9593), .A(n9670), .B(n9578), .ZN(n9751)
         );
  NAND2_X1 U10763 ( .A1(n9751), .A2(n9893), .ZN(n9582) );
  INV_X1 U10764 ( .A(n9579), .ZN(n9580) );
  AOI22_X1 U10765 ( .A1(n4321), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9580), .B2(
        n9897), .ZN(n9581) );
  OAI211_X1 U10766 ( .C1(n9583), .C2(n9884), .A(n9582), .B(n9581), .ZN(n9584)
         );
  AOI21_X1 U10767 ( .B1(n9750), .B2(n9713), .A(n9584), .ZN(n9585) );
  OAI21_X1 U10768 ( .B1(n9754), .B2(n9709), .A(n9585), .ZN(P1_U3269) );
  XNOR2_X1 U10769 ( .A(n9587), .B(n9586), .ZN(n9759) );
  AOI21_X1 U10770 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9591) );
  OAI222_X1 U10771 ( .A1(n9833), .A2(n9626), .B1(n9835), .B2(n9592), .C1(n9842), .C2(n9591), .ZN(n9755) );
  INV_X1 U10772 ( .A(n9604), .ZN(n9595) );
  INV_X1 U10773 ( .A(n9593), .ZN(n9594) );
  AOI211_X1 U10774 ( .C1(n9757), .C2(n9595), .A(n9670), .B(n9594), .ZN(n9756)
         );
  NAND2_X1 U10775 ( .A1(n9756), .A2(n9893), .ZN(n9599) );
  INV_X1 U10776 ( .A(n9596), .ZN(n9597) );
  AOI22_X1 U10777 ( .A1(n4321), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9597), .B2(
        n9897), .ZN(n9598) );
  OAI211_X1 U10778 ( .C1(n9600), .C2(n9884), .A(n9599), .B(n9598), .ZN(n9601)
         );
  AOI21_X1 U10779 ( .B1(n9755), .B2(n9713), .A(n9601), .ZN(n9602) );
  OAI21_X1 U10780 ( .B1(n9759), .B2(n9709), .A(n9602), .ZN(P1_U3270) );
  XNOR2_X1 U10781 ( .A(n9603), .B(n9612), .ZN(n9764) );
  INV_X1 U10782 ( .A(n9627), .ZN(n9605) );
  AOI211_X1 U10783 ( .C1(n9762), .C2(n9605), .A(n9670), .B(n9604), .ZN(n9761)
         );
  NOR2_X1 U10784 ( .A1(n9606), .A2(n9884), .ZN(n9610) );
  OAI22_X1 U10785 ( .A1(n9713), .A2(n9608), .B1(n9607), .B2(n9710), .ZN(n9609)
         );
  AOI211_X1 U10786 ( .C1(n9761), .C2(n9893), .A(n9610), .B(n9609), .ZN(n9619)
         );
  OAI211_X1 U10787 ( .C1(n9613), .C2(n9612), .A(n9611), .B(n9876), .ZN(n9617)
         );
  AOI22_X1 U10788 ( .A1(n9879), .A2(n9615), .B1(n9614), .B2(n9877), .ZN(n9616)
         );
  NAND2_X1 U10789 ( .A1(n9617), .A2(n9616), .ZN(n9760) );
  NAND2_X1 U10790 ( .A1(n9760), .A2(n9713), .ZN(n9618) );
  OAI211_X1 U10791 ( .C1(n9764), .C2(n9709), .A(n9619), .B(n9618), .ZN(
        P1_U3271) );
  XNOR2_X1 U10792 ( .A(n9620), .B(n9623), .ZN(n9769) );
  NOR2_X1 U10793 ( .A1(n9641), .A2(n9640), .ZN(n9639) );
  INV_X1 U10794 ( .A(n9621), .ZN(n9622) );
  NOR2_X1 U10795 ( .A1(n9639), .A2(n9622), .ZN(n9624) );
  XNOR2_X1 U10796 ( .A(n9624), .B(n9623), .ZN(n9625) );
  OAI222_X1 U10797 ( .A1(n9833), .A2(n9663), .B1(n9835), .B2(n9626), .C1(n9842), .C2(n9625), .ZN(n9765) );
  INV_X1 U10798 ( .A(n9644), .ZN(n9628) );
  AOI211_X1 U10799 ( .C1(n9767), .C2(n9628), .A(n9670), .B(n9627), .ZN(n9766)
         );
  NAND2_X1 U10800 ( .A1(n9766), .A2(n9893), .ZN(n9632) );
  INV_X1 U10801 ( .A(n9629), .ZN(n9630) );
  AOI22_X1 U10802 ( .A1(n4321), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9630), .B2(
        n9897), .ZN(n9631) );
  OAI211_X1 U10803 ( .C1(n9633), .C2(n9884), .A(n9632), .B(n9631), .ZN(n9634)
         );
  AOI21_X1 U10804 ( .B1(n9765), .B2(n9713), .A(n9634), .ZN(n9635) );
  OAI21_X1 U10805 ( .B1(n9769), .B2(n9709), .A(n9635), .ZN(P1_U3272) );
  OAI21_X1 U10806 ( .B1(n9637), .B2(n9640), .A(n9636), .ZN(n9638) );
  INV_X1 U10807 ( .A(n9638), .ZN(n9774) );
  AOI21_X1 U10808 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9642) );
  OAI222_X1 U10809 ( .A1(n9833), .A2(n9643), .B1(n9835), .B2(n6260), .C1(n9842), .C2(n9642), .ZN(n9770) );
  AOI211_X1 U10810 ( .C1(n9772), .C2(n9653), .A(n9670), .B(n9644), .ZN(n9771)
         );
  NAND2_X1 U10811 ( .A1(n9771), .A2(n9893), .ZN(n9648) );
  INV_X1 U10812 ( .A(n9645), .ZN(n9646) );
  AOI22_X1 U10813 ( .A1(n4321), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9646), .B2(
        n9897), .ZN(n9647) );
  OAI211_X1 U10814 ( .C1(n9649), .C2(n9884), .A(n9648), .B(n9647), .ZN(n9650)
         );
  AOI21_X1 U10815 ( .B1(n9770), .B2(n9713), .A(n9650), .ZN(n9651) );
  OAI21_X1 U10816 ( .B1(n9774), .B2(n9709), .A(n9651), .ZN(P1_U3273) );
  XNOR2_X1 U10817 ( .A(n9652), .B(n9660), .ZN(n9779) );
  INV_X1 U10818 ( .A(n9653), .ZN(n9654) );
  AOI211_X1 U10819 ( .C1(n9777), .C2(n9668), .A(n9670), .B(n9654), .ZN(n9776)
         );
  NOR2_X1 U10820 ( .A1(n9655), .A2(n9884), .ZN(n9659) );
  OAI22_X1 U10821 ( .A1(n9713), .A2(n9657), .B1(n9656), .B2(n9710), .ZN(n9658)
         );
  AOI211_X1 U10822 ( .C1(n9776), .C2(n9893), .A(n9659), .B(n9658), .ZN(n9666)
         );
  XNOR2_X1 U10823 ( .A(n9661), .B(n9660), .ZN(n9662) );
  OAI222_X1 U10824 ( .A1(n9833), .A2(n9664), .B1(n9835), .B2(n9663), .C1(n9842), .C2(n9662), .ZN(n9775) );
  NAND2_X1 U10825 ( .A1(n9775), .A2(n9713), .ZN(n9665) );
  OAI211_X1 U10826 ( .C1(n9779), .C2(n9709), .A(n9666), .B(n9665), .ZN(
        P1_U3274) );
  XNOR2_X1 U10827 ( .A(n9676), .B(n9667), .ZN(n9784) );
  INV_X1 U10828 ( .A(n9668), .ZN(n9669) );
  AOI211_X1 U10829 ( .C1(n9781), .C2(n9693), .A(n9670), .B(n9669), .ZN(n9780)
         );
  INV_X1 U10830 ( .A(n9671), .ZN(n9672) );
  AOI22_X1 U10831 ( .A1(n4321), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9672), .B2(
        n9897), .ZN(n9673) );
  OAI21_X1 U10832 ( .B1(n4786), .B2(n9884), .A(n9673), .ZN(n9681) );
  AND2_X1 U10833 ( .A1(n9686), .A2(n9674), .ZN(n9677) );
  OAI21_X1 U10834 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9679) );
  AOI222_X1 U10835 ( .A1(n9876), .A2(n9679), .B1(n9703), .B2(n9877), .C1(n9678), .C2(n9879), .ZN(n9783) );
  NOR2_X1 U10836 ( .A1(n9783), .A2(n4321), .ZN(n9680) );
  AOI211_X1 U10837 ( .C1(n9780), .C2(n9893), .A(n9681), .B(n9680), .ZN(n9682)
         );
  OAI21_X1 U10838 ( .B1(n9784), .B2(n9709), .A(n9682), .ZN(P1_U3275) );
  OAI21_X1 U10839 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9815) );
  INV_X1 U10840 ( .A(n9815), .ZN(n9699) );
  OAI211_X1 U10841 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9876), .ZN(n9692)
         );
  AOI22_X1 U10842 ( .A1(n9877), .A2(n9690), .B1(n9689), .B2(n9879), .ZN(n9691)
         );
  NAND2_X1 U10843 ( .A1(n9692), .A2(n9691), .ZN(n9814) );
  OAI211_X1 U10844 ( .C1(n9714), .C2(n9812), .A(n9890), .B(n9693), .ZN(n9811)
         );
  NOR2_X1 U10845 ( .A1(n9811), .A2(n9904), .ZN(n9697) );
  AOI22_X1 U10846 ( .A1(n4321), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9694), .B2(
        n9897), .ZN(n9695) );
  OAI21_X1 U10847 ( .B1(n9812), .B2(n9884), .A(n9695), .ZN(n9696) );
  AOI211_X1 U10848 ( .C1(n9814), .C2(n9713), .A(n9697), .B(n9696), .ZN(n9698)
         );
  OAI21_X1 U10849 ( .B1(n9699), .B2(n9709), .A(n9698), .ZN(P1_U3276) );
  XNOR2_X1 U10850 ( .A(n9700), .B(n9707), .ZN(n9701) );
  NAND2_X1 U10851 ( .A1(n9701), .A2(n9876), .ZN(n9705) );
  AOI22_X1 U10852 ( .A1(n9879), .A2(n9703), .B1(n9702), .B2(n9877), .ZN(n9704)
         );
  NAND2_X1 U10853 ( .A1(n9705), .A2(n9704), .ZN(n9821) );
  INV_X1 U10854 ( .A(n9821), .ZN(n9722) );
  INV_X1 U10855 ( .A(n9706), .ZN(n9817) );
  AND2_X1 U10856 ( .A1(n9708), .A2(n9707), .ZN(n9816) );
  OR3_X1 U10857 ( .A1(n9817), .A2(n9816), .A3(n9709), .ZN(n9721) );
  OAI22_X1 U10858 ( .A1(n9713), .A2(n9712), .B1(n9711), .B2(n9710), .ZN(n9718)
         );
  INV_X1 U10859 ( .A(n9714), .ZN(n9715) );
  OAI211_X1 U10860 ( .C1(n9819), .C2(n9716), .A(n9715), .B(n9890), .ZN(n9818)
         );
  NOR2_X1 U10861 ( .A1(n9818), .A2(n9904), .ZN(n9717) );
  AOI211_X1 U10862 ( .C1(n9901), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9720)
         );
  OAI211_X1 U10863 ( .C1(n4321), .C2(n9722), .A(n9721), .B(n9720), .ZN(
        P1_U3277) );
  OAI211_X1 U10864 ( .C1(n9724), .C2(n9996), .A(n9723), .B(n9725), .ZN(n9785)
         );
  MUX2_X1 U10865 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9785), .S(n10019), .Z(
        P1_U3553) );
  OAI211_X1 U10866 ( .C1(n9727), .C2(n9996), .A(n9726), .B(n9725), .ZN(n9786)
         );
  MUX2_X1 U10867 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9786), .S(n10019), .Z(
        P1_U3552) );
  MUX2_X1 U10868 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9787), .S(n10019), .Z(
        P1_U3551) );
  AOI21_X1 U10869 ( .B1(n9959), .B2(n9735), .A(n9734), .ZN(n9736) );
  OAI211_X1 U10870 ( .C1(n9738), .C2(n9963), .A(n9737), .B(n9736), .ZN(n9788)
         );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9788), .S(n10019), .Z(
        P1_U3550) );
  MUX2_X1 U10872 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9739), .S(n10019), .Z(
        P1_U3549) );
  AOI211_X1 U10873 ( .C1(n9959), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9743)
         );
  OAI21_X1 U10874 ( .B1(n9744), .B2(n9963), .A(n9743), .ZN(n9789) );
  MUX2_X1 U10875 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9789), .S(n10019), .Z(
        P1_U3548) );
  AOI21_X1 U10876 ( .B1(n9959), .B2(n9746), .A(n9745), .ZN(n9747) );
  OAI211_X1 U10877 ( .C1(n9749), .C2(n9963), .A(n9748), .B(n9747), .ZN(n9790)
         );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9790), .S(n10019), .Z(
        P1_U3547) );
  AOI211_X1 U10879 ( .C1(n9959), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9753)
         );
  OAI21_X1 U10880 ( .B1(n9754), .B2(n9963), .A(n9753), .ZN(n9791) );
  MUX2_X1 U10881 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9791), .S(n10019), .Z(
        P1_U3546) );
  AOI211_X1 U10882 ( .C1(n9959), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9758)
         );
  OAI21_X1 U10883 ( .B1(n9759), .B2(n9963), .A(n9758), .ZN(n9792) );
  MUX2_X1 U10884 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9792), .S(n10019), .Z(
        P1_U3545) );
  AOI211_X1 U10885 ( .C1(n9959), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9763)
         );
  OAI21_X1 U10886 ( .B1(n9764), .B2(n9963), .A(n9763), .ZN(n9793) );
  MUX2_X1 U10887 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9793), .S(n10019), .Z(
        P1_U3544) );
  AOI211_X1 U10888 ( .C1(n9959), .C2(n9767), .A(n9766), .B(n9765), .ZN(n9768)
         );
  OAI21_X1 U10889 ( .B1(n9769), .B2(n9963), .A(n9768), .ZN(n9794) );
  MUX2_X1 U10890 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9794), .S(n10019), .Z(
        P1_U3543) );
  AOI211_X1 U10891 ( .C1(n9959), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9773)
         );
  OAI21_X1 U10892 ( .B1(n9774), .B2(n9963), .A(n9773), .ZN(n9795) );
  MUX2_X1 U10893 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9795), .S(n10019), .Z(
        P1_U3542) );
  AOI211_X1 U10894 ( .C1(n9959), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9778)
         );
  OAI21_X1 U10895 ( .B1(n9779), .B2(n9963), .A(n9778), .ZN(n9796) );
  MUX2_X1 U10896 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9796), .S(n10019), .Z(
        P1_U3541) );
  AOI21_X1 U10897 ( .B1(n9959), .B2(n9781), .A(n9780), .ZN(n9782) );
  OAI211_X1 U10898 ( .C1(n9784), .C2(n9963), .A(n9783), .B(n9782), .ZN(n9797)
         );
  MUX2_X1 U10899 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9797), .S(n10019), .Z(
        P1_U3540) );
  MUX2_X1 U10900 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9785), .S(n10004), .Z(
        P1_U3521) );
  MUX2_X1 U10901 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9786), .S(n10004), .Z(
        P1_U3520) );
  MUX2_X1 U10902 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9787), .S(n10004), .Z(
        P1_U3519) );
  MUX2_X1 U10903 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9788), .S(n10004), .Z(
        P1_U3518) );
  MUX2_X1 U10904 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9789), .S(n10004), .Z(
        P1_U3516) );
  MUX2_X1 U10905 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9790), .S(n10004), .Z(
        P1_U3515) );
  MUX2_X1 U10906 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9791), .S(n10004), .Z(
        P1_U3514) );
  MUX2_X1 U10907 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9792), .S(n10004), .Z(
        P1_U3513) );
  MUX2_X1 U10908 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9793), .S(n10004), .Z(
        P1_U3512) );
  MUX2_X1 U10909 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9794), .S(n10004), .Z(
        P1_U3511) );
  MUX2_X1 U10910 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9795), .S(n10004), .Z(
        P1_U3510) );
  MUX2_X1 U10911 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9796), .S(n10004), .Z(
        P1_U3509) );
  MUX2_X1 U10912 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9797), .S(n10004), .Z(
        P1_U3507) );
  NOR4_X1 U10913 ( .A1(n9798), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5288), .A4(
        P1_U3086), .ZN(n9799) );
  AOI21_X1 U10914 ( .B1(n9804), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9799), .ZN(
        n9800) );
  OAI21_X1 U10915 ( .B1(n9801), .B2(n9807), .A(n9800), .ZN(P1_U3324) );
  AOI22_X1 U10916 ( .A1(n4937), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9804), .ZN(n9802) );
  OAI21_X1 U10917 ( .B1(n9803), .B2(n9807), .A(n9802), .ZN(P1_U3325) );
  AOI22_X1 U10918 ( .A1(n9805), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9804), .ZN(n9806) );
  OAI21_X1 U10919 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(P1_U3326) );
  INV_X1 U10920 ( .A(n9809), .ZN(n9810) );
  MUX2_X1 U10921 ( .A(n9810), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U10922 ( .B1(n9812), .B2(n9996), .A(n9811), .ZN(n9813) );
  AOI211_X1 U10923 ( .C1(n9815), .C2(n10000), .A(n9814), .B(n9813), .ZN(n9829)
         );
  AOI22_X1 U10924 ( .A1(n10019), .A2(n9829), .B1(n9450), .B2(n10017), .ZN(
        P1_U3539) );
  NOR3_X1 U10925 ( .A1(n9817), .A2(n9816), .A3(n9963), .ZN(n9822) );
  OAI21_X1 U10926 ( .B1(n9819), .B2(n9996), .A(n9818), .ZN(n9820) );
  NOR3_X1 U10927 ( .A1(n9822), .A2(n9821), .A3(n9820), .ZN(n9830) );
  AOI22_X1 U10928 ( .A1(n10019), .A2(n9830), .B1(n5400), .B2(n10017), .ZN(
        P1_U3538) );
  OAI211_X1 U10929 ( .C1(n9825), .C2(n9996), .A(n9824), .B(n9823), .ZN(n9826)
         );
  AOI21_X1 U10930 ( .B1(n9827), .B2(n10000), .A(n9826), .ZN(n9831) );
  AOI22_X1 U10931 ( .A1(n10019), .A2(n9831), .B1(n5371), .B2(n10017), .ZN(
        P1_U3537) );
  AOI22_X1 U10932 ( .A1(n10004), .A2(n9829), .B1(n9828), .B2(n10002), .ZN(
        P1_U3504) );
  AOI22_X1 U10933 ( .A1(n10004), .A2(n9830), .B1(n5401), .B2(n10002), .ZN(
        P1_U3501) );
  AOI22_X1 U10934 ( .A1(n10004), .A2(n9831), .B1(n5372), .B2(n10002), .ZN(
        P1_U3498) );
  XNOR2_X1 U10935 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10936 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  XNOR2_X1 U10937 ( .A(n9832), .B(n9838), .ZN(n9958) );
  OAI22_X1 U10938 ( .A1(n9836), .A2(n9835), .B1(n9834), .B2(n9833), .ZN(n9846)
         );
  INV_X1 U10939 ( .A(n9837), .ZN(n9844) );
  AOI21_X1 U10940 ( .B1(n9840), .B2(n9839), .A(n4687), .ZN(n9841) );
  AOI211_X1 U10941 ( .C1(n9844), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9845)
         );
  AOI211_X1 U10942 ( .C1(n9847), .C2(n9958), .A(n9846), .B(n9845), .ZN(n9955)
         );
  INV_X1 U10943 ( .A(n9848), .ZN(n9849) );
  AOI22_X1 U10944 ( .A1(n4321), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9849), .B2(
        n9897), .ZN(n9850) );
  OAI21_X1 U10945 ( .B1(n9884), .B2(n9954), .A(n9850), .ZN(n9851) );
  INV_X1 U10946 ( .A(n9851), .ZN(n9858) );
  INV_X1 U10947 ( .A(n9852), .ZN(n9855) );
  INV_X1 U10948 ( .A(n9853), .ZN(n9854) );
  OAI211_X1 U10949 ( .C1(n9954), .C2(n9855), .A(n9854), .B(n9890), .ZN(n9953)
         );
  INV_X1 U10950 ( .A(n9953), .ZN(n9856) );
  AOI22_X1 U10951 ( .A1(n9958), .A2(n9899), .B1(n9893), .B2(n9856), .ZN(n9857)
         );
  OAI211_X1 U10952 ( .C1(n4321), .C2(n9955), .A(n9858), .B(n9857), .ZN(
        P1_U3285) );
  XOR2_X1 U10953 ( .A(n9859), .B(n9867), .Z(n9860) );
  AOI222_X1 U10954 ( .A1(n9861), .A2(n9879), .B1(n9880), .B2(n9877), .C1(n9876), .C2(n9860), .ZN(n9940) );
  INV_X1 U10955 ( .A(n9862), .ZN(n9863) );
  AOI22_X1 U10956 ( .A1(n4321), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9863), .B2(
        n9897), .ZN(n9864) );
  OAI21_X1 U10957 ( .B1(n9884), .B2(n9939), .A(n9864), .ZN(n9865) );
  INV_X1 U10958 ( .A(n9865), .ZN(n9873) );
  XNOR2_X1 U10959 ( .A(n9866), .B(n9867), .ZN(n9943) );
  INV_X1 U10960 ( .A(n9868), .ZN(n9870) );
  OAI211_X1 U10961 ( .C1(n9870), .C2(n9939), .A(n9890), .B(n9869), .ZN(n9938)
         );
  INV_X1 U10962 ( .A(n9938), .ZN(n9871) );
  AOI22_X1 U10963 ( .A1(n9943), .A2(n9894), .B1(n9893), .B2(n9871), .ZN(n9872)
         );
  OAI211_X1 U10964 ( .C1(n4321), .C2(n9940), .A(n9873), .B(n9872), .ZN(
        P1_U3287) );
  XNOR2_X1 U10965 ( .A(n9874), .B(n9887), .ZN(n9875) );
  AOI222_X1 U10966 ( .A1(n9880), .A2(n9879), .B1(n9878), .B2(n9877), .C1(n9876), .C2(n9875), .ZN(n9928) );
  INV_X1 U10967 ( .A(n9881), .ZN(n9882) );
  AOI22_X1 U10968 ( .A1(n4321), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9882), .B2(
        n9897), .ZN(n9883) );
  OAI21_X1 U10969 ( .B1(n9884), .B2(n9927), .A(n9883), .ZN(n9885) );
  INV_X1 U10970 ( .A(n9885), .ZN(n9896) );
  XNOR2_X1 U10971 ( .A(n9886), .B(n9887), .ZN(n9931) );
  INV_X1 U10972 ( .A(n9888), .ZN(n9891) );
  OAI211_X1 U10973 ( .C1(n9927), .C2(n9891), .A(n4779), .B(n9890), .ZN(n9926)
         );
  INV_X1 U10974 ( .A(n9926), .ZN(n9892) );
  AOI22_X1 U10975 ( .A1(n9931), .A2(n9894), .B1(n9893), .B2(n9892), .ZN(n9895)
         );
  OAI211_X1 U10976 ( .C1(n4321), .C2(n9928), .A(n9896), .B(n9895), .ZN(
        P1_U3289) );
  AOI22_X1 U10977 ( .A1(n9897), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n4321), .ZN(n9908) );
  NAND2_X1 U10978 ( .A1(n9899), .A2(n9898), .ZN(n9903) );
  NAND2_X1 U10979 ( .A1(n9901), .A2(n9900), .ZN(n9902) );
  OAI211_X1 U10980 ( .C1(n9905), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9906)
         );
  INV_X1 U10981 ( .A(n9906), .ZN(n9907) );
  OAI211_X1 U10982 ( .C1(n4321), .C2(n9909), .A(n9908), .B(n9907), .ZN(
        P1_U3292) );
  AND2_X1 U10983 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9913), .ZN(P1_U3294) );
  AND2_X1 U10984 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9913), .ZN(P1_U3295) );
  AND2_X1 U10985 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9913), .ZN(P1_U3296) );
  AND2_X1 U10986 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9913), .ZN(P1_U3297) );
  NOR2_X1 U10987 ( .A1(n9912), .A2(n9910), .ZN(P1_U3298) );
  AND2_X1 U10988 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9913), .ZN(P1_U3299) );
  NOR2_X1 U10989 ( .A1(n9912), .A2(n9911), .ZN(P1_U3300) );
  AND2_X1 U10990 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9913), .ZN(P1_U3301) );
  AND2_X1 U10991 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9913), .ZN(P1_U3302) );
  AND2_X1 U10992 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9913), .ZN(P1_U3303) );
  AND2_X1 U10993 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9913), .ZN(P1_U3304) );
  AND2_X1 U10994 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9913), .ZN(P1_U3305) );
  AND2_X1 U10995 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9913), .ZN(P1_U3306) );
  AND2_X1 U10996 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9913), .ZN(P1_U3307) );
  AND2_X1 U10997 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9913), .ZN(P1_U3308) );
  AND2_X1 U10998 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9913), .ZN(P1_U3309) );
  AND2_X1 U10999 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9913), .ZN(P1_U3310) );
  AND2_X1 U11000 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9913), .ZN(P1_U3311) );
  AND2_X1 U11001 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9913), .ZN(P1_U3312) );
  AND2_X1 U11002 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9913), .ZN(P1_U3313) );
  AND2_X1 U11003 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9913), .ZN(P1_U3314) );
  AND2_X1 U11004 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9913), .ZN(P1_U3315) );
  AND2_X1 U11005 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9913), .ZN(P1_U3316) );
  AND2_X1 U11006 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9913), .ZN(P1_U3317) );
  AND2_X1 U11007 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9913), .ZN(P1_U3318) );
  AND2_X1 U11008 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9913), .ZN(P1_U3319) );
  AND2_X1 U11009 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9913), .ZN(P1_U3320) );
  AND2_X1 U11010 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9913), .ZN(P1_U3321) );
  AND2_X1 U11011 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9913), .ZN(P1_U3322) );
  AND2_X1 U11012 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9913), .ZN(P1_U3323) );
  AOI22_X1 U11013 ( .A1(n10004), .A2(n9914), .B1(n4933), .B2(n10002), .ZN(
        P1_U3456) );
  OAI211_X1 U11014 ( .C1(n9917), .C2(n9996), .A(n9916), .B(n9915), .ZN(n9918)
         );
  AOI21_X1 U11015 ( .B1(n9919), .B2(n10000), .A(n9918), .ZN(n10005) );
  AOI22_X1 U11016 ( .A1(n10004), .A2(n10005), .B1(n5023), .B2(n10002), .ZN(
        P1_U3459) );
  OAI21_X1 U11017 ( .B1(n9921), .B2(n9996), .A(n9920), .ZN(n9924) );
  INV_X1 U11018 ( .A(n9922), .ZN(n9923) );
  AOI211_X1 U11019 ( .C1(n10000), .C2(n9925), .A(n9924), .B(n9923), .ZN(n10006) );
  AOI22_X1 U11020 ( .A1(n10004), .A2(n10006), .B1(n5050), .B2(n10002), .ZN(
        P1_U3462) );
  OAI21_X1 U11021 ( .B1(n9927), .B2(n9996), .A(n9926), .ZN(n9930) );
  INV_X1 U11022 ( .A(n9928), .ZN(n9929) );
  AOI211_X1 U11023 ( .C1(n9931), .C2(n10000), .A(n9930), .B(n9929), .ZN(n10007) );
  AOI22_X1 U11024 ( .A1(n10004), .A2(n10007), .B1(n5080), .B2(n10002), .ZN(
        P1_U3465) );
  OAI21_X1 U11025 ( .B1(n9933), .B2(n9996), .A(n9932), .ZN(n9935) );
  AOI211_X1 U11026 ( .C1(n10000), .C2(n9936), .A(n9935), .B(n9934), .ZN(n10008) );
  INV_X1 U11027 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11028 ( .A1(n10004), .A2(n10008), .B1(n9937), .B2(n10002), .ZN(
        P1_U3468) );
  OAI21_X1 U11029 ( .B1(n9939), .B2(n9996), .A(n9938), .ZN(n9942) );
  INV_X1 U11030 ( .A(n9940), .ZN(n9941) );
  AOI211_X1 U11031 ( .C1(n10000), .C2(n9943), .A(n9942), .B(n9941), .ZN(n10009) );
  INV_X1 U11032 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U11033 ( .A1(n10004), .A2(n10009), .B1(n9944), .B2(n10002), .ZN(
        P1_U3471) );
  INV_X1 U11034 ( .A(n9945), .ZN(n9949) );
  NAND2_X1 U11035 ( .A1(n9946), .A2(n9981), .ZN(n9948) );
  OAI211_X1 U11036 ( .C1(n9949), .C2(n9996), .A(n9948), .B(n9947), .ZN(n9950)
         );
  NOR2_X1 U11037 ( .A1(n9951), .A2(n9950), .ZN(n10010) );
  INV_X1 U11038 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U11039 ( .A1(n10004), .A2(n10010), .B1(n9952), .B2(n10002), .ZN(
        P1_U3474) );
  OAI21_X1 U11040 ( .B1(n9954), .B2(n9996), .A(n9953), .ZN(n9957) );
  INV_X1 U11041 ( .A(n9955), .ZN(n9956) );
  AOI211_X1 U11042 ( .C1(n9981), .C2(n9958), .A(n9957), .B(n9956), .ZN(n10011)
         );
  AOI22_X1 U11043 ( .A1(n10004), .A2(n10011), .B1(n5195), .B2(n10002), .ZN(
        P1_U3477) );
  AND2_X1 U11044 ( .A1(n9960), .A2(n9959), .ZN(n9961) );
  NOR2_X1 U11045 ( .A1(n9962), .A2(n9961), .ZN(n9966) );
  OR2_X1 U11046 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  AND3_X1 U11047 ( .A1(n9967), .A2(n9966), .A3(n9965), .ZN(n10012) );
  INV_X1 U11048 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9968) );
  AOI22_X1 U11049 ( .A1(n10004), .A2(n10012), .B1(n9968), .B2(n10002), .ZN(
        P1_U3480) );
  OAI21_X1 U11050 ( .B1(n9970), .B2(n9996), .A(n9969), .ZN(n9972) );
  AOI211_X1 U11051 ( .C1(n10000), .C2(n9973), .A(n9972), .B(n9971), .ZN(n10013) );
  AOI22_X1 U11052 ( .A1(n10004), .A2(n10013), .B1(n9974), .B2(n10002), .ZN(
        P1_U3483) );
  INV_X1 U11053 ( .A(n9975), .ZN(n9980) );
  OAI21_X1 U11054 ( .B1(n9977), .B2(n9996), .A(n9976), .ZN(n9979) );
  AOI211_X1 U11055 ( .C1(n9981), .C2(n9980), .A(n9979), .B(n9978), .ZN(n10014)
         );
  INV_X1 U11056 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11057 ( .A1(n10004), .A2(n10014), .B1(n9982), .B2(n10002), .ZN(
        P1_U3486) );
  OAI211_X1 U11058 ( .C1(n9985), .C2(n9996), .A(n9984), .B(n9983), .ZN(n9986)
         );
  AOI21_X1 U11059 ( .B1(n9987), .B2(n10000), .A(n9986), .ZN(n10015) );
  INV_X1 U11060 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11061 ( .A1(n10004), .A2(n10015), .B1(n9988), .B2(n10002), .ZN(
        P1_U3489) );
  OAI211_X1 U11062 ( .C1(n9991), .C2(n9996), .A(n9990), .B(n9989), .ZN(n9992)
         );
  AOI21_X1 U11063 ( .B1(n9993), .B2(n10000), .A(n9992), .ZN(n10016) );
  INV_X1 U11064 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11065 ( .A1(n10004), .A2(n10016), .B1(n9994), .B2(n10002), .ZN(
        P1_U3492) );
  OAI21_X1 U11066 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n9998) );
  AOI211_X1 U11067 ( .C1(n10001), .C2(n10000), .A(n9999), .B(n9998), .ZN(
        n10018) );
  INV_X1 U11068 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11069 ( .A1(n10004), .A2(n10018), .B1(n10003), .B2(n10002), .ZN(
        P1_U3495) );
  AOI22_X1 U11070 ( .A1(n10019), .A2(n10005), .B1(n5022), .B2(n10017), .ZN(
        P1_U3524) );
  AOI22_X1 U11071 ( .A1(n10019), .A2(n10006), .B1(n5048), .B2(n10017), .ZN(
        P1_U3525) );
  AOI22_X1 U11072 ( .A1(n10019), .A2(n10007), .B1(n6726), .B2(n10017), .ZN(
        P1_U3526) );
  AOI22_X1 U11073 ( .A1(n10019), .A2(n10008), .B1(n6721), .B2(n10017), .ZN(
        P1_U3527) );
  AOI22_X1 U11074 ( .A1(n10019), .A2(n10009), .B1(n6719), .B2(n10017), .ZN(
        P1_U3528) );
  AOI22_X1 U11075 ( .A1(n10019), .A2(n10010), .B1(n6717), .B2(n10017), .ZN(
        P1_U3529) );
  AOI22_X1 U11076 ( .A1(n10019), .A2(n10011), .B1(n6728), .B2(n10017), .ZN(
        P1_U3530) );
  AOI22_X1 U11077 ( .A1(n10019), .A2(n10012), .B1(n6821), .B2(n10017), .ZN(
        P1_U3531) );
  AOI22_X1 U11078 ( .A1(n10019), .A2(n10013), .B1(n6845), .B2(n10017), .ZN(
        P1_U3532) );
  AOI22_X1 U11079 ( .A1(n10019), .A2(n10014), .B1(n6915), .B2(n10017), .ZN(
        P1_U3533) );
  AOI22_X1 U11080 ( .A1(n10019), .A2(n10015), .B1(n7143), .B2(n10017), .ZN(
        P1_U3534) );
  AOI22_X1 U11081 ( .A1(n10019), .A2(n10016), .B1(n7175), .B2(n10017), .ZN(
        P1_U3535) );
  AOI22_X1 U11082 ( .A1(n10019), .A2(n10018), .B1(n7397), .B2(n10017), .ZN(
        P1_U3536) );
  INV_X1 U11083 ( .A(n10029), .ZN(n10022) );
  OAI21_X1 U11084 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10025) );
  AOI222_X1 U11085 ( .A1(n10038), .A2(n10025), .B1(n10024), .B2(n10031), .C1(
        n10023), .C2(n10033), .ZN(n10026) );
  OAI21_X1 U11086 ( .B1(n10038), .B2(n6529), .A(n10026), .ZN(P2_U3226) );
  INV_X1 U11087 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10037) );
  AOI21_X1 U11088 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(n10030) );
  INV_X1 U11089 ( .A(n10030), .ZN(n10035) );
  AOI222_X1 U11090 ( .A1(n10038), .A2(n10035), .B1(n10034), .B2(n10033), .C1(
        n10032), .C2(n10031), .ZN(n10036) );
  OAI21_X1 U11091 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(P2_U3229) );
  INV_X1 U11092 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10044) );
  INV_X1 U11093 ( .A(n10039), .ZN(n10041) );
  AOI211_X1 U11094 ( .C1(n10043), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10082) );
  AOI22_X1 U11095 ( .A1(n10080), .A2(n10044), .B1(n10082), .B2(n10078), .ZN(
        P2_U3396) );
  INV_X1 U11096 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10050) );
  INV_X1 U11097 ( .A(n10045), .ZN(n10049) );
  OAI22_X1 U11098 ( .A1(n10047), .A2(n10074), .B1(n10046), .B2(n10072), .ZN(
        n10048) );
  NOR2_X1 U11099 ( .A1(n10049), .A2(n10048), .ZN(n10084) );
  AOI22_X1 U11100 ( .A1(n10080), .A2(n10050), .B1(n10084), .B2(n10078), .ZN(
        P2_U3405) );
  INV_X1 U11101 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10055) );
  OAI22_X1 U11102 ( .A1(n10052), .A2(n10074), .B1(n10051), .B2(n10072), .ZN(
        n10053) );
  NOR2_X1 U11103 ( .A1(n10054), .A2(n10053), .ZN(n10085) );
  AOI22_X1 U11104 ( .A1(n10080), .A2(n10055), .B1(n10085), .B2(n10078), .ZN(
        P2_U3408) );
  INV_X1 U11105 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10060) );
  OAI22_X1 U11106 ( .A1(n10057), .A2(n10074), .B1(n10056), .B2(n10072), .ZN(
        n10058) );
  NOR2_X1 U11107 ( .A1(n10059), .A2(n10058), .ZN(n10086) );
  AOI22_X1 U11108 ( .A1(n10080), .A2(n10060), .B1(n10086), .B2(n10078), .ZN(
        P2_U3414) );
  OAI22_X1 U11109 ( .A1(n10063), .A2(n10062), .B1(n10061), .B2(n10072), .ZN(
        n10064) );
  NOR2_X1 U11110 ( .A1(n10065), .A2(n10064), .ZN(n10087) );
  AOI22_X1 U11111 ( .A1(n10080), .A2(n10066), .B1(n10087), .B2(n10078), .ZN(
        P2_U3417) );
  INV_X1 U11112 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10071) );
  OAI22_X1 U11113 ( .A1(n10068), .A2(n10074), .B1(n10067), .B2(n10072), .ZN(
        n10069) );
  NOR2_X1 U11114 ( .A1(n10070), .A2(n10069), .ZN(n10089) );
  AOI22_X1 U11115 ( .A1(n10080), .A2(n10071), .B1(n10089), .B2(n10078), .ZN(
        P2_U3420) );
  INV_X1 U11116 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10079) );
  OAI22_X1 U11117 ( .A1(n10075), .A2(n10074), .B1(n10073), .B2(n10072), .ZN(
        n10076) );
  NOR2_X1 U11118 ( .A1(n10077), .A2(n10076), .ZN(n10091) );
  AOI22_X1 U11119 ( .A1(n10080), .A2(n10079), .B1(n10091), .B2(n10078), .ZN(
        P2_U3423) );
  AOI22_X1 U11120 ( .A1(n10092), .A2(n10082), .B1(n10081), .B2(n10090), .ZN(
        P2_U3461) );
  AOI22_X1 U11121 ( .A1(n10092), .A2(n10084), .B1(n10083), .B2(n10090), .ZN(
        P2_U3464) );
  AOI22_X1 U11122 ( .A1(n10092), .A2(n10085), .B1(n6524), .B2(n10090), .ZN(
        P2_U3465) );
  AOI22_X1 U11123 ( .A1(n10092), .A2(n10086), .B1(n6582), .B2(n10090), .ZN(
        P2_U3467) );
  AOI22_X1 U11124 ( .A1(n10092), .A2(n10087), .B1(n6537), .B2(n10090), .ZN(
        P2_U3468) );
  AOI22_X1 U11125 ( .A1(n10092), .A2(n10089), .B1(n10088), .B2(n10090), .ZN(
        P2_U3469) );
  AOI22_X1 U11126 ( .A1(n10092), .A2(n10091), .B1(n6547), .B2(n10090), .ZN(
        P2_U3470) );
  NOR2_X1 U11127 ( .A1(n10094), .A2(n10093), .ZN(n10095) );
  XOR2_X1 U11128 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10095), .Z(ADD_1068_U5) );
  XOR2_X1 U11129 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11130 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10097), .A(n10096), 
        .ZN(n10099) );
  XNOR2_X1 U11131 ( .A(n10099), .B(n10098), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11132 ( .A(n10101), .B(n10100), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11133 ( .A(n10103), .B(n10102), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11134 ( .A(n10105), .B(n10104), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11135 ( .A(n10107), .B(n10106), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11136 ( .A(n10109), .B(n10108), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11137 ( .A(n10111), .B(n10110), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11138 ( .A(n10113), .B(n10112), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11139 ( .A(n10115), .B(n10114), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11140 ( .A(n10117), .B(n10116), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11141 ( .A(n10119), .B(n10118), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11142 ( .A(n10121), .B(n10120), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11143 ( .A(n10123), .B(n10122), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11144 ( .A(n10125), .B(n10124), .ZN(ADD_1068_U50) );
  XOR2_X1 U11145 ( .A(n10127), .B(n10126), .Z(ADD_1068_U54) );
  XOR2_X1 U11146 ( .A(n10129), .B(n10128), .Z(ADD_1068_U53) );
  XNOR2_X1 U11147 ( .A(n10131), .B(n10130), .ZN(ADD_1068_U52) );
  NAND4_X1 U4928 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n8389)
         );
  INV_X2 U4890 ( .A(n8171), .ZN(n8185) );
  NAND2_X1 U6120 ( .A1(n4577), .A2(n4403), .ZN(n8731) );
  OR2_X1 U4826 ( .A1(n8566), .A2(n8588), .ZN(n8614) );
  CLKBUF_X2 U4867 ( .A(n7438), .Z(n7940) );
  NOR2_X1 U4869 ( .A1(n8731), .A2(n8732), .ZN(n8730) );
  NAND2_X1 U4870 ( .A1(n7561), .A2(n5901), .ZN(n7614) );
  OR2_X1 U4898 ( .A1(n5785), .A2(n5763), .ZN(n4463) );
  NAND2_X1 U6119 ( .A1(n8324), .A2(n7929), .ZN(n8223) );
  INV_X1 U6413 ( .A(n5882), .ZN(n4441) );
  NAND2_X2 U9641 ( .A1(n6993), .A2(n4476), .ZN(n4743) );
  OR2_X1 U10096 ( .A1(n5738), .A2(n4939), .ZN(n4940) );
endmodule

