

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2264, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913;

  NOR2_X1 U2299 ( .A1(n3097), .A2(n3096), .ZN(n3104) );
  CLKBUF_X2 U2300 ( .A(n3330), .Z(n3701) );
  AND2_X1 U2301 ( .A1(n3705), .A2(n4848), .ZN(n3330) );
  CLKBUF_X2 U2302 ( .A(n2766), .Z(n2786) );
  CLKBUF_X2 U2303 ( .A(n2766), .Z(n2900) );
  NAND2_X1 U2304 ( .A1(n2666), .A2(n3007), .ZN(n2766) );
  XNOR2_X1 U2305 ( .A(n2661), .B(IR_REG_29__SCAN_IN), .ZN(n3005) );
  NAND2_X1 U2306 ( .A1(n2395), .A2(n2515), .ZN(n2530) );
  INV_X2 U2307 ( .A(n3699), .ZN(n3706) );
  NOR2_X1 U2308 ( .A1(n2530), .A2(IR_REG_22__SCAN_IN), .ZN(n2519) );
  CLKBUF_X2 U2310 ( .A(n2716), .Z(n3585) );
  XNOR2_X1 U2311 ( .A(n2658), .B(n3608), .ZN(n2662) );
  INV_X1 U2312 ( .A(n4909), .ZN(n4526) );
  AND4_X1 U2313 ( .A1(n2550), .A2(n2371), .A3(n2370), .A4(n2369), .ZN(n2264)
         );
  OAI21_X2 U2314 ( .B1(n3176), .B2(n2939), .A(n3856), .ZN(n3275) );
  OAI21_X2 U2315 ( .B1(n3220), .B2(n2938), .A(n3883), .ZN(n3176) );
  AOI21_X2 U2316 ( .B1(n3977), .B2(n4451), .A(n3975), .ZN(n4383) );
  AND2_X2 U2317 ( .A1(n2987), .A2(n3061), .ZN(n4878) );
  INV_X4 U2318 ( .A(n3415), .ZN(n3705) );
  NAND2_X2 U2319 ( .A1(n3041), .A2(n3042), .ZN(n3415) );
  AOI21_X2 U2320 ( .B1(n3482), .B2(n3860), .A(n3865), .ZN(n3970) );
  AND2_X1 U2321 ( .A1(n2424), .A2(n3840), .ZN(n3721) );
  OR2_X1 U2322 ( .A1(n3838), .A2(n3839), .ZN(n2424) );
  OAI21_X1 U2323 ( .B1(n2352), .B2(n2345), .A(n2342), .ZN(n3619) );
  OAI21_X1 U2324 ( .B1(n2431), .B2(n2349), .A(n2347), .ZN(n3617) );
  AND2_X1 U2325 ( .A1(n2363), .A2(n2362), .ZN(n3346) );
  NAND4_X1 U2326 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n2916), .ZN(n4332)
         );
  OAI21_X1 U2327 ( .B1(n3334), .B2(n2365), .A(n2364), .ZN(n2363) );
  NOR2_X1 U2328 ( .A1(n3104), .A2(n3103), .ZN(n3108) );
  BUF_X2 U2329 ( .A(n2904), .Z(n2921) );
  CLKBUF_X1 U2330 ( .A(n3042), .Z(n3217) );
  INV_X2 U2331 ( .A(n4011), .ZN(U4043) );
  CLKBUF_X1 U2332 ( .A(n2706), .Z(n2904) );
  CLKBUF_X3 U2333 ( .A(n2709), .Z(n3017) );
  XNOR2_X1 U2334 ( .A(n2521), .B(IR_REG_24__SCAN_IN), .ZN(n4624) );
  XNOR2_X1 U2335 ( .A(n2518), .B(IR_REG_26__SCAN_IN), .ZN(n4623) );
  OR2_X1 U2336 ( .A1(n2519), .A2(n2645), .ZN(n2524) );
  AND4_X1 U2337 ( .A1(n2368), .A2(n2432), .A3(n2569), .A4(n2367), .ZN(n2600)
         );
  INV_X1 U2338 ( .A(IR_REG_0__SCAN_IN), .ZN(n2432) );
  NOR2_X1 U2339 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2368)
         );
  INV_X1 U2340 ( .A(IR_REG_1__SCAN_IN), .ZN(n2367) );
  NOR2_X1 U2341 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2371)
         );
  NOR2_X1 U2342 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2370)
         );
  NOR2_X1 U2343 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2369)
         );
  NOR2_X1 U2344 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2550)
         );
  NOR2_X2 U2345 ( .A1(n4365), .A2(n3978), .ZN(n4346) );
  NAND2_X1 U2346 ( .A1(n2930), .A2(n3991), .ZN(n3042) );
  NAND2_X1 U2347 ( .A1(n2308), .A2(n2307), .ZN(n4635) );
  NAND2_X1 U2348 ( .A1(n2301), .A2(n2309), .ZN(n2308) );
  NAND2_X1 U2349 ( .A1(n3145), .A2(n2282), .ZN(n2307) );
  INV_X1 U2350 ( .A(n4636), .ZN(n2309) );
  OR2_X1 U2351 ( .A1(n4645), .A2(n4646), .ZN(n2401) );
  INV_X1 U2352 ( .A(n3564), .ZN(n2356) );
  AOI21_X1 U2353 ( .B1(n2426), .B2(n3682), .A(n2360), .ZN(n2359) );
  INV_X1 U2354 ( .A(n3688), .ZN(n2360) );
  NAND2_X1 U2355 ( .A1(n2347), .A2(n2346), .ZN(n2345) );
  INV_X1 U2356 ( .A(n3616), .ZN(n2346) );
  INV_X1 U2357 ( .A(n2498), .ZN(n2497) );
  AND2_X1 U2358 ( .A1(n2267), .A2(n2396), .ZN(n2395) );
  INV_X1 U2359 ( .A(IR_REG_21__SCAN_IN), .ZN(n2396) );
  NOR2_X1 U2360 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2538)
         );
  INV_X1 U2361 ( .A(n4000), .ZN(n3045) );
  NAND2_X1 U2362 ( .A1(n2666), .A2(n2662), .ZN(n2709) );
  NAND2_X1 U2363 ( .A1(n2401), .A2(n2274), .ZN(n2400) );
  OAI22_X1 U2364 ( .A1(n4710), .A2(n4707), .B1(REG2_REG_13__SCAN_IN), .B2(
        n2822), .ZN(n2310) );
  NOR2_X1 U2365 ( .A1(n2310), .A2(n4263), .ZN(n2632) );
  NAND2_X1 U2366 ( .A1(n2319), .A2(n2608), .ZN(n2609) );
  NAND2_X1 U2367 ( .A1(n4268), .A2(n4269), .ZN(n2319) );
  NAND2_X1 U2368 ( .A1(n4284), .A2(n2314), .ZN(n4293) );
  NAND2_X1 U2369 ( .A1(n4291), .A2(n3559), .ZN(n2314) );
  INV_X1 U2370 ( .A(n4785), .ZN(n3918) );
  NOR2_X1 U2371 ( .A1(n4307), .A2(n4883), .ZN(n2438) );
  OR2_X1 U2372 ( .A1(n4734), .A2(n4625), .ZN(n4741) );
  NOR2_X1 U2373 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2494)
         );
  NOR2_X1 U2374 ( .A1(IR_REG_26__SCAN_IN), .A2(n2655), .ZN(n2659) );
  NOR2_X1 U2375 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2516)
         );
  NAND2_X1 U2376 ( .A1(n2310), .A2(n4263), .ZN(n2408) );
  AOI21_X1 U2377 ( .B1(n4310), .B2(n2445), .A(n2443), .ZN(n2442) );
  OR2_X1 U2378 ( .A1(n4310), .A2(n2441), .ZN(n2440) );
  AND2_X1 U2379 ( .A1(n2486), .A2(n2481), .ZN(n2480) );
  NAND2_X1 U2380 ( .A1(n2484), .A2(n2482), .ZN(n2481) );
  INV_X1 U2381 ( .A(n2884), .ZN(n2482) );
  OR2_X1 U2382 ( .A1(n3927), .A2(n2460), .ZN(n2459) );
  INV_X1 U2383 ( .A(n2805), .ZN(n2460) );
  NOR2_X1 U2384 ( .A1(n3652), .A2(n2419), .ZN(n2418) );
  INV_X1 U2385 ( .A(n3798), .ZN(n2419) );
  NAND2_X1 U2386 ( .A1(n3800), .A2(n2283), .ZN(n2341) );
  INV_X1 U2387 ( .A(n3799), .ZN(n2417) );
  OR2_X1 U2388 ( .A1(n3763), .A2(n2418), .ZN(n2416) );
  NOR2_X1 U2389 ( .A1(n2348), .A2(n3616), .ZN(n2344) );
  INV_X1 U2390 ( .A(n2349), .ZN(n2348) );
  INV_X1 U2391 ( .A(n3615), .ZN(n2343) );
  NAND2_X1 U2392 ( .A1(n4245), .A2(n2311), .ZN(n2616) );
  NAND2_X1 U2393 ( .A1(n2312), .A2(REG2_REG_2__SCAN_IN), .ZN(n2311) );
  INV_X1 U2394 ( .A(n2338), .ZN(n2334) );
  NOR2_X1 U2395 ( .A1(n2841), .A2(n2501), .ZN(n2500) );
  INV_X1 U2396 ( .A(n2824), .ZN(n2501) );
  OAI21_X1 U2397 ( .B1(n3310), .B2(n3888), .A(n3890), .ZN(n3394) );
  INV_X1 U2398 ( .A(n2455), .ZN(n2454) );
  OAI21_X1 U2399 ( .B1(n2763), .B2(n2456), .A(n3307), .ZN(n2455) );
  INV_X1 U2400 ( .A(n2765), .ZN(n2456) );
  NAND2_X1 U2401 ( .A1(n3567), .A2(n2947), .ZN(n2380) );
  INV_X1 U2402 ( .A(n3084), .ZN(n3242) );
  XNOR2_X1 U2403 ( .A(n2928), .B(n2927), .ZN(n2930) );
  INV_X1 U2404 ( .A(IR_REG_20__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U2405 ( .A1(n2926), .A2(IR_REG_31__SCAN_IN), .ZN(n2928) );
  INV_X1 U2406 ( .A(IR_REG_6__SCAN_IN), .ZN(n4206) );
  INV_X1 U2407 ( .A(n3332), .ZN(n2364) );
  NAND2_X1 U2408 ( .A1(n2355), .A2(n2356), .ZN(n2349) );
  NAND2_X1 U2409 ( .A1(n2271), .A2(n2356), .ZN(n2347) );
  NAND2_X1 U2410 ( .A1(n3726), .A2(n3682), .ZN(n3729) );
  AND2_X1 U2411 ( .A1(n3720), .A2(n3840), .ZN(n2423) );
  NAND2_X1 U2412 ( .A1(n3459), .A2(n2302), .ZN(n2431) );
  NAND2_X1 U2413 ( .A1(n2358), .A2(n2357), .ZN(n3809) );
  AOI21_X1 U2414 ( .B1(n2359), .B2(n2361), .A(n2293), .ZN(n2357) );
  INV_X1 U2415 ( .A(n3682), .ZN(n2361) );
  AND2_X1 U2416 ( .A1(n3585), .A2(DATAI_24_), .ZN(n3813) );
  INV_X1 U2417 ( .A(n3227), .ZN(n3600) );
  NAND2_X1 U2418 ( .A1(n2528), .A2(n2529), .ZN(n2716) );
  NAND2_X1 U2419 ( .A1(n2535), .A2(n2655), .ZN(n2529) );
  AND2_X1 U2420 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2508)
         );
  AND2_X1 U2421 ( .A1(n3738), .A2(n3735), .ZN(n3409) );
  XNOR2_X1 U2422 ( .A(n3046), .B(n3697), .ZN(n3085) );
  AND2_X1 U2423 ( .A1(n3003), .A2(n4623), .ZN(n2366) );
  OR2_X1 U2424 ( .A1(n2921), .A2(n4327), .ZN(n2668) );
  OR2_X1 U2425 ( .A1(n2921), .A2(n4355), .ZN(n2675) );
  INV_X1 U2426 ( .A(IR_REG_2__SCAN_IN), .ZN(n2557) );
  INV_X1 U2427 ( .A(IR_REG_4__SCAN_IN), .ZN(n4098) );
  OR2_X1 U2428 ( .A1(n3158), .A2(n2574), .ZN(n2338) );
  INV_X1 U2429 ( .A(n4767), .ZN(n2752) );
  OAI21_X1 U2430 ( .B1(n2622), .B2(n4776), .A(n2315), .ZN(n2623) );
  NAND2_X1 U2431 ( .A1(n2400), .A2(REG2_REG_7__SCAN_IN), .ZN(n2315) );
  XNOR2_X1 U2432 ( .A(n2591), .B(n2626), .ZN(n4680) );
  NAND2_X1 U2433 ( .A1(n4671), .A2(n2625), .ZN(n2627) );
  NAND2_X1 U2434 ( .A1(n4692), .A2(n2629), .ZN(n2630) );
  AND3_X1 U2435 ( .A1(n2320), .A2(n2321), .A3(n2306), .ZN(n2603) );
  NAND2_X1 U2436 ( .A1(n2268), .A2(n2322), .ZN(n2321) );
  NOR2_X1 U2437 ( .A1(n2324), .A2(REG1_REG_12__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2438 ( .A1(n4280), .A2(n2305), .ZN(n2325) );
  NAND2_X1 U2439 ( .A1(n2327), .A2(n2305), .ZN(n2326) );
  INV_X1 U2440 ( .A(n2610), .ZN(n2327) );
  OAI21_X1 U2441 ( .B1(n4328), .B2(n3964), .A(n3909), .ZN(n2390) );
  NAND2_X1 U2442 ( .A1(n2466), .A2(n2465), .ZN(n4345) );
  NAND2_X1 U2443 ( .A1(n4390), .A2(n3777), .ZN(n2465) );
  NAND2_X1 U2444 ( .A1(n4362), .A2(n2467), .ZN(n2466) );
  NAND2_X1 U2445 ( .A1(n2468), .A2(n4373), .ZN(n2467) );
  AND2_X1 U2446 ( .A1(n3585), .A2(DATAI_21_), .ZN(n4453) );
  NAND2_X1 U2447 ( .A1(n3551), .A2(n2856), .ZN(n4519) );
  NAND2_X1 U2448 ( .A1(n2825), .A2(n2500), .ZN(n2499) );
  NAND2_X1 U2449 ( .A1(n3481), .A2(n3927), .ZN(n3480) );
  NAND2_X1 U2450 ( .A1(n2732), .A2(n3931), .ZN(n3210) );
  AND2_X1 U2451 ( .A1(n3232), .A2(n2704), .ZN(n3130) );
  NAND2_X1 U2452 ( .A1(n3130), .A2(n3930), .ZN(n3129) );
  NAND2_X1 U2453 ( .A1(n2929), .A2(n3918), .ZN(n4474) );
  NOR2_X1 U2454 ( .A1(n4534), .A2(n2985), .ZN(n2381) );
  AND3_X1 U2455 ( .A1(n2979), .A2(n2978), .A3(n3057), .ZN(n2991) );
  NAND2_X1 U2456 ( .A1(n2965), .A2(n4623), .ZN(n3011) );
  AND3_X1 U2457 ( .A1(n2515), .A2(n2288), .A3(n2395), .ZN(n2527) );
  INV_X1 U2458 ( .A(IR_REG_22__SCAN_IN), .ZN(n2493) );
  NOR2_X1 U2459 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2514)
         );
  NOR2_X1 U2460 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2513)
         );
  INV_X1 U2461 ( .A(n2545), .ZN(n2542) );
  NOR2_X1 U2462 ( .A1(n2575), .A2(IR_REG_5__SCAN_IN), .ZN(n2553) );
  NOR2_X1 U2463 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2560)
         );
  NAND2_X1 U2464 ( .A1(n2412), .A2(IR_REG_1__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U2465 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2412)
         );
  INV_X1 U2466 ( .A(n4625), .ZN(n4005) );
  NAND4_X1 U2467 ( .A1(n2731), .A2(n2730), .A3(n2729), .A4(n2728), .ZN(n4230)
         );
  OR2_X1 U2468 ( .A1(n2900), .A2(n2713), .ZN(n2714) );
  NOR2_X1 U2469 ( .A1(n2712), .A2(n2711), .ZN(n2715) );
  AND2_X1 U2470 ( .A1(n4641), .A2(n2276), .ZN(n2336) );
  NOR2_X1 U2471 ( .A1(n3155), .A2(n2301), .ZN(n4637) );
  NAND2_X1 U2472 ( .A1(n4672), .A2(n4673), .ZN(n4671) );
  XNOR2_X1 U2473 ( .A(n2627), .B(n2626), .ZN(n4678) );
  NAND2_X1 U2474 ( .A1(n4693), .A2(n4694), .ZN(n4692) );
  XNOR2_X1 U2475 ( .A(n2630), .B(n4845), .ZN(n4704) );
  NAND2_X1 U2476 ( .A1(n4704), .A2(REG2_REG_12__SCAN_IN), .ZN(n4702) );
  INV_X1 U2477 ( .A(n2407), .ZN(n2406) );
  NAND2_X1 U2478 ( .A1(n3022), .A2(n4908), .ZN(n4731) );
  AOI21_X1 U2479 ( .B1(n4299), .B2(n4298), .A(n2328), .ZN(n2612) );
  NOR2_X1 U2480 ( .A1(n4303), .A2(n2329), .ZN(n2328) );
  INV_X1 U2481 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2329) );
  AND2_X1 U2482 ( .A1(n3022), .A2(n4002), .ZN(n4726) );
  XNOR2_X1 U2483 ( .A(n2403), .B(n2641), .ZN(n2402) );
  NAND2_X1 U2484 ( .A1(n2405), .A2(n2404), .ZN(n2403) );
  NAND2_X1 U2485 ( .A1(n4627), .A2(REG2_REG_18__SCAN_IN), .ZN(n2404) );
  OR2_X1 U2486 ( .A1(n4310), .A2(n2272), .ZN(n2434) );
  XNOR2_X1 U2487 ( .A(n2382), .B(n3990), .ZN(n3594) );
  OAI211_X1 U2488 ( .C1(n2439), .C2(n2399), .A(n2450), .B(n4888), .ZN(n2398)
         );
  NOR2_X1 U2489 ( .A1(n2530), .A2(n2491), .ZN(n2490) );
  NAND2_X1 U2490 ( .A1(n2657), .A2(n2288), .ZN(n2491) );
  AND2_X1 U2491 ( .A1(n4403), .A2(n2279), .ZN(n2484) );
  AOI21_X1 U2492 ( .B1(n2480), .B2(n2483), .A(n4406), .ZN(n2479) );
  INV_X1 U2493 ( .A(n2484), .ZN(n2483) );
  INV_X1 U2494 ( .A(n3821), .ZN(n3675) );
  AOI22_X1 U2495 ( .A1(n2565), .A2(n4249), .B1(n2312), .B2(REG1_REG_2__SCAN_IN), .ZN(n2567) );
  NOR2_X1 U2496 ( .A1(n3028), .A2(n2617), .ZN(n2618) );
  NOR2_X1 U2497 ( .A1(n2451), .A2(n2291), .ZN(n2447) );
  INV_X1 U2498 ( .A(n4316), .ZN(n2446) );
  NOR2_X1 U2499 ( .A1(n4383), .A2(n3980), .ZN(n4365) );
  AOI21_X1 U2500 ( .B1(n2479), .B2(n2477), .A(n2476), .ZN(n2475) );
  INV_X1 U2501 ( .A(n3921), .ZN(n2476) );
  INV_X1 U2502 ( .A(n2480), .ZN(n2477) );
  INV_X1 U2503 ( .A(n2479), .ZN(n2478) );
  AND2_X1 U2504 ( .A1(n2899), .A2(n2933), .ZN(n4431) );
  AND2_X1 U2505 ( .A1(REG3_REG_20__SCAN_IN), .A2(n2664), .ZN(n2876) );
  NAND2_X1 U2506 ( .A1(n2394), .A2(n2393), .ZN(n4468) );
  INV_X1 U2507 ( .A(n3899), .ZN(n2393) );
  INV_X1 U2508 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U2509 ( .A1(n2458), .A2(n2457), .ZN(n3429) );
  AOI21_X1 U2510 ( .B1(n2269), .B2(n2460), .A(n2296), .ZN(n2457) );
  INV_X1 U2511 ( .A(n2718), .ZN(n2489) );
  NOR2_X1 U2512 ( .A1(n4339), .A2(n3713), .ZN(n2984) );
  OR3_X1 U2513 ( .A1(n3777), .A2(n3813), .A3(n2385), .ZN(n2384) );
  AOI21_X1 U2514 ( .B1(n4485), .B2(n2875), .A(n2874), .ZN(n4473) );
  NOR2_X1 U2515 ( .A1(n3831), .A2(n4499), .ZN(n2374) );
  XNOR2_X1 U2516 ( .A(n2414), .B(n3707), .ZN(n3187) );
  NAND2_X1 U2517 ( .A1(n3106), .A2(n2415), .ZN(n2414) );
  NAND2_X1 U2518 ( .A1(n3093), .A2(n3105), .ZN(n2415) );
  INV_X1 U2519 ( .A(n4312), .ZN(n3713) );
  OR2_X1 U2520 ( .A1(n3041), .A2(n3048), .ZN(n2503) );
  OR2_X1 U2521 ( .A1(n3532), .A2(n3533), .ZN(n2355) );
  OAI22_X1 U2522 ( .A1(n2270), .A2(n2354), .B1(n3460), .B2(n3531), .ZN(n2353)
         );
  INV_X1 U2523 ( .A(n3532), .ZN(n2354) );
  AND2_X1 U2524 ( .A1(n2806), .A2(REG3_REG_12__SCAN_IN), .ZN(n2815) );
  AND2_X1 U2525 ( .A1(n2815), .A2(REG3_REG_13__SCAN_IN), .ZN(n2826) );
  AOI21_X1 U2526 ( .B1(n2340), .B2(n4897), .A(n3670), .ZN(n3671) );
  NAND2_X1 U2527 ( .A1(n2341), .A2(n2416), .ZN(n2340) );
  AND2_X1 U2528 ( .A1(n2280), .A2(n2339), .ZN(n3094) );
  XNOR2_X1 U2529 ( .A(n3092), .B(n3697), .ZN(n3095) );
  NAND2_X1 U2530 ( .A1(n3800), .A2(n3799), .ZN(n2420) );
  NAND2_X1 U2531 ( .A1(n2826), .A2(REG3_REG_14__SCAN_IN), .ZN(n2833) );
  INV_X1 U2532 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2832) );
  OR2_X1 U2533 ( .A1(n2833), .A2(n2832), .ZN(n2842) );
  AOI21_X1 U2534 ( .B1(n2347), .B2(n2344), .A(n2343), .ZN(n2342) );
  NOR2_X1 U2535 ( .A1(n4785), .A2(n4005), .ZN(n4000) );
  OR2_X1 U2536 ( .A1(n2709), .A2(n2690), .ZN(n2691) );
  OR2_X1 U2537 ( .A1(n2766), .A2(n2689), .ZN(n2692) );
  NAND2_X1 U2538 ( .A1(n2920), .A2(REG2_REG_0__SCAN_IN), .ZN(n2701) );
  OAI21_X1 U2539 ( .B1(n4253), .B2(REG2_REG_2__SCAN_IN), .A(n2313), .ZN(n4247)
         );
  NAND2_X1 U2540 ( .A1(n4253), .A2(REG2_REG_2__SCAN_IN), .ZN(n2313) );
  NAND2_X1 U2541 ( .A1(n4246), .A2(n4247), .ZN(n4245) );
  INV_X1 U2542 ( .A(IR_REG_3__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U2543 ( .A(n2618), .B(n4630), .ZN(n3145) );
  NOR2_X1 U2544 ( .A1(n4635), .A2(n2292), .ZN(n2621) );
  AOI21_X1 U2545 ( .B1(n2336), .B2(n2334), .A(n2275), .ZN(n2333) );
  INV_X1 U2546 ( .A(n2336), .ZN(n2335) );
  OR2_X1 U2547 ( .A1(n4698), .A2(n4699), .ZN(n2323) );
  AND2_X1 U2548 ( .A1(n2408), .A2(REG2_REG_14__SCAN_IN), .ZN(n2407) );
  NOR2_X1 U2549 ( .A1(n2407), .A2(n2632), .ZN(n4273) );
  OR2_X1 U2550 ( .A1(n4273), .A2(n4272), .ZN(n4270) );
  INV_X1 U2551 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4184) );
  AND2_X1 U2552 ( .A1(n4270), .A2(n2634), .ZN(n2636) );
  NAND2_X1 U2553 ( .A1(n4283), .A2(n4285), .ZN(n4284) );
  AND2_X1 U2554 ( .A1(n3585), .A2(n2534), .ZN(n2650) );
  INV_X1 U2555 ( .A(n2447), .ZN(n2441) );
  NAND2_X1 U2556 ( .A1(n2444), .A2(n2448), .ZN(n2443) );
  NAND2_X1 U2557 ( .A1(n2451), .A2(n2291), .ZN(n2448) );
  NAND2_X1 U2558 ( .A1(n2447), .A2(n2446), .ZN(n2444) );
  NOR2_X1 U2559 ( .A1(n3957), .A2(n2446), .ZN(n2445) );
  OAI21_X1 U2560 ( .B1(n4346), .B2(n3963), .A(n3960), .ZN(n4330) );
  INV_X1 U2561 ( .A(n4337), .ZN(n4329) );
  INV_X1 U2562 ( .A(n2461), .ZN(n4338) );
  OAI21_X1 U2563 ( .B1(n4345), .B2(n2463), .A(n2462), .ZN(n2461) );
  NAND2_X1 U2564 ( .A1(n2464), .A2(n4359), .ZN(n2462) );
  NOR2_X1 U2565 ( .A1(n2464), .A2(n4359), .ZN(n2463) );
  OR3_X1 U2566 ( .A1(n2683), .A2(n4181), .A3(n3844), .ZN(n2671) );
  INV_X1 U2567 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4181) );
  AOI21_X1 U2568 ( .B1(n4368), .B2(n4393), .A(n2909), .ZN(n4362) );
  NAND2_X1 U2569 ( .A1(n2474), .A2(n2472), .ZN(n4399) );
  AOI21_X1 U2570 ( .B1(n2475), .B2(n2478), .A(n2473), .ZN(n2472) );
  NAND2_X1 U2571 ( .A1(n4473), .A2(n2475), .ZN(n2474) );
  INV_X1 U2572 ( .A(n3920), .ZN(n2473) );
  NAND2_X1 U2573 ( .A1(n3585), .A2(DATAI_23_), .ZN(n4413) );
  NAND2_X1 U2574 ( .A1(n2893), .A2(REG3_REG_22__SCAN_IN), .ZN(n2901) );
  AND2_X1 U2575 ( .A1(n2876), .A2(REG3_REG_21__SCAN_IN), .ZN(n2893) );
  AND2_X1 U2576 ( .A1(n2485), .A2(n2279), .ZN(n4449) );
  NAND2_X1 U2577 ( .A1(n4473), .A2(n2884), .ZN(n2485) );
  AND4_X1 U2578 ( .A1(n2883), .A2(n2882), .A3(n2881), .A4(n2880), .ZN(n4457)
         );
  INV_X1 U2579 ( .A(n2391), .ZN(n4451) );
  OAI21_X1 U2580 ( .B1(n4468), .B2(n3949), .A(n2392), .ZN(n2391) );
  NOR2_X1 U2581 ( .A1(n2857), .A2(n3832), .ZN(n2869) );
  NOR2_X1 U2582 ( .A1(n2842), .A2(n4184), .ZN(n2851) );
  OAI21_X1 U2583 ( .B1(n2825), .B2(n2497), .A(n2495), .ZN(n3551) );
  AND2_X1 U2584 ( .A1(n2496), .A2(n2850), .ZN(n2495) );
  OR2_X1 U2585 ( .A1(n2497), .A2(n2500), .ZN(n2496) );
  INV_X1 U2586 ( .A(n3628), .ZN(n3791) );
  AND2_X1 U2587 ( .A1(n2502), .A2(n2840), .ZN(n2498) );
  NAND2_X1 U2588 ( .A1(n2825), .A2(n2824), .ZN(n3448) );
  NOR2_X2 U2589 ( .A1(n3970), .A2(n3943), .ZN(n3519) );
  NAND2_X1 U2590 ( .A1(n3394), .A2(n3859), .ZN(n2945) );
  OR2_X1 U2591 ( .A1(n2775), .A2(n2774), .ZN(n2787) );
  INV_X1 U2592 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4065) );
  AOI21_X1 U2593 ( .B1(n2454), .B2(n2456), .A(n2287), .ZN(n2453) );
  INV_X1 U2594 ( .A(n3371), .ZN(n3314) );
  NAND2_X1 U2595 ( .A1(n2944), .A2(n3854), .ZN(n3310) );
  NOR2_X1 U2596 ( .A1(n2755), .A2(n2754), .ZN(n2767) );
  NAND2_X1 U2597 ( .A1(n2372), .A2(n2942), .ZN(n4778) );
  INV_X1 U2598 ( .A(n4777), .ZN(n2372) );
  NAND2_X1 U2599 ( .A1(n2764), .A2(n2763), .ZN(n4782) );
  NAND2_X1 U2600 ( .A1(n2470), .A2(n2469), .ZN(n3274) );
  AOI21_X1 U2601 ( .B1(n2744), .B2(n2471), .A(n2278), .ZN(n2469) );
  INV_X1 U2602 ( .A(n2733), .ZN(n2471) );
  AND2_X1 U2603 ( .A1(n3879), .A2(n3883), .ZN(n3219) );
  AND2_X1 U2604 ( .A1(n4908), .A2(n3060), .ZN(n4493) );
  NAND2_X1 U2605 ( .A1(n2935), .A2(n3870), .ZN(n3929) );
  OAI21_X1 U2606 ( .B1(n2716), .B2(n4232), .A(n2696), .ZN(n2703) );
  NAND2_X1 U2607 ( .A1(n2716), .A2(n2695), .ZN(n2696) );
  INV_X1 U2608 ( .A(n4794), .ZN(n4509) );
  NAND2_X1 U2609 ( .A1(n3234), .A2(n3872), .ZN(n2387) );
  INV_X1 U2610 ( .A(n3929), .ZN(n3234) );
  INV_X1 U2611 ( .A(n4493), .ZN(n4799) );
  AND2_X1 U2612 ( .A1(n4005), .A2(n3073), .ZN(n3061) );
  NAND2_X1 U2613 ( .A1(n2443), .A2(n4874), .ZN(n2435) );
  AND2_X1 U2614 ( .A1(n2445), .A2(n4874), .ZN(n2436) );
  INV_X1 U2615 ( .A(n3912), .ZN(n4534) );
  AND2_X1 U2616 ( .A1(n4626), .A2(n3061), .ZN(n4794) );
  NAND2_X1 U2617 ( .A1(n3585), .A2(DATAI_27_), .ZN(n4340) );
  NOR3_X1 U2618 ( .A1(n4421), .A2(n3777), .A3(n3813), .ZN(n4375) );
  NOR2_X1 U2619 ( .A1(n4421), .A2(n3813), .ZN(n4391) );
  OR2_X1 U2620 ( .A1(n4562), .A2(n4419), .ZN(n4421) );
  AND2_X1 U2621 ( .A1(n4508), .A2(n2300), .ZN(n4460) );
  NAND2_X1 U2622 ( .A1(n4508), .A2(n4510), .ZN(n4507) );
  NAND2_X1 U2623 ( .A1(n4508), .A2(n2374), .ZN(n4501) );
  NOR2_X1 U2624 ( .A1(n4879), .A2(n3802), .ZN(n4508) );
  NAND2_X1 U2625 ( .A1(n2379), .A2(n2378), .ZN(n2377) );
  NOR2_X1 U2626 ( .A1(n3544), .A2(n4860), .ZN(n2378) );
  INV_X1 U2627 ( .A(n2380), .ZN(n2379) );
  INV_X1 U2628 ( .A(n3570), .ZN(n3567) );
  NOR3_X1 U2629 ( .A1(n3477), .A2(n3544), .A3(n3463), .ZN(n3454) );
  NOR2_X1 U2630 ( .A1(n3477), .A2(n3463), .ZN(n3442) );
  OR2_X1 U2631 ( .A1(n3476), .A2(n3484), .ZN(n3477) );
  INV_X1 U2632 ( .A(n3740), .ZN(n3391) );
  AND2_X1 U2633 ( .A1(n4812), .A2(n3314), .ZN(n3392) );
  INV_X1 U2634 ( .A(n3276), .ZN(n3282) );
  NAND2_X1 U2635 ( .A1(n3283), .A2(n3282), .ZN(n4777) );
  OR2_X1 U2636 ( .A1(n3169), .A2(n3600), .ZN(n3226) );
  NOR2_X1 U2637 ( .A1(n3226), .A2(n3202), .ZN(n3283) );
  AND2_X1 U2638 ( .A1(n2703), .A2(n3084), .ZN(n3241) );
  INV_X1 U2639 ( .A(n4878), .ZN(n4848) );
  INV_X1 U2640 ( .A(n4624), .ZN(n2980) );
  AND2_X1 U2641 ( .A1(n3041), .A2(n3012), .ZN(n3074) );
  NAND2_X1 U2642 ( .A1(n3607), .A2(IR_REG_31__SCAN_IN), .ZN(n2658) );
  INV_X1 U2643 ( .A(IR_REG_28__SCAN_IN), .ZN(n2647) );
  INV_X1 U2644 ( .A(IR_REG_26__SCAN_IN), .ZN(n2526) );
  INV_X1 U2645 ( .A(IR_REG_27__SCAN_IN), .ZN(n2643) );
  XNOR2_X1 U2646 ( .A(n2524), .B(n2523), .ZN(n3999) );
  CLKBUF_X1 U2647 ( .A(n2930), .Z(n2987) );
  NOR2_X1 U2648 ( .A1(n2430), .A2(IR_REG_19__SCAN_IN), .ZN(n2429) );
  INV_X1 U2649 ( .A(n2541), .ZN(n2430) );
  NAND2_X1 U2650 ( .A1(n2549), .A2(n2537), .ZN(n2605) );
  OR2_X1 U2651 ( .A1(n2589), .A2(IR_REG_9__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U2652 ( .A1(n2560), .A2(n2557), .ZN(n2566) );
  NAND2_X1 U2653 ( .A1(n3334), .A2(n2365), .ZN(n2362) );
  INV_X1 U2654 ( .A(n4340), .ZN(n4331) );
  NAND2_X1 U2655 ( .A1(n2424), .A2(n2423), .ZN(n3719) );
  INV_X1 U2656 ( .A(n4413), .ZN(n4419) );
  NAND2_X1 U2657 ( .A1(n2422), .A2(n2421), .ZN(n3712) );
  AOI21_X1 U2658 ( .B1(n2423), .B2(n3839), .A(n3704), .ZN(n2421) );
  INV_X1 U2659 ( .A(n2703), .ZN(n3243) );
  NAND2_X1 U2660 ( .A1(n2431), .A2(n3460), .ZN(n3534) );
  AND2_X1 U2661 ( .A1(n2351), .A2(n2350), .ZN(n3565) );
  INV_X1 U2662 ( .A(n2353), .ZN(n2350) );
  NAND2_X1 U2663 ( .A1(n2352), .A2(n2355), .ZN(n2351) );
  NAND2_X1 U2664 ( .A1(n2427), .A2(n2504), .ZN(n3820) );
  NAND2_X1 U2665 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  NAND2_X1 U2666 ( .A1(n2420), .A2(n3798), .ZN(n3830) );
  AND2_X1 U2667 ( .A1(n3113), .A2(n3112), .ZN(n4906) );
  INV_X1 U2668 ( .A(n4896), .ZN(n4867) );
  NAND4_X1 U2669 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .ZN(n4350)
         );
  OR2_X1 U2670 ( .A1(n3017), .A2(n2673), .ZN(n2674) );
  INV_X1 U2671 ( .A(n4457), .ZN(n4494) );
  CLKBUF_X1 U2672 ( .A(n3040), .Z(n4231) );
  AND2_X1 U2673 ( .A1(n2651), .A2(n2650), .ZN(n3022) );
  AND2_X1 U2674 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4234)
         );
  XNOR2_X1 U2675 ( .A(n2573), .B(n3158), .ZN(n3146) );
  AND2_X1 U2676 ( .A1(n3145), .A2(REG2_REG_4__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U2677 ( .A1(n2573), .A2(n2338), .ZN(n2337) );
  INV_X1 U2678 ( .A(n2316), .ZN(n4657) );
  NAND2_X1 U2679 ( .A1(n3125), .A2(n2624), .ZN(n4672) );
  NAND2_X1 U2680 ( .A1(n4677), .A2(n2628), .ZN(n4693) );
  NAND2_X1 U2681 ( .A1(n4679), .A2(n2592), .ZN(n4688) );
  INV_X1 U2682 ( .A(n2323), .ZN(n4697) );
  NAND2_X1 U2683 ( .A1(n4702), .A2(n2631), .ZN(n4710) );
  NAND2_X1 U2684 ( .A1(n4258), .A2(n2604), .ZN(n4268) );
  XNOR2_X1 U2685 ( .A(n2636), .B(n2635), .ZN(n4722) );
  XNOR2_X1 U2686 ( .A(n2609), .B(n2635), .ZN(n4727) );
  AND2_X1 U2687 ( .A1(n2962), .A2(n2299), .ZN(n2388) );
  XNOR2_X1 U2688 ( .A(n2390), .B(n2451), .ZN(n2389) );
  NAND2_X1 U2689 ( .A1(n4460), .A2(n4428), .ZN(n4562) );
  OR2_X1 U2690 ( .A1(n2266), .A2(n3791), .ZN(n4879) );
  NAND2_X1 U2691 ( .A1(n2499), .A2(n2840), .ZN(n3504) );
  NAND2_X1 U2692 ( .A1(n2499), .A2(n2498), .ZN(n4876) );
  NAND2_X1 U2693 ( .A1(n3480), .A2(n2805), .ZN(n3384) );
  NOR2_X1 U2694 ( .A1(n4778), .A2(n3355), .ZN(n4812) );
  NAND2_X1 U2695 ( .A1(n3210), .A2(n2733), .ZN(n3175) );
  NAND2_X1 U2696 ( .A1(n3129), .A2(n2718), .ZN(n3159) );
  INV_X1 U2697 ( .A(n4833), .ZN(n4910) );
  AND2_X1 U2698 ( .A1(n4526), .A2(n3218), .ZN(n4825) );
  AND2_X1 U2699 ( .A1(n2981), .A2(n2980), .ZN(n3013) );
  NAND2_X1 U2700 ( .A1(n3011), .A2(n3074), .ZN(n4634) );
  NAND2_X1 U2701 ( .A1(n2660), .A2(IR_REG_31__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U2702 ( .A1(n2527), .A2(n2659), .ZN(n2660) );
  NAND2_X1 U2703 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2518) );
  XNOR2_X1 U2704 ( .A(n2522), .B(IR_REG_25__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U2705 ( .A1(n2516), .A2(n2493), .ZN(n2492) );
  XNOR2_X1 U2706 ( .A(n2531), .B(IR_REG_22__SCAN_IN), .ZN(n4625) );
  XNOR2_X1 U2707 ( .A(n2533), .B(IR_REG_21__SCAN_IN), .ZN(n3991) );
  OR2_X1 U2708 ( .A1(n2556), .A2(n2555), .ZN(n4767) );
  NAND2_X1 U2709 ( .A1(n2411), .A2(n2410), .ZN(n2562) );
  NAND2_X1 U2710 ( .A1(n2367), .A2(IR_REG_31__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U2711 ( .A1(n2337), .A2(n2336), .ZN(n4640) );
  NAND2_X1 U2712 ( .A1(n2409), .A2(n2408), .ZN(n4264) );
  AOI21_X1 U2713 ( .B1(n2405), .B2(n4297), .A(n4296), .ZN(n4302) );
  AOI21_X1 U2714 ( .B1(n2402), .B2(n4703), .A(n2303), .ZN(n2511) );
  OAI21_X1 U2715 ( .B1(n3594), .B2(n4833), .A(n3593), .ZN(U3260) );
  NAND2_X1 U2716 ( .A1(n2437), .A2(n2449), .ZN(n2996) );
  NAND2_X1 U2717 ( .A1(n4883), .A2(n2992), .ZN(n2449) );
  NAND2_X1 U2718 ( .A1(n2398), .A2(n2397), .ZN(n2990) );
  NAND2_X1 U2719 ( .A1(n4886), .A2(n2983), .ZN(n2397) );
  NAND3_X2 U2720 ( .A1(n2286), .A2(n2723), .A3(n2722), .ZN(n3105) );
  OAI21_X1 U2721 ( .B1(n2389), .B2(n4513), .A(n2388), .ZN(n4307) );
  OR2_X1 U2722 ( .A1(n3477), .A2(n2377), .ZN(n2266) );
  INV_X2 U2723 ( .A(n3093), .ZN(n3699) );
  XNOR2_X1 U2724 ( .A(n2558), .B(n2557), .ZN(n4253) );
  INV_X1 U2725 ( .A(n4253), .ZN(n2312) );
  AND4_X1 U2726 ( .A1(n2538), .A2(n2514), .A3(n2513), .A4(n2512), .ZN(n2267)
         );
  OR2_X1 U2727 ( .A1(n2599), .A2(n4845), .ZN(n2268) );
  AND2_X1 U2728 ( .A1(n2459), .A2(n2814), .ZN(n2269) );
  AND2_X1 U2729 ( .A1(n3460), .A2(n3531), .ZN(n2270) );
  OR2_X1 U2730 ( .A1(n2353), .A2(n2298), .ZN(n2271) );
  INV_X1 U2731 ( .A(n4390), .ZN(n2468) );
  NAND4_X1 U2732 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(n4370)
         );
  INV_X1 U2733 ( .A(n4370), .ZN(n2464) );
  INV_X1 U2734 ( .A(n3971), .ZN(n2392) );
  OR2_X1 U2735 ( .A1(n2441), .A2(n2439), .ZN(n2272) );
  AND2_X1 U2736 ( .A1(n2374), .A2(n4890), .ZN(n2273) );
  INV_X1 U2737 ( .A(n4359), .ZN(n2385) );
  INV_X1 U2738 ( .A(n3333), .ZN(n2365) );
  INV_X1 U2739 ( .A(IR_REG_31__SCAN_IN), .ZN(n2645) );
  OR2_X1 U2740 ( .A1(n3040), .A2(n2703), .ZN(n2935) );
  OR2_X1 U2741 ( .A1(n2621), .A2(n4767), .ZN(n2274) );
  INV_X1 U2742 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U2743 ( .A1(n2366), .A2(n4624), .ZN(n3041) );
  NAND2_X1 U2744 ( .A1(n2562), .A2(n2561), .ZN(n4236) );
  OR2_X1 U2745 ( .A1(n4293), .A2(n4292), .ZN(n2405) );
  AND2_X1 U2746 ( .A1(n2743), .A2(REG1_REG_5__SCAN_IN), .ZN(n2275) );
  NAND2_X1 U2747 ( .A1(n3158), .A2(n2574), .ZN(n2276) );
  NAND2_X1 U2748 ( .A1(n3692), .A2(n2510), .ZN(n3838) );
  AND2_X1 U2749 ( .A1(n4348), .A2(n4347), .ZN(n2277) );
  AND2_X1 U2750 ( .A1(n4229), .A2(n3202), .ZN(n2278) );
  NAND2_X1 U2751 ( .A1(n4494), .A2(n4479), .ZN(n2279) );
  OR2_X1 U2752 ( .A1(n3140), .A2(n3699), .ZN(n2280) );
  OAI21_X1 U2753 ( .B1(n3497), .B2(n2502), .A(n3966), .ZN(n3552) );
  INV_X1 U2754 ( .A(n3552), .ZN(n2394) );
  OR2_X1 U2755 ( .A1(n2530), .A2(n2492), .ZN(n2281) );
  NOR2_X1 U2756 ( .A1(n4636), .A2(n2726), .ZN(n2282) );
  NOR2_X1 U2757 ( .A1(n3763), .A2(n2417), .ZN(n2283) );
  NOR2_X1 U2758 ( .A1(n4281), .A2(n4280), .ZN(n2284) );
  AND2_X1 U2759 ( .A1(n2440), .A2(n2442), .ZN(n2399) );
  AND2_X1 U2760 ( .A1(n3190), .A2(n3191), .ZN(n2285) );
  AND2_X1 U2761 ( .A1(n2720), .A2(n2719), .ZN(n2286) );
  NAND2_X1 U2762 ( .A1(n3306), .A2(n2782), .ZN(n2287) );
  INV_X1 U2763 ( .A(n2426), .ZN(n2425) );
  NAND2_X1 U2764 ( .A1(n3675), .A2(n2504), .ZN(n2426) );
  AND2_X1 U2765 ( .A1(n2516), .A2(n2494), .ZN(n2288) );
  AND2_X1 U2766 ( .A1(n2438), .A2(n2435), .ZN(n2289) );
  NAND2_X1 U2767 ( .A1(n2515), .A2(n2267), .ZN(n2532) );
  AND2_X1 U2768 ( .A1(n2420), .A2(n2418), .ZN(n2290) );
  AND2_X1 U2769 ( .A1(n3852), .A2(n3966), .ZN(n3503) );
  INV_X1 U2770 ( .A(n3503), .ZN(n2502) );
  INV_X1 U2771 ( .A(n3544), .ZN(n3441) );
  AND2_X1 U2772 ( .A1(n4332), .A2(n3713), .ZN(n2291) );
  OAI21_X1 U2773 ( .B1(n3783), .B2(n3633), .A(n2509), .ZN(n3800) );
  NAND2_X1 U2774 ( .A1(n4508), .A2(n2273), .ZN(n2375) );
  AND2_X1 U2775 ( .A1(n2743), .A2(REG2_REG_5__SCAN_IN), .ZN(n2292) );
  XOR2_X1 U2776 ( .A(n3687), .B(n3707), .Z(n2293) );
  AND2_X1 U2777 ( .A1(n2323), .A2(n2268), .ZN(n2294) );
  INV_X1 U2778 ( .A(n3957), .ZN(n2451) );
  OR2_X1 U2779 ( .A1(n4223), .A2(n3544), .ZN(n2295) );
  NOR3_X1 U2780 ( .A1(n4421), .A2(n2384), .A3(n4331), .ZN(n2386) );
  INV_X1 U2781 ( .A(n2383), .ZN(n4544) );
  NOR2_X1 U2782 ( .A1(n4421), .A2(n2384), .ZN(n2383) );
  NOR2_X1 U2783 ( .A1(n4224), .A2(n3463), .ZN(n2296) );
  NAND4_X1 U2784 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(n4390)
         );
  NOR2_X1 U2785 ( .A1(n2406), .A2(n2632), .ZN(n2297) );
  INV_X1 U2786 ( .A(DATAI_0_), .ZN(n2373) );
  NAND2_X1 U2787 ( .A1(n4782), .A2(n2765), .ZN(n3291) );
  AND2_X1 U2788 ( .A1(n3540), .A2(n3539), .ZN(n2298) );
  OR2_X1 U2789 ( .A1(n3586), .A2(n3851), .ZN(n2299) );
  INV_X1 U2790 ( .A(n2376), .ZN(n3524) );
  NOR3_X1 U2791 ( .A1(n3477), .A2(n2380), .A3(n3544), .ZN(n2376) );
  INV_X1 U2792 ( .A(n4890), .ZN(n4479) );
  NAND2_X1 U2793 ( .A1(n3585), .A2(DATAI_20_), .ZN(n4890) );
  AND2_X1 U2794 ( .A1(n2273), .A2(n4458), .ZN(n2300) );
  INV_X1 U2795 ( .A(n4885), .ZN(n4883) );
  INV_X1 U2796 ( .A(n4888), .ZN(n4886) );
  INV_X1 U2797 ( .A(n4874), .ZN(n2439) );
  NAND2_X1 U2798 ( .A1(n2642), .A2(IR_REG_31__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U2799 ( .A1(n3929), .A2(n3233), .ZN(n3232) );
  INV_X1 U2800 ( .A(n3777), .ZN(n4373) );
  AND2_X1 U2801 ( .A1(n2619), .A2(n4630), .ZN(n2301) );
  NAND2_X1 U2802 ( .A1(n3421), .A2(n3420), .ZN(n2302) );
  NAND2_X1 U2803 ( .A1(n2653), .A2(n2505), .ZN(n2303) );
  INV_X1 U2804 ( .A(n4711), .ZN(n2324) );
  AND2_X1 U2805 ( .A1(n2337), .A2(n2276), .ZN(n2304) );
  OR2_X1 U2806 ( .A1(n3001), .A2(REG1_REG_17__SCAN_IN), .ZN(n2305) );
  OR2_X1 U2807 ( .A1(n2822), .A2(REG1_REG_13__SCAN_IN), .ZN(n2306) );
  OAI211_X1 U2808 ( .C1(n2400), .C2(n2318), .A(n2317), .B(n4703), .ZN(n2316)
         );
  NAND2_X1 U2809 ( .A1(n2400), .A2(n2318), .ZN(n2317) );
  INV_X1 U2810 ( .A(n4655), .ZN(n2318) );
  NAND3_X1 U2811 ( .A1(n2268), .A2(n4711), .A3(n4698), .ZN(n2320) );
  XNOR2_X1 U2812 ( .A(n2599), .B(n4845), .ZN(n4698) );
  OAI21_X1 U2813 ( .B1(n4728), .B2(n2326), .A(n2325), .ZN(n4299) );
  NOR2_X1 U2814 ( .A1(n4728), .A2(n2610), .ZN(n4281) );
  NAND2_X1 U2815 ( .A1(n2331), .A2(n2330), .ZN(n2591) );
  OR2_X1 U2816 ( .A1(n4668), .A2(n4664), .ZN(n2330) );
  NAND2_X1 U2817 ( .A1(n2332), .A2(n4665), .ZN(n2331) );
  NAND2_X1 U2818 ( .A1(n4668), .A2(n4664), .ZN(n2332) );
  NOR2_X1 U2819 ( .A1(n3121), .A2(n2588), .ZN(n4668) );
  OAI21_X1 U2820 ( .B1(n2573), .B2(n2335), .A(n2333), .ZN(n2578) );
  OAI21_X1 U2821 ( .B1(n3095), .B2(n3094), .A(n3102), .ZN(n3096) );
  NAND2_X1 U2822 ( .A1(n3330), .A2(n3089), .ZN(n2339) );
  INV_X1 U2823 ( .A(n2431), .ZN(n2352) );
  NAND2_X1 U2824 ( .A1(n2427), .A2(n2359), .ZN(n2358) );
  NAND2_X1 U2825 ( .A1(n2427), .A2(n2425), .ZN(n3726) );
  AOI21_X2 U2826 ( .B1(n3253), .B2(n3252), .A(n3251), .ZN(n3334) );
  INV_X2 U2827 ( .A(n2536), .ZN(n2515) );
  NAND3_X1 U2828 ( .A1(n2264), .A2(n2600), .A3(n2413), .ZN(n2536) );
  MUX2_X1 U2829 ( .A(n2432), .B(n2373), .S(n2716), .Z(n3084) );
  INV_X1 U2830 ( .A(n2375), .ZN(n4478) );
  NAND2_X1 U2831 ( .A1(n2984), .A2(n2381), .ZN(n2382) );
  NAND2_X1 U2832 ( .A1(n2984), .A2(n3914), .ZN(n4532) );
  INV_X1 U2833 ( .A(n2382), .ZN(n4531) );
  INV_X1 U2834 ( .A(n2386), .ZN(n4339) );
  NAND2_X1 U2835 ( .A1(n2387), .A2(n2935), .ZN(n3132) );
  OAI21_X1 U2836 ( .B1(n3872), .B2(n3234), .A(n2387), .ZN(n3238) );
  NOR2_X2 U2837 ( .A1(n4330), .A2(n4329), .ZN(n4328) );
  NAND2_X1 U2838 ( .A1(n2945), .A2(n3863), .ZN(n3482) );
  OR2_X1 U2839 ( .A1(n3049), .A2(n3084), .ZN(n3036) );
  AOI211_X2 U2840 ( .C1(n4493), .C2(n4321), .A(n4320), .B(n4319), .ZN(n4538)
         );
  INV_X1 U2841 ( .A(n2401), .ZN(n4644) );
  NOR2_X1 U2842 ( .A1(n2400), .A2(REG2_REG_7__SCAN_IN), .ZN(n2622) );
  XNOR2_X1 U2843 ( .A(n2621), .B(n4767), .ZN(n4645) );
  INV_X1 U2844 ( .A(n2632), .ZN(n2409) );
  INV_X1 U2845 ( .A(IR_REG_13__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U2846 ( .A1(n3838), .A2(n2423), .ZN(n2422) );
  INV_X1 U2847 ( .A(n3671), .ZN(n2427) );
  NOR2_X2 U2848 ( .A1(n3597), .A2(n2285), .ZN(n3253) );
  NOR2_X1 U2849 ( .A1(n3596), .A2(n2428), .ZN(n3597) );
  OR2_X1 U2850 ( .A1(n3599), .A2(n3595), .ZN(n2428) );
  NAND2_X1 U2851 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  NAND2_X1 U2852 ( .A1(n2542), .A2(n2429), .ZN(n2926) );
  NAND3_X1 U2853 ( .A1(n2549), .A2(n2537), .A3(n2506), .ZN(n2547) );
  INV_X1 U2854 ( .A(n2547), .ZN(n2540) );
  AND2_X2 U2855 ( .A1(n2662), .A2(n3005), .ZN(n2707) );
  NAND3_X1 U2856 ( .A1(n2289), .A2(n2434), .A3(n2433), .ZN(n2437) );
  NAND2_X1 U2857 ( .A1(n4310), .A2(n2436), .ZN(n2433) );
  INV_X1 U2858 ( .A(n4307), .ZN(n2450) );
  NAND2_X1 U2859 ( .A1(n2452), .A2(n2453), .ZN(n2784) );
  NAND2_X1 U2860 ( .A1(n2764), .A2(n2454), .ZN(n2452) );
  NAND2_X1 U2861 ( .A1(n3481), .A2(n2269), .ZN(n2458) );
  NAND3_X1 U2862 ( .A1(n2732), .A2(n2744), .A3(n3931), .ZN(n2470) );
  NOR2_X1 U2863 ( .A1(n4431), .A2(n4404), .ZN(n2486) );
  NAND3_X1 U2864 ( .A1(n2488), .A2(n2725), .A3(n2487), .ZN(n3208) );
  NAND2_X1 U2865 ( .A1(n2724), .A2(n2489), .ZN(n2487) );
  NAND3_X1 U2866 ( .A1(n3130), .A2(n2724), .A3(n3930), .ZN(n2488) );
  INV_X1 U2867 ( .A(n2490), .ZN(n3607) );
  XNOR2_X1 U2868 ( .A(n2623), .B(n2586), .ZN(n3126) );
  NAND2_X1 U2869 ( .A1(n3689), .A2(n3810), .ZN(n3773) );
  AOI22_X1 U2870 ( .A1(n3049), .A2(n3093), .B1(n3242), .B2(n3705), .ZN(n3053)
         );
  NAND4_X2 U2871 ( .A1(n2702), .A2(n2701), .A3(n2700), .A4(n2699), .ZN(n3049)
         );
  NAND2_X1 U2872 ( .A1(n3005), .A2(n3007), .ZN(n2706) );
  INV_X1 U2873 ( .A(n3005), .ZN(n2666) );
  INV_X1 U2874 ( .A(n4621), .ZN(n2988) );
  INV_X1 U2875 ( .A(n4585), .ZN(n2993) );
  AND2_X1 U2876 ( .A1(n3076), .A2(n4838), .ZN(n4891) );
  INV_X2 U2877 ( .A(n4836), .ZN(n4909) );
  INV_X1 U2878 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2774) );
  OR2_X1 U2879 ( .A1(n3673), .A2(n3672), .ZN(n2504) );
  OR2_X1 U2880 ( .A1(n4731), .A2(n3918), .ZN(n2505) );
  NAND2_X1 U2881 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U2882 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2507) );
  AND2_X1 U2883 ( .A1(n3632), .A2(n3787), .ZN(n2509) );
  OR2_X1 U2884 ( .A1(n3773), .A2(n3774), .ZN(n2510) );
  XNOR2_X1 U2885 ( .A(n2552), .B(IR_REG_10__SCAN_IN), .ZN(n4676) );
  INV_X1 U2886 ( .A(n2766), .ZN(n2920) );
  INV_X1 U2887 ( .A(n2635), .ZN(n4873) );
  INV_X1 U2888 ( .A(IR_REG_19__SCAN_IN), .ZN(n2512) );
  OR2_X1 U2889 ( .A1(n3140), .A2(n3415), .ZN(n3090) );
  AND2_X1 U2890 ( .A1(n2616), .A2(n4631), .ZN(n2617) );
  INV_X1 U2891 ( .A(n3341), .ZN(n3342) );
  AOI22_X1 U2892 ( .A1(n4224), .A2(n3701), .B1(n3706), .B2(n3463), .ZN(n3531)
         );
  INV_X1 U2893 ( .A(n3411), .ZN(n3412) );
  INV_X1 U2894 ( .A(n4676), .ZN(n2626) );
  NAND2_X1 U2895 ( .A1(n2823), .A2(n2295), .ZN(n2825) );
  INV_X1 U2896 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2797) );
  INV_X1 U2897 ( .A(n4789), .ZN(n2763) );
  INV_X1 U2898 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4165) );
  OR2_X1 U2899 ( .A1(n2535), .A2(n2508), .ZN(n2528) );
  AND2_X1 U2900 ( .A1(n3621), .A2(n3620), .ZN(n4864) );
  NOR2_X1 U2901 ( .A1(n2706), .A2(n2705), .ZN(n2712) );
  NOR2_X1 U2902 ( .A1(n2585), .A2(n2586), .ZN(n2588) );
  OAI22_X1 U2903 ( .A1(n4688), .A2(n2594), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4686), .ZN(n2599) );
  NAND2_X1 U2904 ( .A1(n2540), .A2(n2507), .ZN(n2545) );
  NAND2_X1 U2905 ( .A1(n2902), .A2(REG3_REG_24__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U2906 ( .A1(n2851), .A2(REG3_REG_17__SCAN_IN), .ZN(n2857) );
  OR2_X1 U2907 ( .A1(n4857), .A2(n3567), .ZN(n3864) );
  NOR2_X1 U2908 ( .A1(n2798), .A2(n2797), .ZN(n2806) );
  AND3_X1 U2909 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2734) );
  AND2_X1 U2910 ( .A1(n3585), .A2(DATAI_25_), .ZN(n3777) );
  INV_X1 U2911 ( .A(n2642), .ZN(n2644) );
  OR2_X1 U2912 ( .A1(n2580), .A2(n2551), .ZN(n2589) );
  NOR2_X1 U2913 ( .A1(n2671), .A2(n4108), .ZN(n2911) );
  NOR2_X1 U2914 ( .A1(n2901), .A2(n4165), .ZN(n2902) );
  OAI21_X1 U2915 ( .B1(n3346), .B2(n3345), .A(n3344), .ZN(n3368) );
  NAND2_X1 U2916 ( .A1(n3053), .A2(n2503), .ZN(n3081) );
  AOI21_X1 U2917 ( .B1(n4725), .B2(ADDR_REG_18__SCAN_IN), .A(n4294), .ZN(n4295) );
  AND2_X1 U2918 ( .A1(n4314), .A2(n3907), .ZN(n4337) );
  NAND2_X1 U2919 ( .A1(n3585), .A2(DATAI_26_), .ZN(n4359) );
  NAND2_X1 U2920 ( .A1(n3585), .A2(DATAI_22_), .ZN(n4428) );
  AND2_X1 U2921 ( .A1(n4625), .A2(n3991), .ZN(n3060) );
  OR2_X1 U2922 ( .A1(n2787), .A2(n4065), .ZN(n2798) );
  INV_X1 U2923 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2754) );
  INV_X1 U2924 ( .A(n4795), .ZN(n4471) );
  INV_X1 U2925 ( .A(n3011), .ZN(n2982) );
  INV_X1 U2926 ( .A(n4453), .ZN(n4458) );
  INV_X1 U2927 ( .A(n3478), .ZN(n3484) );
  INV_X1 U2928 ( .A(n4791), .ZN(n4513) );
  INV_X1 U2929 ( .A(IR_REG_23__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U2930 ( .A1(n2536), .A2(IR_REG_31__SCAN_IN), .ZN(n2549) );
  OR2_X1 U2931 ( .A1(n2665), .A2(n2911), .ZN(n4327) );
  OAI22_X1 U2932 ( .A1(n3088), .A2(n3087), .B1(n3086), .B2(n3085), .ZN(n3097)
         );
  OR2_X1 U2933 ( .A1(n3017), .A2(n4591), .ZN(n2667) );
  AND4_X1 U2934 ( .A1(n2908), .A2(n2907), .A3(n2906), .A4(n2905), .ZN(n4382)
         );
  NAND2_X1 U2935 ( .A1(n3126), .A2(REG2_REG_8__SCAN_IN), .ZN(n3125) );
  AND2_X1 U2936 ( .A1(n3022), .A2(n2649), .ZN(n4703) );
  INV_X1 U2937 ( .A(n4295), .ZN(n4296) );
  AND2_X1 U2938 ( .A1(n3074), .A2(n3073), .ZN(n3075) );
  NAND2_X1 U2939 ( .A1(n2960), .A2(n2959), .ZN(n4791) );
  INV_X1 U2940 ( .A(n4305), .ZN(n2994) );
  AOI21_X1 U2941 ( .B1(n2982), .B2(n3014), .A(n3013), .ZN(n3058) );
  NAND2_X1 U2942 ( .A1(n4474), .A2(n4741), .ZN(n4874) );
  INV_X1 U2943 ( .A(n4741), .ZN(n4853) );
  INV_X1 U2944 ( .A(IR_REG_30__SCAN_IN), .ZN(n3608) );
  AND2_X1 U2945 ( .A1(n2607), .A2(n2606), .ZN(n4275) );
  AND2_X1 U2946 ( .A1(n2652), .A2(n2651), .ZN(n4725) );
  NAND2_X1 U2947 ( .A1(n3072), .A2(n3065), .ZN(n4896) );
  OR2_X1 U2948 ( .A1(n3041), .A2(n2997), .ZN(n4011) );
  INV_X1 U2949 ( .A(n4382), .ZN(n4435) );
  INV_X1 U2950 ( .A(n4703), .ZN(n4719) );
  INV_X1 U2951 ( .A(n4726), .ZN(n4714) );
  NAND2_X1 U2952 ( .A1(n4836), .A2(n3240), .ZN(n4833) );
  NAND2_X2 U2953 ( .A1(n3075), .A2(n4853), .ZN(n4838) );
  NAND2_X1 U2954 ( .A1(n4526), .A2(n4783), .ZN(n4524) );
  NAND2_X1 U2955 ( .A1(n3216), .A2(n4838), .ZN(n4836) );
  NAND2_X1 U2956 ( .A1(n4885), .A2(n4878), .ZN(n4585) );
  AND2_X2 U2957 ( .A1(n2991), .A2(n3058), .ZN(n4885) );
  NAND2_X1 U2958 ( .A1(n2994), .A2(n2988), .ZN(n2989) );
  AND3_X1 U2959 ( .A1(n4882), .A2(n4881), .A3(n4880), .ZN(n4887) );
  NAND2_X1 U2960 ( .A1(n4888), .A2(n4878), .ZN(n4621) );
  AND2_X1 U2961 ( .A1(n4809), .A2(n4808), .ZN(n4811) );
  AND2_X2 U2962 ( .A1(n2991), .A2(n3215), .ZN(n4888) );
  AND2_X1 U2963 ( .A1(n3999), .A2(STATE_REG_SCAN_IN), .ZN(n3012) );
  XNOR2_X1 U2964 ( .A(n2648), .B(n2647), .ZN(n4908) );
  INV_X1 U2965 ( .A(n4686), .ZN(n4830) );
  INV_X1 U2966 ( .A(n4654), .ZN(n4776) );
  NAND2_X1 U2967 ( .A1(n2654), .A2(n2511), .ZN(U3259) );
  INV_X2 U2968 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2969 ( .A(n2527), .ZN(n2517) );
  NAND2_X1 U2970 ( .A1(n2524), .A2(n2523), .ZN(n2520) );
  NAND2_X1 U2971 ( .A1(n2520), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U2972 ( .A1(n2281), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  INV_X1 U2973 ( .A(n3074), .ZN(n3059) );
  INV_X1 U2974 ( .A(n3999), .ZN(n2525) );
  NAND2_X1 U2975 ( .A1(n2525), .A2(STATE_REG_SCAN_IN), .ZN(n4632) );
  NAND2_X1 U2976 ( .A1(n3059), .A2(n4632), .ZN(n2651) );
  NAND2_X1 U2977 ( .A1(n2527), .A2(n2526), .ZN(n2642) );
  NAND2_X1 U2978 ( .A1(n2647), .A2(n2643), .ZN(n2655) );
  NAND2_X1 U2979 ( .A1(n2530), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U2980 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U2981 ( .A1(n3999), .A2(n3060), .ZN(n2534) );
  XNOR2_X1 U2982 ( .A(n2535), .B(n2643), .ZN(n4002) );
  INV_X1 U2983 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4577) );
  NAND2_X1 U2984 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2537) );
  INV_X1 U2985 ( .A(n2538), .ZN(n2539) );
  NAND2_X1 U2986 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U2987 ( .A1(n2543), .A2(IR_REG_19__SCAN_IN), .ZN(n2544) );
  AND2_X2 U2988 ( .A1(n2926), .A2(n2544), .ZN(n4785) );
  MUX2_X1 U2989 ( .A(REG1_REG_19__SCAN_IN), .B(n4577), .S(n4785), .Z(n2613) );
  XNOR2_X1 U2990 ( .A(n2545), .B(IR_REG_18__SCAN_IN), .ZN(n4303) );
  XNOR2_X1 U2991 ( .A(n4303), .B(REG1_REG_18__SCAN_IN), .ZN(n4298) );
  INV_X1 U2992 ( .A(IR_REG_17__SCAN_IN), .ZN(n2546) );
  XNOR2_X1 U2993 ( .A(n2547), .B(n2546), .ZN(n3001) );
  OR2_X1 U2994 ( .A1(n2605), .A2(IR_REG_15__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U2995 ( .A1(n2607), .A2(IR_REG_31__SCAN_IN), .ZN(n2548) );
  XNOR2_X1 U2996 ( .A(n2548), .B(IR_REG_16__SCAN_IN), .ZN(n2635) );
  XNOR2_X1 U2997 ( .A(n2549), .B(IR_REG_14__SCAN_IN), .ZN(n4628) );
  INV_X1 U2998 ( .A(n2600), .ZN(n2575) );
  NAND2_X1 U2999 ( .A1(n2553), .A2(n4206), .ZN(n2580) );
  INV_X1 U3000 ( .A(n2550), .ZN(n2551) );
  NAND2_X1 U3001 ( .A1(n2593), .A2(IR_REG_31__SCAN_IN), .ZN(n2552) );
  NOR2_X1 U3002 ( .A1(n2553), .A2(n2645), .ZN(n2554) );
  MUX2_X1 U3003 ( .A(n2645), .B(n2554), .S(IR_REG_6__SCAN_IN), .Z(n2556) );
  INV_X1 U3004 ( .A(n2580), .ZN(n2555) );
  OR2_X1 U3005 ( .A1(n2560), .A2(n2645), .ZN(n2558) );
  INV_X1 U3006 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2559) );
  XNOR2_X1 U3007 ( .A(n4253), .B(n2559), .ZN(n4248) );
  INV_X1 U3008 ( .A(n4248), .ZN(n2565) );
  INV_X1 U3009 ( .A(n2560), .ZN(n2561) );
  INV_X1 U3010 ( .A(n4236), .ZN(n4232) );
  NAND2_X1 U3011 ( .A1(n4232), .A2(REG1_REG_1__SCAN_IN), .ZN(n2564) );
  INV_X1 U3012 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U3013 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n4237) );
  AOI21_X1 U3014 ( .B1(n4236), .B2(n4745), .A(n4237), .ZN(n2563) );
  NAND2_X1 U3015 ( .A1(n2564), .A2(n2563), .ZN(n4240) );
  NAND2_X1 U3016 ( .A1(n4240), .A2(n2564), .ZN(n4249) );
  NAND2_X1 U3017 ( .A1(n2566), .A2(IR_REG_31__SCAN_IN), .ZN(n2570) );
  XNOR2_X1 U3018 ( .A(n2570), .B(IR_REG_3__SCAN_IN), .ZN(n4631) );
  XNOR2_X1 U3019 ( .A(n2567), .B(n4631), .ZN(n3027) );
  INV_X1 U3020 ( .A(n2567), .ZN(n2568) );
  AOI22_X1 U3021 ( .A1(n3027), .A2(REG1_REG_3__SCAN_IN), .B1(n4631), .B2(n2568), .ZN(n2573) );
  NAND2_X1 U3022 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  NAND2_X1 U3023 ( .A1(n2571), .A2(IR_REG_31__SCAN_IN), .ZN(n2572) );
  XNOR2_X1 U3024 ( .A(n2572), .B(n4098), .ZN(n3158) );
  INV_X1 U3025 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U3026 ( .A1(n2575), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  XNOR2_X1 U3027 ( .A(n2576), .B(IR_REG_5__SCAN_IN), .ZN(n2743) );
  INV_X1 U3028 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2577) );
  INV_X1 U3029 ( .A(n2743), .ZN(n4765) );
  AOI22_X1 U3030 ( .A1(n2743), .A2(REG1_REG_5__SCAN_IN), .B1(n2577), .B2(n4765), .ZN(n4641) );
  NAND2_X1 U3031 ( .A1(n2752), .A2(n2578), .ZN(n2579) );
  XOR2_X1 U3032 ( .A(n2578), .B(n2752), .Z(n4650) );
  NAND2_X1 U3033 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U3034 ( .A1(n2579), .A2(n4649), .ZN(n4660) );
  NAND2_X1 U3035 ( .A1(n2580), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  XNOR2_X1 U3036 ( .A(n2582), .B(IR_REG_7__SCAN_IN), .ZN(n4654) );
  INV_X1 U3037 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4810) );
  NOR2_X1 U3038 ( .A1(n4776), .A2(n4810), .ZN(n4658) );
  OAI22_X1 U3039 ( .A1(n4660), .A2(n4658), .B1(n4654), .B2(REG1_REG_7__SCAN_IN), .ZN(n2585) );
  INV_X1 U3040 ( .A(IR_REG_7__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U3041 ( .A1(n2582), .A2(n2581), .ZN(n2583) );
  NAND2_X1 U3042 ( .A1(n2583), .A2(IR_REG_31__SCAN_IN), .ZN(n2584) );
  XNOR2_X1 U3043 ( .A(n2584), .B(IR_REG_8__SCAN_IN), .ZN(n4629) );
  INV_X1 U3044 ( .A(n4629), .ZN(n2586) );
  INV_X1 U3045 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4817) );
  AOI21_X1 U3046 ( .B1(n2586), .B2(n2585), .A(n2588), .ZN(n2587) );
  INV_X1 U3047 ( .A(n2587), .ZN(n3122) );
  NOR2_X1 U3048 ( .A1(n4817), .A2(n3122), .ZN(n3121) );
  INV_X1 U3049 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U3050 ( .A1(n2589), .A2(IR_REG_31__SCAN_IN), .ZN(n2590) );
  XNOR2_X1 U3051 ( .A(n2590), .B(IR_REG_9__SCAN_IN), .ZN(n4665) );
  INV_X1 U3052 ( .A(n4665), .ZN(n4820) );
  NAND2_X1 U3053 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U3054 ( .A1(n2591), .A2(n4676), .ZN(n2592) );
  OAI21_X1 U3055 ( .B1(n2593), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2596) );
  XNOR2_X1 U3056 ( .A(n2596), .B(IR_REG_11__SCAN_IN), .ZN(n4686) );
  AND2_X1 U3057 ( .A1(n4686), .A2(REG1_REG_11__SCAN_IN), .ZN(n2594) );
  INV_X1 U3058 ( .A(IR_REG_11__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U3059 ( .A1(n2596), .A2(n2595), .ZN(n2597) );
  NAND2_X1 U3060 ( .A1(n2597), .A2(IR_REG_31__SCAN_IN), .ZN(n2598) );
  XNOR2_X1 U3061 ( .A(n2598), .B(IR_REG_12__SCAN_IN), .ZN(n2813) );
  INV_X1 U3062 ( .A(n2813), .ZN(n4845) );
  INV_X1 U3063 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4699) );
  AND2_X1 U3064 ( .A1(n2264), .A2(n2600), .ZN(n2601) );
  OR2_X1 U3065 ( .A1(n2601), .A2(n2645), .ZN(n2602) );
  XNOR2_X1 U3066 ( .A(n2602), .B(IR_REG_13__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U3067 ( .A1(n2822), .A2(REG1_REG_13__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U3068 ( .A1(n4628), .A2(n2603), .ZN(n2604) );
  XOR2_X1 U3069 ( .A(n4628), .B(n2603), .Z(n4259) );
  NAND2_X1 U3070 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4259), .ZN(n4258) );
  NAND2_X1 U3071 ( .A1(n2605), .A2(IR_REG_15__SCAN_IN), .ZN(n2606) );
  INV_X1 U3072 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3579) );
  XNOR2_X1 U3073 ( .A(n4275), .B(n3579), .ZN(n4269) );
  NAND2_X1 U3074 ( .A1(n4275), .A2(REG1_REG_15__SCAN_IN), .ZN(n2608) );
  NOR2_X1 U3075 ( .A1(n2635), .A2(n2609), .ZN(n2610) );
  NOR2_X1 U3076 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4727), .ZN(n4728) );
  INV_X1 U3077 ( .A(n3001), .ZN(n4291) );
  INV_X1 U3078 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2611) );
  OAI21_X1 U3079 ( .B1(n4291), .B2(n2611), .A(n2305), .ZN(n4280) );
  INV_X1 U3080 ( .A(n4303), .ZN(n4627) );
  XNOR2_X1 U3081 ( .A(n2613), .B(n2612), .ZN(n2614) );
  NAND2_X1 U3082 ( .A1(n4726), .A2(n2614), .ZN(n2654) );
  NAND2_X1 U3083 ( .A1(n4686), .A2(REG2_REG_11__SCAN_IN), .ZN(n2629) );
  INV_X1 U3084 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4837) );
  AOI22_X1 U3085 ( .A1(n4686), .A2(REG2_REG_11__SCAN_IN), .B1(n4837), .B2(
        n4830), .ZN(n4694) );
  INV_X1 U3086 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U3087 ( .A1(n4665), .A2(REG2_REG_9__SCAN_IN), .B1(n3316), .B2(n4820), .ZN(n4673) );
  INV_X1 U3088 ( .A(n3158), .ZN(n4630) );
  XNOR2_X1 U3089 ( .A(n4236), .B(REG2_REG_1__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U3090 ( .A1(n4235), .A2(n4234), .ZN(n4233) );
  NAND2_X1 U3091 ( .A1(n4232), .A2(REG2_REG_1__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U3092 ( .A1(n4233), .A2(n2615), .ZN(n4246) );
  XNOR2_X1 U3093 ( .A(n2616), .B(n4631), .ZN(n3029) );
  INV_X1 U3094 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3030) );
  NOR2_X1 U3095 ( .A1(n3029), .A2(n3030), .ZN(n3028) );
  INV_X1 U3096 ( .A(n2618), .ZN(n2619) );
  NAND2_X1 U3097 ( .A1(n2743), .A2(REG2_REG_5__SCAN_IN), .ZN(n2620) );
  OAI21_X1 U3098 ( .B1(n2743), .B2(REG2_REG_5__SCAN_IN), .A(n2620), .ZN(n4636)
         );
  INV_X1 U3099 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4646) );
  INV_X1 U3100 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U3101 ( .A1(n2623), .A2(n4629), .ZN(n2624) );
  NAND2_X1 U3102 ( .A1(n4665), .A2(REG2_REG_9__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3103 ( .A1(n2627), .A2(n4676), .ZN(n2628) );
  NAND2_X1 U3104 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U3105 ( .A1(n2813), .A2(n2630), .ZN(n2631) );
  INV_X1 U3106 ( .A(n2822), .ZN(n4847) );
  INV_X1 U3107 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4708) );
  NOR2_X1 U3108 ( .A1(n4847), .A2(n4708), .ZN(n4707) );
  INV_X1 U3109 ( .A(n4628), .ZN(n4263) );
  INV_X1 U3110 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U3111 ( .A1(n4275), .A2(REG2_REG_15__SCAN_IN), .ZN(n2634) );
  OR2_X1 U3112 ( .A1(n4275), .A2(REG2_REG_15__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3113 ( .A1(n2634), .A2(n2633), .ZN(n4272) );
  NAND2_X1 U3114 ( .A1(n2636), .A2(n4873), .ZN(n2637) );
  INV_X1 U3115 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U3116 ( .A1(n4722), .A2(n4720), .ZN(n4721) );
  NAND2_X1 U3117 ( .A1(n2637), .A2(n4721), .ZN(n4283) );
  INV_X1 U3118 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3559) );
  XNOR2_X1 U3119 ( .A(n3001), .B(n3559), .ZN(n4285) );
  INV_X1 U3120 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2639) );
  NOR2_X1 U3121 ( .A1(n4627), .A2(n2639), .ZN(n2638) );
  AOI21_X1 U3122 ( .B1(n2639), .B2(n4627), .A(n2638), .ZN(n4292) );
  INV_X1 U3123 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2640) );
  MUX2_X1 U3124 ( .A(n2640), .B(REG2_REG_19__SCAN_IN), .S(n4785), .Z(n2641) );
  AND2_X1 U3125 ( .A1(n2644), .A2(n2643), .ZN(n2646) );
  OR2_X1 U3126 ( .A1(n2646), .A2(n2645), .ZN(n2648) );
  NOR2_X1 U3127 ( .A1(n4908), .A2(n4002), .ZN(n2649) );
  INV_X1 U3128 ( .A(n2650), .ZN(n2652) );
  AND2_X1 U3129 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3757) );
  AOI21_X1 U3130 ( .B1(n4725), .B2(ADDR_REG_19__SCAN_IN), .A(n3757), .ZN(n2653) );
  INV_X1 U3131 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2983) );
  INV_X1 U3132 ( .A(IR_REG_29__SCAN_IN), .ZN(n2656) );
  AND2_X1 U3133 ( .A1(n2656), .A2(n2659), .ZN(n2657) );
  NAND2_X1 U3134 ( .A1(n2931), .A2(REG1_REG_27__SCAN_IN), .ZN(n2670) );
  INV_X1 U3135 ( .A(n2662), .ZN(n3007) );
  INV_X1 U3136 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2663) );
  OR2_X1 U3137 ( .A1(n2786), .A2(n2663), .ZN(n2669) );
  NAND2_X1 U3138 ( .A1(n2734), .A2(REG3_REG_6__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U3139 ( .A1(n2767), .A2(REG3_REG_8__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3140 ( .A1(n2869), .A2(REG3_REG_19__SCAN_IN), .ZN(n2877) );
  INV_X1 U3141 ( .A(n2877), .ZN(n2664) );
  INV_X1 U3142 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3844) );
  INV_X1 U3143 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4108) );
  AND2_X1 U3144 ( .A1(n2671), .A2(n4108), .ZN(n2665) );
  INV_X1 U3145 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4591) );
  INV_X1 U3146 ( .A(n4350), .ZN(n4313) );
  NAND2_X1 U3147 ( .A1(n2931), .A2(REG1_REG_26__SCAN_IN), .ZN(n2677) );
  INV_X1 U31480 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4356) );
  OR2_X1 U31490 ( .A1(n2786), .A2(n4356), .ZN(n2676) );
  OAI21_X1 U3150 ( .B1(n2683), .B2(n4181), .A(n3844), .ZN(n2672) );
  NAND2_X1 U3151 ( .A1(n2672), .A2(n2671), .ZN(n4355) );
  INV_X1 U3152 ( .A(REG0_REG_26__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3153 ( .A1(n2931), .A2(REG1_REG_25__SCAN_IN), .ZN(n2681) );
  INV_X1 U3154 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4377) );
  OR2_X1 U3155 ( .A1(n2786), .A2(n4377), .ZN(n2680) );
  XNOR2_X1 U3156 ( .A(n2683), .B(n4181), .ZN(n4376) );
  OR2_X1 U3157 ( .A1(n2921), .A2(n4376), .ZN(n2679) );
  INV_X1 U3158 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4596) );
  OR2_X1 U3159 ( .A1(n3017), .A2(n4596), .ZN(n2678) );
  NAND2_X1 U3160 ( .A1(n2931), .A2(REG1_REG_24__SCAN_IN), .ZN(n2687) );
  INV_X1 U3161 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4396) );
  OR2_X1 U3162 ( .A1(n2900), .A2(n4396), .ZN(n2686) );
  OR2_X1 U3163 ( .A1(n2902), .A2(REG3_REG_24__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3164 ( .A1(n2683), .A2(n2682), .ZN(n4395) );
  OR2_X1 U3165 ( .A1(n2921), .A2(n4395), .ZN(n2685) );
  INV_X1 U3166 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4600) );
  OR2_X1 U3167 ( .A1(n3017), .A2(n4600), .ZN(n2684) );
  NAND4_X1 U3168 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2684), .ZN(n4416)
         );
  INV_X1 U3169 ( .A(n4416), .ZN(n4368) );
  INV_X1 U3170 ( .A(n3813), .ZN(n4393) );
  INV_X1 U3171 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2688) );
  OR2_X1 U3172 ( .A1(n2706), .A2(n2688), .ZN(n2694) );
  NAND2_X1 U3173 ( .A1(n2707), .A2(REG1_REG_1__SCAN_IN), .ZN(n2693) );
  INV_X1 U3174 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2689) );
  INV_X1 U3175 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2690) );
  NAND4_X1 U3176 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(n3040)
         );
  INV_X1 U3177 ( .A(DATAI_1_), .ZN(n2695) );
  NAND2_X1 U3178 ( .A1(n3040), .A2(n2703), .ZN(n3870) );
  INV_X1 U3179 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2697) );
  OR2_X1 U3180 ( .A1(n2706), .A2(n2697), .ZN(n2702) );
  INV_X1 U3181 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2698) );
  OR2_X1 U3182 ( .A1(n2709), .A2(n2698), .ZN(n2700) );
  NAND2_X1 U3183 ( .A1(n2707), .A2(REG1_REG_0__SCAN_IN), .ZN(n2699) );
  AND2_X1 U3184 ( .A1(n3049), .A2(n3242), .ZN(n3233) );
  NAND2_X1 U3185 ( .A1(n4231), .A2(n3243), .ZN(n2704) );
  INV_X1 U3186 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2705) );
  INV_X1 U3187 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U3188 ( .A1(n2707), .A2(REG1_REG_2__SCAN_IN), .ZN(n2708) );
  OAI21_X1 U3189 ( .B1(n2710), .B2(n2709), .A(n2708), .ZN(n2711) );
  NAND2_X2 U3190 ( .A1(n2715), .A2(n2714), .ZN(n3089) );
  INV_X1 U3191 ( .A(DATAI_2_), .ZN(n2717) );
  MUX2_X1 U3192 ( .A(n4253), .B(n2717), .S(n2716), .Z(n3140) );
  OR2_X1 U3193 ( .A1(n3089), .A2(n3140), .ZN(n3873) );
  NAND2_X1 U3194 ( .A1(n3089), .A2(n3140), .ZN(n3876) );
  NAND2_X1 U3195 ( .A1(n3873), .A2(n3876), .ZN(n3930) );
  INV_X1 U3196 ( .A(n3140), .ZN(n3133) );
  OR2_X1 U3197 ( .A1(n3089), .A2(n3133), .ZN(n2718) );
  OR2_X1 U3198 ( .A1(n2904), .A2(REG3_REG_3__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3199 ( .A1(n2707), .A2(REG1_REG_3__SCAN_IN), .ZN(n2719) );
  INV_X1 U3200 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2721) );
  OR2_X1 U3201 ( .A1(n3017), .A2(n2721), .ZN(n2723) );
  OR2_X1 U3202 ( .A1(n2786), .A2(n3030), .ZN(n2722) );
  MUX2_X1 U3203 ( .A(n4631), .B(DATAI_3_), .S(n2716), .Z(n3171) );
  NAND2_X1 U3204 ( .A1(n3105), .A2(n3171), .ZN(n2724) );
  OR2_X1 U3205 ( .A1(n3105), .A2(n3171), .ZN(n2725) );
  INV_X1 U3206 ( .A(n3208), .ZN(n2732) );
  NAND2_X1 U3207 ( .A1(n2707), .A2(REG1_REG_4__SCAN_IN), .ZN(n2731) );
  INV_X1 U3208 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2726) );
  OR2_X1 U3209 ( .A1(n2786), .A2(n2726), .ZN(n2730) );
  XNOR2_X1 U32100 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(
        n3604) );
  OR2_X1 U32110 ( .A1(n2904), .A2(n3604), .ZN(n2729) );
  INV_X1 U32120 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2727) );
  OR2_X1 U32130 ( .A1(n3017), .A2(n2727), .ZN(n2728) );
  INV_X1 U32140 ( .A(DATAI_4_), .ZN(n4145) );
  MUX2_X1 U32150 ( .A(n3158), .B(n4145), .S(n3585), .Z(n3227) );
  OR2_X1 U32160 ( .A1(n4230), .A2(n3227), .ZN(n3879) );
  NAND2_X1 U32170 ( .A1(n4230), .A2(n3227), .ZN(n3883) );
  INV_X1 U32180 ( .A(n3219), .ZN(n3931) );
  NAND2_X1 U32190 ( .A1(n4230), .A2(n3600), .ZN(n2733) );
  NAND2_X1 U32200 ( .A1(n2707), .A2(REG1_REG_5__SCAN_IN), .ZN(n2742) );
  INV_X1 U32210 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3267) );
  OR2_X1 U32220 ( .A1(n2786), .A2(n3267), .ZN(n2741) );
  INV_X1 U32230 ( .A(n2734), .ZN(n2745) );
  INV_X1 U32240 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U32250 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2735) );
  NAND2_X1 U32260 ( .A1(n2736), .A2(n2735), .ZN(n2737) );
  NAND2_X1 U32270 ( .A1(n2745), .A2(n2737), .ZN(n3266) );
  OR2_X1 U32280 ( .A1(n2921), .A2(n3266), .ZN(n2740) );
  INV_X1 U32290 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2738) );
  OR2_X1 U32300 ( .A1(n3017), .A2(n2738), .ZN(n2739) );
  NAND4_X1 U32310 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .ZN(n4229)
         );
  MUX2_X1 U32320 ( .A(n2743), .B(DATAI_5_), .S(n3585), .Z(n3202) );
  OR2_X1 U32330 ( .A1(n4229), .A2(n3202), .ZN(n2744) );
  NAND2_X1 U32340 ( .A1(n2707), .A2(REG1_REG_6__SCAN_IN), .ZN(n2751) );
  OR2_X1 U32350 ( .A1(n2786), .A2(n4646), .ZN(n2750) );
  INV_X1 U32360 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U32370 ( .A1(n2745), .A2(n3256), .ZN(n2746) );
  AND2_X1 U32380 ( .A1(n2746), .A2(n2755), .ZN(n4768) );
  INV_X1 U32390 ( .A(n4768), .ZN(n3259) );
  OR2_X1 U32400 ( .A1(n2921), .A2(n3259), .ZN(n2749) );
  INV_X1 U32410 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2747) );
  OR2_X1 U32420 ( .A1(n3017), .A2(n2747), .ZN(n2748) );
  NAND4_X1 U32430 ( .A1(n2751), .A2(n2750), .A3(n2749), .A4(n2748), .ZN(n4796)
         );
  MUX2_X1 U32440 ( .A(n2752), .B(DATAI_6_), .S(n3585), .Z(n3276) );
  AND2_X1 U32450 ( .A1(n4796), .A2(n3276), .ZN(n2753) );
  OAI22_X1 U32460 ( .A1(n3274), .A2(n2753), .B1(n3276), .B2(n4796), .ZN(n4780)
         );
  INV_X1 U32470 ( .A(n4780), .ZN(n2764) );
  NAND2_X1 U32480 ( .A1(n2931), .A2(REG1_REG_7__SCAN_IN), .ZN(n2761) );
  OR2_X1 U32490 ( .A1(n2786), .A2(n4653), .ZN(n2760) );
  AND2_X1 U32500 ( .A1(n2755), .A2(n2754), .ZN(n2756) );
  OR2_X1 U32510 ( .A1(n2756), .A2(n2767), .ZN(n4803) );
  OR2_X1 U32520 ( .A1(n2921), .A2(n4803), .ZN(n2759) );
  INV_X1 U32530 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2757) );
  OR2_X1 U32540 ( .A1(n3017), .A2(n2757), .ZN(n2758) );
  NAND4_X1 U32550 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n4228)
         );
  MUX2_X1 U32560 ( .A(n4654), .B(DATAI_7_), .S(n3585), .Z(n4793) );
  NAND2_X1 U32570 ( .A1(n4228), .A2(n4793), .ZN(n2765) );
  OR2_X1 U32580 ( .A1(n4228), .A2(n4793), .ZN(n2762) );
  NAND2_X1 U32590 ( .A1(n2765), .A2(n2762), .ZN(n4789) );
  NAND2_X1 U32600 ( .A1(n2931), .A2(REG1_REG_8__SCAN_IN), .ZN(n2773) );
  INV_X1 U32610 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3301) );
  OR2_X1 U32620 ( .A1(n2786), .A2(n3301), .ZN(n2772) );
  OR2_X1 U32630 ( .A1(n2767), .A2(REG3_REG_8__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U32640 ( .A1(n2775), .A2(n2768), .ZN(n3359) );
  OR2_X1 U32650 ( .A1(n2921), .A2(n3359), .ZN(n2771) );
  INV_X1 U32660 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2769) );
  OR2_X1 U32670 ( .A1(n3017), .A2(n2769), .ZN(n2770) );
  NAND4_X1 U32680 ( .A1(n2773), .A2(n2772), .A3(n2771), .A4(n2770), .ZN(n4786)
         );
  MUX2_X1 U32690 ( .A(n4629), .B(DATAI_8_), .S(n3585), .Z(n3355) );
  OR2_X1 U32700 ( .A1(n4786), .A2(n3355), .ZN(n3307) );
  NAND2_X1 U32710 ( .A1(n4786), .A2(n3355), .ZN(n3306) );
  NAND2_X1 U32720 ( .A1(n2931), .A2(REG1_REG_9__SCAN_IN), .ZN(n2781) );
  OR2_X1 U32730 ( .A1(n2786), .A2(n3316), .ZN(n2780) );
  NAND2_X1 U32740 ( .A1(n2775), .A2(n2774), .ZN(n2776) );
  NAND2_X1 U32750 ( .A1(n2787), .A2(n2776), .ZN(n3374) );
  OR2_X1 U32760 ( .A1(n2921), .A2(n3374), .ZN(n2779) );
  INV_X1 U32770 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2777) );
  OR2_X1 U32780 ( .A1(n3017), .A2(n2777), .ZN(n2778) );
  NAND4_X1 U32790 ( .A1(n2781), .A2(n2780), .A3(n2779), .A4(n2778), .ZN(n4227)
         );
  MUX2_X1 U32800 ( .A(n4665), .B(DATAI_9_), .S(n3585), .Z(n3371) );
  NAND2_X1 U32810 ( .A1(n4227), .A2(n3371), .ZN(n2782) );
  OR2_X1 U32820 ( .A1(n4227), .A2(n3371), .ZN(n2783) );
  NAND2_X1 U32830 ( .A1(n2784), .A2(n2783), .ZN(n3393) );
  NAND2_X1 U32840 ( .A1(n2931), .A2(REG1_REG_10__SCAN_IN), .ZN(n2793) );
  INV_X1 U32850 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2785) );
  OR2_X1 U32860 ( .A1(n2786), .A2(n2785), .ZN(n2792) );
  NAND2_X1 U32870 ( .A1(n2787), .A2(n4065), .ZN(n2788) );
  AND2_X1 U32880 ( .A1(n2798), .A2(n2788), .ZN(n4822) );
  INV_X1 U32890 ( .A(n4822), .ZN(n3741) );
  OR2_X1 U32900 ( .A1(n2921), .A2(n3741), .ZN(n2791) );
  INV_X1 U32910 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2789) );
  OR2_X1 U32920 ( .A1(n3017), .A2(n2789), .ZN(n2790) );
  NAND4_X1 U32930 ( .A1(n2793), .A2(n2792), .A3(n2791), .A4(n2790), .ZN(n4226)
         );
  MUX2_X1 U32940 ( .A(n4676), .B(DATAI_10_), .S(n3585), .Z(n3740) );
  NOR2_X1 U32950 ( .A1(n4226), .A2(n3740), .ZN(n2795) );
  NAND2_X1 U32960 ( .A1(n4226), .A2(n3740), .ZN(n2794) );
  OAI21_X1 U32970 ( .B1(n3393), .B2(n2795), .A(n2794), .ZN(n2796) );
  INV_X1 U32980 ( .A(n2796), .ZN(n3481) );
  NAND2_X1 U32990 ( .A1(n2931), .A2(REG1_REG_11__SCAN_IN), .ZN(n2803) );
  OR2_X1 U33000 ( .A1(n2900), .A2(n4837), .ZN(n2802) );
  AND2_X1 U33010 ( .A1(n2798), .A2(n2797), .ZN(n2799) );
  OR2_X1 U33020 ( .A1(n2799), .A2(n2806), .ZN(n4839) );
  OR2_X1 U33030 ( .A1(n2921), .A2(n4839), .ZN(n2801) );
  INV_X1 U33040 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3491) );
  OR2_X1 U33050 ( .A1(n3017), .A2(n3491), .ZN(n2800) );
  NAND4_X1 U33060 ( .A1(n2803), .A2(n2802), .A3(n2801), .A4(n2800), .ZN(n4225)
         );
  INV_X1 U33070 ( .A(DATAI_11_), .ZN(n2804) );
  MUX2_X1 U33080 ( .A(n4830), .B(n2804), .S(n3585), .Z(n3478) );
  OR2_X1 U33090 ( .A1(n4225), .A2(n3478), .ZN(n3378) );
  NAND2_X1 U33100 ( .A1(n4225), .A2(n3478), .ZN(n3380) );
  NAND2_X1 U33110 ( .A1(n3378), .A2(n3380), .ZN(n3927) );
  OR2_X1 U33120 ( .A1(n4225), .A2(n3484), .ZN(n2805) );
  NAND2_X1 U33130 ( .A1(n2931), .A2(REG1_REG_12__SCAN_IN), .ZN(n2812) );
  INV_X1 U33140 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3386) );
  OR2_X1 U33150 ( .A1(n2786), .A2(n3386), .ZN(n2811) );
  NOR2_X1 U33160 ( .A1(n2806), .A2(REG3_REG_12__SCAN_IN), .ZN(n2807) );
  OR2_X1 U33170 ( .A1(n2815), .A2(n2807), .ZN(n3466) );
  OR2_X1 U33180 ( .A1(n2921), .A2(n3466), .ZN(n2810) );
  INV_X1 U33190 ( .A(REG0_REG_12__SCAN_IN), .ZN(n2808) );
  OR2_X1 U33200 ( .A1(n3017), .A2(n2808), .ZN(n2809) );
  NAND4_X1 U33210 ( .A1(n2812), .A2(n2811), .A3(n2810), .A4(n2809), .ZN(n4224)
         );
  MUX2_X1 U33220 ( .A(n2813), .B(DATAI_12_), .S(n3585), .Z(n3463) );
  NAND2_X1 U33230 ( .A1(n4224), .A2(n3463), .ZN(n2814) );
  INV_X1 U33240 ( .A(n3429), .ZN(n2823) );
  NAND2_X1 U33250 ( .A1(n2931), .A2(REG1_REG_13__SCAN_IN), .ZN(n2821) );
  OR2_X1 U33260 ( .A1(n2786), .A2(n4708), .ZN(n2820) );
  NOR2_X1 U33270 ( .A1(n2815), .A2(REG3_REG_13__SCAN_IN), .ZN(n2816) );
  OR2_X1 U33280 ( .A1(n2826), .A2(n2816), .ZN(n3547) );
  OR2_X1 U33290 ( .A1(n2921), .A2(n3547), .ZN(n2819) );
  INV_X1 U33300 ( .A(REG0_REG_13__SCAN_IN), .ZN(n2817) );
  OR2_X1 U33310 ( .A1(n3017), .A2(n2817), .ZN(n2818) );
  NAND4_X1 U33320 ( .A1(n2821), .A2(n2820), .A3(n2819), .A4(n2818), .ZN(n4223)
         );
  MUX2_X1 U33330 ( .A(n2822), .B(DATAI_13_), .S(n3585), .Z(n3544) );
  NAND2_X1 U33340 ( .A1(n4223), .A2(n3544), .ZN(n2824) );
  NAND2_X1 U33350 ( .A1(n2931), .A2(REG1_REG_14__SCAN_IN), .ZN(n2831) );
  OR2_X1 U33360 ( .A1(n2900), .A2(n4265), .ZN(n2830) );
  OR2_X1 U33370 ( .A1(n2826), .A2(REG3_REG_14__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U33380 ( .A1(n2833), .A2(n2827), .ZN(n3573) );
  OR2_X1 U33390 ( .A1(n2921), .A2(n3573), .ZN(n2829) );
  INV_X1 U33400 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3509) );
  OR2_X1 U33410 ( .A1(n3017), .A2(n3509), .ZN(n2828) );
  NAND4_X1 U33420 ( .A1(n2831), .A2(n2830), .A3(n2829), .A4(n2828), .ZN(n4857)
         );
  MUX2_X1 U33430 ( .A(n4628), .B(DATAI_14_), .S(n3585), .Z(n3570) );
  NAND2_X1 U33440 ( .A1(n4857), .A2(n3567), .ZN(n3867) );
  NAND2_X1 U33450 ( .A1(n3864), .A2(n3867), .ZN(n3943) );
  NAND2_X1 U33460 ( .A1(n2931), .A2(REG1_REG_15__SCAN_IN), .ZN(n2838) );
  INV_X1 U33470 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3526) );
  OR2_X1 U33480 ( .A1(n2786), .A2(n3526), .ZN(n2837) );
  NAND2_X1 U33490 ( .A1(n2833), .A2(n2832), .ZN(n2834) );
  NAND2_X1 U33500 ( .A1(n2842), .A2(n2834), .ZN(n4871) );
  OR2_X1 U33510 ( .A1(n2921), .A2(n4871), .ZN(n2836) );
  INV_X1 U33520 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3582) );
  OR2_X1 U3353 ( .A1(n3017), .A2(n3582), .ZN(n2835) );
  NAND4_X1 U33540 ( .A1(n2838), .A2(n2837), .A3(n2836), .A4(n2835), .ZN(n4012)
         );
  MUX2_X1 U3355 ( .A(n4275), .B(DATAI_15_), .S(n3585), .Z(n4860) );
  NAND2_X1 U3356 ( .A1(n4012), .A2(n4860), .ZN(n2839) );
  NAND2_X1 U3357 ( .A1(n3943), .A2(n2839), .ZN(n2841) );
  NOR2_X1 U3358 ( .A1(n4857), .A2(n3570), .ZN(n3515) );
  INV_X1 U3359 ( .A(n4012), .ZN(n3496) );
  INV_X1 U3360 ( .A(n4860), .ZN(n3525) );
  AOI22_X1 U3361 ( .A1(n3515), .A2(n2839), .B1(n3496), .B2(n3525), .ZN(n2840)
         );
  NAND2_X1 U3362 ( .A1(n2931), .A2(REG1_REG_16__SCAN_IN), .ZN(n2849) );
  OR2_X1 U3363 ( .A1(n2900), .A2(n4720), .ZN(n2848) );
  NAND2_X1 U3364 ( .A1(n2842), .A2(n4184), .ZN(n2844) );
  INV_X1 U3365 ( .A(n2851), .ZN(n2843) );
  NAND2_X1 U3366 ( .A1(n2844), .A2(n2843), .ZN(n3794) );
  OR2_X1 U3367 ( .A1(n2904), .A2(n3794), .ZN(n2847) );
  INV_X1 U3368 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2845) );
  OR2_X1 U3369 ( .A1(n3017), .A2(n2845), .ZN(n2846) );
  NAND4_X1 U3370 ( .A1(n2849), .A2(n2848), .A3(n2847), .A4(n2846), .ZN(n4858)
         );
  INV_X1 U3371 ( .A(DATAI_16_), .ZN(n4872) );
  MUX2_X1 U3372 ( .A(n4873), .B(n4872), .S(n3585), .Z(n3628) );
  OR2_X1 U3373 ( .A1(n4858), .A2(n3628), .ZN(n3852) );
  NAND2_X1 U3374 ( .A1(n4858), .A2(n3628), .ZN(n3966) );
  NAND2_X1 U3375 ( .A1(n4858), .A2(n3791), .ZN(n2850) );
  NAND2_X1 U3376 ( .A1(n2931), .A2(REG1_REG_17__SCAN_IN), .ZN(n2855) );
  OR2_X1 U3377 ( .A1(n2900), .A2(n3559), .ZN(n2854) );
  OAI21_X1 U3378 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2851), .A(n2857), .ZN(n3805) );
  OR2_X1 U3379 ( .A1(n2921), .A2(n3805), .ZN(n2853) );
  INV_X1 U3380 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4619) );
  OR2_X1 U3381 ( .A1(n3017), .A2(n4619), .ZN(n2852) );
  NAND4_X1 U3382 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .ZN(n4517)
         );
  MUX2_X1 U3383 ( .A(n3001), .B(DATAI_17_), .S(n3585), .Z(n3802) );
  OR2_X1 U3384 ( .A1(n4517), .A2(n3802), .ZN(n2856) );
  NAND2_X1 U3385 ( .A1(n2931), .A2(REG1_REG_18__SCAN_IN), .ZN(n2864) );
  OR2_X1 U3386 ( .A1(n2900), .A2(n2639), .ZN(n2863) );
  INV_X1 U3387 ( .A(n2857), .ZN(n2859) );
  INV_X1 U3388 ( .A(n2869), .ZN(n2858) );
  OAI21_X1 U3389 ( .B1(REG3_REG_18__SCAN_IN), .B2(n2859), .A(n2858), .ZN(n4525) );
  OR2_X1 U3390 ( .A1(n2921), .A2(n4525), .ZN(n2862) );
  INV_X1 U3391 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2860) );
  OR2_X1 U3392 ( .A1(n3017), .A2(n2860), .ZN(n2861) );
  NAND4_X1 U3393 ( .A1(n2864), .A2(n2863), .A3(n2862), .A4(n2861), .ZN(n4495)
         );
  INV_X1 U3394 ( .A(DATAI_18_), .ZN(n2865) );
  MUX2_X1 U3395 ( .A(n4303), .B(n2865), .S(n3585), .Z(n4510) );
  OR2_X1 U3396 ( .A1(n4495), .A2(n4510), .ZN(n4490) );
  INV_X1 U3397 ( .A(n4490), .ZN(n2866) );
  AND2_X1 U3398 ( .A1(n4495), .A2(n4510), .ZN(n4489) );
  NOR2_X1 U3399 ( .A1(n2866), .A2(n4489), .ZN(n4523) );
  INV_X1 U3400 ( .A(n4523), .ZN(n3946) );
  NAND2_X1 U3401 ( .A1(n4517), .A2(n3802), .ZN(n4518) );
  AND2_X1 U3402 ( .A1(n3946), .A2(n4518), .ZN(n2867) );
  NAND2_X1 U3403 ( .A1(n4519), .A2(n2867), .ZN(n4520) );
  INV_X1 U3404 ( .A(n4510), .ZN(n3831) );
  OR2_X1 U3405 ( .A1(n4495), .A2(n3831), .ZN(n2868) );
  NAND2_X1 U3406 ( .A1(n4520), .A2(n2868), .ZN(n4485) );
  NAND2_X1 U3407 ( .A1(n2931), .A2(REG1_REG_19__SCAN_IN), .ZN(n2873) );
  OR2_X1 U3408 ( .A1(n2786), .A2(n2640), .ZN(n2872) );
  OAI21_X1 U3409 ( .B1(REG3_REG_19__SCAN_IN), .B2(n2869), .A(n2877), .ZN(n3758) );
  OR2_X1 U3410 ( .A1(n2904), .A2(n3758), .ZN(n2871) );
  INV_X1 U3411 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4614) );
  OR2_X1 U3412 ( .A1(n3017), .A2(n4614), .ZN(n2870) );
  NAND4_X1 U3413 ( .A1(n2873), .A2(n2872), .A3(n2871), .A4(n2870), .ZN(n4901)
         );
  MUX2_X1 U3414 ( .A(n4785), .B(DATAI_19_), .S(n3585), .Z(n4499) );
  NAND2_X1 U3415 ( .A1(n4901), .A2(n4499), .ZN(n2875) );
  NOR2_X1 U3416 ( .A1(n4901), .A2(n4499), .ZN(n2874) );
  NAND2_X1 U3417 ( .A1(n2931), .A2(REG1_REG_20__SCAN_IN), .ZN(n2883) );
  INV_X1 U3418 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4480) );
  OR2_X1 U3419 ( .A1(n2900), .A2(n4480), .ZN(n2882) );
  INV_X1 U3420 ( .A(n2876), .ZN(n2886) );
  INV_X1 U3421 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U3422 ( .A1(n4087), .A2(n2877), .ZN(n2878) );
  NAND2_X1 U3423 ( .A1(n2886), .A2(n2878), .ZN(n4905) );
  OR2_X1 U3424 ( .A1(n2921), .A2(n4905), .ZN(n2881) );
  INV_X1 U3425 ( .A(REG0_REG_20__SCAN_IN), .ZN(n2879) );
  OR2_X1 U3426 ( .A1(n3017), .A2(n2879), .ZN(n2880) );
  NAND2_X1 U3427 ( .A1(n4457), .A2(n4890), .ZN(n2884) );
  NAND2_X1 U3428 ( .A1(n2931), .A2(REG1_REG_21__SCAN_IN), .ZN(n2892) );
  INV_X1 U3429 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4462) );
  OR2_X1 U3430 ( .A1(n2900), .A2(n4462), .ZN(n2891) );
  INV_X1 U3431 ( .A(n2893), .ZN(n2888) );
  INV_X1 U3432 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2885) );
  NAND2_X1 U3433 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  NAND2_X1 U3434 ( .A1(n2888), .A2(n2887), .ZN(n4461) );
  OR2_X1 U3435 ( .A1(n2921), .A2(n4461), .ZN(n2890) );
  INV_X1 U3436 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4609) );
  OR2_X1 U3437 ( .A1(n3017), .A2(n4609), .ZN(n2889) );
  NAND4_X1 U3438 ( .A1(n2892), .A2(n2891), .A3(n2890), .A4(n2889), .ZN(n4889)
         );
  NAND2_X1 U3439 ( .A1(n4889), .A2(n4453), .ZN(n4403) );
  NAND2_X1 U3440 ( .A1(n2931), .A2(REG1_REG_22__SCAN_IN), .ZN(n2898) );
  INV_X1 U3441 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4443) );
  OR2_X1 U3442 ( .A1(n2786), .A2(n4443), .ZN(n2897) );
  OAI21_X1 U3443 ( .B1(n2893), .B2(REG3_REG_22__SCAN_IN), .A(n2901), .ZN(n4442) );
  OR2_X1 U3444 ( .A1(n2921), .A2(n4442), .ZN(n2896) );
  INV_X1 U3445 ( .A(REG0_REG_22__SCAN_IN), .ZN(n2894) );
  OR2_X1 U3446 ( .A1(n3017), .A2(n2894), .ZN(n2895) );
  NAND4_X1 U3447 ( .A1(n2898), .A2(n2897), .A3(n2896), .A4(n2895), .ZN(n4454)
         );
  AND2_X1 U3448 ( .A1(n4454), .A2(n4428), .ZN(n2956) );
  INV_X1 U3449 ( .A(n2956), .ZN(n2899) );
  OR2_X1 U3450 ( .A1(n4454), .A2(n4428), .ZN(n2933) );
  NOR2_X1 U3451 ( .A1(n4889), .A2(n4453), .ZN(n4404) );
  INV_X1 U3452 ( .A(n4454), .ZN(n4414) );
  NOR2_X1 U3453 ( .A1(n4414), .A2(n4428), .ZN(n4406) );
  NAND2_X1 U3454 ( .A1(n2931), .A2(REG1_REG_23__SCAN_IN), .ZN(n2908) );
  INV_X1 U3455 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4423) );
  OR2_X1 U3456 ( .A1(n2900), .A2(n4423), .ZN(n2907) );
  AND2_X1 U3457 ( .A1(n2901), .A2(n4165), .ZN(n2903) );
  OR2_X1 U34580 ( .A1(n2903), .A2(n2902), .ZN(n4422) );
  OR2_X1 U34590 ( .A1(n2904), .A2(n4422), .ZN(n2906) );
  INV_X1 U3460 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4604) );
  OR2_X1 U3461 ( .A1(n3017), .A2(n4604), .ZN(n2905) );
  NAND2_X1 U3462 ( .A1(n4382), .A2(n4413), .ZN(n3921) );
  NAND2_X1 U3463 ( .A1(n4435), .A2(n4419), .ZN(n3920) );
  AOI21_X1 U3464 ( .B1(n3813), .B2(n4416), .A(n4399), .ZN(n2909) );
  OAI21_X1 U3465 ( .B1(n4331), .B2(n4350), .A(n4338), .ZN(n2910) );
  OAI21_X1 U3466 ( .B1(n4313), .B2(n4340), .A(n2910), .ZN(n4310) );
  NAND2_X1 U34670 ( .A1(n2931), .A2(REG1_REG_28__SCAN_IN), .ZN(n2919) );
  INV_X1 U3468 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4323) );
  OR2_X1 U34690 ( .A1(n2786), .A2(n4323), .ZN(n2918) );
  NAND2_X1 U3470 ( .A1(n2911), .A2(REG3_REG_28__SCAN_IN), .ZN(n4304) );
  INV_X1 U34710 ( .A(n2911), .ZN(n2913) );
  INV_X1 U3472 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2912) );
  NAND2_X1 U34730 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  NAND2_X1 U3474 ( .A1(n4304), .A2(n2914), .ZN(n4322) );
  OR2_X1 U34750 ( .A1(n2921), .A2(n4322), .ZN(n2917) );
  INV_X1 U3476 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2915) );
  OR2_X1 U34770 ( .A1(n3017), .A2(n2915), .ZN(n2916) );
  NAND2_X1 U3478 ( .A1(n3585), .A2(DATAI_28_), .ZN(n4312) );
  OR2_X1 U34790 ( .A1(n4332), .A2(n4312), .ZN(n2958) );
  NAND2_X1 U3480 ( .A1(n4332), .A2(n4312), .ZN(n3909) );
  NAND2_X1 U34810 ( .A1(n2958), .A2(n3909), .ZN(n4316) );
  NAND2_X1 U3482 ( .A1(n2931), .A2(REG1_REG_29__SCAN_IN), .ZN(n2925) );
  NAND2_X1 U34830 ( .A1(n2920), .A2(REG2_REG_29__SCAN_IN), .ZN(n2924) );
  OR2_X1 U3484 ( .A1(n2921), .A2(n4304), .ZN(n2923) );
  OR2_X1 U34850 ( .A1(n3017), .A2(n2983), .ZN(n2922) );
  NAND4_X1 U3486 ( .A1(n2925), .A2(n2924), .A3(n2923), .A4(n2922), .ZN(n4321)
         );
  NAND2_X1 U34870 ( .A1(n3585), .A2(DATAI_29_), .ZN(n3914) );
  XNOR2_X1 U3488 ( .A(n4321), .B(n3914), .ZN(n3957) );
  XNOR2_X1 U34890 ( .A(n3217), .B(n4625), .ZN(n2929) );
  NAND2_X1 U3490 ( .A1(n2987), .A2(n4785), .ZN(n4734) );
  INV_X1 U34910 ( .A(n3017), .ZN(n2932) );
  AOI222_X1 U3492 ( .A1(n2920), .A2(REG2_REG_30__SCAN_IN), .B1(n2932), .B2(
        REG0_REG_30__SCAN_IN), .C1(n2931), .C2(REG1_REG_30__SCAN_IN), .ZN(
        n3851) );
  INV_X1 U34930 ( .A(B_REG_SCAN_IN), .ZN(n4004) );
  OAI21_X1 U3494 ( .B1(n4004), .B2(n4002), .A(n4493), .ZN(n3586) );
  INV_X1 U34950 ( .A(n2933), .ZN(n4410) );
  OR2_X1 U3496 ( .A1(n4889), .A2(n4458), .ZN(n4408) );
  INV_X1 U34970 ( .A(n4408), .ZN(n2934) );
  NOR2_X1 U3498 ( .A1(n4410), .A2(n2934), .ZN(n3977) );
  INV_X1 U34990 ( .A(n4499), .ZN(n3755) );
  AND2_X1 U3500 ( .A1(n4901), .A2(n3755), .ZN(n3941) );
  NOR2_X1 U35010 ( .A1(n4489), .A2(n3941), .ZN(n2955) );
  INV_X1 U3502 ( .A(n3802), .ZN(n3557) );
  NAND2_X1 U35030 ( .A1(n4517), .A2(n3557), .ZN(n4488) );
  NAND2_X1 U3504 ( .A1(n2955), .A2(n4488), .ZN(n3899) );
  INV_X1 U35050 ( .A(n3036), .ZN(n3872) );
  INV_X1 U35060 ( .A(n3930), .ZN(n3131) );
  NAND2_X1 U35070 ( .A1(n3132), .A2(n3131), .ZN(n2936) );
  NAND2_X1 U35080 ( .A1(n2936), .A2(n3873), .ZN(n3161) );
  INV_X1 U35090 ( .A(n3171), .ZN(n2937) );
  OR2_X1 U35100 ( .A1(n3105), .A2(n2937), .ZN(n3878) );
  NAND2_X1 U35110 ( .A1(n3105), .A2(n2937), .ZN(n3875) );
  NAND2_X1 U35120 ( .A1(n3878), .A2(n3875), .ZN(n3928) );
  INV_X1 U35130 ( .A(n3928), .ZN(n3162) );
  NAND2_X1 U35140 ( .A1(n3161), .A2(n3162), .ZN(n3160) );
  NAND2_X1 U35150 ( .A1(n3160), .A2(n3878), .ZN(n3220) );
  INV_X1 U35160 ( .A(n3879), .ZN(n2938) );
  INV_X1 U35170 ( .A(n3202), .ZN(n2940) );
  NAND2_X1 U35180 ( .A1(n4229), .A2(n2940), .ZN(n3881) );
  INV_X1 U35190 ( .A(n3881), .ZN(n2939) );
  OR2_X1 U35200 ( .A1(n4229), .A2(n2940), .ZN(n3856) );
  NAND2_X1 U35210 ( .A1(n4796), .A2(n3282), .ZN(n3882) );
  NAND2_X1 U35220 ( .A1(n3275), .A2(n3882), .ZN(n4788) );
  OR2_X1 U35230 ( .A1(n4796), .A2(n3282), .ZN(n4787) );
  INV_X1 U35240 ( .A(n4793), .ZN(n2942) );
  OR2_X1 U35250 ( .A1(n4228), .A2(n2942), .ZN(n2941) );
  AND2_X1 U35260 ( .A1(n4787), .A2(n2941), .ZN(n3886) );
  NAND2_X1 U35270 ( .A1(n4788), .A2(n3886), .ZN(n2943) );
  NAND2_X1 U35280 ( .A1(n4228), .A2(n2942), .ZN(n3853) );
  NAND2_X1 U35290 ( .A1(n2943), .A2(n3853), .ZN(n3292) );
  INV_X1 U35300 ( .A(n3355), .ZN(n3299) );
  OR2_X1 U35310 ( .A1(n4786), .A2(n3299), .ZN(n3889) );
  NAND2_X1 U35320 ( .A1(n3292), .A2(n3889), .ZN(n2944) );
  NAND2_X1 U35330 ( .A1(n4786), .A2(n3299), .ZN(n3854) );
  NAND2_X1 U35340 ( .A1(n4227), .A2(n3314), .ZN(n3855) );
  INV_X1 U35350 ( .A(n3855), .ZN(n3888) );
  OR2_X1 U35360 ( .A1(n4227), .A2(n3314), .ZN(n3890) );
  NAND2_X1 U35370 ( .A1(n4226), .A2(n3391), .ZN(n3859) );
  OR2_X1 U35380 ( .A1(n4226), .A2(n3391), .ZN(n3863) );
  INV_X1 U35390 ( .A(n3463), .ZN(n2947) );
  NAND2_X1 U35400 ( .A1(n4224), .A2(n2947), .ZN(n3430) );
  NAND2_X1 U35410 ( .A1(n4223), .A2(n3441), .ZN(n2946) );
  AND2_X1 U35420 ( .A1(n3430), .A2(n2946), .ZN(n2949) );
  AND2_X1 U35430 ( .A1(n2949), .A2(n3380), .ZN(n3860) );
  OR2_X1 U35440 ( .A1(n4224), .A2(n2947), .ZN(n3432) );
  NAND2_X1 U35450 ( .A1(n3378), .A2(n3432), .ZN(n2948) );
  NAND2_X1 U35460 ( .A1(n2949), .A2(n2948), .ZN(n2951) );
  OR2_X1 U35470 ( .A1(n4223), .A2(n3441), .ZN(n2950) );
  NAND2_X1 U35480 ( .A1(n2951), .A2(n2950), .ZN(n3865) );
  INV_X1 U35490 ( .A(n3864), .ZN(n3518) );
  OR2_X1 U35500 ( .A1(n4012), .A2(n3525), .ZN(n3869) );
  NAND2_X1 U35510 ( .A1(n4012), .A2(n3525), .ZN(n3868) );
  NAND2_X1 U35520 ( .A1(n3869), .A2(n3868), .ZN(n3938) );
  NOR3_X1 U35530 ( .A1(n3519), .A2(n3518), .A3(n3938), .ZN(n2953) );
  INV_X1 U35540 ( .A(n3868), .ZN(n2952) );
  NOR2_X1 U35550 ( .A1(n2953), .A2(n2952), .ZN(n3497) );
  NOR2_X1 U35560 ( .A1(n4457), .A2(n4479), .ZN(n3949) );
  OR2_X1 U35570 ( .A1(n4517), .A2(n3557), .ZN(n4486) );
  NAND2_X1 U35580 ( .A1(n4490), .A2(n4486), .ZN(n2954) );
  NOR2_X1 U35590 ( .A1(n4901), .A2(n3755), .ZN(n3940) );
  AOI21_X1 U35600 ( .B1(n2955), .B2(n2954), .A(n3940), .ZN(n4467) );
  NAND2_X1 U35610 ( .A1(n4457), .A2(n4479), .ZN(n3947) );
  AOI21_X1 U35620 ( .B1(n4467), .B2(n3947), .A(n3949), .ZN(n3971) );
  NAND2_X1 U35630 ( .A1(n4889), .A2(n4458), .ZN(n3951) );
  NOR2_X1 U35640 ( .A1(n4382), .A2(n4419), .ZN(n2957) );
  NOR2_X1 U35650 ( .A1(n2957), .A2(n2956), .ZN(n3903) );
  OAI21_X1 U35660 ( .B1(n4410), .B2(n3951), .A(n3903), .ZN(n3975) );
  NAND2_X1 U35670 ( .A1(n4382), .A2(n4419), .ZN(n4384) );
  NAND2_X1 U35680 ( .A1(n4368), .A2(n3813), .ZN(n3944) );
  NAND2_X1 U35690 ( .A1(n4384), .A2(n3944), .ZN(n3980) );
  NAND2_X1 U35700 ( .A1(n4416), .A2(n4393), .ZN(n4363) );
  NAND2_X1 U35710 ( .A1(n4390), .A2(n4373), .ZN(n3942) );
  NAND2_X1 U35720 ( .A1(n4363), .A2(n3942), .ZN(n3978) );
  OR2_X1 U35730 ( .A1(n4390), .A2(n4373), .ZN(n4348) );
  OR2_X1 U35740 ( .A1(n4370), .A2(n4359), .ZN(n3950) );
  NAND2_X1 U35750 ( .A1(n4348), .A2(n3950), .ZN(n3963) );
  NAND2_X1 U35760 ( .A1(n4370), .A2(n4359), .ZN(n3960) );
  OR2_X1 U35770 ( .A1(n4350), .A2(n4340), .ZN(n4314) );
  NAND2_X1 U35780 ( .A1(n4350), .A2(n4340), .ZN(n3907) );
  NAND2_X1 U35790 ( .A1(n4314), .A2(n2958), .ZN(n3964) );
  INV_X1 U35800 ( .A(n2987), .ZN(n4626) );
  NAND2_X1 U35810 ( .A1(n4626), .A2(n3991), .ZN(n2960) );
  OR2_X1 U3582 ( .A1(n3918), .A2(n4005), .ZN(n2959) );
  INV_X1 U3583 ( .A(n3060), .ZN(n2961) );
  NOR2_X2 U3584 ( .A1(n4908), .A2(n2961), .ZN(n4795) );
  INV_X1 U3585 ( .A(n3914), .ZN(n2985) );
  INV_X1 U3586 ( .A(n3991), .ZN(n3073) );
  AOI22_X1 U3587 ( .A1(n4332), .A2(n4795), .B1(n2985), .B2(n4794), .ZN(n2962)
         );
  NOR2_X1 U3588 ( .A1(n4741), .A2(n3991), .ZN(n2963) );
  NAND2_X1 U3589 ( .A1(n2987), .A2(n3918), .ZN(n3062) );
  NAND2_X1 U3590 ( .A1(n3062), .A2(n3060), .ZN(n3066) );
  NAND2_X1 U3591 ( .A1(n3074), .A2(n3066), .ZN(n3211) );
  NOR2_X1 U3592 ( .A1(n2963), .A2(n3211), .ZN(n2979) );
  INV_X1 U3593 ( .A(n3003), .ZN(n2967) );
  NAND2_X1 U3594 ( .A1(n2980), .A2(n2967), .ZN(n2964) );
  MUX2_X1 U3595 ( .A(n2980), .B(n2964), .S(B_REG_SCAN_IN), .Z(n2965) );
  INV_X1 U3596 ( .A(D_REG_1__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3597 ( .A1(n2982), .A2(n2966), .ZN(n3212) );
  INV_X1 U3598 ( .A(n4623), .ZN(n2981) );
  NAND2_X1 U3599 ( .A1(n2981), .A2(n2967), .ZN(n3056) );
  NAND2_X1 U3600 ( .A1(n3212), .A2(n3056), .ZN(n2978) );
  NOR4_X1 U3601 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2971) );
  NOR4_X1 U3602 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2970) );
  NOR4_X1 U3603 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2969) );
  NOR4_X1 U3604 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2968) );
  NAND4_X1 U3605 ( .A1(n2971), .A2(n2970), .A3(n2969), .A4(n2968), .ZN(n2977)
         );
  NOR2_X1 U3606 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_30__SCAN_IN), .ZN(n2975)
         );
  NOR4_X1 U3607 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2974) );
  NOR4_X1 U3608 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2973) );
  NOR4_X1 U3609 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2972) );
  NAND4_X1 U3610 ( .A1(n2975), .A2(n2974), .A3(n2973), .A4(n2972), .ZN(n2976)
         );
  OAI21_X1 U3611 ( .B1(n2977), .B2(n2976), .A(n2982), .ZN(n3057) );
  INV_X1 U3612 ( .A(D_REG_0__SCAN_IN), .ZN(n3014) );
  INV_X1 U3613 ( .A(n3058), .ZN(n3215) );
  NAND2_X1 U3614 ( .A1(n3241), .A2(n3140), .ZN(n3170) );
  OR2_X1 U3615 ( .A1(n3170), .A2(n3171), .ZN(n3169) );
  NAND2_X1 U3616 ( .A1(n3392), .A2(n3391), .ZN(n3476) );
  INV_X1 U3617 ( .A(n2984), .ZN(n4311) );
  NAND2_X1 U3618 ( .A1(n4311), .A2(n2985), .ZN(n2986) );
  NAND2_X1 U3619 ( .A1(n4532), .A2(n2986), .ZN(n4305) );
  NAND2_X1 U3620 ( .A1(n2990), .A2(n2989), .ZN(U3515) );
  INV_X1 U3621 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U3622 ( .A1(n2994), .A2(n2993), .ZN(n2995) );
  NAND2_X1 U3623 ( .A1(n2996), .A2(n2995), .ZN(U3547) );
  INV_X1 U3624 ( .A(n3012), .ZN(n2997) );
  MUX2_X1 U3625 ( .A(n4236), .B(n2695), .S(U3149), .Z(n2998) );
  INV_X1 U3626 ( .A(n2998), .ZN(U3351) );
  INV_X1 U3627 ( .A(DATAI_15_), .ZN(n4017) );
  NAND2_X1 U3628 ( .A1(n4275), .A2(STATE_REG_SCAN_IN), .ZN(n2999) );
  OAI21_X1 U3629 ( .B1(STATE_REG_SCAN_IN), .B2(n4017), .A(n2999), .ZN(U3337)
         );
  INV_X1 U3630 ( .A(DATAI_21_), .ZN(n4110) );
  NAND2_X1 U3631 ( .A1(n3991), .A2(STATE_REG_SCAN_IN), .ZN(n3000) );
  OAI21_X1 U3632 ( .B1(STATE_REG_SCAN_IN), .B2(n4110), .A(n3000), .ZN(U3331)
         );
  INV_X1 U3633 ( .A(DATAI_17_), .ZN(n4132) );
  NAND2_X1 U3634 ( .A1(n3001), .A2(STATE_REG_SCAN_IN), .ZN(n3002) );
  OAI21_X1 U3635 ( .B1(STATE_REG_SCAN_IN), .B2(n4132), .A(n3002), .ZN(U3335)
         );
  INV_X1 U3636 ( .A(DATAI_25_), .ZN(n4123) );
  NAND2_X1 U3637 ( .A1(n3003), .A2(STATE_REG_SCAN_IN), .ZN(n3004) );
  OAI21_X1 U3638 ( .B1(STATE_REG_SCAN_IN), .B2(n4123), .A(n3004), .ZN(U3327)
         );
  INV_X1 U3639 ( .A(DATAI_29_), .ZN(n4115) );
  NAND2_X1 U3640 ( .A1(n3005), .A2(STATE_REG_SCAN_IN), .ZN(n3006) );
  OAI21_X1 U3641 ( .B1(STATE_REG_SCAN_IN), .B2(n4115), .A(n3006), .ZN(U3323)
         );
  INV_X1 U3642 ( .A(DATAI_30_), .ZN(n3009) );
  NAND2_X1 U3643 ( .A1(n3007), .A2(STATE_REG_SCAN_IN), .ZN(n3008) );
  OAI21_X1 U3644 ( .B1(STATE_REG_SCAN_IN), .B2(n3009), .A(n3008), .ZN(U3322)
         );
  INV_X1 U3645 ( .A(DATAI_27_), .ZN(n4119) );
  INV_X1 U3646 ( .A(n4002), .ZN(n3020) );
  NAND2_X1 U3647 ( .A1(n3020), .A2(STATE_REG_SCAN_IN), .ZN(n3010) );
  OAI21_X1 U3648 ( .B1(STATE_REG_SCAN_IN), .B2(n4119), .A(n3010), .ZN(U3325)
         );
  AOI22_X1 U3649 ( .A1(n4634), .A2(n3014), .B1(n3013), .B2(n3012), .ZN(U3458)
         );
  INV_X1 U3650 ( .A(n4634), .ZN(n3016) );
  NAND2_X1 U3651 ( .A1(n3016), .A2(n3056), .ZN(n3015) );
  OAI21_X1 U3652 ( .B1(n3016), .B2(n2966), .A(n3015), .ZN(U3459) );
  NOR2_X1 U3653 ( .A1(n4725), .A2(U4043), .ZN(U3148) );
  AOI222_X1 U3654 ( .A1(n2920), .A2(REG2_REG_31__SCAN_IN), .B1(n2932), .B2(
        REG0_REG_31__SCAN_IN), .C1(n2707), .C2(REG1_REG_31__SCAN_IN), .ZN(
        n3987) );
  NAND2_X1 U3655 ( .A1(n4011), .A2(DATAO_REG_31__SCAN_IN), .ZN(n3018) );
  OAI21_X1 U3656 ( .B1(n3987), .B2(n4011), .A(n3018), .ZN(U3581) );
  INV_X1 U3657 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U3658 ( .A1(n4002), .A2(REG2_REG_0__SCAN_IN), .ZN(n3019) );
  NOR2_X1 U3659 ( .A1(n4908), .A2(n3019), .ZN(n3152) );
  OAI21_X1 U3660 ( .B1(REG1_REG_0__SCAN_IN), .B2(n3020), .A(n3152), .ZN(n3021)
         );
  MUX2_X1 U3661 ( .A(n3021), .B(n3152), .S(IR_REG_0__SCAN_IN), .Z(n3026) );
  INV_X1 U3662 ( .A(n3022), .ZN(n3025) );
  AOI22_X1 U3663 ( .A1(n4725), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3024) );
  INV_X1 U3664 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3048) );
  NAND3_X1 U3665 ( .A1(n4726), .A2(IR_REG_0__SCAN_IN), .A3(n3048), .ZN(n3023)
         );
  OAI211_X1 U3666 ( .C1(n3026), .C2(n3025), .A(n3024), .B(n3023), .ZN(U3240)
         );
  INV_X1 U3667 ( .A(n4631), .ZN(n3035) );
  XOR2_X1 U3668 ( .A(REG1_REG_3__SCAN_IN), .B(n3027), .Z(n3032) );
  AOI211_X1 U3669 ( .C1(n3030), .C2(n3029), .A(n3028), .B(n4719), .ZN(n3031)
         );
  AOI21_X1 U3670 ( .B1(n4726), .B2(n3032), .A(n3031), .ZN(n3034) );
  INV_X1 U3671 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U3672 ( .A1(STATE_REG_SCAN_IN), .A2(n4752), .ZN(n3114) );
  AOI21_X1 U3673 ( .B1(n4725), .B2(ADDR_REG_3__SCAN_IN), .A(n3114), .ZN(n3033)
         );
  OAI211_X1 U3674 ( .C1(n3035), .C2(n4731), .A(n3034), .B(n3033), .ZN(U3243)
         );
  NAND2_X1 U3675 ( .A1(n3049), .A2(n3084), .ZN(n3871) );
  NAND2_X1 U3676 ( .A1(n3036), .A2(n3871), .ZN(n4736) );
  INV_X1 U3677 ( .A(n3061), .ZN(n3037) );
  NOR2_X1 U3678 ( .A1(n3084), .A2(n3037), .ZN(n4735) );
  INV_X1 U3679 ( .A(n4231), .ZN(n3136) );
  INV_X1 U3680 ( .A(n4474), .ZN(n3483) );
  OAI21_X1 U3681 ( .B1(n3483), .B2(n4791), .A(n4736), .ZN(n3038) );
  OAI21_X1 U3682 ( .B1(n3136), .B2(n4799), .A(n3038), .ZN(n4733) );
  AOI211_X1 U3683 ( .C1(n4853), .C2(n4736), .A(n4735), .B(n4733), .ZN(n4732)
         );
  NAND2_X1 U3684 ( .A1(n4883), .A2(REG1_REG_0__SCAN_IN), .ZN(n3039) );
  OAI21_X1 U3685 ( .B1(n4732), .B2(n4883), .A(n3039), .ZN(U3518) );
  INV_X1 U3686 ( .A(n3042), .ZN(n3063) );
  AND2_X2 U3687 ( .A1(n3063), .A2(n3041), .ZN(n3093) );
  NAND2_X1 U3688 ( .A1(n3040), .A2(n3093), .ZN(n3044) );
  NAND2_X1 U3689 ( .A1(n3243), .A2(n3705), .ZN(n3043) );
  NAND2_X1 U3690 ( .A1(n3044), .A2(n3043), .ZN(n3046) );
  NAND2_X4 U3691 ( .A1(n3217), .A2(n3045), .ZN(n3707) );
  NOR2_X1 U3692 ( .A1(n2703), .A2(n3699), .ZN(n3047) );
  AOI21_X1 U3693 ( .B1(n3040), .B2(n3330), .A(n3047), .ZN(n3086) );
  XNOR2_X1 U3694 ( .A(n3085), .B(n3086), .ZN(n3088) );
  NAND2_X1 U3695 ( .A1(n3049), .A2(n3330), .ZN(n3052) );
  NOR2_X1 U3696 ( .A1(n3041), .A2(n2432), .ZN(n3050) );
  AOI21_X1 U3697 ( .B1(n3242), .B2(n3093), .A(n3050), .ZN(n3051) );
  NAND2_X1 U3698 ( .A1(n3052), .A2(n3051), .ZN(n3080) );
  NAND2_X1 U3699 ( .A1(n3081), .A2(n3080), .ZN(n3055) );
  INV_X2 U3700 ( .A(n3707), .ZN(n3697) );
  NAND2_X1 U3701 ( .A1(n3053), .A2(n3697), .ZN(n3054) );
  AND2_X1 U3702 ( .A1(n3055), .A2(n3054), .ZN(n3087) );
  XNOR2_X1 U3703 ( .A(n3088), .B(n3087), .ZN(n3079) );
  AND2_X1 U3704 ( .A1(n3057), .A2(n3056), .ZN(n3214) );
  NAND3_X1 U3705 ( .A1(n3214), .A2(n3058), .A3(n3212), .ZN(n3070) );
  NOR2_X1 U3706 ( .A1(n3070), .A2(n3059), .ZN(n3072) );
  AOI21_X1 U3707 ( .B1(n3062), .B2(n3061), .A(n3060), .ZN(n3065) );
  NAND3_X1 U3708 ( .A1(n3074), .A2(n3063), .A3(n4000), .ZN(n3068) );
  NOR2_X1 U3709 ( .A1(n3070), .A2(n3068), .ZN(n3064) );
  INV_X1 U3710 ( .A(n4908), .ZN(n3149) );
  AND2_X2 U3711 ( .A1(n3064), .A2(n3149), .ZN(n4902) );
  AND2_X2 U3712 ( .A1(n3064), .A2(n4908), .ZN(n4859) );
  AOI22_X1 U3713 ( .A1(n4902), .A2(n3049), .B1(n4859), .B2(n3089), .ZN(n3078)
         );
  NAND2_X1 U3714 ( .A1(n3070), .A2(n3065), .ZN(n3067) );
  NAND2_X1 U3715 ( .A1(n3067), .A2(n3066), .ZN(n3110) );
  INV_X1 U3716 ( .A(n3110), .ZN(n3071) );
  OAI21_X1 U3717 ( .B1(U3149), .B2(n4509), .A(n3068), .ZN(n3069) );
  NAND2_X1 U3718 ( .A1(n3070), .A2(n3069), .ZN(n3111) );
  NAND3_X1 U3719 ( .A1(n3071), .A2(n3074), .A3(n3111), .ZN(n3098) );
  NAND2_X1 U3720 ( .A1(n3072), .A2(n4794), .ZN(n3076) );
  AOI22_X1 U3721 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3098), .B1(n3843), .B2(n3243), .ZN(n3077) );
  OAI211_X1 U3722 ( .C1(n3079), .C2(n4896), .A(n3078), .B(n3077), .ZN(U3219)
         );
  XOR2_X1 U3723 ( .A(n3081), .B(n3080), .Z(n3148) );
  NAND2_X1 U3724 ( .A1(n3148), .A2(n4867), .ZN(n3083) );
  AOI22_X1 U3725 ( .A1(n3098), .A2(REG3_REG_0__SCAN_IN), .B1(n4859), .B2(n4231), .ZN(n3082) );
  OAI211_X1 U3726 ( .C1(n4891), .C2(n3084), .A(n3083), .B(n3082), .ZN(U3229)
         );
  NAND2_X1 U3727 ( .A1(n3089), .A2(n3093), .ZN(n3091) );
  NAND2_X1 U3728 ( .A1(n3091), .A2(n3090), .ZN(n3092) );
  NAND2_X1 U3729 ( .A1(n3095), .A2(n3094), .ZN(n3102) );
  AOI21_X1 U3730 ( .B1(n3097), .B2(n3096), .A(n3104), .ZN(n3101) );
  AOI22_X1 U3731 ( .A1(n4859), .A2(n3105), .B1(n4902), .B2(n4231), .ZN(n3100)
         );
  AOI22_X1 U3732 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3098), .B1(n3843), .B2(n3133), .ZN(n3099) );
  OAI211_X1 U3733 ( .C1(n3101), .C2(n4896), .A(n3100), .B(n3099), .ZN(U3234)
         );
  INV_X1 U3734 ( .A(n3102), .ZN(n3103) );
  AOI22_X1 U3735 ( .A1(n3105), .A2(n3701), .B1(n3706), .B2(n3171), .ZN(n3185)
         );
  NAND2_X1 U3736 ( .A1(n3171), .A2(n3705), .ZN(n3106) );
  XOR2_X1 U3737 ( .A(n3185), .B(n3187), .Z(n3107) );
  NOR2_X2 U3738 ( .A1(n3108), .A2(n3107), .ZN(n3596) );
  AOI21_X1 U3739 ( .B1(n3108), .B2(n3107), .A(n3596), .ZN(n3119) );
  INV_X1 U3740 ( .A(n3041), .ZN(n3109) );
  OAI21_X1 U3741 ( .B1(n3110), .B2(n3109), .A(STATE_REG_SCAN_IN), .ZN(n3113)
         );
  AND2_X1 U3742 ( .A1(n3111), .A2(n4632), .ZN(n3112) );
  AOI22_X1 U3743 ( .A1(n3171), .A2(n3843), .B1(n4859), .B2(n4230), .ZN(n3116)
         );
  AOI21_X1 U3744 ( .B1(n4902), .B2(n3089), .A(n3114), .ZN(n3115) );
  OAI211_X1 U3745 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4906), .A(n3116), .B(n3115), 
        .ZN(n3117) );
  INV_X1 U3746 ( .A(n3117), .ZN(n3118) );
  OAI21_X1 U3747 ( .B1(n3119), .B2(n4896), .A(n3118), .ZN(U3215) );
  INV_X1 U3748 ( .A(n4731), .ZN(n4276) );
  INV_X1 U3749 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4169) );
  NOR2_X1 U3750 ( .A1(STATE_REG_SCAN_IN), .A2(n4169), .ZN(n3356) );
  AOI21_X1 U3751 ( .B1(n4725), .B2(ADDR_REG_8__SCAN_IN), .A(n3356), .ZN(n3120)
         );
  INV_X1 U3752 ( .A(n3120), .ZN(n3124) );
  AOI211_X1 U3753 ( .C1(n4817), .C2(n3122), .A(n3121), .B(n4714), .ZN(n3123)
         );
  AOI211_X1 U3754 ( .C1(n4276), .C2(n4629), .A(n3124), .B(n3123), .ZN(n3128)
         );
  OAI211_X1 U3755 ( .C1(n3126), .C2(REG2_REG_8__SCAN_IN), .A(n4703), .B(n3125), 
        .ZN(n3127) );
  NAND2_X1 U3756 ( .A1(n3128), .A2(n3127), .ZN(U3248) );
  OAI21_X1 U3757 ( .B1(n3130), .B2(n3930), .A(n3129), .ZN(n4748) );
  XNOR2_X1 U3758 ( .A(n3132), .B(n3131), .ZN(n3138) );
  NAND2_X1 U3759 ( .A1(n4748), .A2(n3483), .ZN(n3135) );
  AOI22_X1 U3760 ( .A1(n4493), .A2(n3105), .B1(n3133), .B2(n4794), .ZN(n3134)
         );
  OAI211_X1 U3761 ( .C1(n3136), .C2(n4471), .A(n3135), .B(n3134), .ZN(n3137)
         );
  AOI21_X1 U3762 ( .B1(n3138), .B2(n4791), .A(n3137), .ZN(n4751) );
  INV_X1 U3763 ( .A(n4751), .ZN(n3139) );
  AOI21_X1 U3764 ( .B1(n4853), .B2(n4748), .A(n3139), .ZN(n3144) );
  OR2_X1 U3765 ( .A1(n3241), .A2(n3140), .ZN(n3141) );
  AND2_X1 U3766 ( .A1(n3170), .A2(n3141), .ZN(n4747) );
  AOI22_X1 U3767 ( .A1(n2993), .A2(n4747), .B1(REG1_REG_2__SCAN_IN), .B2(n4883), .ZN(n3142) );
  OAI21_X1 U3768 ( .B1(n3144), .B2(n4883), .A(n3142), .ZN(U3520) );
  AOI22_X1 U3769 ( .A1(n2988), .A2(n4747), .B1(REG0_REG_2__SCAN_IN), .B2(n4886), .ZN(n3143) );
  OAI21_X1 U3770 ( .B1(n3144), .B2(n4886), .A(n3143), .ZN(U3471) );
  INV_X1 U3771 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4193) );
  NOR2_X1 U3772 ( .A1(STATE_REG_SCAN_IN), .A2(n4193), .ZN(n3601) );
  OAI21_X1 U3773 ( .B1(REG2_REG_4__SCAN_IN), .B2(n3145), .A(n4703), .ZN(n3154)
         );
  XNOR2_X1 U3774 ( .A(REG1_REG_4__SCAN_IN), .B(n3146), .ZN(n3147) );
  NAND2_X1 U3775 ( .A1(n4726), .A2(n3147), .ZN(n3153) );
  NAND2_X1 U3776 ( .A1(n3148), .A2(n4002), .ZN(n3150) );
  OAI211_X1 U3777 ( .C1(n4234), .C2(n4002), .A(n3150), .B(n3149), .ZN(n3151)
         );
  OAI211_X1 U3778 ( .C1(IR_REG_0__SCAN_IN), .C2(n3152), .A(n3151), .B(U4043), 
        .ZN(n4257) );
  OAI211_X1 U3779 ( .C1(n3155), .C2(n3154), .A(n3153), .B(n4257), .ZN(n3156)
         );
  AOI211_X1 U3780 ( .C1(n4725), .C2(ADDR_REG_4__SCAN_IN), .A(n3601), .B(n3156), 
        .ZN(n3157) );
  OAI21_X1 U3781 ( .B1(n3158), .B2(n4731), .A(n3157), .ZN(U3244) );
  XNOR2_X1 U3782 ( .A(n3159), .B(n3928), .ZN(n4754) );
  INV_X1 U3783 ( .A(n3089), .ZN(n3166) );
  OAI21_X1 U3784 ( .B1(n3162), .B2(n3161), .A(n3160), .ZN(n3163) );
  NAND2_X1 U3785 ( .A1(n3163), .A2(n4791), .ZN(n3165) );
  AOI22_X1 U3786 ( .A1(n4493), .A2(n4230), .B1(n4794), .B2(n3171), .ZN(n3164)
         );
  OAI211_X1 U3787 ( .C1(n3166), .C2(n4471), .A(n3165), .B(n3164), .ZN(n3167)
         );
  AOI21_X1 U3788 ( .B1(n3483), .B2(n4754), .A(n3167), .ZN(n4757) );
  INV_X1 U3789 ( .A(n4757), .ZN(n3168) );
  AOI21_X1 U3790 ( .B1(n4853), .B2(n4754), .A(n3168), .ZN(n3174) );
  INV_X1 U3791 ( .A(n3169), .ZN(n3228) );
  AOI21_X1 U3792 ( .B1(n3171), .B2(n3170), .A(n3228), .ZN(n4753) );
  AOI22_X1 U3793 ( .A1(n4753), .A2(n2988), .B1(REG0_REG_3__SCAN_IN), .B2(n4886), .ZN(n3172) );
  OAI21_X1 U3794 ( .B1(n3174), .B2(n4886), .A(n3172), .ZN(U3473) );
  AOI22_X1 U3795 ( .A1(n4753), .A2(n2993), .B1(REG1_REG_3__SCAN_IN), .B2(n4883), .ZN(n3173) );
  OAI21_X1 U3796 ( .B1(n3174), .B2(n4883), .A(n3173), .ZN(U3521) );
  NAND2_X1 U3797 ( .A1(n3856), .A2(n3881), .ZN(n3925) );
  XOR2_X1 U3798 ( .A(n3175), .B(n3925), .Z(n3263) );
  XOR2_X1 U3799 ( .A(n3925), .B(n3176), .Z(n3179) );
  AOI22_X1 U3800 ( .A1(n4230), .A2(n4795), .B1(n3202), .B2(n4794), .ZN(n3178)
         );
  NAND2_X1 U3801 ( .A1(n4796), .A2(n4493), .ZN(n3177) );
  OAI211_X1 U3802 ( .C1(n3179), .C2(n4513), .A(n3178), .B(n3177), .ZN(n3265)
         );
  AOI21_X1 U3803 ( .B1(n3263), .B2(n4874), .A(n3265), .ZN(n3182) );
  AOI21_X1 U3804 ( .B1(n3202), .B2(n3226), .A(n3283), .ZN(n3270) );
  AOI22_X1 U3805 ( .A1(n3270), .A2(n2993), .B1(REG1_REG_5__SCAN_IN), .B2(n4883), .ZN(n3180) );
  OAI21_X1 U3806 ( .B1(n3182), .B2(n4883), .A(n3180), .ZN(U3523) );
  AOI22_X1 U3807 ( .A1(n3270), .A2(n2988), .B1(REG0_REG_5__SCAN_IN), .B2(n4886), .ZN(n3181) );
  OAI21_X1 U3808 ( .B1(n3182), .B2(n4886), .A(n3181), .ZN(U3477) );
  NOR2_X1 U3809 ( .A1(n3227), .A2(n3699), .ZN(n3183) );
  AOI21_X1 U3810 ( .B1(n4230), .B2(n3701), .A(n3183), .ZN(n3188) );
  INV_X1 U3811 ( .A(n3188), .ZN(n3191) );
  AOI22_X1 U3812 ( .A1(n4230), .A2(n3093), .B1(n3705), .B2(n3600), .ZN(n3184)
         );
  XNOR2_X1 U3813 ( .A(n3184), .B(n3707), .ZN(n3189) );
  INV_X1 U3814 ( .A(n3189), .ZN(n3190) );
  INV_X1 U3815 ( .A(n3185), .ZN(n3186) );
  NOR2_X1 U3816 ( .A1(n3187), .A2(n3186), .ZN(n3595) );
  XNOR2_X1 U3817 ( .A(n3189), .B(n3188), .ZN(n3599) );
  NAND2_X1 U3818 ( .A1(n4229), .A2(n3706), .ZN(n3193) );
  NAND2_X1 U3819 ( .A1(n3202), .A2(n3705), .ZN(n3192) );
  NAND2_X1 U3820 ( .A1(n3193), .A2(n3192), .ZN(n3194) );
  XNOR2_X1 U3821 ( .A(n3194), .B(n3697), .ZN(n3199) );
  INV_X1 U3822 ( .A(n3199), .ZN(n3197) );
  AND2_X1 U3823 ( .A1(n3202), .A2(n3706), .ZN(n3195) );
  AOI21_X1 U3824 ( .B1(n4229), .B2(n3701), .A(n3195), .ZN(n3198) );
  INV_X1 U3825 ( .A(n3198), .ZN(n3196) );
  NAND2_X1 U3826 ( .A1(n3197), .A2(n3196), .ZN(n3252) );
  INV_X1 U3827 ( .A(n3252), .ZN(n3200) );
  AND2_X1 U3828 ( .A1(n3199), .A2(n3198), .ZN(n3251) );
  NOR2_X1 U3829 ( .A1(n3200), .A2(n3251), .ZN(n3201) );
  XNOR2_X1 U3830 ( .A(n3253), .B(n3201), .ZN(n3206) );
  INV_X2 U3831 ( .A(n4891), .ZN(n3843) );
  AOI22_X1 U3832 ( .A1(n3202), .A2(n3843), .B1(n4902), .B2(n4230), .ZN(n3204)
         );
  AND2_X1 U3833 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4638) );
  AOI21_X1 U3834 ( .B1(n4859), .B2(n4796), .A(n4638), .ZN(n3203) );
  OAI211_X1 U3835 ( .C1(n4906), .C2(n3266), .A(n3204), .B(n3203), .ZN(n3205)
         );
  AOI21_X1 U3836 ( .B1(n3206), .B2(n4867), .A(n3205), .ZN(n3207) );
  INV_X1 U3837 ( .A(n3207), .ZN(U3224) );
  NAND2_X1 U3838 ( .A1(n3208), .A2(n3219), .ZN(n3209) );
  NAND2_X1 U3839 ( .A1(n3210), .A2(n3209), .ZN(n4758) );
  INV_X1 U3840 ( .A(n3211), .ZN(n3213) );
  NAND4_X1 U3841 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3216)
         );
  OR2_X1 U3842 ( .A1(n3217), .A2(n3918), .ZN(n3264) );
  INV_X1 U3843 ( .A(n3264), .ZN(n3218) );
  INV_X1 U3844 ( .A(n4825), .ZN(n4834) );
  XNOR2_X1 U3845 ( .A(n3220), .B(n3219), .ZN(n3224) );
  AOI22_X1 U3846 ( .A1(n3105), .A2(n4795), .B1(n3600), .B2(n4794), .ZN(n3222)
         );
  NAND2_X1 U3847 ( .A1(n4229), .A2(n4493), .ZN(n3221) );
  OAI211_X1 U3848 ( .C1(n4758), .C2(n4474), .A(n3222), .B(n3221), .ZN(n3223)
         );
  AOI21_X1 U3849 ( .B1(n3224), .B2(n4791), .A(n3223), .ZN(n3225) );
  INV_X1 U3850 ( .A(n3225), .ZN(n4760) );
  OAI211_X1 U3851 ( .C1(n3228), .C2(n3227), .A(n4878), .B(n3226), .ZN(n4759)
         );
  OAI22_X1 U3852 ( .A1(n4759), .A2(n4785), .B1(n4838), .B2(n3604), .ZN(n3229)
         );
  OAI21_X1 U3853 ( .B1(n4760), .B2(n3229), .A(n4526), .ZN(n3231) );
  NAND2_X1 U3854 ( .A1(n4909), .A2(REG2_REG_4__SCAN_IN), .ZN(n3230) );
  OAI211_X1 U3855 ( .C1(n4758), .C2(n4834), .A(n3231), .B(n3230), .ZN(U3286)
         );
  OAI21_X1 U3856 ( .B1(n3929), .B2(n3233), .A(n3232), .ZN(n4742) );
  NAND2_X1 U3857 ( .A1(n3049), .A2(n4795), .ZN(n3236) );
  NAND2_X1 U3858 ( .A1(n3089), .A2(n4493), .ZN(n3235) );
  OAI211_X1 U3859 ( .C1(n4509), .C2(n2703), .A(n3236), .B(n3235), .ZN(n3237)
         );
  AOI21_X1 U3860 ( .B1(n3238), .B2(n4791), .A(n3237), .ZN(n3239) );
  OAI21_X1 U3861 ( .B1(n4474), .B2(n4742), .A(n3239), .ZN(n4744) );
  INV_X1 U3862 ( .A(n4744), .ZN(n3250) );
  INV_X1 U3863 ( .A(n4742), .ZN(n3248) );
  AND2_X1 U3864 ( .A1(n4878), .A2(n3918), .ZN(n3240) );
  INV_X1 U3865 ( .A(n3241), .ZN(n3245) );
  NAND2_X1 U3866 ( .A1(n3243), .A2(n3242), .ZN(n3244) );
  NAND2_X1 U3867 ( .A1(n3245), .A2(n3244), .ZN(n4740) );
  INV_X1 U3868 ( .A(n4838), .ZN(n4821) );
  AOI22_X1 U3869 ( .A1(n4909), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4821), .ZN(n3246) );
  OAI21_X1 U3870 ( .B1(n4833), .B2(n4740), .A(n3246), .ZN(n3247) );
  AOI21_X1 U3871 ( .B1(n3248), .B2(n4825), .A(n3247), .ZN(n3249) );
  OAI21_X1 U3872 ( .B1(n3250), .B2(n4909), .A(n3249), .ZN(U3289) );
  AOI22_X1 U3873 ( .A1(n4796), .A2(n3706), .B1(n3705), .B2(n3276), .ZN(n3254)
         );
  XNOR2_X1 U3874 ( .A(n3254), .B(n3707), .ZN(n3332) );
  AOI22_X1 U3875 ( .A1(n4796), .A2(n3701), .B1(n3706), .B2(n3276), .ZN(n3333)
         );
  XNOR2_X1 U3876 ( .A(n3332), .B(n3333), .ZN(n3255) );
  XNOR2_X1 U3877 ( .A(n3334), .B(n3255), .ZN(n3261) );
  AOI22_X1 U3878 ( .A1(n3276), .A2(n3843), .B1(n4902), .B2(n4229), .ZN(n3258)
         );
  NOR2_X1 U3879 ( .A1(STATE_REG_SCAN_IN), .A2(n3256), .ZN(n4647) );
  AOI21_X1 U3880 ( .B1(n4859), .B2(n4228), .A(n4647), .ZN(n3257) );
  OAI211_X1 U3881 ( .C1(n4906), .C2(n3259), .A(n3258), .B(n3257), .ZN(n3260)
         );
  AOI21_X1 U3882 ( .B1(n3261), .B2(n4867), .A(n3260), .ZN(n3262) );
  INV_X1 U3883 ( .A(n3262), .ZN(U3236) );
  INV_X1 U3884 ( .A(n3263), .ZN(n3273) );
  NAND2_X1 U3885 ( .A1(n4474), .A2(n3264), .ZN(n4783) );
  NAND2_X1 U3886 ( .A1(n3265), .A2(n4836), .ZN(n3272) );
  NOR2_X1 U3887 ( .A1(n3266), .A2(n4838), .ZN(n3269) );
  NOR2_X1 U3888 ( .A1(n4836), .A2(n3267), .ZN(n3268) );
  AOI211_X1 U3889 ( .C1(n3270), .C2(n4910), .A(n3269), .B(n3268), .ZN(n3271)
         );
  OAI211_X1 U3890 ( .C1(n3273), .C2(n4524), .A(n3272), .B(n3271), .ZN(U3285)
         );
  NAND2_X1 U3891 ( .A1(n4787), .A2(n3882), .ZN(n3936) );
  XOR2_X1 U3892 ( .A(n3274), .B(n3936), .Z(n4771) );
  INV_X1 U3893 ( .A(n4771), .ZN(n3281) );
  XNOR2_X1 U3894 ( .A(n3275), .B(n3936), .ZN(n3279) );
  AOI22_X1 U3895 ( .A1(n4228), .A2(n4493), .B1(n3276), .B2(n4794), .ZN(n3278)
         );
  NAND2_X1 U3896 ( .A1(n4229), .A2(n4795), .ZN(n3277) );
  OAI211_X1 U3897 ( .C1(n3279), .C2(n4513), .A(n3278), .B(n3277), .ZN(n3280)
         );
  AOI21_X1 U3898 ( .B1(n3483), .B2(n4771), .A(n3280), .ZN(n4774) );
  OAI21_X1 U3899 ( .B1(n4741), .B2(n3281), .A(n4774), .ZN(n3289) );
  OR2_X1 U3900 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  NAND2_X1 U3901 ( .A1(n4777), .A2(n3284), .ZN(n4769) );
  OAI22_X1 U3902 ( .A1(n4769), .A2(n4621), .B1(n4888), .B2(n2747), .ZN(n3285)
         );
  AOI21_X1 U3903 ( .B1(n3289), .B2(n4888), .A(n3285), .ZN(n3286) );
  INV_X1 U3904 ( .A(n3286), .ZN(U3479) );
  INV_X1 U3905 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3287) );
  OAI22_X1 U3906 ( .A1(n4769), .A2(n4585), .B1(n4885), .B2(n3287), .ZN(n3288)
         );
  AOI21_X1 U3907 ( .B1(n3289), .B2(n4885), .A(n3288), .ZN(n3290) );
  INV_X1 U3908 ( .A(n3290), .ZN(U3524) );
  NAND2_X1 U3909 ( .A1(n3889), .A2(n3854), .ZN(n3926) );
  XNOR2_X1 U3910 ( .A(n3291), .B(n3926), .ZN(n3298) );
  XNOR2_X1 U3911 ( .A(n3292), .B(n3926), .ZN(n3296) );
  INV_X1 U3912 ( .A(n4227), .ZN(n3294) );
  AOI22_X1 U3913 ( .A1(n4228), .A2(n4795), .B1(n3355), .B2(n4794), .ZN(n3293)
         );
  OAI21_X1 U3914 ( .B1(n3294), .B2(n4799), .A(n3293), .ZN(n3295) );
  AOI21_X1 U3915 ( .B1(n3296), .B2(n4791), .A(n3295), .ZN(n3297) );
  OAI21_X1 U3916 ( .B1(n3298), .B2(n4474), .A(n3297), .ZN(n4814) );
  INV_X1 U3917 ( .A(n4814), .ZN(n3305) );
  INV_X1 U3918 ( .A(n3298), .ZN(n4816) );
  INV_X1 U3919 ( .A(n4778), .ZN(n3300) );
  NOR2_X1 U3920 ( .A1(n3300), .A2(n3299), .ZN(n4813) );
  NOR3_X1 U3921 ( .A1(n4813), .A2(n4812), .A3(n4833), .ZN(n3303) );
  OAI22_X1 U3922 ( .A1(n4526), .A2(n3301), .B1(n3359), .B2(n4838), .ZN(n3302)
         );
  AOI211_X1 U3923 ( .C1(n4816), .C2(n4825), .A(n3303), .B(n3302), .ZN(n3304)
         );
  OAI21_X1 U3924 ( .B1(n3305), .B2(n4909), .A(n3304), .ZN(U3282) );
  INV_X1 U3925 ( .A(n3306), .ZN(n3308) );
  OAI21_X1 U3926 ( .B1(n3291), .B2(n3308), .A(n3307), .ZN(n3309) );
  NAND2_X1 U3927 ( .A1(n3890), .A2(n3855), .ZN(n3937) );
  XNOR2_X1 U3928 ( .A(n3309), .B(n3937), .ZN(n3322) );
  INV_X1 U3929 ( .A(n3322), .ZN(n3320) );
  INV_X1 U3930 ( .A(n4226), .ZN(n3487) );
  XNOR2_X1 U3931 ( .A(n3310), .B(n3937), .ZN(n3311) );
  NAND2_X1 U3932 ( .A1(n3311), .A2(n4791), .ZN(n3313) );
  AOI22_X1 U3933 ( .A1(n4786), .A2(n4795), .B1(n4794), .B2(n3371), .ZN(n3312)
         );
  OAI211_X1 U3934 ( .C1(n3487), .C2(n4799), .A(n3313), .B(n3312), .ZN(n3321)
         );
  NOR2_X1 U3935 ( .A1(n4812), .A2(n3314), .ZN(n3315) );
  OR2_X1 U3936 ( .A1(n3392), .A2(n3315), .ZN(n3323) );
  NOR2_X1 U3937 ( .A1(n3323), .A2(n4833), .ZN(n3318) );
  OAI22_X1 U3938 ( .A1(n3374), .A2(n4838), .B1(n3316), .B2(n4526), .ZN(n3317)
         );
  AOI211_X1 U3939 ( .C1(n3321), .C2(n4526), .A(n3318), .B(n3317), .ZN(n3319)
         );
  OAI21_X1 U3940 ( .B1(n3320), .B2(n4524), .A(n3319), .ZN(U3281) );
  AOI21_X1 U3941 ( .B1(n4874), .B2(n3322), .A(n3321), .ZN(n3328) );
  INV_X1 U3942 ( .A(n3323), .ZN(n3325) );
  AOI22_X1 U3943 ( .A1(n3325), .A2(n2988), .B1(REG0_REG_9__SCAN_IN), .B2(n4886), .ZN(n3324) );
  OAI21_X1 U3944 ( .B1(n3328), .B2(n4886), .A(n3324), .ZN(U3485) );
  NAND2_X1 U3945 ( .A1(n4883), .A2(REG1_REG_9__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U3946 ( .A1(n3325), .A2(n2993), .ZN(n3326) );
  OAI211_X1 U3947 ( .C1(n3328), .C2(n4883), .A(n3327), .B(n3326), .ZN(U3527)
         );
  AOI22_X1 U3948 ( .A1(n4228), .A2(n3706), .B1(n3705), .B2(n4793), .ZN(n3329)
         );
  XNOR2_X1 U3949 ( .A(n3329), .B(n3707), .ZN(n3340) );
  AND2_X1 U3950 ( .A1(n4793), .A2(n3706), .ZN(n3331) );
  AOI21_X1 U3951 ( .B1(n4228), .B2(n3701), .A(n3331), .ZN(n3341) );
  XNOR2_X1 U3952 ( .A(n3340), .B(n3341), .ZN(n3345) );
  XOR2_X1 U3953 ( .A(n3345), .B(n3346), .Z(n3338) );
  AOI22_X1 U3954 ( .A1(n4793), .A2(n3843), .B1(n4902), .B2(n4796), .ZN(n3336)
         );
  NOR2_X1 U3955 ( .A1(STATE_REG_SCAN_IN), .A2(n2754), .ZN(n4656) );
  AOI21_X1 U3956 ( .B1(n4859), .B2(n4786), .A(n4656), .ZN(n3335) );
  OAI211_X1 U3957 ( .C1(n4906), .C2(n4803), .A(n3336), .B(n3335), .ZN(n3337)
         );
  AOI21_X1 U3958 ( .B1(n3338), .B2(n4867), .A(n3337), .ZN(n3339) );
  INV_X1 U3959 ( .A(n3339), .ZN(U3210) );
  INV_X1 U3960 ( .A(n3340), .ZN(n3343) );
  NAND2_X1 U3961 ( .A1(n3343), .A2(n3342), .ZN(n3344) );
  NAND2_X1 U3962 ( .A1(n4786), .A2(n3706), .ZN(n3348) );
  NAND2_X1 U3963 ( .A1(n3355), .A2(n3705), .ZN(n3347) );
  NAND2_X1 U3964 ( .A1(n3348), .A2(n3347), .ZN(n3349) );
  XNOR2_X1 U3965 ( .A(n3349), .B(n3697), .ZN(n3352) );
  AND2_X1 U3966 ( .A1(n3355), .A2(n3706), .ZN(n3350) );
  AOI21_X1 U3967 ( .B1(n4786), .B2(n3701), .A(n3350), .ZN(n3351) );
  NOR2_X1 U3968 ( .A1(n3352), .A2(n3351), .ZN(n3367) );
  INV_X1 U3969 ( .A(n3367), .ZN(n3353) );
  NAND2_X1 U3970 ( .A1(n3352), .A2(n3351), .ZN(n3366) );
  NAND2_X1 U3971 ( .A1(n3353), .A2(n3366), .ZN(n3354) );
  XNOR2_X1 U3972 ( .A(n3368), .B(n3354), .ZN(n3361) );
  AOI22_X1 U3973 ( .A1(n3355), .A2(n3843), .B1(n4859), .B2(n4227), .ZN(n3358)
         );
  AOI21_X1 U3974 ( .B1(n4902), .B2(n4228), .A(n3356), .ZN(n3357) );
  OAI211_X1 U3975 ( .C1(n4906), .C2(n3359), .A(n3358), .B(n3357), .ZN(n3360)
         );
  AOI21_X1 U3976 ( .B1(n3361), .B2(n4867), .A(n3360), .ZN(n3362) );
  INV_X1 U3977 ( .A(n3362), .ZN(U3218) );
  NAND2_X1 U3978 ( .A1(n4227), .A2(n3706), .ZN(n3364) );
  NAND2_X1 U3979 ( .A1(n3371), .A2(n3705), .ZN(n3363) );
  NAND2_X1 U3980 ( .A1(n3364), .A2(n3363), .ZN(n3365) );
  XNOR2_X1 U3981 ( .A(n3365), .B(n3707), .ZN(n3406) );
  AOI22_X1 U3982 ( .A1(n4227), .A2(n3701), .B1(n3706), .B2(n3371), .ZN(n3407)
         );
  XNOR2_X1 U3983 ( .A(n3406), .B(n3407), .ZN(n3370) );
  OAI21_X1 U3984 ( .B1(n3368), .B2(n3367), .A(n3366), .ZN(n3369) );
  NAND2_X1 U3985 ( .A1(n3369), .A2(n3370), .ZN(n3736) );
  OAI21_X1 U3986 ( .B1(n3370), .B2(n3369), .A(n3736), .ZN(n3376) );
  AOI22_X1 U3987 ( .A1(n3371), .A2(n3843), .B1(n4902), .B2(n4786), .ZN(n3373)
         );
  NOR2_X1 U3988 ( .A1(STATE_REG_SCAN_IN), .A2(n2774), .ZN(n4669) );
  AOI21_X1 U3989 ( .B1(n4859), .B2(n4226), .A(n4669), .ZN(n3372) );
  OAI211_X1 U3990 ( .C1(n4906), .C2(n3374), .A(n3373), .B(n3372), .ZN(n3375)
         );
  AOI21_X1 U3991 ( .B1(n3376), .B2(n4867), .A(n3375), .ZN(n3377) );
  INV_X1 U3992 ( .A(n3377), .ZN(U3228) );
  NAND2_X1 U3993 ( .A1(n3432), .A2(n3430), .ZN(n3923) );
  INV_X1 U3994 ( .A(n3378), .ZN(n3379) );
  AOI21_X1 U3995 ( .B1(n3482), .B2(n3380), .A(n3379), .ZN(n3433) );
  XOR2_X1 U3996 ( .A(n3923), .B(n3433), .Z(n3383) );
  AOI22_X1 U3997 ( .A1(n4223), .A2(n4493), .B1(n4794), .B2(n3463), .ZN(n3382)
         );
  NAND2_X1 U3998 ( .A1(n4225), .A2(n4795), .ZN(n3381) );
  OAI211_X1 U3999 ( .C1(n3383), .C2(n4513), .A(n3382), .B(n3381), .ZN(n3470)
         );
  INV_X1 U4000 ( .A(n3470), .ZN(n3390) );
  XNOR2_X1 U4001 ( .A(n3384), .B(n3923), .ZN(n3471) );
  INV_X1 U4002 ( .A(n4524), .ZN(n4446) );
  AND2_X1 U4003 ( .A1(n3477), .A2(n3463), .ZN(n3385) );
  OR2_X1 U4004 ( .A1(n3385), .A2(n3442), .ZN(n3475) );
  NOR2_X1 U4005 ( .A1(n3475), .A2(n4833), .ZN(n3388) );
  OAI22_X1 U4006 ( .A1(n4526), .A2(n3386), .B1(n3466), .B2(n4838), .ZN(n3387)
         );
  AOI211_X1 U4007 ( .C1(n3471), .C2(n4446), .A(n3388), .B(n3387), .ZN(n3389)
         );
  OAI21_X1 U4008 ( .B1(n3390), .B2(n4909), .A(n3389), .ZN(U3278) );
  OAI21_X1 U4009 ( .B1(n3392), .B2(n3391), .A(n3476), .ZN(n4823) );
  NAND2_X1 U4010 ( .A1(n3863), .A2(n3859), .ZN(n3922) );
  XNOR2_X1 U4011 ( .A(n3393), .B(n3922), .ZN(n4826) );
  XNOR2_X1 U4012 ( .A(n3394), .B(n3922), .ZN(n3397) );
  AOI22_X1 U4013 ( .A1(n4225), .A2(n4493), .B1(n4794), .B2(n3740), .ZN(n3396)
         );
  NAND2_X1 U4014 ( .A1(n4227), .A2(n4795), .ZN(n3395) );
  OAI211_X1 U4015 ( .C1(n3397), .C2(n4513), .A(n3396), .B(n3395), .ZN(n3398)
         );
  AOI21_X1 U4016 ( .B1(n3483), .B2(n4826), .A(n3398), .ZN(n4829) );
  INV_X1 U4017 ( .A(n4829), .ZN(n3399) );
  AOI21_X1 U4018 ( .B1(n4853), .B2(n4826), .A(n3399), .ZN(n3401) );
  MUX2_X1 U4019 ( .A(n2789), .B(n3401), .S(n4888), .Z(n3400) );
  OAI21_X1 U4020 ( .B1(n4823), .B2(n4621), .A(n3400), .ZN(U3487) );
  INV_X1 U4021 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3402) );
  MUX2_X1 U4022 ( .A(n3402), .B(n3401), .S(n4885), .Z(n3403) );
  OAI21_X1 U4023 ( .B1(n4823), .B2(n4585), .A(n3403), .ZN(U3528) );
  AND2_X1 U4024 ( .A1(n3740), .A2(n3706), .ZN(n3404) );
  AOI21_X1 U4025 ( .B1(n4226), .B2(n3701), .A(n3404), .ZN(n3411) );
  AOI22_X1 U4026 ( .A1(n4226), .A2(n3706), .B1(n3705), .B2(n3740), .ZN(n3405)
         );
  XNOR2_X1 U4027 ( .A(n3405), .B(n3707), .ZN(n3410) );
  XOR2_X1 U4028 ( .A(n3411), .B(n3410), .Z(n3738) );
  INV_X1 U4029 ( .A(n3406), .ZN(n3408) );
  NAND2_X1 U4030 ( .A1(n3408), .A2(n3407), .ZN(n3735) );
  NAND2_X1 U4031 ( .A1(n3736), .A2(n3409), .ZN(n3737) );
  INV_X1 U4032 ( .A(n3410), .ZN(n3413) );
  NAND2_X1 U4033 ( .A1(n3737), .A2(n3414), .ZN(n3459) );
  NAND2_X1 U4034 ( .A1(n4225), .A2(n3706), .ZN(n3417) );
  OR2_X1 U4035 ( .A1(n3478), .A2(n3415), .ZN(n3416) );
  NAND2_X1 U4036 ( .A1(n3417), .A2(n3416), .ZN(n3418) );
  XNOR2_X1 U4037 ( .A(n3418), .B(n3697), .ZN(n3421) );
  NOR2_X1 U4038 ( .A1(n3478), .A2(n3699), .ZN(n3419) );
  AOI21_X1 U4039 ( .B1(n4225), .B2(n3701), .A(n3419), .ZN(n3420) );
  OR2_X1 U4040 ( .A1(n3421), .A2(n3420), .ZN(n3460) );
  NAND2_X1 U4041 ( .A1(n2302), .A2(n3460), .ZN(n3422) );
  XNOR2_X1 U4042 ( .A(n3459), .B(n3422), .ZN(n3426) );
  AOI22_X1 U40430 ( .A1(n3484), .A2(n3843), .B1(n4902), .B2(n4226), .ZN(n3424)
         );
  AND2_X1 U4044 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4690) );
  AOI21_X1 U4045 ( .B1(n4859), .B2(n4224), .A(n4690), .ZN(n3423) );
  OAI211_X1 U4046 ( .C1(n4906), .C2(n4839), .A(n3424), .B(n3423), .ZN(n3425)
         );
  AOI21_X1 U4047 ( .B1(n3426), .B2(n4867), .A(n3425), .ZN(n3427) );
  INV_X1 U4048 ( .A(n3427), .ZN(U3233) );
  XNOR2_X1 U4049 ( .A(n4223), .B(n3441), .ZN(n3956) );
  INV_X1 U4050 ( .A(n3956), .ZN(n3428) );
  XNOR2_X1 U4051 ( .A(n3429), .B(n3428), .ZN(n3439) );
  INV_X1 U4052 ( .A(n3430), .ZN(n3431) );
  AOI21_X1 U4053 ( .B1(n3433), .B2(n3432), .A(n3431), .ZN(n3434) );
  XOR2_X1 U4054 ( .A(n3956), .B(n3434), .Z(n3437) );
  INV_X1 U4055 ( .A(n4857), .ZN(n3568) );
  AOI22_X1 U4056 ( .A1(n4224), .A2(n4795), .B1(n3544), .B2(n4794), .ZN(n3435)
         );
  OAI21_X1 U4057 ( .B1(n3568), .B2(n4799), .A(n3435), .ZN(n3436) );
  AOI21_X1 U4058 ( .B1(n3437), .B2(n4791), .A(n3436), .ZN(n3438) );
  OAI21_X1 U4059 ( .B1(n3439), .B2(n4474), .A(n3438), .ZN(n4850) );
  INV_X1 U4060 ( .A(n4850), .ZN(n3446) );
  INV_X1 U4061 ( .A(n3439), .ZN(n4852) );
  INV_X1 U4062 ( .A(n3454), .ZN(n3440) );
  OAI21_X1 U4063 ( .B1(n3442), .B2(n3441), .A(n3440), .ZN(n4849) );
  NOR2_X1 U4064 ( .A1(n4849), .A2(n4833), .ZN(n3444) );
  OAI22_X1 U4065 ( .A1(n4526), .A2(n4708), .B1(n3547), .B2(n4838), .ZN(n3443)
         );
  AOI211_X1 U4066 ( .C1(n4852), .C2(n4825), .A(n3444), .B(n3443), .ZN(n3445)
         );
  OAI21_X1 U4067 ( .B1(n3446), .B2(n4909), .A(n3445), .ZN(U3277) );
  INV_X1 U4068 ( .A(n3448), .ZN(n3450) );
  INV_X1 U4069 ( .A(n3943), .ZN(n3447) );
  NOR2_X1 U4070 ( .A1(n3448), .A2(n3447), .ZN(n3516) );
  INV_X1 U4071 ( .A(n3516), .ZN(n3449) );
  OAI21_X1 U4072 ( .B1(n3450), .B2(n3943), .A(n3449), .ZN(n3508) );
  INV_X1 U4073 ( .A(n3508), .ZN(n3458) );
  AOI21_X1 U4074 ( .B1(n3970), .B2(n3943), .A(n3519), .ZN(n3453) );
  OAI22_X1 U4075 ( .A1(n3496), .A2(n4799), .B1(n3567), .B2(n4509), .ZN(n3451)
         );
  AOI21_X1 U4076 ( .B1(n4795), .B2(n4223), .A(n3451), .ZN(n3452) );
  OAI21_X1 U4077 ( .B1(n3453), .B2(n4513), .A(n3452), .ZN(n3507) );
  OAI21_X1 U4078 ( .B1(n3454), .B2(n3567), .A(n3524), .ZN(n3514) );
  NOR2_X1 U4079 ( .A1(n3514), .A2(n4833), .ZN(n3456) );
  OAI22_X1 U4080 ( .A1(n4526), .A2(n4265), .B1(n3573), .B2(n4838), .ZN(n3455)
         );
  AOI211_X1 U4081 ( .C1(n3507), .C2(n4836), .A(n3456), .B(n3455), .ZN(n3457)
         );
  OAI21_X1 U4082 ( .B1(n3458), .B2(n4524), .A(n3457), .ZN(U3276) );
  AOI22_X1 U4083 ( .A1(n4224), .A2(n3706), .B1(n3705), .B2(n3463), .ZN(n3461)
         );
  XOR2_X1 U4084 ( .A(n3707), .B(n3461), .Z(n3532) );
  INV_X1 U4085 ( .A(n3531), .ZN(n3533) );
  XNOR2_X1 U4086 ( .A(n3532), .B(n3533), .ZN(n3462) );
  XNOR2_X1 U4087 ( .A(n3534), .B(n3462), .ZN(n3468) );
  AOI22_X1 U4088 ( .A1(n3463), .A2(n3843), .B1(n4902), .B2(n4225), .ZN(n3465)
         );
  INV_X1 U4089 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4179) );
  NOR2_X1 U4090 ( .A1(STATE_REG_SCAN_IN), .A2(n4179), .ZN(n4700) );
  AOI21_X1 U4091 ( .B1(n4859), .B2(n4223), .A(n4700), .ZN(n3464) );
  OAI211_X1 U4092 ( .C1(n4906), .C2(n3466), .A(n3465), .B(n3464), .ZN(n3467)
         );
  AOI21_X1 U4093 ( .B1(n3468), .B2(n4867), .A(n3467), .ZN(n3469) );
  INV_X1 U4094 ( .A(n3469), .ZN(U3221) );
  AOI21_X1 U4095 ( .B1(n4874), .B2(n3471), .A(n3470), .ZN(n3473) );
  MUX2_X1 U4096 ( .A(n2808), .B(n3473), .S(n4888), .Z(n3472) );
  OAI21_X1 U4097 ( .B1(n3475), .B2(n4621), .A(n3472), .ZN(U3491) );
  MUX2_X1 U4098 ( .A(n4699), .B(n3473), .S(n4885), .Z(n3474) );
  OAI21_X1 U4099 ( .B1(n3475), .B2(n4585), .A(n3474), .ZN(U3530) );
  INV_X1 U4100 ( .A(n3476), .ZN(n3479) );
  OAI21_X1 U4101 ( .B1(n3479), .B2(n3478), .A(n3477), .ZN(n4832) );
  OAI21_X1 U4102 ( .B1(n3481), .B2(n3927), .A(n3480), .ZN(n4831) );
  XOR2_X1 U4103 ( .A(n3482), .B(n3927), .Z(n3489) );
  NAND2_X1 U4104 ( .A1(n4831), .A2(n3483), .ZN(n3486) );
  AOI22_X1 U4105 ( .A1(n4224), .A2(n4493), .B1(n4794), .B2(n3484), .ZN(n3485)
         );
  OAI211_X1 U4106 ( .C1(n3487), .C2(n4471), .A(n3486), .B(n3485), .ZN(n3488)
         );
  AOI21_X1 U4107 ( .B1(n3489), .B2(n4791), .A(n3488), .ZN(n4843) );
  INV_X1 U4108 ( .A(n4843), .ZN(n3490) );
  AOI21_X1 U4109 ( .B1(n4853), .B2(n4831), .A(n3490), .ZN(n3493) );
  MUX2_X1 U4110 ( .A(n3491), .B(n3493), .S(n4888), .Z(n3492) );
  OAI21_X1 U4111 ( .B1(n4832), .B2(n4621), .A(n3492), .ZN(U3489) );
  INV_X1 U4112 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3494) );
  MUX2_X1 U4113 ( .A(n3494), .B(n3493), .S(n4885), .Z(n3495) );
  OAI21_X1 U4114 ( .B1(n4585), .B2(n4832), .A(n3495), .ZN(U3529) );
  OAI22_X1 U4115 ( .A1(n3496), .A2(n4471), .B1(n3628), .B2(n4509), .ZN(n3500)
         );
  XNOR2_X1 U4116 ( .A(n3497), .B(n2502), .ZN(n3498) );
  NOR2_X1 U4117 ( .A1(n3498), .A2(n4513), .ZN(n3499) );
  AOI211_X1 U4118 ( .C1(n4493), .C2(n4517), .A(n3500), .B(n3499), .ZN(n4882)
         );
  NAND2_X1 U4119 ( .A1(n2266), .A2(n3791), .ZN(n4877) );
  AND3_X1 U4120 ( .A1(n4879), .A2(n4910), .A3(n4877), .ZN(n3502) );
  OAI22_X1 U4121 ( .A1(n4526), .A2(n4720), .B1(n3794), .B2(n4838), .ZN(n3501)
         );
  NOR2_X1 U4122 ( .A1(n3502), .A2(n3501), .ZN(n3506) );
  NAND2_X1 U4123 ( .A1(n3504), .A2(n3503), .ZN(n4875) );
  NAND3_X1 U4124 ( .A1(n4876), .A2(n4875), .A3(n4446), .ZN(n3505) );
  OAI211_X1 U4125 ( .C1(n4882), .C2(n4909), .A(n3506), .B(n3505), .ZN(U3274)
         );
  AOI21_X1 U4126 ( .B1(n3508), .B2(n4874), .A(n3507), .ZN(n3511) );
  MUX2_X1 U4127 ( .A(n3509), .B(n3511), .S(n4888), .Z(n3510) );
  OAI21_X1 U4128 ( .B1(n3514), .B2(n4621), .A(n3510), .ZN(U3495) );
  INV_X1 U4129 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3512) );
  MUX2_X1 U4130 ( .A(n3512), .B(n3511), .S(n4885), .Z(n3513) );
  OAI21_X1 U4131 ( .B1(n4585), .B2(n3514), .A(n3513), .ZN(U3532) );
  NOR2_X1 U4132 ( .A1(n3516), .A2(n3515), .ZN(n3517) );
  XOR2_X1 U4133 ( .A(n3938), .B(n3517), .Z(n3578) );
  INV_X1 U4134 ( .A(n3578), .ZN(n3530) );
  NOR2_X1 U4135 ( .A1(n3519), .A2(n3518), .ZN(n3520) );
  XNOR2_X1 U4136 ( .A(n3520), .B(n3938), .ZN(n3521) );
  NAND2_X1 U4137 ( .A1(n3521), .A2(n4791), .ZN(n3523) );
  AOI22_X1 U4138 ( .A1(n4858), .A2(n4493), .B1(n4794), .B2(n4860), .ZN(n3522)
         );
  OAI211_X1 U4139 ( .C1(n3568), .C2(n4471), .A(n3523), .B(n3522), .ZN(n3577)
         );
  OAI21_X1 U4140 ( .B1(n2376), .B2(n3525), .A(n2266), .ZN(n3584) );
  NOR2_X1 U4141 ( .A1(n3584), .A2(n4833), .ZN(n3528) );
  OAI22_X1 U4142 ( .A1(n4526), .A2(n3526), .B1(n4871), .B2(n4838), .ZN(n3527)
         );
  AOI211_X1 U4143 ( .C1(n3577), .C2(n4836), .A(n3528), .B(n3527), .ZN(n3529)
         );
  OAI21_X1 U4144 ( .B1(n3530), .B2(n4524), .A(n3529), .ZN(U3275) );
  NAND2_X1 U4145 ( .A1(n4223), .A2(n3706), .ZN(n3536) );
  NAND2_X1 U4146 ( .A1(n3544), .A2(n3705), .ZN(n3535) );
  NAND2_X1 U4147 ( .A1(n3536), .A2(n3535), .ZN(n3537) );
  XNOR2_X1 U4148 ( .A(n3537), .B(n3697), .ZN(n3542) );
  INV_X1 U4149 ( .A(n3542), .ZN(n3540) );
  AND2_X1 U4150 ( .A1(n3544), .A2(n3706), .ZN(n3538) );
  AOI21_X1 U4151 ( .B1(n4223), .B2(n3701), .A(n3538), .ZN(n3541) );
  INV_X1 U4152 ( .A(n3541), .ZN(n3539) );
  AND2_X1 U4153 ( .A1(n3542), .A2(n3541), .ZN(n3564) );
  NOR2_X1 U4154 ( .A1(n2298), .A2(n3564), .ZN(n3543) );
  XNOR2_X1 U4155 ( .A(n3565), .B(n3543), .ZN(n3549) );
  AOI22_X1 U4156 ( .A1(n3544), .A2(n3843), .B1(n4902), .B2(n4224), .ZN(n3546)
         );
  INV_X1 U4157 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4200) );
  NOR2_X1 U4158 ( .A1(STATE_REG_SCAN_IN), .A2(n4200), .ZN(n4716) );
  AOI21_X1 U4159 ( .B1(n4859), .B2(n4857), .A(n4716), .ZN(n3545) );
  OAI211_X1 U4160 ( .C1(n4906), .C2(n3547), .A(n3546), .B(n3545), .ZN(n3548)
         );
  AOI21_X1 U4161 ( .B1(n3549), .B2(n4867), .A(n3548), .ZN(n3550) );
  INV_X1 U4162 ( .A(n3550), .ZN(U3231) );
  NAND2_X1 U4163 ( .A1(n4486), .A2(n4488), .ZN(n3945) );
  XOR2_X1 U4164 ( .A(n3945), .B(n3551), .Z(n4583) );
  INV_X1 U4165 ( .A(n4583), .ZN(n3563) );
  XNOR2_X1 U4166 ( .A(n2394), .B(n3945), .ZN(n3555) );
  INV_X1 U4167 ( .A(n4495), .ZN(n3753) );
  OAI22_X1 U4168 ( .A1(n3753), .A2(n4799), .B1(n4509), .B2(n3557), .ZN(n3553)
         );
  AOI21_X1 U4169 ( .B1(n4795), .B2(n4858), .A(n3553), .ZN(n3554) );
  OAI21_X1 U4170 ( .B1(n3555), .B2(n4513), .A(n3554), .ZN(n4582) );
  INV_X1 U4171 ( .A(n4879), .ZN(n3558) );
  INV_X1 U4172 ( .A(n4508), .ZN(n3556) );
  OAI21_X1 U4173 ( .B1(n3558), .B2(n3557), .A(n3556), .ZN(n4622) );
  NOR2_X1 U4174 ( .A1(n4622), .A2(n4833), .ZN(n3561) );
  OAI22_X1 U4175 ( .A1(n4526), .A2(n3559), .B1(n3805), .B2(n4838), .ZN(n3560)
         );
  AOI211_X1 U4176 ( .C1(n4582), .C2(n4836), .A(n3561), .B(n3560), .ZN(n3562)
         );
  OAI21_X1 U4177 ( .B1(n4524), .B2(n3563), .A(n3562), .ZN(U3273) );
  AOI22_X1 U4178 ( .A1(n4857), .A2(n3706), .B1(n3705), .B2(n3570), .ZN(n3566)
         );
  XOR2_X1 U4179 ( .A(n3707), .B(n3566), .Z(n3615) );
  INV_X1 U4180 ( .A(n3701), .ZN(n3677) );
  OAI22_X1 U4181 ( .A1(n3568), .A2(n3677), .B1(n3699), .B2(n3567), .ZN(n3616)
         );
  XNOR2_X1 U4182 ( .A(n3615), .B(n3616), .ZN(n3569) );
  XNOR2_X1 U4183 ( .A(n3617), .B(n3569), .ZN(n3575) );
  AOI22_X1 U4184 ( .A1(n3570), .A2(n3843), .B1(n4902), .B2(n4223), .ZN(n3572)
         );
  AND2_X1 U4185 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4260) );
  AOI21_X1 U4186 ( .B1(n4859), .B2(n4012), .A(n4260), .ZN(n3571) );
  OAI211_X1 U4187 ( .C1(n4906), .C2(n3573), .A(n3572), .B(n3571), .ZN(n3574)
         );
  AOI21_X1 U4188 ( .B1(n3575), .B2(n4867), .A(n3574), .ZN(n3576) );
  INV_X1 U4189 ( .A(n3576), .ZN(U3212) );
  AOI21_X1 U4190 ( .B1(n3578), .B2(n4874), .A(n3577), .ZN(n3581) );
  MUX2_X1 U4191 ( .A(n3579), .B(n3581), .S(n4885), .Z(n3580) );
  OAI21_X1 U4192 ( .B1(n4585), .B2(n3584), .A(n3580), .ZN(U3533) );
  MUX2_X1 U4193 ( .A(n3582), .B(n3581), .S(n4888), .Z(n3583) );
  OAI21_X1 U4194 ( .B1(n3584), .B2(n4621), .A(n3583), .ZN(U3497) );
  AND2_X1 U4195 ( .A1(n3585), .A2(DATAI_31_), .ZN(n3990) );
  NAND2_X1 U4196 ( .A1(n3585), .A2(DATAI_30_), .ZN(n3912) );
  NOR2_X1 U4197 ( .A1(n3987), .A2(n3586), .ZN(n4533) );
  AOI21_X1 U4198 ( .B1(n3990), .B2(n4794), .A(n4533), .ZN(n3591) );
  NOR2_X1 U4199 ( .A1(n3591), .A2(n4886), .ZN(n3587) );
  AOI21_X1 U4200 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4886), .A(n3587), .ZN(n3588) );
  OAI21_X1 U4201 ( .B1(n3594), .B2(n4621), .A(n3588), .ZN(U3517) );
  NOR2_X1 U4202 ( .A1(n3591), .A2(n4883), .ZN(n3589) );
  AOI21_X1 U4203 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4883), .A(n3589), .ZN(n3590) );
  OAI21_X1 U4204 ( .B1(n3594), .B2(n4585), .A(n3590), .ZN(U3549) );
  NOR2_X1 U4205 ( .A1(n3591), .A2(n4909), .ZN(n3592) );
  AOI21_X1 U4206 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4909), .A(n3592), .ZN(n3593) );
  OR2_X1 U4207 ( .A1(n3596), .A2(n3595), .ZN(n3598) );
  AOI211_X1 U4208 ( .C1(n3599), .C2(n3598), .A(n4896), .B(n3597), .ZN(n3606)
         );
  AOI22_X1 U4209 ( .A1(n3600), .A2(n3843), .B1(n4859), .B2(n4229), .ZN(n3603)
         );
  AOI21_X1 U4210 ( .B1(n4902), .B2(n3105), .A(n3601), .ZN(n3602) );
  OAI211_X1 U4211 ( .C1(n4906), .C2(n3604), .A(n3603), .B(n3602), .ZN(n3605)
         );
  OR2_X1 U4212 ( .A1(n3606), .A2(n3605), .ZN(U3227) );
  NAND3_X1 U4213 ( .A1(n3608), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3610) );
  INV_X1 U4214 ( .A(DATAI_31_), .ZN(n3609) );
  OAI22_X1 U4215 ( .A1(n3607), .A2(n3610), .B1(STATE_REG_SCAN_IN), .B2(n3609), 
        .ZN(U3321) );
  NAND2_X1 U4216 ( .A1(n4370), .A2(n3706), .ZN(n3612) );
  OR2_X1 U4217 ( .A1(n4359), .A2(n3415), .ZN(n3611) );
  NAND2_X1 U4218 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  XNOR2_X1 U4219 ( .A(n3613), .B(n3697), .ZN(n3694) );
  NOR2_X1 U4220 ( .A1(n4359), .A2(n3699), .ZN(n3614) );
  AOI21_X1 U4221 ( .B1(n4370), .B2(n3701), .A(n3614), .ZN(n3693) );
  NOR2_X1 U4222 ( .A1(n3694), .A2(n3693), .ZN(n3839) );
  NAND2_X1 U4223 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  NAND2_X1 U4224 ( .A1(n3619), .A2(n3618), .ZN(n3783) );
  NAND2_X1 U4225 ( .A1(n4012), .A2(n3701), .ZN(n3621) );
  NAND2_X1 U4226 ( .A1(n4860), .A2(n3706), .ZN(n3620) );
  NAND2_X1 U4227 ( .A1(n4012), .A2(n3706), .ZN(n3623) );
  NAND2_X1 U4228 ( .A1(n4860), .A2(n3705), .ZN(n3622) );
  NAND2_X1 U4229 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  XNOR2_X1 U4230 ( .A(n3624), .B(n3697), .ZN(n4865) );
  NAND2_X1 U4231 ( .A1(n4858), .A2(n3706), .ZN(n3626) );
  OR2_X1 U4232 ( .A1(n3628), .A2(n3415), .ZN(n3625) );
  NAND2_X1 U4233 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  XNOR2_X1 U4234 ( .A(n3627), .B(n3697), .ZN(n3631) );
  NOR2_X1 U4235 ( .A1(n3628), .A2(n3699), .ZN(n3629) );
  AOI21_X1 U4236 ( .B1(n4858), .B2(n3701), .A(n3629), .ZN(n3630) );
  OR2_X1 U4237 ( .A1(n3631), .A2(n3630), .ZN(n3788) );
  OAI21_X1 U4238 ( .B1(n4864), .B2(n4865), .A(n3788), .ZN(n3633) );
  NAND3_X1 U4239 ( .A1(n3788), .A2(n4864), .A3(n4865), .ZN(n3632) );
  NAND2_X1 U4240 ( .A1(n3631), .A2(n3630), .ZN(n3787) );
  NAND2_X1 U4241 ( .A1(n4517), .A2(n3706), .ZN(n3635) );
  NAND2_X1 U4242 ( .A1(n3802), .A2(n3705), .ZN(n3634) );
  NAND2_X1 U4243 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  XNOR2_X1 U4244 ( .A(n3636), .B(n3707), .ZN(n3639) );
  NAND2_X1 U4245 ( .A1(n4517), .A2(n3701), .ZN(n3638) );
  NAND2_X1 U4246 ( .A1(n3802), .A2(n3706), .ZN(n3637) );
  NAND2_X1 U4247 ( .A1(n3638), .A2(n3637), .ZN(n3640) );
  NAND2_X1 U4248 ( .A1(n3639), .A2(n3640), .ZN(n3799) );
  INV_X1 U4249 ( .A(n3639), .ZN(n3642) );
  INV_X1 U4250 ( .A(n3640), .ZN(n3641) );
  NAND2_X1 U4251 ( .A1(n3642), .A2(n3641), .ZN(n3798) );
  NAND2_X1 U4252 ( .A1(n4495), .A2(n3706), .ZN(n3644) );
  OR2_X1 U4253 ( .A1(n4510), .A2(n3415), .ZN(n3643) );
  NAND2_X1 U4254 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  XNOR2_X1 U4255 ( .A(n3645), .B(n3707), .ZN(n3827) );
  NAND2_X1 U4256 ( .A1(n4495), .A2(n3701), .ZN(n3647) );
  OR2_X1 U4257 ( .A1(n4510), .A2(n3699), .ZN(n3646) );
  NAND2_X1 U4258 ( .A1(n3647), .A2(n3646), .ZN(n3828) );
  NOR2_X1 U4259 ( .A1(n3827), .A2(n3828), .ZN(n3746) );
  NAND2_X1 U4260 ( .A1(n4901), .A2(n3706), .ZN(n3649) );
  NAND2_X1 U4261 ( .A1(n4499), .A2(n3705), .ZN(n3648) );
  NAND2_X1 U4262 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  XNOR2_X1 U4263 ( .A(n3650), .B(n3697), .ZN(n3655) );
  AND2_X1 U4264 ( .A1(n4499), .A2(n3706), .ZN(n3651) );
  AOI21_X1 U4265 ( .B1(n4901), .B2(n3701), .A(n3651), .ZN(n3654) );
  NAND2_X1 U4266 ( .A1(n3655), .A2(n3654), .ZN(n3653) );
  INV_X1 U4267 ( .A(n3653), .ZN(n3657) );
  OR2_X1 U4268 ( .A1(n3746), .A2(n3657), .ZN(n3652) );
  OAI21_X1 U4269 ( .B1(n3655), .B2(n3654), .A(n3653), .ZN(n3751) );
  INV_X1 U4270 ( .A(n3751), .ZN(n3656) );
  NAND2_X1 U4271 ( .A1(n3827), .A2(n3828), .ZN(n3747) );
  AND2_X1 U4272 ( .A1(n3656), .A2(n3747), .ZN(n3748) );
  NOR2_X1 U4273 ( .A1(n3657), .A2(n3748), .ZN(n3763) );
  OAI22_X1 U4274 ( .A1(n4457), .A2(n3699), .B1(n3415), .B2(n4890), .ZN(n3658)
         );
  XNOR2_X1 U4275 ( .A(n3658), .B(n3697), .ZN(n3669) );
  INV_X1 U4276 ( .A(n3669), .ZN(n3662) );
  OR2_X1 U4277 ( .A1(n4457), .A2(n3677), .ZN(n3660) );
  OR2_X1 U4278 ( .A1(n4890), .A2(n3699), .ZN(n3659) );
  AND2_X1 U4279 ( .A1(n3660), .A2(n3659), .ZN(n3668) );
  INV_X1 U4280 ( .A(n3668), .ZN(n3661) );
  NAND2_X1 U4281 ( .A1(n3662), .A2(n3661), .ZN(n4897) );
  NAND2_X1 U4282 ( .A1(n4889), .A2(n3701), .ZN(n3664) );
  NAND2_X1 U4283 ( .A1(n4453), .A2(n3706), .ZN(n3663) );
  NAND2_X1 U4284 ( .A1(n3664), .A2(n3663), .ZN(n3764) );
  NAND2_X1 U4285 ( .A1(n4889), .A2(n3706), .ZN(n3666) );
  NAND2_X1 U4286 ( .A1(n4453), .A2(n3705), .ZN(n3665) );
  NAND2_X1 U4287 ( .A1(n3666), .A2(n3665), .ZN(n3667) );
  XNOR2_X1 U4288 ( .A(n3667), .B(n3707), .ZN(n3765) );
  NAND2_X1 U4289 ( .A1(n3669), .A2(n3668), .ZN(n4894) );
  OAI21_X1 U4290 ( .B1(n3764), .B2(n3765), .A(n4894), .ZN(n3670) );
  INV_X1 U4291 ( .A(n3765), .ZN(n3673) );
  INV_X1 U4292 ( .A(n3764), .ZN(n3672) );
  OAI22_X1 U4293 ( .A1(n4414), .A2(n3699), .B1(n3415), .B2(n4428), .ZN(n3674)
         );
  XNOR2_X1 U4294 ( .A(n3674), .B(n3707), .ZN(n3681) );
  OAI22_X1 U4295 ( .A1(n4414), .A2(n3677), .B1(n3699), .B2(n4428), .ZN(n3680)
         );
  XNOR2_X1 U4296 ( .A(n3681), .B(n3680), .ZN(n3821) );
  OAI22_X1 U4297 ( .A1(n4382), .A2(n3699), .B1(n3415), .B2(n4413), .ZN(n3676)
         );
  XNOR2_X1 U4298 ( .A(n3676), .B(n3707), .ZN(n3684) );
  OR2_X1 U4299 ( .A1(n4382), .A2(n3677), .ZN(n3679) );
  OR2_X1 U4300 ( .A1(n4413), .A2(n3699), .ZN(n3678) );
  NAND2_X1 U4301 ( .A1(n3679), .A2(n3678), .ZN(n3683) );
  XNOR2_X1 U4302 ( .A(n3684), .B(n3683), .ZN(n3727) );
  NOR2_X1 U4303 ( .A1(n3681), .A2(n3680), .ZN(n3728) );
  NOR2_X1 U4304 ( .A1(n3727), .A2(n3728), .ZN(n3682) );
  NAND2_X1 U4305 ( .A1(n3684), .A2(n3683), .ZN(n3688) );
  NAND2_X1 U4306 ( .A1(n4416), .A2(n3706), .ZN(n3686) );
  NAND2_X1 U4307 ( .A1(n3813), .A2(n3705), .ZN(n3685) );
  NAND2_X1 U4308 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  AOI22_X1 U4309 ( .A1(n4416), .A2(n3701), .B1(n3706), .B2(n3813), .ZN(n3812)
         );
  NAND2_X1 U4310 ( .A1(n3809), .A2(n3812), .ZN(n3689) );
  NAND3_X1 U4311 ( .A1(n3729), .A2(n2293), .A3(n3688), .ZN(n3810) );
  OAI22_X1 U4312 ( .A1(n2468), .A2(n3699), .B1(n3415), .B2(n4373), .ZN(n3690)
         );
  XOR2_X1 U4313 ( .A(n3707), .B(n3690), .Z(n3774) );
  AOI22_X1 U4314 ( .A1(n4390), .A2(n3701), .B1(n3706), .B2(n3777), .ZN(n3775)
         );
  AOI21_X1 U4315 ( .B1(n3773), .B2(n3774), .A(n3775), .ZN(n3691) );
  INV_X1 U4316 ( .A(n3691), .ZN(n3692) );
  NAND2_X1 U4317 ( .A1(n3694), .A2(n3693), .ZN(n3840) );
  NAND2_X1 U4318 ( .A1(n4350), .A2(n3706), .ZN(n3696) );
  OR2_X1 U4319 ( .A1(n4340), .A2(n3415), .ZN(n3695) );
  NAND2_X1 U4320 ( .A1(n3696), .A2(n3695), .ZN(n3698) );
  XNOR2_X1 U4321 ( .A(n3698), .B(n3697), .ZN(n3703) );
  NOR2_X1 U4322 ( .A1(n4340), .A2(n3699), .ZN(n3700) );
  AOI21_X1 U4323 ( .B1(n4350), .B2(n3701), .A(n3700), .ZN(n3702) );
  NOR2_X1 U4324 ( .A1(n3703), .A2(n3702), .ZN(n3704) );
  AOI21_X1 U4325 ( .B1(n3703), .B2(n3702), .A(n3704), .ZN(n3720) );
  AOI22_X1 U4326 ( .A1(n4332), .A2(n3706), .B1(n3705), .B2(n3713), .ZN(n3710)
         );
  AOI22_X1 U4327 ( .A1(n4332), .A2(n3701), .B1(n3706), .B2(n3713), .ZN(n3708)
         );
  XNOR2_X1 U4328 ( .A(n3708), .B(n3707), .ZN(n3709) );
  XOR2_X1 U4329 ( .A(n3710), .B(n3709), .Z(n3711) );
  XNOR2_X1 U4330 ( .A(n3712), .B(n3711), .ZN(n3718) );
  AOI22_X1 U4331 ( .A1(n3713), .A2(n3843), .B1(n4859), .B2(n4321), .ZN(n3715)
         );
  AOI22_X1 U4332 ( .A1(n4902), .A2(n4350), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3714) );
  OAI211_X1 U4333 ( .C1(n4906), .C2(n4322), .A(n3715), .B(n3714), .ZN(n3716)
         );
  INV_X1 U4334 ( .A(n3716), .ZN(n3717) );
  OAI21_X1 U4335 ( .B1(n3718), .B2(n4896), .A(n3717), .ZN(U3217) );
  OAI211_X1 U4336 ( .C1(n3721), .C2(n3720), .A(n3719), .B(n4867), .ZN(n3725)
         );
  AOI22_X1 U4337 ( .A1(n4902), .A2(n4370), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3724) );
  AOI22_X1 U4338 ( .A1(n4331), .A2(n3843), .B1(n4859), .B2(n4332), .ZN(n3723)
         );
  OR2_X1 U4339 ( .A1(n4906), .A2(n4327), .ZN(n3722) );
  NAND4_X1 U4340 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(U3211)
         );
  INV_X1 U4341 ( .A(n3726), .ZN(n3819) );
  OAI21_X1 U4342 ( .B1(n3819), .B2(n3728), .A(n3727), .ZN(n3730) );
  NAND3_X1 U4343 ( .A1(n3730), .A2(n4867), .A3(n3729), .ZN(n3734) );
  AOI22_X1 U4344 ( .A1(n4902), .A2(n4454), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3733) );
  AOI22_X1 U4345 ( .A1(n4419), .A2(n3843), .B1(n4859), .B2(n4416), .ZN(n3732)
         );
  OR2_X1 U4346 ( .A1(n4906), .A2(n4422), .ZN(n3731) );
  NAND4_X1 U4347 ( .A1(n3734), .A2(n3733), .A3(n3732), .A4(n3731), .ZN(U3213)
         );
  AND2_X1 U4348 ( .A1(n3736), .A2(n3735), .ZN(n3739) );
  OAI211_X1 U4349 ( .C1(n3739), .C2(n3738), .A(n4867), .B(n3737), .ZN(n3745)
         );
  NOR2_X1 U4350 ( .A1(STATE_REG_SCAN_IN), .A2(n4065), .ZN(n4684) );
  AOI21_X1 U4351 ( .B1(n4859), .B2(n4225), .A(n4684), .ZN(n3744) );
  AOI22_X1 U4352 ( .A1(n3740), .A2(n3843), .B1(n4902), .B2(n4227), .ZN(n3743)
         );
  OR2_X1 U4353 ( .A1(n4906), .A2(n3741), .ZN(n3742) );
  NAND4_X1 U4354 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(U3214)
         );
  OR2_X1 U4355 ( .A1(n3830), .A2(n3746), .ZN(n3749) );
  NAND2_X1 U4356 ( .A1(n3749), .A2(n3747), .ZN(n3752) );
  AND2_X1 U4357 ( .A1(n3749), .A2(n3748), .ZN(n3750) );
  AOI21_X1 U4358 ( .B1(n3752), .B2(n3751), .A(n3750), .ZN(n3762) );
  INV_X1 U4359 ( .A(n4902), .ZN(n3754) );
  OAI22_X1 U4360 ( .A1(n4891), .A2(n3755), .B1(n3754), .B2(n3753), .ZN(n3756)
         );
  AOI211_X1 U4361 ( .C1(n4859), .C2(n4494), .A(n3757), .B(n3756), .ZN(n3761)
         );
  INV_X1 U4362 ( .A(n4906), .ZN(n3759) );
  INV_X1 U4363 ( .A(n3758), .ZN(n4502) );
  NAND2_X1 U4364 ( .A1(n3759), .A2(n4502), .ZN(n3760) );
  OAI211_X1 U4365 ( .C1(n3762), .C2(n4896), .A(n3761), .B(n3760), .ZN(U3216)
         );
  OR2_X1 U4366 ( .A1(n2290), .A2(n3763), .ZN(n4893) );
  NAND2_X1 U4367 ( .A1(n4893), .A2(n4894), .ZN(n4892) );
  NAND2_X1 U4368 ( .A1(n4892), .A2(n4897), .ZN(n3767) );
  XNOR2_X1 U4369 ( .A(n3765), .B(n3764), .ZN(n3766) );
  XNOR2_X1 U4370 ( .A(n3767), .B(n3766), .ZN(n3771) );
  AOI22_X1 U4371 ( .A1(n4453), .A2(n3843), .B1(n4859), .B2(n4454), .ZN(n3769)
         );
  AOI22_X1 U4372 ( .A1(n4902), .A2(n4494), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3768) );
  OAI211_X1 U4373 ( .C1(n4906), .C2(n4461), .A(n3769), .B(n3768), .ZN(n3770)
         );
  AOI21_X1 U4374 ( .B1(n3771), .B2(n4867), .A(n3770), .ZN(n3772) );
  INV_X1 U4375 ( .A(n3772), .ZN(U3220) );
  XOR2_X1 U4376 ( .A(n3775), .B(n3774), .Z(n3776) );
  XNOR2_X1 U4377 ( .A(n3773), .B(n3776), .ZN(n3781) );
  AOI22_X1 U4378 ( .A1(n3777), .A2(n3843), .B1(n4859), .B2(n4370), .ZN(n3779)
         );
  AOI22_X1 U4379 ( .A1(n4902), .A2(n4416), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3778) );
  OAI211_X1 U4380 ( .C1(n4906), .C2(n4376), .A(n3779), .B(n3778), .ZN(n3780)
         );
  AOI21_X1 U4381 ( .B1(n3781), .B2(n4867), .A(n3780), .ZN(n3782) );
  INV_X1 U4382 ( .A(n3782), .ZN(U3222) );
  INV_X1 U4383 ( .A(n4864), .ZN(n3784) );
  NOR2_X1 U4384 ( .A1(n3783), .A2(n3784), .ZN(n3786) );
  INV_X1 U4385 ( .A(n3783), .ZN(n3785) );
  OAI22_X1 U4386 ( .A1(n3786), .A2(n4865), .B1(n3785), .B2(n4864), .ZN(n3790)
         );
  NAND2_X1 U4387 ( .A1(n3788), .A2(n3787), .ZN(n3789) );
  XNOR2_X1 U4388 ( .A(n3790), .B(n3789), .ZN(n3796) );
  AOI22_X1 U4389 ( .A1(n3791), .A2(n3843), .B1(n4859), .B2(n4517), .ZN(n3793)
         );
  NOR2_X1 U4390 ( .A1(STATE_REG_SCAN_IN), .A2(n4184), .ZN(n4724) );
  AOI21_X1 U4391 ( .B1(n4902), .B2(n4012), .A(n4724), .ZN(n3792) );
  OAI211_X1 U4392 ( .C1(n4906), .C2(n3794), .A(n3793), .B(n3792), .ZN(n3795)
         );
  AOI21_X1 U4393 ( .B1(n3796), .B2(n4867), .A(n3795), .ZN(n3797) );
  INV_X1 U4394 ( .A(n3797), .ZN(U3223) );
  NAND2_X1 U4395 ( .A1(n3799), .A2(n3798), .ZN(n3801) );
  XOR2_X1 U4396 ( .A(n3801), .B(n3800), .Z(n3807) );
  AOI22_X1 U4397 ( .A1(n3802), .A2(n3843), .B1(n4859), .B2(n4495), .ZN(n3804)
         );
  INV_X1 U4398 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4188) );
  NOR2_X1 U4399 ( .A1(STATE_REG_SCAN_IN), .A2(n4188), .ZN(n4287) );
  AOI21_X1 U4400 ( .B1(n4902), .B2(n4858), .A(n4287), .ZN(n3803) );
  OAI211_X1 U4401 ( .C1(n4906), .C2(n3805), .A(n3804), .B(n3803), .ZN(n3806)
         );
  AOI21_X1 U4402 ( .B1(n3807), .B2(n4867), .A(n3806), .ZN(n3808) );
  INV_X1 U4403 ( .A(n3808), .ZN(U3225) );
  NAND2_X1 U4404 ( .A1(n3809), .A2(n3810), .ZN(n3811) );
  XOR2_X1 U4405 ( .A(n3812), .B(n3811), .Z(n3817) );
  AOI22_X1 U4406 ( .A1(n3813), .A2(n3843), .B1(n4859), .B2(n4390), .ZN(n3815)
         );
  AOI22_X1 U4407 ( .A1(n4902), .A2(n4435), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3814) );
  OAI211_X1 U4408 ( .C1(n4906), .C2(n4395), .A(n3815), .B(n3814), .ZN(n3816)
         );
  AOI21_X1 U4409 ( .B1(n3817), .B2(n4867), .A(n3816), .ZN(n3818) );
  INV_X1 U4410 ( .A(n3818), .ZN(U3226) );
  AOI21_X1 U4411 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n3826) );
  INV_X1 U4412 ( .A(n4428), .ZN(n4440) );
  AOI22_X1 U4413 ( .A1(n4859), .A2(n4435), .B1(n3843), .B2(n4440), .ZN(n3823)
         );
  AOI22_X1 U4414 ( .A1(n4902), .A2(n4889), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3822) );
  OAI211_X1 U4415 ( .C1(n4906), .C2(n4442), .A(n3823), .B(n3822), .ZN(n3824)
         );
  INV_X1 U4416 ( .A(n3824), .ZN(n3825) );
  OAI21_X1 U4417 ( .B1(n3826), .B2(n4896), .A(n3825), .ZN(U3232) );
  XOR2_X1 U4418 ( .A(n3828), .B(n3827), .Z(n3829) );
  XNOR2_X1 U4419 ( .A(n3830), .B(n3829), .ZN(n3836) );
  AOI22_X1 U4420 ( .A1(n3831), .A2(n3843), .B1(n4859), .B2(n4901), .ZN(n3834)
         );
  NOR2_X1 U4421 ( .A1(STATE_REG_SCAN_IN), .A2(n3832), .ZN(n4294) );
  AOI21_X1 U4422 ( .B1(n4902), .B2(n4517), .A(n4294), .ZN(n3833) );
  OAI211_X1 U4423 ( .C1(n4906), .C2(n4525), .A(n3834), .B(n3833), .ZN(n3835)
         );
  AOI21_X1 U4424 ( .B1(n3836), .B2(n4867), .A(n3835), .ZN(n3837) );
  INV_X1 U4425 ( .A(n3837), .ZN(U3235) );
  INV_X1 U4426 ( .A(n3839), .ZN(n3841) );
  NAND2_X1 U4427 ( .A1(n3841), .A2(n3840), .ZN(n3842) );
  XNOR2_X1 U4428 ( .A(n3838), .B(n3842), .ZN(n3849) );
  AOI22_X1 U4429 ( .A1(n2385), .A2(n3843), .B1(n4859), .B2(n4350), .ZN(n3847)
         );
  NOR2_X1 U4430 ( .A1(n3844), .A2(STATE_REG_SCAN_IN), .ZN(n3845) );
  AOI21_X1 U4431 ( .B1(n4902), .B2(n4390), .A(n3845), .ZN(n3846) );
  OAI211_X1 U4432 ( .C1(n4906), .C2(n4355), .A(n3847), .B(n3846), .ZN(n3848)
         );
  AOI21_X1 U4433 ( .B1(n3849), .B2(n4867), .A(n3848), .ZN(n3850) );
  INV_X1 U4434 ( .A(n3850), .ZN(U3237) );
  INV_X1 U4435 ( .A(n3851), .ZN(n4010) );
  AOI22_X1 U4436 ( .A1(n4010), .A2(n3912), .B1(n3987), .B2(n3990), .ZN(n3919)
         );
  INV_X1 U4437 ( .A(n3951), .ZN(n4409) );
  INV_X1 U4438 ( .A(n3852), .ZN(n3974) );
  NAND3_X1 U4439 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n3885) );
  INV_X1 U4440 ( .A(n3885), .ZN(n3858) );
  INV_X1 U4441 ( .A(n3856), .ZN(n3857) );
  NAND3_X1 U4442 ( .A1(n3858), .A2(n3857), .A3(n3882), .ZN(n3862) );
  AND2_X1 U4443 ( .A1(n3860), .A2(n3859), .ZN(n3892) );
  INV_X1 U4444 ( .A(n3892), .ZN(n3861) );
  AOI21_X1 U4445 ( .B1(n3863), .B2(n3862), .A(n3861), .ZN(n3866) );
  NAND2_X1 U4446 ( .A1(n3864), .A2(n3869), .ZN(n3965) );
  NOR3_X1 U4447 ( .A1(n3866), .A2(n3965), .A3(n3865), .ZN(n3898) );
  NAND2_X1 U4448 ( .A1(n3868), .A2(n3867), .ZN(n3891) );
  NAND2_X1 U4449 ( .A1(n3891), .A2(n3869), .ZN(n3967) );
  INV_X1 U4450 ( .A(n3967), .ZN(n3897) );
  OAI211_X1 U4451 ( .C1(n3872), .C2(n3991), .A(n3871), .B(n3870), .ZN(n3874)
         );
  NAND3_X1 U4452 ( .A1(n3874), .A2(n3873), .A3(n2935), .ZN(n3877) );
  NAND3_X1 U4453 ( .A1(n3877), .A2(n3876), .A3(n3875), .ZN(n3880) );
  NAND3_X1 U4454 ( .A1(n3880), .A2(n3879), .A3(n3878), .ZN(n3884) );
  NAND4_X1 U4455 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3887)
         );
  AOI21_X1 U4456 ( .B1(n3887), .B2(n3886), .A(n3885), .ZN(n3895) );
  AOI21_X1 U4457 ( .B1(n3890), .B2(n3889), .A(n3888), .ZN(n3894) );
  INV_X1 U4458 ( .A(n3891), .ZN(n3893) );
  OAI211_X1 U4459 ( .C1(n3895), .C2(n3894), .A(n3893), .B(n3892), .ZN(n3896)
         );
  OAI21_X1 U4460 ( .B1(n3898), .B2(n3897), .A(n3896), .ZN(n3900) );
  NOR2_X1 U4461 ( .A1(n3949), .A2(n3899), .ZN(n3973) );
  OAI211_X1 U4462 ( .C1(n3974), .C2(n3900), .A(n3966), .B(n3973), .ZN(n3901)
         );
  OAI221_X1 U4463 ( .B1(n4409), .B2(n2392), .C1(n4409), .C2(n3901), .A(n3977), 
        .ZN(n3902) );
  AOI21_X1 U4464 ( .B1(n3903), .B2(n3902), .A(n3980), .ZN(n3905) );
  INV_X1 U4465 ( .A(n3963), .ZN(n3904) );
  OAI21_X1 U4466 ( .B1(n3905), .B2(n3978), .A(n3904), .ZN(n3906) );
  NAND4_X1 U4467 ( .A1(n3919), .A2(n3907), .A3(n3960), .A4(n3906), .ZN(n3917)
         );
  NAND2_X1 U4468 ( .A1(n4321), .A2(n3914), .ZN(n3908) );
  AND2_X1 U4469 ( .A1(n3909), .A2(n3908), .ZN(n3961) );
  INV_X1 U4470 ( .A(n3961), .ZN(n3916) );
  NOR2_X1 U4471 ( .A1(n3987), .A2(n3990), .ZN(n3910) );
  NOR2_X1 U4472 ( .A1(n3919), .A2(n3910), .ZN(n3915) );
  INV_X1 U4473 ( .A(n3910), .ZN(n3911) );
  OAI21_X1 U4474 ( .B1(n3912), .B2(n4010), .A(n3911), .ZN(n3939) );
  INV_X1 U4475 ( .A(n3939), .ZN(n3913) );
  OAI21_X1 U4476 ( .B1(n4321), .B2(n3914), .A(n3913), .ZN(n3962) );
  AOI21_X1 U4477 ( .B1(n3961), .B2(n3964), .A(n3962), .ZN(n3985) );
  OAI22_X1 U4478 ( .A1(n3917), .A2(n3916), .B1(n3915), .B2(n3985), .ZN(n3998)
         );
  NAND2_X1 U4479 ( .A1(n3998), .A2(n3918), .ZN(n3996) );
  INV_X1 U4480 ( .A(n3919), .ZN(n3989) );
  NAND2_X1 U4481 ( .A1(n3921), .A2(n3920), .ZN(n4411) );
  INV_X1 U4482 ( .A(n4411), .ZN(n3924) );
  NOR4_X1 U4483 ( .A1(n3989), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3935)
         );
  NOR2_X1 U4484 ( .A1(n4329), .A2(n2502), .ZN(n3934) );
  NOR4_X1 U4485 ( .A1(n2763), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3933)
         );
  NOR4_X1 U4486 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3932)
         );
  NAND4_X1 U4487 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3959)
         );
  NOR4_X1 U4488 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3955)
         );
  OR2_X1 U4489 ( .A1(n3941), .A2(n3940), .ZN(n4491) );
  NAND2_X1 U4490 ( .A1(n4348), .A2(n3942), .ZN(n4366) );
  NOR4_X1 U4491 ( .A1(n3943), .A2(n4491), .A3(n4366), .A4(n4736), .ZN(n3954)
         );
  NAND2_X1 U4492 ( .A1(n3944), .A2(n4363), .ZN(n4400) );
  NOR4_X1 U4493 ( .A1(n3946), .A2(n4400), .A3(n4316), .A4(n3945), .ZN(n3953)
         );
  INV_X1 U4494 ( .A(n4431), .ZN(n4438) );
  INV_X1 U4495 ( .A(n3947), .ZN(n3948) );
  OR2_X1 U4496 ( .A1(n3949), .A2(n3948), .ZN(n4472) );
  NAND2_X1 U4497 ( .A1(n3950), .A2(n3960), .ZN(n4349) );
  NAND2_X1 U4498 ( .A1(n4408), .A2(n3951), .ZN(n4450) );
  NOR4_X1 U4499 ( .A1(n4438), .A2(n4472), .A3(n4349), .A4(n4450), .ZN(n3952)
         );
  NAND4_X1 U4500 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3958)
         );
  NOR4_X1 U4501 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3993)
         );
  NAND3_X1 U4502 ( .A1(n4337), .A2(n3961), .A3(n3960), .ZN(n3984) );
  NOR3_X1 U4503 ( .A1(n3964), .A2(n3963), .A3(n3962), .ZN(n3983) );
  INV_X1 U4504 ( .A(n3965), .ZN(n3969) );
  NAND2_X1 U4505 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  AOI21_X1 U4506 ( .B1(n3970), .B2(n3969), .A(n3968), .ZN(n3972) );
  AOI221_X1 U4507 ( .B1(n3974), .B2(n3973), .C1(n3972), .C2(n3973), .A(n3971), 
        .ZN(n3976) );
  AOI21_X1 U4508 ( .B1(n3977), .B2(n3976), .A(n3975), .ZN(n3981) );
  INV_X1 U4509 ( .A(n3978), .ZN(n3979) );
  OAI21_X1 U4510 ( .B1(n3981), .B2(n3980), .A(n3979), .ZN(n3982) );
  AOI22_X1 U4511 ( .A1(n3985), .A2(n3984), .B1(n3983), .B2(n3982), .ZN(n3986)
         );
  AOI21_X1 U4512 ( .B1(n3987), .B2(n4534), .A(n3986), .ZN(n3988) );
  AOI21_X1 U4513 ( .B1(n3990), .B2(n3989), .A(n3988), .ZN(n3992) );
  MUX2_X1 U4514 ( .A(n3993), .B(n3992), .S(n3991), .Z(n3994) );
  XNOR2_X1 U4515 ( .A(n3994), .B(n4785), .ZN(n3995) );
  MUX2_X1 U4516 ( .A(n3996), .B(n3995), .S(n4626), .Z(n3997) );
  OAI21_X1 U4517 ( .B1(n3998), .B2(n4734), .A(n3997), .ZN(n4008) );
  INV_X1 U4518 ( .A(n4632), .ZN(n4007) );
  NAND3_X1 U4519 ( .A1(n4000), .A2(STATE_REG_SCAN_IN), .A3(n3999), .ZN(n4001)
         );
  NOR4_X1 U4520 ( .A1(n3699), .A2(n4908), .A3(n4002), .A4(n4001), .ZN(n4003)
         );
  AOI211_X1 U4521 ( .C1(n4007), .C2(n4005), .A(n4004), .B(n4003), .ZN(n4006)
         );
  AOI21_X1 U4522 ( .B1(n4008), .B2(n4007), .A(n4006), .ZN(n4009) );
  INV_X1 U4523 ( .A(n4009), .ZN(U3239) );
  MUX2_X1 U4524 ( .A(DATAO_REG_30__SCAN_IN), .B(n4010), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4525 ( .A(DATAO_REG_29__SCAN_IN), .B(n4321), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4526 ( .A(DATAO_REG_28__SCAN_IN), .B(n4332), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4527 ( .A(DATAO_REG_27__SCAN_IN), .B(n4350), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4528 ( .A(DATAO_REG_26__SCAN_IN), .B(n4370), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4529 ( .A(DATAO_REG_25__SCAN_IN), .B(n4390), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4530 ( .A(DATAO_REG_24__SCAN_IN), .B(n4416), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4531 ( .A(DATAO_REG_23__SCAN_IN), .B(n4435), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4532 ( .A(DATAO_REG_22__SCAN_IN), .B(n4454), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4533 ( .A(DATAO_REG_21__SCAN_IN), .B(n4889), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4534 ( .A(DATAO_REG_20__SCAN_IN), .B(n4494), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4535 ( .A(DATAO_REG_19__SCAN_IN), .B(n4901), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4536 ( .A(DATAO_REG_18__SCAN_IN), .B(n4495), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4537 ( .A(DATAO_REG_17__SCAN_IN), .B(n4517), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4538 ( .A(DATAO_REG_16__SCAN_IN), .B(n4858), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4539 ( .A(DATAO_REG_15__SCAN_IN), .B(n4012), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4540 ( .A(DATAO_REG_14__SCAN_IN), .B(n4857), .S(U4043), .Z(n4222)
         );
  XNOR2_X1 U4541 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n4220) );
  INV_X1 U4542 ( .A(keyinput_50), .ZN(n4085) );
  INV_X1 U4543 ( .A(keyinput_49), .ZN(n4083) );
  INV_X1 U4544 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4190) );
  OAI22_X1 U4545 ( .A1(n4184), .A2(keyinput_46), .B1(keyinput_47), .B2(
        REG3_REG_5__SCAN_IN), .ZN(n4013) );
  AOI221_X1 U4546 ( .B1(n4184), .B2(keyinput_46), .C1(REG3_REG_5__SCAN_IN), 
        .C2(keyinput_47), .A(n4013), .ZN(n4080) );
  INV_X1 U4547 ( .A(keyinput_45), .ZN(n4078) );
  INV_X1 U4548 ( .A(keyinput_44), .ZN(n4076) );
  INV_X1 U4549 ( .A(keyinput_43), .ZN(n4074) );
  AOI22_X1 U4550 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_35), .B1(n4108), 
        .B2(keyinput_34), .ZN(n4014) );
  OAI221_X1 U4551 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_35), .C1(n4108), 
        .C2(keyinput_34), .A(n4014), .ZN(n4062) );
  INV_X1 U4552 ( .A(DATAI_3_), .ZN(n4155) );
  INV_X1 U4553 ( .A(DATAI_14_), .ZN(n4016) );
  OAI22_X1 U4554 ( .A1(n4017), .A2(keyinput_16), .B1(n4016), .B2(keyinput_17), 
        .ZN(n4015) );
  AOI221_X1 U4555 ( .B1(n4017), .B2(keyinput_16), .C1(keyinput_17), .C2(n4016), 
        .A(n4015), .ZN(n4042) );
  INV_X1 U4556 ( .A(keyinput_15), .ZN(n4038) );
  INV_X1 U4557 ( .A(keyinput_4), .ZN(n4024) );
  INV_X1 U4558 ( .A(DATAI_28_), .ZN(n4907) );
  INV_X1 U4559 ( .A(keyinput_3), .ZN(n4022) );
  INV_X1 U4560 ( .A(keyinput_2), .ZN(n4020) );
  AOI22_X1 U4561 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n4018) );
  OAI221_X1 U4562 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n4018), .ZN(n4019) );
  AOI221_X1 U4563 ( .B1(DATAI_29_), .B2(keyinput_2), .C1(n4115), .C2(n4020), 
        .A(n4019), .ZN(n4021) );
  AOI221_X1 U4564 ( .B1(DATAI_28_), .B2(keyinput_3), .C1(n4907), .C2(n4022), 
        .A(n4021), .ZN(n4023) );
  AOI221_X1 U4565 ( .B1(DATAI_27_), .B2(keyinput_4), .C1(n4119), .C2(n4024), 
        .A(n4023), .ZN(n4030) );
  XNOR2_X1 U4566 ( .A(DATAI_22_), .B(keyinput_9), .ZN(n4029) );
  AOI22_X1 U4567 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(n4123), .B2(keyinput_6), .ZN(n4025) );
  OAI221_X1 U4568 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n4123), .C2(
        keyinput_6), .A(n4025), .ZN(n4028) );
  INV_X1 U4569 ( .A(DATAI_23_), .ZN(n4633) );
  AOI22_X1 U4570 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(n4633), .B2(keyinput_8), .ZN(n4026) );
  OAI221_X1 U4571 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(n4633), .C2(
        keyinput_8), .A(n4026), .ZN(n4027) );
  NOR4_X1 U4572 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4036)
         );
  INV_X1 U4573 ( .A(DATAI_20_), .ZN(n4111) );
  AOI22_X1 U4574 ( .A1(n4111), .A2(keyinput_11), .B1(n4110), .B2(keyinput_10), 
        .ZN(n4031) );
  OAI221_X1 U4575 ( .B1(n4111), .B2(keyinput_11), .C1(n4110), .C2(keyinput_10), 
        .A(n4031), .ZN(n4035) );
  OAI22_X1 U4576 ( .A1(n4132), .A2(keyinput_14), .B1(DATAI_18_), .B2(
        keyinput_13), .ZN(n4032) );
  AOI221_X1 U4577 ( .B1(n4132), .B2(keyinput_14), .C1(keyinput_13), .C2(
        DATAI_18_), .A(n4032), .ZN(n4034) );
  XNOR2_X1 U4578 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n4033) );
  OAI211_X1 U4579 ( .C1(n4036), .C2(n4035), .A(n4034), .B(n4033), .ZN(n4037)
         );
  OAI221_X1 U4580 ( .B1(DATAI_16_), .B2(n4038), .C1(n4872), .C2(keyinput_15), 
        .A(n4037), .ZN(n4041) );
  AOI22_X1 U4581 ( .A1(DATAI_13_), .A2(keyinput_18), .B1(DATAI_12_), .B2(
        keyinput_19), .ZN(n4039) );
  OAI221_X1 U4582 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(DATAI_12_), .C2(
        keyinput_19), .A(n4039), .ZN(n4040) );
  AOI21_X1 U4583 ( .B1(n4042), .B2(n4041), .A(n4040), .ZN(n4049) );
  AOI22_X1 U4584 ( .A1(DATAI_10_), .A2(keyinput_21), .B1(n2804), .B2(
        keyinput_20), .ZN(n4043) );
  OAI221_X1 U4585 ( .B1(DATAI_10_), .B2(keyinput_21), .C1(n2804), .C2(
        keyinput_20), .A(n4043), .ZN(n4048) );
  OAI22_X1 U4586 ( .A1(DATAI_7_), .A2(keyinput_24), .B1(DATAI_6_), .B2(
        keyinput_25), .ZN(n4044) );
  AOI221_X1 U4587 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(keyinput_25), .C2(
        DATAI_6_), .A(n4044), .ZN(n4047) );
  OAI22_X1 U4588 ( .A1(DATAI_8_), .A2(keyinput_23), .B1(DATAI_4_), .B2(
        keyinput_27), .ZN(n4045) );
  AOI221_X1 U4589 ( .B1(DATAI_8_), .B2(keyinput_23), .C1(keyinput_27), .C2(
        DATAI_4_), .A(n4045), .ZN(n4046) );
  OAI211_X1 U4590 ( .C1(n4049), .C2(n4048), .A(n4047), .B(n4046), .ZN(n4052)
         );
  INV_X1 U4591 ( .A(DATAI_5_), .ZN(n4764) );
  INV_X1 U4592 ( .A(DATAI_9_), .ZN(n4819) );
  AOI22_X1 U4593 ( .A1(n4764), .A2(keyinput_26), .B1(n4819), .B2(keyinput_22), 
        .ZN(n4050) );
  OAI221_X1 U4594 ( .B1(n4764), .B2(keyinput_26), .C1(n4819), .C2(keyinput_22), 
        .A(n4050), .ZN(n4051) );
  OAI22_X1 U4595 ( .A1(keyinput_28), .A2(n4155), .B1(n4052), .B2(n4051), .ZN(
        n4053) );
  AOI21_X1 U4596 ( .B1(keyinput_28), .B2(n4155), .A(n4053), .ZN(n4060) );
  AOI22_X1 U4597 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_32), .B1(n2754), .B2(
        keyinput_33), .ZN(n4054) );
  OAI221_X1 U4598 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_32), .C1(n2754), .C2(
        keyinput_33), .A(n4054), .ZN(n4059) );
  XNOR2_X1 U4599 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n4058) );
  XOR2_X1 U4600 ( .A(DATAI_0_), .B(keyinput_31), .Z(n4056) );
  XNOR2_X1 U4601 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n4055) );
  NAND2_X1 U4602 ( .A1(n4056), .A2(n4055), .ZN(n4057) );
  NOR4_X1 U4603 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4061)
         );
  OAI22_X1 U4604 ( .A1(keyinput_36), .A2(n4165), .B1(n4062), .B2(n4061), .ZN(
        n4063) );
  AOI21_X1 U4605 ( .B1(keyinput_36), .B2(n4165), .A(n4063), .ZN(n4067) );
  AOI22_X1 U4606 ( .A1(n4065), .A2(keyinput_37), .B1(n4752), .B2(keyinput_38), 
        .ZN(n4064) );
  OAI221_X1 U4607 ( .B1(n4065), .B2(keyinput_37), .C1(n4752), .C2(keyinput_38), 
        .A(n4064), .ZN(n4066) );
  OR2_X1 U4608 ( .A1(n4067), .A2(n4066), .ZN(n4072) );
  OAI22_X1 U4609 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_41), .B1(keyinput_39), .B2(REG3_REG_19__SCAN_IN), .ZN(n4068) );
  AOI221_X1 U4610 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_41), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_39), .A(n4068), .ZN(n4071) );
  XNOR2_X1 U4611 ( .A(keyinput_40), .B(REG3_REG_28__SCAN_IN), .ZN(n4070) );
  XNOR2_X1 U4612 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n4069) );
  NAND4_X1 U4613 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4073)
         );
  OAI221_X1 U4614 ( .B1(REG3_REG_21__SCAN_IN), .B2(n4074), .C1(n2885), .C2(
        keyinput_43), .A(n4073), .ZN(n4075) );
  OAI221_X1 U4615 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_44), .C1(n4179), 
        .C2(n4076), .A(n4075), .ZN(n4077) );
  OAI221_X1 U4616 ( .B1(REG3_REG_25__SCAN_IN), .B2(n4078), .C1(n4181), .C2(
        keyinput_45), .A(n4077), .ZN(n4079) );
  OAI211_X1 U4617 ( .C1(REG3_REG_17__SCAN_IN), .C2(keyinput_48), .A(n4080), 
        .B(n4079), .ZN(n4081) );
  AOI21_X1 U4618 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_48), .A(n4081), 
        .ZN(n4082) );
  AOI221_X1 U4619 ( .B1(REG3_REG_24__SCAN_IN), .B2(n4083), .C1(n4190), .C2(
        keyinput_49), .A(n4082), .ZN(n4084) );
  AOI221_X1 U4620 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_50), .C1(n4193), 
        .C2(n4085), .A(n4084), .ZN(n4089) );
  AOI22_X1 U4621 ( .A1(n2697), .A2(keyinput_52), .B1(n4087), .B2(keyinput_53), 
        .ZN(n4086) );
  OAI221_X1 U4622 ( .B1(n2697), .B2(keyinput_52), .C1(n4087), .C2(keyinput_53), 
        .A(n4086), .ZN(n4088) );
  AOI211_X1 U4623 ( .C1(n2774), .C2(keyinput_51), .A(n4089), .B(n4088), .ZN(
        n4090) );
  OAI21_X1 U4624 ( .B1(n2774), .B2(keyinput_51), .A(n4090), .ZN(n4097) );
  XNOR2_X1 U4625 ( .A(keyinput_54), .B(n4200), .ZN(n4096) );
  AOI22_X1 U4626 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_57), .B1(n2367), .B2(
        keyinput_56), .ZN(n4091) );
  OAI221_X1 U4627 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_57), .C1(n2367), .C2(
        keyinput_56), .A(n4091), .ZN(n4095) );
  XNOR2_X1 U4628 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .ZN(n4093) );
  XNOR2_X1 U4629 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n4092) );
  NAND2_X1 U4630 ( .A1(n4093), .A2(n4092), .ZN(n4094) );
  AOI211_X1 U4631 ( .C1(n4097), .C2(n4096), .A(n4095), .B(n4094), .ZN(n4102)
         );
  AND2_X1 U4632 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_61), .ZN(n4101) );
  XNOR2_X1 U4633 ( .A(n4098), .B(keyinput_59), .ZN(n4100) );
  XNOR2_X1 U4634 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4099) );
  NOR4_X1 U4635 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4103)
         );
  OAI21_X1 U4636 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_61), .A(n4103), .ZN(
        n4219) );
  INV_X1 U4637 ( .A(keyinput_118), .ZN(n4199) );
  OAI22_X1 U4638 ( .A1(n2697), .A2(keyinput_116), .B1(keyinput_115), .B2(
        REG3_REG_9__SCAN_IN), .ZN(n4104) );
  AOI221_X1 U4639 ( .B1(n2697), .B2(keyinput_116), .C1(REG3_REG_9__SCAN_IN), 
        .C2(keyinput_115), .A(n4104), .ZN(n4196) );
  INV_X1 U4640 ( .A(keyinput_114), .ZN(n4194) );
  INV_X1 U4641 ( .A(keyinput_113), .ZN(n4191) );
  INV_X1 U4642 ( .A(keyinput_109), .ZN(n4182) );
  INV_X1 U4643 ( .A(keyinput_108), .ZN(n4178) );
  INV_X1 U4644 ( .A(keyinput_107), .ZN(n4176) );
  OAI22_X1 U4645 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_102), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_101), .ZN(n4105) );
  AOI221_X1 U4646 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_102), .C1(
        keyinput_101), .C2(REG3_REG_10__SCAN_IN), .A(n4105), .ZN(n4174) );
  INV_X1 U4647 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4648 ( .A1(n4108), .A2(keyinput_98), .B1(n4107), .B2(keyinput_99), 
        .ZN(n4106) );
  OAI221_X1 U4649 ( .B1(n4108), .B2(keyinput_98), .C1(n4107), .C2(keyinput_99), 
        .A(n4106), .ZN(n4167) );
  INV_X1 U4650 ( .A(keyinput_92), .ZN(n4154) );
  AOI22_X1 U4651 ( .A1(n4111), .A2(keyinput_75), .B1(n4110), .B2(keyinput_74), 
        .ZN(n4109) );
  OAI221_X1 U4652 ( .B1(n4111), .B2(keyinput_75), .C1(n4110), .C2(keyinput_74), 
        .A(n4109), .ZN(n4130) );
  INV_X1 U4653 ( .A(keyinput_68), .ZN(n4120) );
  INV_X1 U4654 ( .A(keyinput_67), .ZN(n4117) );
  INV_X1 U4655 ( .A(keyinput_66), .ZN(n4114) );
  AOI22_X1 U4656 ( .A1(DATAI_31_), .A2(keyinput_64), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n4112) );
  OAI221_X1 U4657 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(DATAI_30_), .C2(
        keyinput_65), .A(n4112), .ZN(n4113) );
  AOI221_X1 U4658 ( .B1(DATAI_29_), .B2(keyinput_66), .C1(n4115), .C2(n4114), 
        .A(n4113), .ZN(n4116) );
  AOI221_X1 U4659 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(n4907), .C2(n4117), 
        .A(n4116), .ZN(n4118) );
  AOI221_X1 U4660 ( .B1(DATAI_27_), .B2(n4120), .C1(n4119), .C2(keyinput_68), 
        .A(n4118), .ZN(n4127) );
  XNOR2_X1 U4661 ( .A(DATAI_22_), .B(keyinput_73), .ZN(n4126) );
  AOI22_X1 U4662 ( .A1(DATAI_23_), .A2(keyinput_72), .B1(DATAI_26_), .B2(
        keyinput_69), .ZN(n4121) );
  OAI221_X1 U4663 ( .B1(DATAI_23_), .B2(keyinput_72), .C1(DATAI_26_), .C2(
        keyinput_69), .A(n4121), .ZN(n4125) );
  AOI22_X1 U4664 ( .A1(DATAI_24_), .A2(keyinput_71), .B1(n4123), .B2(
        keyinput_70), .ZN(n4122) );
  OAI221_X1 U4665 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(n4123), .C2(
        keyinput_70), .A(n4122), .ZN(n4124) );
  NOR4_X1 U4666 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4129)
         );
  NAND2_X1 U4667 ( .A1(keyinput_76), .A2(DATAI_19_), .ZN(n4128) );
  OAI221_X1 U4668 ( .B1(n4130), .B2(n4129), .C1(keyinput_76), .C2(DATAI_19_), 
        .A(n4128), .ZN(n4134) );
  AOI22_X1 U4669 ( .A1(DATAI_18_), .A2(keyinput_77), .B1(n4132), .B2(
        keyinput_78), .ZN(n4131) );
  OAI221_X1 U4670 ( .B1(DATAI_18_), .B2(keyinput_77), .C1(n4132), .C2(
        keyinput_78), .A(n4131), .ZN(n4133) );
  OAI22_X1 U4671 ( .A1(n4134), .A2(n4133), .B1(keyinput_79), .B2(DATAI_16_), 
        .ZN(n4135) );
  AOI21_X1 U4672 ( .B1(keyinput_79), .B2(DATAI_16_), .A(n4135), .ZN(n4143) );
  INV_X1 U4673 ( .A(DATAI_12_), .ZN(n4844) );
  OAI22_X1 U4674 ( .A1(n4844), .A2(keyinput_83), .B1(keyinput_82), .B2(
        DATAI_13_), .ZN(n4136) );
  AOI221_X1 U4675 ( .B1(n4844), .B2(keyinput_83), .C1(DATAI_13_), .C2(
        keyinput_82), .A(n4136), .ZN(n4142) );
  AOI22_X1 U4676 ( .A1(DATAI_14_), .A2(keyinput_81), .B1(DATAI_15_), .B2(
        keyinput_80), .ZN(n4137) );
  OAI221_X1 U4677 ( .B1(DATAI_14_), .B2(keyinput_81), .C1(DATAI_15_), .C2(
        keyinput_80), .A(n4137), .ZN(n4141) );
  INV_X1 U4678 ( .A(DATAI_10_), .ZN(n4139) );
  AOI22_X1 U4679 ( .A1(n4139), .A2(keyinput_85), .B1(n2804), .B2(keyinput_84), 
        .ZN(n4138) );
  OAI221_X1 U4680 ( .B1(n4139), .B2(keyinput_85), .C1(n2804), .C2(keyinput_84), 
        .A(n4138), .ZN(n4140) );
  AOI221_X1 U4681 ( .B1(n4143), .B2(n4142), .C1(n4141), .C2(n4142), .A(n4140), 
        .ZN(n4152) );
  INV_X1 U4682 ( .A(DATAI_6_), .ZN(n4766) );
  AOI22_X1 U4683 ( .A1(n4766), .A2(keyinput_89), .B1(keyinput_91), .B2(n4145), 
        .ZN(n4144) );
  OAI221_X1 U4684 ( .B1(n4766), .B2(keyinput_89), .C1(n4145), .C2(keyinput_91), 
        .A(n4144), .ZN(n4151) );
  INV_X1 U4685 ( .A(DATAI_8_), .ZN(n4147) );
  AOI22_X1 U4686 ( .A1(n4764), .A2(keyinput_90), .B1(n4147), .B2(keyinput_87), 
        .ZN(n4146) );
  OAI221_X1 U4687 ( .B1(n4764), .B2(keyinput_90), .C1(n4147), .C2(keyinput_87), 
        .A(n4146), .ZN(n4150) );
  INV_X1 U4688 ( .A(DATAI_7_), .ZN(n4775) );
  AOI22_X1 U4689 ( .A1(n4775), .A2(keyinput_88), .B1(n4819), .B2(keyinput_86), 
        .ZN(n4148) );
  OAI221_X1 U4690 ( .B1(n4775), .B2(keyinput_88), .C1(n4819), .C2(keyinput_86), 
        .A(n4148), .ZN(n4149) );
  NOR4_X1 U4691 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4153)
         );
  AOI221_X1 U4692 ( .B1(DATAI_3_), .B2(keyinput_92), .C1(n4155), .C2(n4154), 
        .A(n4153), .ZN(n4163) );
  AOI22_X1 U4693 ( .A1(n2373), .A2(keyinput_95), .B1(U3149), .B2(keyinput_96), 
        .ZN(n4156) );
  OAI221_X1 U4694 ( .B1(n2373), .B2(keyinput_95), .C1(U3149), .C2(keyinput_96), 
        .A(n4156), .ZN(n4157) );
  INV_X1 U4695 ( .A(n4157), .ZN(n4161) );
  XNOR2_X1 U4696 ( .A(keyinput_97), .B(REG3_REG_7__SCAN_IN), .ZN(n4160) );
  XOR2_X1 U4697 ( .A(DATAI_1_), .B(keyinput_94), .Z(n4159) );
  XNOR2_X1 U4698 ( .A(DATAI_2_), .B(keyinput_93), .ZN(n4158) );
  NAND4_X1 U4699 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4162)
         );
  NOR2_X1 U4700 ( .A1(n4163), .A2(n4162), .ZN(n4166) );
  NAND2_X1 U4701 ( .A1(n4165), .A2(keyinput_100), .ZN(n4164) );
  OAI221_X1 U4702 ( .B1(n4167), .B2(n4166), .C1(n4165), .C2(keyinput_100), .A(
        n4164), .ZN(n4173) );
  AOI22_X1 U4703 ( .A1(n2912), .A2(keyinput_104), .B1(n4169), .B2(keyinput_105), .ZN(n4168) );
  OAI221_X1 U4704 ( .B1(n2912), .B2(keyinput_104), .C1(n4169), .C2(
        keyinput_105), .A(n4168), .ZN(n4172) );
  AOI22_X1 U4705 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_106), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_103), .ZN(n4170) );
  OAI221_X1 U4706 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_106), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_103), .A(n4170), .ZN(n4171) );
  AOI211_X1 U4707 ( .C1(n4174), .C2(n4173), .A(n4172), .B(n4171), .ZN(n4175)
         );
  AOI221_X1 U4708 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_107), .C1(n2885), 
        .C2(n4176), .A(n4175), .ZN(n4177) );
  AOI221_X1 U4709 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_108), .C1(n4179), 
        .C2(n4178), .A(n4177), .ZN(n4180) );
  AOI221_X1 U4710 ( .B1(REG3_REG_25__SCAN_IN), .B2(n4182), .C1(n4181), .C2(
        keyinput_109), .A(n4180), .ZN(n4186) );
  AOI22_X1 U4711 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_111), .B1(n4184), 
        .B2(keyinput_110), .ZN(n4183) );
  OAI221_X1 U4712 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_111), .C1(n4184), 
        .C2(keyinput_110), .A(n4183), .ZN(n4185) );
  AOI211_X1 U4713 ( .C1(n4188), .C2(keyinput_112), .A(n4186), .B(n4185), .ZN(
        n4187) );
  OAI21_X1 U4714 ( .B1(n4188), .B2(keyinput_112), .A(n4187), .ZN(n4189) );
  OAI221_X1 U4715 ( .B1(REG3_REG_24__SCAN_IN), .B2(n4191), .C1(n4190), .C2(
        keyinput_113), .A(n4189), .ZN(n4192) );
  OAI221_X1 U4716 ( .B1(REG3_REG_4__SCAN_IN), .B2(n4194), .C1(n4193), .C2(
        keyinput_114), .A(n4192), .ZN(n4195) );
  OAI211_X1 U4717 ( .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_117), .A(n4196), 
        .B(n4195), .ZN(n4197) );
  AOI21_X1 U4718 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_117), .A(n4197), 
        .ZN(n4198) );
  AOI221_X1 U4719 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_118), .C1(n4200), 
        .C2(n4199), .A(n4198), .ZN(n4205) );
  AOI22_X1 U4720 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_122), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_121), .ZN(n4201) );
  OAI221_X1 U4721 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_122), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_121), .A(n4201), .ZN(n4204) );
  AOI22_X1 U4722 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput_120), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_119), .ZN(n4202) );
  OAI221_X1 U4723 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_120), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_119), .A(n4202), .ZN(n4203) );
  NOR3_X1 U4724 ( .A1(n4205), .A2(n4204), .A3(n4203), .ZN(n4213) );
  XNOR2_X1 U4725 ( .A(n4206), .B(keyinput_125), .ZN(n4209) );
  XNOR2_X1 U4726 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_124), .ZN(n4208) );
  XNOR2_X1 U4727 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n4207) );
  NAND3_X1 U4728 ( .A1(n4209), .A2(n4208), .A3(n4207), .ZN(n4212) );
  INV_X1 U4729 ( .A(keyinput_126), .ZN(n4210) );
  MUX2_X1 U4730 ( .A(keyinput_126), .B(n4210), .S(IR_REG_7__SCAN_IN), .Z(n4211) );
  OAI21_X1 U4731 ( .B1(n4213), .B2(n4212), .A(n4211), .ZN(n4215) );
  AOI21_X1 U4732 ( .B1(n4215), .B2(keyinput_127), .A(IR_REG_8__SCAN_IN), .ZN(
        n4217) );
  INV_X1 U4733 ( .A(keyinput_127), .ZN(n4214) );
  AOI21_X1 U4734 ( .B1(n4215), .B2(n4214), .A(keyinput_63), .ZN(n4216) );
  AOI22_X1 U4735 ( .A1(keyinput_63), .A2(n4217), .B1(IR_REG_8__SCAN_IN), .B2(
        n4216), .ZN(n4218) );
  AOI21_X1 U4736 ( .B1(n4220), .B2(n4219), .A(n4218), .ZN(n4221) );
  XOR2_X1 U4737 ( .A(n4222), .B(n4221), .Z(U3564) );
  MUX2_X1 U4738 ( .A(DATAO_REG_13__SCAN_IN), .B(n4223), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4739 ( .A(DATAO_REG_12__SCAN_IN), .B(n4224), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4740 ( .A(DATAO_REG_11__SCAN_IN), .B(n4225), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4741 ( .A(DATAO_REG_10__SCAN_IN), .B(n4226), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4742 ( .A(DATAO_REG_9__SCAN_IN), .B(n4227), .S(U4043), .Z(U3559) );
  MUX2_X1 U4743 ( .A(DATAO_REG_8__SCAN_IN), .B(n4786), .S(U4043), .Z(U3558) );
  MUX2_X1 U4744 ( .A(DATAO_REG_7__SCAN_IN), .B(n4228), .S(U4043), .Z(U3557) );
  MUX2_X1 U4745 ( .A(DATAO_REG_6__SCAN_IN), .B(n4796), .S(U4043), .Z(U3556) );
  MUX2_X1 U4746 ( .A(DATAO_REG_5__SCAN_IN), .B(n4229), .S(U4043), .Z(U3555) );
  MUX2_X1 U4747 ( .A(DATAO_REG_4__SCAN_IN), .B(n4230), .S(U4043), .Z(U3554) );
  MUX2_X1 U4748 ( .A(DATAO_REG_3__SCAN_IN), .B(n3105), .S(U4043), .Z(U3553) );
  MUX2_X1 U4749 ( .A(DATAO_REG_2__SCAN_IN), .B(n3089), .S(U4043), .Z(U3552) );
  MUX2_X1 U4750 ( .A(DATAO_REG_1__SCAN_IN), .B(n4231), .S(U4043), .Z(U3551) );
  MUX2_X1 U4751 ( .A(DATAO_REG_0__SCAN_IN), .B(n3049), .S(U4043), .Z(U3550) );
  NAND2_X1 U4752 ( .A1(n4276), .A2(n4232), .ZN(n4244) );
  OAI211_X1 U4753 ( .C1(n4235), .C2(n4234), .A(n4703), .B(n4233), .ZN(n4243)
         );
  AOI22_X1 U4754 ( .A1(n4725), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4242) );
  MUX2_X1 U4755 ( .A(REG1_REG_1__SCAN_IN), .B(n4745), .S(n4236), .Z(n4238) );
  NAND2_X1 U4756 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  NAND3_X1 U4757 ( .A1(n4726), .A2(n4240), .A3(n4239), .ZN(n4241) );
  NAND4_X1 U4758 ( .A1(n4244), .A2(n4243), .A3(n4242), .A4(n4241), .ZN(U3241)
         );
  AOI22_X1 U4759 ( .A1(n4725), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4256) );
  OAI211_X1 U4760 ( .C1(n4247), .C2(n4246), .A(n4703), .B(n4245), .ZN(n4252)
         );
  XNOR2_X1 U4761 ( .A(n4249), .B(n4248), .ZN(n4250) );
  NAND2_X1 U4762 ( .A1(n4726), .A2(n4250), .ZN(n4251) );
  AND2_X1 U4763 ( .A1(n4252), .A2(n4251), .ZN(n4255) );
  OR2_X1 U4764 ( .A1(n4731), .A2(n4253), .ZN(n4254) );
  NAND4_X1 U4765 ( .A1(n4257), .A2(n4256), .A3(n4255), .A4(n4254), .ZN(U3242)
         );
  OAI211_X1 U4766 ( .C1(n4259), .C2(REG1_REG_14__SCAN_IN), .A(n4726), .B(n4258), .ZN(n4262) );
  AOI21_X1 U4767 ( .B1(n4725), .B2(ADDR_REG_14__SCAN_IN), .A(n4260), .ZN(n4261) );
  OAI211_X1 U4768 ( .C1(n4731), .C2(n4263), .A(n4262), .B(n4261), .ZN(n4267)
         );
  AOI211_X1 U4769 ( .C1(n4265), .C2(n4264), .A(n2297), .B(n4719), .ZN(n4266)
         );
  OR2_X1 U4770 ( .A1(n4267), .A2(n4266), .ZN(U3254) );
  XNOR2_X1 U4771 ( .A(n4269), .B(n4268), .ZN(n4279) );
  AND2_X1 U4772 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4856) );
  INV_X1 U4773 ( .A(n4270), .ZN(n4271) );
  AOI211_X1 U4774 ( .C1(n4273), .C2(n4272), .A(n4271), .B(n4719), .ZN(n4274)
         );
  AOI211_X1 U4775 ( .C1(n4725), .C2(ADDR_REG_15__SCAN_IN), .A(n4856), .B(n4274), .ZN(n4278) );
  NAND2_X1 U4776 ( .A1(n4276), .A2(n4275), .ZN(n4277) );
  OAI211_X1 U4777 ( .C1(n4714), .C2(n4279), .A(n4278), .B(n4277), .ZN(U3255)
         );
  AOI21_X1 U4778 ( .B1(n4281), .B2(n4280), .A(n2284), .ZN(n4282) );
  OR2_X1 U4779 ( .A1(n4282), .A2(n4714), .ZN(n4290) );
  AOI221_X1 U4780 ( .B1(n4285), .B2(n4284), .C1(n4283), .C2(n4284), .A(n4719), 
        .ZN(n4286) );
  OR2_X1 U4781 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  AOI21_X1 U4782 ( .B1(n4725), .B2(ADDR_REG_17__SCAN_IN), .A(n4288), .ZN(n4289) );
  OAI211_X1 U4783 ( .C1(n4291), .C2(n4731), .A(n4290), .B(n4289), .ZN(U3257)
         );
  AOI21_X1 U4784 ( .B1(n4293), .B2(n4292), .A(n4719), .ZN(n4297) );
  XOR2_X1 U4785 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND2_X1 U4786 ( .A1(n4726), .A2(n4300), .ZN(n4301) );
  OAI211_X1 U4787 ( .C1(n4303), .C2(n4731), .A(n4302), .B(n4301), .ZN(U3258)
         );
  OAI22_X1 U4788 ( .A1(n4305), .A2(n4833), .B1(n4304), .B2(n4838), .ZN(n4306)
         );
  OAI21_X1 U4789 ( .B1(n4307), .B2(n4306), .A(n4526), .ZN(n4309) );
  NAND2_X1 U4790 ( .A1(n4909), .A2(REG2_REG_29__SCAN_IN), .ZN(n4308) );
  OAI211_X1 U4791 ( .C1(n2399), .C2(n4524), .A(n4309), .B(n4308), .ZN(U3354)
         );
  XNOR2_X1 U4792 ( .A(n4310), .B(n4316), .ZN(n4539) );
  OAI211_X1 U4793 ( .C1(n2386), .C2(n4312), .A(n4311), .B(n4878), .ZN(n4537)
         );
  OAI22_X1 U4794 ( .A1(n4313), .A2(n4471), .B1(n4509), .B2(n4312), .ZN(n4320)
         );
  INV_X1 U4795 ( .A(n4328), .ZN(n4315) );
  NAND2_X1 U4796 ( .A1(n4315), .A2(n4314), .ZN(n4317) );
  XNOR2_X1 U4797 ( .A(n4317), .B(n4316), .ZN(n4318) );
  NOR2_X1 U4798 ( .A1(n4318), .A2(n4513), .ZN(n4319) );
  OAI21_X1 U4799 ( .B1(n4785), .B2(n4537), .A(n4538), .ZN(n4325) );
  OAI22_X1 U4800 ( .A1(n4836), .A2(n4323), .B1(n4322), .B2(n4838), .ZN(n4324)
         );
  AOI21_X1 U4801 ( .B1(n4325), .B2(n4836), .A(n4324), .ZN(n4326) );
  OAI21_X1 U4802 ( .B1(n4539), .B2(n4524), .A(n4326), .ZN(U3262) );
  INV_X1 U4803 ( .A(n4327), .ZN(n4336) );
  AOI21_X1 U4804 ( .B1(n4330), .B2(n4329), .A(n4328), .ZN(n4335) );
  AOI22_X1 U4805 ( .A1(n4370), .A2(n4795), .B1(n4331), .B2(n4794), .ZN(n4334)
         );
  NAND2_X1 U4806 ( .A1(n4332), .A2(n4493), .ZN(n4333) );
  OAI211_X1 U4807 ( .C1(n4335), .C2(n4513), .A(n4334), .B(n4333), .ZN(n4540)
         );
  AOI21_X1 U4808 ( .B1(n4336), .B2(n4821), .A(n4540), .ZN(n4344) );
  XNOR2_X1 U4809 ( .A(n4338), .B(n4337), .ZN(n4541) );
  NAND2_X1 U4810 ( .A1(n4541), .A2(n4446), .ZN(n4343) );
  OAI21_X1 U4811 ( .B1(n2383), .B2(n4340), .A(n4339), .ZN(n4593) );
  INV_X1 U4812 ( .A(n4593), .ZN(n4341) );
  AOI22_X1 U4813 ( .A1(n4341), .A2(n4910), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4909), .ZN(n4342) );
  OAI211_X1 U4814 ( .C1(n4909), .C2(n4344), .A(n4343), .B(n4342), .ZN(U3263)
         );
  XNOR2_X1 U4815 ( .A(n4345), .B(n4349), .ZN(n4548) );
  INV_X1 U4816 ( .A(n4346), .ZN(n4347) );
  XNOR2_X1 U4817 ( .A(n2277), .B(n4349), .ZN(n4354) );
  NAND2_X1 U4818 ( .A1(n4350), .A2(n4493), .ZN(n4352) );
  NAND2_X1 U4819 ( .A1(n4390), .A2(n4795), .ZN(n4351) );
  OAI211_X1 U4820 ( .C1(n4509), .C2(n4359), .A(n4352), .B(n4351), .ZN(n4353)
         );
  AOI21_X1 U4821 ( .B1(n4354), .B2(n4791), .A(n4353), .ZN(n4547) );
  INV_X1 U4822 ( .A(n4547), .ZN(n4358) );
  OAI22_X1 U4823 ( .A1(n4836), .A2(n4356), .B1(n4355), .B2(n4838), .ZN(n4357)
         );
  AOI21_X1 U4824 ( .B1(n4358), .B2(n4836), .A(n4357), .ZN(n4361) );
  OR2_X1 U4825 ( .A1(n4375), .A2(n4359), .ZN(n4545) );
  NAND3_X1 U4826 ( .A1(n4545), .A2(n4544), .A3(n4910), .ZN(n4360) );
  OAI211_X1 U4827 ( .C1(n4548), .C2(n4524), .A(n4361), .B(n4360), .ZN(U3264)
         );
  XOR2_X1 U4828 ( .A(n4366), .B(n4362), .Z(n4550) );
  INV_X1 U4829 ( .A(n4550), .ZN(n4381) );
  INV_X1 U4830 ( .A(n4363), .ZN(n4364) );
  NOR2_X1 U4831 ( .A1(n4365), .A2(n4364), .ZN(n4367) );
  XNOR2_X1 U4832 ( .A(n4367), .B(n4366), .ZN(n4372) );
  OAI22_X1 U4833 ( .A1(n4368), .A2(n4471), .B1(n4373), .B2(n4509), .ZN(n4369)
         );
  AOI21_X1 U4834 ( .B1(n4493), .B2(n4370), .A(n4369), .ZN(n4371) );
  OAI21_X1 U4835 ( .B1(n4372), .B2(n4513), .A(n4371), .ZN(n4549) );
  NOR2_X1 U4836 ( .A1(n4391), .A2(n4373), .ZN(n4374) );
  OR2_X1 U4837 ( .A1(n4375), .A2(n4374), .ZN(n4598) );
  NOR2_X1 U4838 ( .A1(n4598), .A2(n4833), .ZN(n4379) );
  OAI22_X1 U4839 ( .A1(n4526), .A2(n4377), .B1(n4376), .B2(n4838), .ZN(n4378)
         );
  AOI211_X1 U4840 ( .C1(n4549), .C2(n4836), .A(n4379), .B(n4378), .ZN(n4380)
         );
  OAI21_X1 U4841 ( .B1(n4381), .B2(n4524), .A(n4380), .ZN(U3265) );
  OAI22_X1 U4842 ( .A1(n4382), .A2(n4471), .B1(n4509), .B2(n4393), .ZN(n4389)
         );
  INV_X1 U4843 ( .A(n4383), .ZN(n4385) );
  NAND2_X1 U4844 ( .A1(n4385), .A2(n4384), .ZN(n4386) );
  XNOR2_X1 U4845 ( .A(n4386), .B(n4400), .ZN(n4387) );
  NOR2_X1 U4846 ( .A1(n4387), .A2(n4513), .ZN(n4388) );
  AOI211_X1 U4847 ( .C1(n4493), .C2(n4390), .A(n4389), .B(n4388), .ZN(n4553)
         );
  INV_X1 U4848 ( .A(n4421), .ZN(n4394) );
  INV_X1 U4849 ( .A(n4391), .ZN(n4392) );
  OAI21_X1 U4850 ( .B1(n4394), .B2(n4393), .A(n4392), .ZN(n4602) );
  INV_X1 U4851 ( .A(n4602), .ZN(n4398) );
  OAI22_X1 U4852 ( .A1(n4836), .A2(n4396), .B1(n4395), .B2(n4838), .ZN(n4397)
         );
  AOI21_X1 U4853 ( .B1(n4398), .B2(n4910), .A(n4397), .ZN(n4402) );
  XOR2_X1 U4854 ( .A(n4400), .B(n4399), .Z(n4555) );
  NAND2_X1 U4855 ( .A1(n4555), .A2(n4446), .ZN(n4401) );
  OAI211_X1 U4856 ( .C1(n4553), .C2(n4909), .A(n4402), .B(n4401), .ZN(U3266)
         );
  OAI21_X1 U4857 ( .B1(n4449), .B2(n4404), .A(n4403), .ZN(n4439) );
  INV_X1 U4858 ( .A(n4439), .ZN(n4405) );
  NOR2_X1 U4859 ( .A1(n4405), .A2(n4431), .ZN(n4436) );
  NOR2_X1 U4860 ( .A1(n4436), .A2(n4406), .ZN(n4407) );
  XOR2_X1 U4861 ( .A(n4411), .B(n4407), .Z(n4559) );
  INV_X1 U4862 ( .A(n4559), .ZN(n4427) );
  OAI21_X1 U4863 ( .B1(n4451), .B2(n4409), .A(n4408), .ZN(n4430) );
  AOI21_X1 U4864 ( .B1(n4430), .B2(n4431), .A(n4410), .ZN(n4412) );
  XNOR2_X1 U4865 ( .A(n4412), .B(n4411), .ZN(n4418) );
  OAI22_X1 U4866 ( .A1(n4414), .A2(n4471), .B1(n4509), .B2(n4413), .ZN(n4415)
         );
  AOI21_X1 U4867 ( .B1(n4493), .B2(n4416), .A(n4415), .ZN(n4417) );
  OAI21_X1 U4868 ( .B1(n4418), .B2(n4513), .A(n4417), .ZN(n4558) );
  NAND2_X1 U4869 ( .A1(n4562), .A2(n4419), .ZN(n4420) );
  NAND2_X1 U4870 ( .A1(n4421), .A2(n4420), .ZN(n4606) );
  NOR2_X1 U4871 ( .A1(n4606), .A2(n4833), .ZN(n4425) );
  OAI22_X1 U4872 ( .A1(n4526), .A2(n4423), .B1(n4422), .B2(n4838), .ZN(n4424)
         );
  AOI211_X1 U4873 ( .C1(n4558), .C2(n4836), .A(n4425), .B(n4424), .ZN(n4426)
         );
  OAI21_X1 U4874 ( .B1(n4427), .B2(n4524), .A(n4426), .ZN(U3267) );
  INV_X1 U4875 ( .A(n4889), .ZN(n4429) );
  OAI22_X1 U4876 ( .A1(n4429), .A2(n4471), .B1(n4428), .B2(n4509), .ZN(n4434)
         );
  XOR2_X1 U4877 ( .A(n4431), .B(n4430), .Z(n4432) );
  NOR2_X1 U4878 ( .A1(n4432), .A2(n4513), .ZN(n4433) );
  AOI211_X1 U4879 ( .C1(n4493), .C2(n4435), .A(n4434), .B(n4433), .ZN(n4565)
         );
  INV_X1 U4880 ( .A(n4436), .ZN(n4437) );
  OAI21_X1 U4881 ( .B1(n4439), .B2(n4438), .A(n4437), .ZN(n4566) );
  INV_X1 U4882 ( .A(n4566), .ZN(n4447) );
  INV_X1 U4883 ( .A(n4460), .ZN(n4441) );
  NAND2_X1 U4884 ( .A1(n4441), .A2(n4440), .ZN(n4563) );
  AND3_X1 U4885 ( .A1(n4563), .A2(n4910), .A3(n4562), .ZN(n4445) );
  OAI22_X1 U4886 ( .A1(n4526), .A2(n4443), .B1(n4442), .B2(n4838), .ZN(n4444)
         );
  AOI211_X1 U4887 ( .C1(n4447), .C2(n4446), .A(n4445), .B(n4444), .ZN(n4448)
         );
  OAI21_X1 U4888 ( .B1(n4909), .B2(n4565), .A(n4448), .ZN(U3268) );
  XNOR2_X1 U4889 ( .A(n4449), .B(n4450), .ZN(n4568) );
  INV_X1 U4890 ( .A(n4568), .ZN(n4466) );
  XNOR2_X1 U4891 ( .A(n4451), .B(n4450), .ZN(n4452) );
  NAND2_X1 U4892 ( .A1(n4452), .A2(n4791), .ZN(n4456) );
  AOI22_X1 U4893 ( .A1(n4454), .A2(n4493), .B1(n4794), .B2(n4453), .ZN(n4455)
         );
  OAI211_X1 U4894 ( .C1(n4457), .C2(n4471), .A(n4456), .B(n4455), .ZN(n4567)
         );
  NOR2_X1 U4895 ( .A1(n4478), .A2(n4458), .ZN(n4459) );
  OR2_X1 U4896 ( .A1(n4460), .A2(n4459), .ZN(n4611) );
  NOR2_X1 U4897 ( .A1(n4611), .A2(n4833), .ZN(n4464) );
  OAI22_X1 U4898 ( .A1(n4526), .A2(n4462), .B1(n4461), .B2(n4838), .ZN(n4463)
         );
  AOI211_X1 U4899 ( .C1(n4567), .C2(n4836), .A(n4464), .B(n4463), .ZN(n4465)
         );
  OAI21_X1 U4900 ( .B1(n4466), .B2(n4524), .A(n4465), .ZN(U3269) );
  NAND2_X1 U4901 ( .A1(n4468), .A2(n4467), .ZN(n4469) );
  XOR2_X1 U4902 ( .A(n4469), .B(n4472), .Z(n4477) );
  INV_X1 U4903 ( .A(n4901), .ZN(n4511) );
  AOI22_X1 U4904 ( .A1(n4889), .A2(n4493), .B1(n4479), .B2(n4794), .ZN(n4470)
         );
  OAI21_X1 U4905 ( .B1(n4511), .B2(n4471), .A(n4470), .ZN(n4476) );
  XNOR2_X1 U4906 ( .A(n4473), .B(n4472), .ZN(n4574) );
  NOR2_X1 U4907 ( .A1(n4574), .A2(n4474), .ZN(n4475) );
  AOI211_X1 U4908 ( .C1(n4477), .C2(n4791), .A(n4476), .B(n4475), .ZN(n4573)
         );
  INV_X1 U4909 ( .A(n4574), .ZN(n4483) );
  NAND2_X1 U4910 ( .A1(n4501), .A2(n4479), .ZN(n4571) );
  AND3_X1 U4911 ( .A1(n2375), .A2(n4910), .A3(n4571), .ZN(n4482) );
  OAI22_X1 U4912 ( .A1(n4526), .A2(n4480), .B1(n4905), .B2(n4838), .ZN(n4481)
         );
  AOI211_X1 U4913 ( .C1(n4483), .C2(n4825), .A(n4482), .B(n4481), .ZN(n4484)
         );
  OAI21_X1 U4914 ( .B1(n4573), .B2(n4909), .A(n4484), .ZN(U3270) );
  XNOR2_X1 U4915 ( .A(n4485), .B(n4491), .ZN(n4576) );
  INV_X1 U4916 ( .A(n4576), .ZN(n4506) );
  INV_X1 U4917 ( .A(n4486), .ZN(n4487) );
  AOI21_X1 U4918 ( .B1(n2394), .B2(n4488), .A(n4487), .ZN(n4512) );
  AOI21_X1 U4919 ( .B1(n4512), .B2(n4490), .A(n4489), .ZN(n4492) );
  XNOR2_X1 U4920 ( .A(n4492), .B(n4491), .ZN(n4498) );
  AOI22_X1 U4921 ( .A1(n4494), .A2(n4493), .B1(n4499), .B2(n4794), .ZN(n4497)
         );
  NAND2_X1 U4922 ( .A1(n4495), .A2(n4795), .ZN(n4496) );
  OAI211_X1 U4923 ( .C1(n4498), .C2(n4513), .A(n4497), .B(n4496), .ZN(n4575)
         );
  NAND2_X1 U4924 ( .A1(n4507), .A2(n4499), .ZN(n4500) );
  NAND2_X1 U4925 ( .A1(n4501), .A2(n4500), .ZN(n4616) );
  AOI22_X1 U4926 ( .A1(n4909), .A2(REG2_REG_19__SCAN_IN), .B1(n4502), .B2(
        n4821), .ZN(n4503) );
  OAI21_X1 U4927 ( .B1(n4616), .B2(n4833), .A(n4503), .ZN(n4504) );
  AOI21_X1 U4928 ( .B1(n4575), .B2(n4836), .A(n4504), .ZN(n4505) );
  OAI21_X1 U4929 ( .B1(n4506), .B2(n4524), .A(n4505), .ZN(U3271) );
  OAI211_X1 U4930 ( .C1(n4508), .C2(n4510), .A(n4507), .B(n4878), .ZN(n4579)
         );
  OAI22_X1 U4931 ( .A1(n4511), .A2(n4799), .B1(n4510), .B2(n4509), .ZN(n4516)
         );
  XNOR2_X1 U4932 ( .A(n4512), .B(n4523), .ZN(n4514) );
  NOR2_X1 U4933 ( .A1(n4514), .A2(n4513), .ZN(n4515) );
  AOI211_X1 U4934 ( .C1(n4795), .C2(n4517), .A(n4516), .B(n4515), .ZN(n4580)
         );
  OAI21_X1 U4935 ( .B1(n4785), .B2(n4579), .A(n4580), .ZN(n4529) );
  NAND2_X1 U4936 ( .A1(n4519), .A2(n4518), .ZN(n4522) );
  INV_X1 U4937 ( .A(n4520), .ZN(n4521) );
  AOI21_X1 U4938 ( .B1(n4523), .B2(n4522), .A(n4521), .ZN(n4581) );
  NOR2_X1 U4939 ( .A1(n4581), .A2(n4524), .ZN(n4528) );
  OAI22_X1 U4940 ( .A1(n4526), .A2(n2639), .B1(n4525), .B2(n4838), .ZN(n4527)
         );
  AOI211_X1 U4941 ( .C1(n4529), .C2(n4526), .A(n4528), .B(n4527), .ZN(n4530)
         );
  INV_X1 U4942 ( .A(n4530), .ZN(U3272) );
  AOI21_X1 U4943 ( .B1(n4534), .B2(n4532), .A(n4531), .ZN(n4911) );
  INV_X1 U4944 ( .A(n4911), .ZN(n4588) );
  INV_X1 U4945 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4535) );
  AOI21_X1 U4946 ( .B1(n4534), .B2(n4794), .A(n4533), .ZN(n4913) );
  MUX2_X1 U4947 ( .A(n4535), .B(n4913), .S(n4885), .Z(n4536) );
  OAI21_X1 U4948 ( .B1(n4588), .B2(n4585), .A(n4536), .ZN(U3548) );
  OAI211_X1 U4949 ( .C1(n4539), .C2(n2439), .A(n4538), .B(n4537), .ZN(n4589)
         );
  MUX2_X1 U4950 ( .A(REG1_REG_28__SCAN_IN), .B(n4589), .S(n4885), .Z(U3546) );
  INV_X1 U4951 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4542) );
  AOI21_X1 U4952 ( .B1(n4541), .B2(n4874), .A(n4540), .ZN(n4590) );
  MUX2_X1 U4953 ( .A(n4542), .B(n4590), .S(n4885), .Z(n4543) );
  OAI21_X1 U4954 ( .B1(n4585), .B2(n4593), .A(n4543), .ZN(U3545) );
  NAND3_X1 U4955 ( .A1(n4545), .A2(n4544), .A3(n4878), .ZN(n4546) );
  OAI211_X1 U4956 ( .C1(n4548), .C2(n2439), .A(n4547), .B(n4546), .ZN(n4594)
         );
  MUX2_X1 U4957 ( .A(REG1_REG_26__SCAN_IN), .B(n4594), .S(n4885), .Z(U3544) );
  INV_X1 U4958 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4551) );
  AOI21_X1 U4959 ( .B1(n4550), .B2(n4874), .A(n4549), .ZN(n4595) );
  MUX2_X1 U4960 ( .A(n4551), .B(n4595), .S(n4885), .Z(n4552) );
  OAI21_X1 U4961 ( .B1(n4585), .B2(n4598), .A(n4552), .ZN(U3543) );
  INV_X1 U4962 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4556) );
  INV_X1 U4963 ( .A(n4553), .ZN(n4554) );
  AOI21_X1 U4964 ( .B1(n4555), .B2(n4874), .A(n4554), .ZN(n4599) );
  MUX2_X1 U4965 ( .A(n4556), .B(n4599), .S(n4885), .Z(n4557) );
  OAI21_X1 U4966 ( .B1(n4585), .B2(n4602), .A(n4557), .ZN(U3542) );
  INV_X1 U4967 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4560) );
  AOI21_X1 U4968 ( .B1(n4559), .B2(n4874), .A(n4558), .ZN(n4603) );
  MUX2_X1 U4969 ( .A(n4560), .B(n4603), .S(n4885), .Z(n4561) );
  OAI21_X1 U4970 ( .B1(n4585), .B2(n4606), .A(n4561), .ZN(U3541) );
  NAND3_X1 U4971 ( .A1(n4563), .A2(n4878), .A3(n4562), .ZN(n4564) );
  OAI211_X1 U4972 ( .C1(n4566), .C2(n2439), .A(n4565), .B(n4564), .ZN(n4607)
         );
  MUX2_X1 U4973 ( .A(REG1_REG_22__SCAN_IN), .B(n4607), .S(n4885), .Z(U3540) );
  INV_X1 U4974 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4569) );
  AOI21_X1 U4975 ( .B1(n4568), .B2(n4874), .A(n4567), .ZN(n4608) );
  MUX2_X1 U4976 ( .A(n4569), .B(n4608), .S(n4885), .Z(n4570) );
  OAI21_X1 U4977 ( .B1(n4585), .B2(n4611), .A(n4570), .ZN(U3539) );
  NAND3_X1 U4978 ( .A1(n2375), .A2(n4571), .A3(n4878), .ZN(n4572) );
  OAI211_X1 U4979 ( .C1(n4574), .C2(n4741), .A(n4573), .B(n4572), .ZN(n4612)
         );
  MUX2_X1 U4980 ( .A(REG1_REG_20__SCAN_IN), .B(n4612), .S(n4885), .Z(U3538) );
  AOI21_X1 U4981 ( .B1(n4874), .B2(n4576), .A(n4575), .ZN(n4613) );
  MUX2_X1 U4982 ( .A(n4577), .B(n4613), .S(n4885), .Z(n4578) );
  OAI21_X1 U4983 ( .B1(n4585), .B2(n4616), .A(n4578), .ZN(U3537) );
  OAI211_X1 U4984 ( .C1(n2439), .C2(n4581), .A(n4580), .B(n4579), .ZN(n4617)
         );
  MUX2_X1 U4985 ( .A(REG1_REG_18__SCAN_IN), .B(n4617), .S(n4885), .Z(U3536) );
  AOI21_X1 U4986 ( .B1(n4583), .B2(n4874), .A(n4582), .ZN(n4618) );
  MUX2_X1 U4987 ( .A(n2611), .B(n4618), .S(n4885), .Z(n4584) );
  OAI21_X1 U4988 ( .B1(n4585), .B2(n4622), .A(n4584), .ZN(U3535) );
  INV_X1 U4989 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4586) );
  MUX2_X1 U4990 ( .A(n4586), .B(n4913), .S(n4888), .Z(n4587) );
  OAI21_X1 U4991 ( .B1(n4588), .B2(n4621), .A(n4587), .ZN(U3516) );
  MUX2_X1 U4992 ( .A(REG0_REG_28__SCAN_IN), .B(n4589), .S(n4888), .Z(U3514) );
  MUX2_X1 U4993 ( .A(n4591), .B(n4590), .S(n4888), .Z(n4592) );
  OAI21_X1 U4994 ( .B1(n4593), .B2(n4621), .A(n4592), .ZN(U3513) );
  MUX2_X1 U4995 ( .A(REG0_REG_26__SCAN_IN), .B(n4594), .S(n4888), .Z(U3512) );
  MUX2_X1 U4996 ( .A(n4596), .B(n4595), .S(n4888), .Z(n4597) );
  OAI21_X1 U4997 ( .B1(n4598), .B2(n4621), .A(n4597), .ZN(U3511) );
  MUX2_X1 U4998 ( .A(n4600), .B(n4599), .S(n4888), .Z(n4601) );
  OAI21_X1 U4999 ( .B1(n4602), .B2(n4621), .A(n4601), .ZN(U3510) );
  MUX2_X1 U5000 ( .A(n4604), .B(n4603), .S(n4888), .Z(n4605) );
  OAI21_X1 U5001 ( .B1(n4606), .B2(n4621), .A(n4605), .ZN(U3509) );
  MUX2_X1 U5002 ( .A(REG0_REG_22__SCAN_IN), .B(n4607), .S(n4888), .Z(U3508) );
  MUX2_X1 U5003 ( .A(n4609), .B(n4608), .S(n4888), .Z(n4610) );
  OAI21_X1 U5004 ( .B1(n4611), .B2(n4621), .A(n4610), .ZN(U3507) );
  MUX2_X1 U5005 ( .A(REG0_REG_20__SCAN_IN), .B(n4612), .S(n4888), .Z(U3506) );
  MUX2_X1 U5006 ( .A(n4614), .B(n4613), .S(n4888), .Z(n4615) );
  OAI21_X1 U5007 ( .B1(n4616), .B2(n4621), .A(n4615), .ZN(U3505) );
  MUX2_X1 U5008 ( .A(REG0_REG_18__SCAN_IN), .B(n4617), .S(n4888), .Z(U3503) );
  MUX2_X1 U5009 ( .A(n4619), .B(n4618), .S(n4888), .Z(n4620) );
  OAI21_X1 U5010 ( .B1(n4622), .B2(n4621), .A(n4620), .ZN(U3501) );
  MUX2_X1 U5011 ( .A(n4623), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5012 ( .A(n4624), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5013 ( .A(n4625), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5014 ( .A(DATAI_20_), .B(n4626), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5015 ( .A(DATAI_19_), .B(n4785), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5016 ( .A(n4627), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5017 ( .A(DATAI_14_), .B(n4628), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5018 ( .A(n4676), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5019 ( .A(DATAI_8_), .B(n4629), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5020 ( .A(DATAI_4_), .B(n4630), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5021 ( .A(DATAI_3_), .B(n4631), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5022 ( .A(n2312), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  OAI21_X1 U5023 ( .B1(STATE_REG_SCAN_IN), .B2(n4633), .A(n4632), .ZN(U3329)
         );
  AND2_X1 U5024 ( .A1(D_REG_2__SCAN_IN), .A2(n4634), .ZN(U3320) );
  AND2_X1 U5025 ( .A1(D_REG_3__SCAN_IN), .A2(n4634), .ZN(U3319) );
  AND2_X1 U5026 ( .A1(D_REG_4__SCAN_IN), .A2(n4634), .ZN(U3318) );
  AND2_X1 U5027 ( .A1(D_REG_5__SCAN_IN), .A2(n4634), .ZN(U3317) );
  AND2_X1 U5028 ( .A1(D_REG_6__SCAN_IN), .A2(n4634), .ZN(U3316) );
  AND2_X1 U5029 ( .A1(D_REG_7__SCAN_IN), .A2(n4634), .ZN(U3315) );
  AND2_X1 U5030 ( .A1(D_REG_8__SCAN_IN), .A2(n4634), .ZN(U3314) );
  AND2_X1 U5031 ( .A1(D_REG_9__SCAN_IN), .A2(n4634), .ZN(U3313) );
  AND2_X1 U5032 ( .A1(D_REG_10__SCAN_IN), .A2(n4634), .ZN(U3312) );
  AND2_X1 U5033 ( .A1(D_REG_11__SCAN_IN), .A2(n4634), .ZN(U3311) );
  AND2_X1 U5034 ( .A1(D_REG_12__SCAN_IN), .A2(n4634), .ZN(U3310) );
  AND2_X1 U5035 ( .A1(D_REG_13__SCAN_IN), .A2(n4634), .ZN(U3309) );
  AND2_X1 U5036 ( .A1(D_REG_14__SCAN_IN), .A2(n4634), .ZN(U3308) );
  AND2_X1 U5037 ( .A1(D_REG_15__SCAN_IN), .A2(n4634), .ZN(U3307) );
  AND2_X1 U5038 ( .A1(D_REG_16__SCAN_IN), .A2(n4634), .ZN(U3306) );
  AND2_X1 U5039 ( .A1(D_REG_17__SCAN_IN), .A2(n4634), .ZN(U3305) );
  AND2_X1 U5040 ( .A1(D_REG_18__SCAN_IN), .A2(n4634), .ZN(U3304) );
  AND2_X1 U5041 ( .A1(D_REG_19__SCAN_IN), .A2(n4634), .ZN(U3303) );
  AND2_X1 U5042 ( .A1(D_REG_20__SCAN_IN), .A2(n4634), .ZN(U3302) );
  AND2_X1 U5043 ( .A1(D_REG_21__SCAN_IN), .A2(n4634), .ZN(U3301) );
  AND2_X1 U5044 ( .A1(D_REG_22__SCAN_IN), .A2(n4634), .ZN(U3300) );
  AND2_X1 U5045 ( .A1(D_REG_23__SCAN_IN), .A2(n4634), .ZN(U3299) );
  AND2_X1 U5046 ( .A1(D_REG_24__SCAN_IN), .A2(n4634), .ZN(U3298) );
  AND2_X1 U5047 ( .A1(D_REG_25__SCAN_IN), .A2(n4634), .ZN(U3297) );
  AND2_X1 U5048 ( .A1(D_REG_26__SCAN_IN), .A2(n4634), .ZN(U3296) );
  AND2_X1 U5049 ( .A1(D_REG_27__SCAN_IN), .A2(n4634), .ZN(U3295) );
  AND2_X1 U5050 ( .A1(D_REG_28__SCAN_IN), .A2(n4634), .ZN(U3294) );
  AND2_X1 U5051 ( .A1(D_REG_29__SCAN_IN), .A2(n4634), .ZN(U3293) );
  AND2_X1 U5052 ( .A1(D_REG_30__SCAN_IN), .A2(n4634), .ZN(U3292) );
  AND2_X1 U5053 ( .A1(D_REG_31__SCAN_IN), .A2(n4634), .ZN(U3291) );
  AOI211_X1 U5054 ( .C1(n4637), .C2(n4636), .A(n4635), .B(n4719), .ZN(n4639)
         );
  AOI211_X1 U5055 ( .C1(n4725), .C2(ADDR_REG_5__SCAN_IN), .A(n4639), .B(n4638), 
        .ZN(n4643) );
  OAI211_X1 U5056 ( .C1(n4641), .C2(n2304), .A(n4726), .B(n4640), .ZN(n4642)
         );
  OAI211_X1 U5057 ( .C1(n4731), .C2(n4765), .A(n4643), .B(n4642), .ZN(U3245)
         );
  AOI211_X1 U5058 ( .C1(n4646), .C2(n4645), .A(n4644), .B(n4719), .ZN(n4648)
         );
  AOI211_X1 U5059 ( .C1(n4725), .C2(ADDR_REG_6__SCAN_IN), .A(n4648), .B(n4647), 
        .ZN(n4652) );
  OAI211_X1 U5060 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4650), .A(n4726), .B(n4649), 
        .ZN(n4651) );
  OAI211_X1 U5061 ( .C1(n4731), .C2(n4767), .A(n4652), .B(n4651), .ZN(U3246)
         );
  AOI22_X1 U5062 ( .A1(n4654), .A2(n4653), .B1(REG2_REG_7__SCAN_IN), .B2(n4776), .ZN(n4655) );
  AOI211_X1 U5063 ( .C1(n4725), .C2(ADDR_REG_7__SCAN_IN), .A(n4657), .B(n4656), 
        .ZN(n4663) );
  AOI21_X1 U5064 ( .B1(n4776), .B2(n4810), .A(n4658), .ZN(n4661) );
  AOI21_X1 U5065 ( .B1(n4661), .B2(n4660), .A(n4714), .ZN(n4659) );
  OAI21_X1 U5066 ( .B1(n4661), .B2(n4660), .A(n4659), .ZN(n4662) );
  OAI211_X1 U5067 ( .C1(n4731), .C2(n4776), .A(n4663), .B(n4662), .ZN(U3247)
         );
  AOI22_X1 U5068 ( .A1(n4665), .A2(n4664), .B1(REG1_REG_9__SCAN_IN), .B2(n4820), .ZN(n4667) );
  OAI21_X1 U5069 ( .B1(n4668), .B2(n4667), .A(n4726), .ZN(n4666) );
  AOI21_X1 U5070 ( .B1(n4668), .B2(n4667), .A(n4666), .ZN(n4670) );
  AOI211_X1 U5071 ( .C1(n4725), .C2(ADDR_REG_9__SCAN_IN), .A(n4670), .B(n4669), 
        .ZN(n4675) );
  OAI211_X1 U5072 ( .C1(n4673), .C2(n4672), .A(n4703), .B(n4671), .ZN(n4674)
         );
  OAI211_X1 U5073 ( .C1(n4731), .C2(n4820), .A(n4675), .B(n4674), .ZN(U3249)
         );
  OAI211_X1 U5074 ( .C1(n4678), .C2(REG2_REG_10__SCAN_IN), .A(n4677), .B(n4703), .ZN(n4682) );
  OAI211_X1 U5075 ( .C1(n4680), .C2(REG1_REG_10__SCAN_IN), .A(n4726), .B(n4679), .ZN(n4681) );
  OAI211_X1 U5076 ( .C1(n4731), .C2(n2626), .A(n4682), .B(n4681), .ZN(n4683)
         );
  AOI211_X1 U5077 ( .C1(n4725), .C2(ADDR_REG_10__SCAN_IN), .A(n4684), .B(n4683), .ZN(n4685) );
  INV_X1 U5078 ( .A(n4685), .ZN(U3250) );
  AOI22_X1 U5079 ( .A1(n4686), .A2(REG1_REG_11__SCAN_IN), .B1(n3494), .B2(
        n4830), .ZN(n4689) );
  OAI21_X1 U5080 ( .B1(n4689), .B2(n4688), .A(n4726), .ZN(n4687) );
  AOI21_X1 U5081 ( .B1(n4689), .B2(n4688), .A(n4687), .ZN(n4691) );
  AOI211_X1 U5082 ( .C1(n4725), .C2(ADDR_REG_11__SCAN_IN), .A(n4691), .B(n4690), .ZN(n4696) );
  OAI211_X1 U5083 ( .C1(n4694), .C2(n4693), .A(n4703), .B(n4692), .ZN(n4695)
         );
  OAI211_X1 U5084 ( .C1(n4731), .C2(n4830), .A(n4696), .B(n4695), .ZN(U3251)
         );
  AOI211_X1 U5085 ( .C1(n4699), .C2(n4698), .A(n4697), .B(n4714), .ZN(n4701)
         );
  AOI211_X1 U5086 ( .C1(n4725), .C2(ADDR_REG_12__SCAN_IN), .A(n4701), .B(n4700), .ZN(n4706) );
  OAI211_X1 U5087 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4704), .A(n4703), .B(n4702), .ZN(n4705) );
  OAI211_X1 U5088 ( .C1(n4731), .C2(n4845), .A(n4706), .B(n4705), .ZN(U3252)
         );
  AOI21_X1 U5089 ( .B1(n4847), .B2(n4708), .A(n4707), .ZN(n4709) );
  XNOR2_X1 U5090 ( .A(n4710), .B(n4709), .ZN(n4718) );
  NAND2_X1 U5091 ( .A1(n4711), .A2(n2306), .ZN(n4712) );
  XNOR2_X1 U5092 ( .A(n2294), .B(n4712), .ZN(n4713) );
  OAI22_X1 U5093 ( .A1(n4847), .A2(n4731), .B1(n4714), .B2(n4713), .ZN(n4715)
         );
  AOI211_X1 U5094 ( .C1(n4725), .C2(ADDR_REG_13__SCAN_IN), .A(n4716), .B(n4715), .ZN(n4717) );
  OAI21_X1 U5095 ( .B1(n4718), .B2(n4719), .A(n4717), .ZN(U3253) );
  AOI221_X1 U5096 ( .B1(n4722), .B2(n4721), .C1(n4720), .C2(n4721), .A(n4719), 
        .ZN(n4723) );
  AOI211_X1 U5097 ( .C1(n4725), .C2(ADDR_REG_16__SCAN_IN), .A(n4724), .B(n4723), .ZN(n4730) );
  OAI221_X1 U5098 ( .B1(n4728), .B2(REG1_REG_16__SCAN_IN), .C1(n4728), .C2(
        n4727), .A(n4726), .ZN(n4729) );
  OAI211_X1 U5099 ( .C1(n4731), .C2(n4873), .A(n4730), .B(n4729), .ZN(U3256)
         );
  AOI22_X1 U5100 ( .A1(STATE_REG_SCAN_IN), .A2(n2432), .B1(n2373), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5101 ( .A1(n4888), .A2(n4732), .B1(n2698), .B2(n4886), .ZN(U3467)
         );
  AOI21_X1 U5102 ( .B1(n4735), .B2(n4734), .A(n4733), .ZN(n4739) );
  AOI22_X1 U5103 ( .A1(n4736), .A2(n4825), .B1(REG3_REG_0__SCAN_IN), .B2(n4821), .ZN(n4737) );
  OAI221_X1 U5104 ( .B1(n4909), .B2(n4739), .C1(n4836), .C2(n4738), .A(n4737), 
        .ZN(U3290) );
  OAI22_X1 U5105 ( .A1(n4742), .A2(n4741), .B1(n4848), .B2(n4740), .ZN(n4743)
         );
  NOR2_X1 U5106 ( .A1(n4744), .A2(n4743), .ZN(n4746) );
  AOI22_X1 U5107 ( .A1(n4885), .A2(n4746), .B1(n4745), .B2(n4883), .ZN(U3519)
         );
  AOI22_X1 U5108 ( .A1(n4888), .A2(n4746), .B1(n2690), .B2(n4886), .ZN(U3469)
         );
  AOI22_X1 U5109 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4909), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4821), .ZN(n4750) );
  AOI22_X1 U5110 ( .A1(n4748), .A2(n4825), .B1(n4910), .B2(n4747), .ZN(n4749)
         );
  OAI211_X1 U5111 ( .C1(n4909), .C2(n4751), .A(n4750), .B(n4749), .ZN(U3288)
         );
  AOI22_X1 U5112 ( .A1(n4909), .A2(REG2_REG_3__SCAN_IN), .B1(n4821), .B2(n4752), .ZN(n4756) );
  AOI22_X1 U5113 ( .A1(n4754), .A2(n4825), .B1(n4910), .B2(n4753), .ZN(n4755)
         );
  OAI211_X1 U5114 ( .C1(n4909), .C2(n4757), .A(n4756), .B(n4755), .ZN(U3287)
         );
  INV_X1 U5115 ( .A(n4758), .ZN(n4762) );
  INV_X1 U5116 ( .A(n4759), .ZN(n4761) );
  AOI211_X1 U5117 ( .C1(n4762), .C2(n4853), .A(n4761), .B(n4760), .ZN(n4763)
         );
  AOI22_X1 U5118 ( .A1(n4885), .A2(n4763), .B1(n2574), .B2(n4883), .ZN(U3522)
         );
  AOI22_X1 U5119 ( .A1(n4888), .A2(n4763), .B1(n2727), .B2(n4886), .ZN(U3475)
         );
  AOI22_X1 U5120 ( .A1(STATE_REG_SCAN_IN), .A2(n4765), .B1(n4764), .B2(U3149), 
        .ZN(U3347) );
  AOI22_X1 U5121 ( .A1(STATE_REG_SCAN_IN), .A2(n4767), .B1(n4766), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5122 ( .A1(n4768), .A2(n4821), .B1(REG2_REG_6__SCAN_IN), .B2(n4909), .ZN(n4773) );
  INV_X1 U5123 ( .A(n4769), .ZN(n4770) );
  AOI22_X1 U5124 ( .A1(n4771), .A2(n4825), .B1(n4910), .B2(n4770), .ZN(n4772)
         );
  OAI211_X1 U5125 ( .C1(n4909), .C2(n4774), .A(n4773), .B(n4772), .ZN(U3284)
         );
  AOI22_X1 U5126 ( .A1(STATE_REG_SCAN_IN), .A2(n4776), .B1(n4775), .B2(U3149), 
        .ZN(U3345) );
  AOI21_X1 U5127 ( .B1(n4777), .B2(n4793), .A(n4848), .ZN(n4779) );
  NAND2_X1 U5128 ( .A1(n4779), .A2(n4778), .ZN(n4805) );
  NAND2_X1 U5129 ( .A1(n4780), .A2(n4789), .ZN(n4781) );
  AND2_X1 U5130 ( .A1(n4782), .A2(n4781), .ZN(n4807) );
  NAND2_X1 U5131 ( .A1(n4807), .A2(n4783), .ZN(n4784) );
  OAI211_X1 U5132 ( .C1(n4785), .C2(n4805), .A(n4784), .B(n4836), .ZN(n4801)
         );
  INV_X1 U5133 ( .A(n4786), .ZN(n4800) );
  NAND2_X1 U5134 ( .A1(n4788), .A2(n4787), .ZN(n4790) );
  XNOR2_X1 U5135 ( .A(n4790), .B(n4789), .ZN(n4792) );
  NAND2_X1 U5136 ( .A1(n4792), .A2(n4791), .ZN(n4798) );
  AOI22_X1 U5137 ( .A1(n4796), .A2(n4795), .B1(n4794), .B2(n4793), .ZN(n4797)
         );
  OAI211_X1 U5138 ( .C1(n4800), .C2(n4799), .A(n4798), .B(n4797), .ZN(n4804)
         );
  OAI22_X1 U5139 ( .A1(n4801), .A2(n4804), .B1(REG2_REG_7__SCAN_IN), .B2(n4836), .ZN(n4802) );
  OAI21_X1 U5140 ( .B1(n4803), .B2(n4838), .A(n4802), .ZN(U3283) );
  INV_X1 U5141 ( .A(n4804), .ZN(n4809) );
  INV_X1 U5142 ( .A(n4805), .ZN(n4806) );
  AOI21_X1 U5143 ( .B1(n4807), .B2(n4874), .A(n4806), .ZN(n4808) );
  AOI22_X1 U5144 ( .A1(n4885), .A2(n4811), .B1(n4810), .B2(n4883), .ZN(U3525)
         );
  AOI22_X1 U5145 ( .A1(n4888), .A2(n4811), .B1(n2757), .B2(n4886), .ZN(U3481)
         );
  NOR3_X1 U5146 ( .A1(n4813), .A2(n4812), .A3(n4848), .ZN(n4815) );
  AOI211_X1 U5147 ( .C1(n4816), .C2(n4853), .A(n4815), .B(n4814), .ZN(n4818)
         );
  AOI22_X1 U5148 ( .A1(n4885), .A2(n4818), .B1(n4817), .B2(n4883), .ZN(U3526)
         );
  AOI22_X1 U5149 ( .A1(n4888), .A2(n4818), .B1(n2769), .B2(n4886), .ZN(U3483)
         );
  AOI22_X1 U5150 ( .A1(STATE_REG_SCAN_IN), .A2(n4820), .B1(n4819), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5151 ( .A1(n4822), .A2(n4821), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4909), .ZN(n4828) );
  INV_X1 U5152 ( .A(n4823), .ZN(n4824) );
  AOI22_X1 U5153 ( .A1(n4826), .A2(n4825), .B1(n4910), .B2(n4824), .ZN(n4827)
         );
  OAI211_X1 U5154 ( .C1(n4909), .C2(n4829), .A(n4828), .B(n4827), .ZN(U3280)
         );
  AOI22_X1 U5155 ( .A1(STATE_REG_SCAN_IN), .A2(n4830), .B1(n2804), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5156 ( .A(n4831), .ZN(n4835) );
  OAI22_X1 U5157 ( .A1(n4835), .A2(n4834), .B1(n4833), .B2(n4832), .ZN(n4841)
         );
  OAI22_X1 U5158 ( .A1(n4839), .A2(n4838), .B1(n4837), .B2(n4836), .ZN(n4840)
         );
  NOR2_X1 U5159 ( .A1(n4841), .A2(n4840), .ZN(n4842) );
  OAI21_X1 U5160 ( .B1(n4843), .B2(n4909), .A(n4842), .ZN(U3279) );
  AOI22_X1 U5161 ( .A1(STATE_REG_SCAN_IN), .A2(n4845), .B1(n4844), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5162 ( .A(DATAI_13_), .ZN(n4846) );
  AOI22_X1 U5163 ( .A1(STATE_REG_SCAN_IN), .A2(n4847), .B1(n4846), .B2(U3149), 
        .ZN(U3339) );
  NOR2_X1 U5164 ( .A1(n4849), .A2(n4848), .ZN(n4851) );
  AOI211_X1 U5165 ( .C1(n4853), .C2(n4852), .A(n4851), .B(n4850), .ZN(n4855)
         );
  INV_X1 U5166 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U5167 ( .A1(n4885), .A2(n4855), .B1(n4854), .B2(n4883), .ZN(U3531)
         );
  AOI22_X1 U5168 ( .A1(n4888), .A2(n4855), .B1(n2817), .B2(n4886), .ZN(U3493)
         );
  AOI21_X1 U5169 ( .B1(n4902), .B2(n4857), .A(n4856), .ZN(n4863) );
  NAND2_X1 U5170 ( .A1(n4859), .A2(n4858), .ZN(n4862) );
  NAND2_X1 U5171 ( .A1(n3843), .A2(n4860), .ZN(n4861) );
  AND3_X1 U5172 ( .A1(n4863), .A2(n4862), .A3(n4861), .ZN(n4870) );
  XNOR2_X1 U5173 ( .A(n4865), .B(n4864), .ZN(n4866) );
  XNOR2_X1 U5174 ( .A(n3783), .B(n4866), .ZN(n4868) );
  NAND2_X1 U5175 ( .A1(n4868), .A2(n4867), .ZN(n4869) );
  OAI211_X1 U5176 ( .C1(n4906), .C2(n4871), .A(n4870), .B(n4869), .ZN(U3238)
         );
  AOI22_X1 U5177 ( .A1(STATE_REG_SCAN_IN), .A2(n4873), .B1(n4872), .B2(U3149), 
        .ZN(U3336) );
  NAND3_X1 U5178 ( .A1(n4876), .A2(n4875), .A3(n4874), .ZN(n4881) );
  NAND3_X1 U5179 ( .A1(n4879), .A2(n4878), .A3(n4877), .ZN(n4880) );
  INV_X1 U5180 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U5181 ( .A1(n4885), .A2(n4887), .B1(n4884), .B2(n4883), .ZN(U3534)
         );
  AOI22_X1 U5182 ( .A1(n4888), .A2(n4887), .B1(n2845), .B2(n4886), .ZN(U3499)
         );
  AOI22_X1 U5183 ( .A1(n4859), .A2(n4889), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4904) );
  NOR2_X1 U5184 ( .A1(n4891), .A2(n4890), .ZN(n4900) );
  INV_X1 U5185 ( .A(n4892), .ZN(n4898) );
  AOI21_X1 U5186 ( .B1(n4897), .B2(n4894), .A(n4893), .ZN(n4895) );
  AOI211_X1 U5187 ( .C1(n4898), .C2(n4897), .A(n4896), .B(n4895), .ZN(n4899)
         );
  AOI211_X1 U5188 ( .C1(n4902), .C2(n4901), .A(n4900), .B(n4899), .ZN(n4903)
         );
  OAI211_X1 U5189 ( .C1(n4906), .C2(n4905), .A(n4904), .B(n4903), .ZN(U3230)
         );
  AOI22_X1 U5190 ( .A1(STATE_REG_SCAN_IN), .A2(n4908), .B1(n4907), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5191 ( .A1(n4911), .A2(n4910), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4909), .ZN(n4912) );
  OAI21_X1 U5192 ( .B1(n4909), .B2(n4913), .A(n4912), .ZN(U3261) );
  CLKBUF_X1 U2309 ( .A(n2707), .Z(n2931) );
endmodule

