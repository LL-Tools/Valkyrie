

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698;

  AOI211_X1 U4910 ( .C1(n8070), .C2(n8002), .A(n9920), .B(n8001), .ZN(n8003)
         );
  OR2_X1 U4911 ( .A1(n7101), .A2(n7078), .ZN(n9672) );
  NAND2_X1 U4912 ( .A1(n7101), .A2(n9659), .ZN(n9643) );
  BUF_X2 U4913 ( .A(n9794), .Z(n4580) );
  OAI21_X1 U4914 ( .B1(n6099), .B2(n6098), .A(n6097), .ZN(n6102) );
  CLKBUF_X1 U4915 ( .A(n9735), .Z(n4426) );
  XNOR2_X1 U4916 ( .A(n5702), .B(n5715), .ZN(n8305) );
  OR2_X1 U4917 ( .A1(n6804), .A2(n9269), .ZN(n6824) );
  BUF_X1 U4918 ( .A(n8364), .Z(n8394) );
  NAND2_X1 U4919 ( .A1(n6174), .A2(n6179), .ZN(n8915) );
  NOR2_X1 U4920 ( .A1(n6564), .A2(n6563), .ZN(n9152) );
  INV_X1 U4921 ( .A(n5842), .ZN(n6010) );
  CLKBUF_X2 U4922 ( .A(n7520), .Z(n8381) );
  AND2_X2 U4923 ( .A1(n6525), .A2(n6524), .ZN(n7021) );
  INV_X1 U4924 ( .A(n7672), .ZN(n5051) );
  NOR2_X2 U4925 ( .A1(n9592), .A2(n7811), .ZN(n7060) );
  INV_X1 U4926 ( .A(n6399), .ZN(n6947) );
  INV_X1 U4927 ( .A(n6488), .ZN(n6778) );
  INV_X2 U4928 ( .A(n6650), .ZN(n7103) );
  NAND4_X1 U4929 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n7009)
         );
  CLKBUF_X2 U4930 ( .A(n6520), .Z(n4408) );
  AND2_X1 U4931 ( .A1(n7648), .A2(n7156), .ZN(n6373) );
  INV_X2 U4932 ( .A(n6091), .ZN(n5844) );
  CLKBUF_X3 U4933 ( .A(n6944), .Z(n4427) );
  INV_X1 U4934 ( .A(n6463), .ZN(n6384) );
  AND2_X1 U4935 ( .A1(n8336), .A2(n6327), .ZN(n6427) );
  AND3_X1 U4936 ( .A1(n5225), .A2(n5224), .A3(n5223), .ZN(n7409) );
  AND2_X2 U4937 ( .A1(n6351), .A2(n6361), .ZN(n9522) );
  NAND2_X1 U4938 ( .A1(n5107), .A2(n5108), .ZN(n5257) );
  CLKBUF_X2 U4939 ( .A(n5302), .Z(n7161) );
  NOR2_X1 U4940 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4793) );
  INV_X1 U4941 ( .A(n6537), .ZN(n6933) );
  OAI21_X1 U4942 ( .B1(n4451), .B2(n4841), .A(n9758), .ZN(n4840) );
  NOR2_X1 U4943 ( .A1(n5192), .A2(n5172), .ZN(n6239) );
  AND2_X1 U4944 ( .A1(n8652), .A2(n5970), .ZN(n5971) );
  AOI22_X1 U4945 ( .A1(n8698), .A2(n8697), .B1(n6047), .B2(n6046), .ZN(n6049)
         );
  AND2_X1 U4946 ( .A1(n9276), .A2(n6674), .ZN(n9127) );
  NAND2_X1 U4947 ( .A1(n6358), .A2(n6356), .ZN(n6944) );
  OR2_X1 U4948 ( .A1(n9183), .A2(n9257), .ZN(n7995) );
  NOR2_X1 U4949 ( .A1(n10225), .A2(n7009), .ZN(n7057) );
  INV_X1 U4950 ( .A(n6121), .ZN(n7521) );
  INV_X1 U4951 ( .A(n10311), .ZN(n7573) );
  AND2_X1 U4952 ( .A1(n4869), .A2(n8702), .ZN(n5974) );
  OR2_X1 U4953 ( .A1(n6632), .A2(n10500), .ZN(n6660) );
  INV_X1 U4954 ( .A(n6906), .ZN(n8318) );
  NAND2_X1 U4955 ( .A1(n8001), .A2(n4487), .ZN(n9918) );
  INV_X1 U4956 ( .A(n4421), .ZN(n6777) );
  INV_X1 U4957 ( .A(n6086), .ZN(n5848) );
  XNOR2_X1 U4958 ( .A(n4704), .B(n8757), .ZN(n5125) );
  OAI21_X1 U4959 ( .B1(n8785), .B2(n6215), .A(n6243), .ZN(n8774) );
  OAI21_X1 U4960 ( .B1(n5811), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U4961 ( .A1(n9731), .A2(n5059), .ZN(n7077) );
  AND2_X2 U4962 ( .A1(n9483), .A2(n9490), .ZN(n9736) );
  OAI21_X1 U4963 ( .B1(n5028), .B2(n5027), .A(n5024), .ZN(n5702) );
  NAND2_X2 U4964 ( .A1(n5842), .A2(n5841), .ZN(n5243) );
  OAI22_X1 U4965 ( .A1(n8756), .A2(n8853), .B1(n8755), .B2(n10256), .ZN(n8958)
         );
  AOI211_X1 U4966 ( .C1(n7788), .C2(n7787), .A(n9340), .B(n7786), .ZN(n7789)
         );
  NOR2_X1 U4967 ( .A1(n6546), .A2(n6545), .ZN(n9257) );
  INV_X1 U4968 ( .A(n9926), .ZN(n9930) );
  XNOR2_X1 U4969 ( .A(n5406), .B(n5424), .ZN(n7201) );
  INV_X1 U4970 ( .A(n10282), .ZN(n10296) );
  OAI211_X1 U4971 ( .C1(n9479), .C2(n7993), .A(n9478), .B(n9523), .ZN(n9582)
         );
  INV_X1 U4972 ( .A(n7021), .ZN(n9591) );
  AND2_X1 U4973 ( .A1(n7097), .A2(n7096), .ZN(n10067) );
  CLKBUF_X3 U4974 ( .A(n6386), .Z(n4429) );
  INV_X1 U4975 ( .A(n5243), .ZN(n5621) );
  AND2_X1 U4976 ( .A1(n8408), .A2(n5229), .ZN(n4404) );
  NAND2_X2 U4977 ( .A1(n8539), .A2(n8380), .ZN(n8427) );
  NAND2_X2 U4978 ( .A1(n5071), .A2(n5069), .ZN(n8539) );
  AND2_X1 U4979 ( .A1(n9451), .A2(n7837), .ZN(n6356) );
  NAND2_X1 U4980 ( .A1(n5243), .A2(n6393), .ZN(n4405) );
  NAND2_X1 U4981 ( .A1(n5243), .A2(n6393), .ZN(n4406) );
  NAND2_X1 U4982 ( .A1(n5243), .A2(n6393), .ZN(n6104) );
  INV_X1 U4983 ( .A(n6104), .ZN(n5622) );
  NAND2_X2 U4984 ( .A1(n7758), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U4985 ( .A1(n8061), .A2(n4718), .ZN(n4717) );
  AND2_X2 U4986 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8061) );
  INV_X2 U4987 ( .A(n6114), .ZN(n7385) );
  NAND2_X2 U4988 ( .A1(n7976), .A2(n7062), .ZN(n8025) );
  AND3_X4 U4989 ( .A1(n6453), .A2(n6452), .A3(n6451), .ZN(n7637) );
  NOR2_X2 U4990 ( .A1(n7755), .A2(n4787), .ZN(n7953) );
  NOR2_X2 U4991 ( .A1(n7757), .A2(n7756), .ZN(n7755) );
  NAND2_X2 U4992 ( .A1(n4920), .A2(n4919), .ZN(n9741) );
  NAND2_X2 U4993 ( .A1(n9804), .A2(n9411), .ZN(n9788) );
  NAND2_X2 U4994 ( .A1(n8311), .A2(n6324), .ZN(n6463) );
  BUF_X4 U4995 ( .A(n5621), .Z(n4407) );
  AOI21_X2 U4996 ( .B1(n7007), .B2(n4418), .A(n6357), .ZN(n6379) );
  AOI21_X2 U4997 ( .B1(n4630), .B2(n9988), .A(n4627), .ZN(n9964) );
  AOI21_X2 U4998 ( .B1(n5755), .B2(n5754), .A(n5753), .ZN(n5770) );
  XNOR2_X2 U4999 ( .A(n7118), .B(n9475), .ZN(n9665) );
  INV_X1 U5000 ( .A(n8482), .ZN(n9102) );
  NAND2_X2 U5001 ( .A1(n5481), .A2(n5480), .ZN(n8482) );
  OAI22_X2 U5002 ( .A1(n8285), .A2(n8286), .B1(n6036), .B2(n7208), .ZN(n8627)
         );
  AOI22_X2 U5003 ( .A1(n8248), .A2(n8249), .B1(n6035), .B2(n6034), .ZN(n8285)
         );
  XNOR2_X2 U5004 ( .A(n6390), .B(n6389), .ZN(n7218) );
  NAND2_X1 U5005 ( .A1(n6929), .A2(n6928), .ZN(n9321) );
  NAND2_X1 U5006 ( .A1(n5120), .A2(n5123), .ZN(n6083) );
  CLKBUF_X1 U5008 ( .A(n9752), .Z(n4611) );
  NAND2_X1 U5009 ( .A1(n9856), .A2(n9868), .ZN(n9837) );
  OR2_X1 U5010 ( .A1(n5834), .A2(n5116), .ZN(n5115) );
  NAND2_X1 U5011 ( .A1(n8797), .A2(n6201), .ZN(n8829) );
  NAND2_X1 U5012 ( .A1(n6745), .A2(n6744), .ZN(n10020) );
  NAND2_X1 U5013 ( .A1(n5636), .A2(n5635), .ZN(n5662) );
  NAND2_X1 U5014 ( .A1(n9370), .A2(n9380), .ZN(n9460) );
  NAND2_X2 U5015 ( .A1(n6155), .A2(n6156), .ZN(n8345) );
  INV_X1 U5016 ( .A(n9863), .ZN(n9921) );
  INV_X2 U5017 ( .A(n10252), .ZN(n4409) );
  INV_X1 U5018 ( .A(n7917), .ZN(n7914) );
  INV_X2 U5019 ( .A(n10285), .ZN(n7894) );
  INV_X1 U5020 ( .A(n8604), .ZN(n8554) );
  INV_X1 U5021 ( .A(n10275), .ZN(n7930) );
  INV_X1 U5022 ( .A(n10276), .ZN(n7617) );
  INV_X4 U5023 ( .A(n6241), .ZN(n6237) );
  BUF_X1 U5024 ( .A(n6358), .Z(n7156) );
  AND3_X1 U5025 ( .A1(n5262), .A2(n5261), .A3(n5260), .ZN(n10302) );
  BUF_X2 U5026 ( .A(n6488), .Z(n6930) );
  BUF_X1 U5027 ( .A(n7751), .Z(n4428) );
  XNOR2_X1 U5028 ( .A(n6083), .B(n6242), .ZN(n8742) );
  AND2_X1 U5029 ( .A1(n4938), .A2(n4939), .ZN(n7055) );
  NAND2_X1 U5030 ( .A1(n5835), .A2(n6245), .ZN(n8785) );
  NAND2_X1 U5031 ( .A1(n8947), .A2(n8599), .ZN(n6272) );
  CLKBUF_X1 U5032 ( .A(n9819), .Z(n4413) );
  AOI21_X1 U5033 ( .B1(n4837), .B2(n4687), .A(n4692), .ZN(n4691) );
  NAND2_X1 U5034 ( .A1(n6897), .A2(n6896), .ZN(n9961) );
  NAND2_X1 U5035 ( .A1(n6181), .A2(n6180), .ZN(n8898) );
  NAND2_X1 U5036 ( .A1(n9054), .A2(n8816), .ZN(n6201) );
  OR2_X1 U5037 ( .A1(n8998), .A2(n8893), .ZN(n6174) );
  NAND2_X1 U5038 ( .A1(n8025), .A2(n7063), .ZN(n8115) );
  XNOR2_X1 U5039 ( .A(n5662), .B(n5637), .ZN(n7991) );
  NAND2_X2 U5040 ( .A1(n9359), .A2(n9347), .ZN(n9452) );
  NAND2_X1 U5041 ( .A1(n5428), .A2(n5420), .ZN(n5405) );
  AND2_X1 U5042 ( .A1(n5017), .A2(n6358), .ZN(n6418) );
  BUF_X2 U5043 ( .A(n5291), .Z(n6091) );
  INV_X1 U5044 ( .A(n9527), .ZN(n5016) );
  NAND2_X1 U5045 ( .A1(n5270), .A2(n5319), .ZN(n7166) );
  INV_X2 U5046 ( .A(n5302), .ZN(n5277) );
  INV_X4 U5047 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5048 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6718) );
  OAI21_X1 U5049 ( .B1(n8955), .B2(n9011), .A(n4612), .ZN(n8957) );
  NAND2_X1 U5050 ( .A1(n4698), .A2(n4697), .ZN(n10073) );
  AOI21_X1 U5051 ( .B1(n9956), .B2(n10241), .A(n4699), .ZN(n4698) );
  OR2_X1 U5052 ( .A1(n7055), .A2(n9475), .ZN(n5188) );
  NAND2_X1 U5053 ( .A1(n7055), .A2(n9475), .ZN(n7135) );
  OR3_X1 U5054 ( .A1(n9972), .A2(n9971), .A3(n9970), .ZN(n10076) );
  MUX2_X1 U5055 ( .A(n10068), .B(P1_REG0_REG_30__SCAN_IN), .S(n7144), .Z(
        n10069) );
  NAND2_X1 U5056 ( .A1(n5032), .A2(n4459), .ZN(n9639) );
  OR2_X1 U5057 ( .A1(n9661), .A2(n9660), .ZN(n9662) );
  NAND2_X1 U5058 ( .A1(n4543), .A2(n10002), .ZN(n9942) );
  OAI21_X1 U5059 ( .B1(n6193), .B2(n6194), .A(n6192), .ZN(n6200) );
  AND2_X1 U5060 ( .A1(n9945), .A2(n9585), .ZN(n4412) );
  AND2_X1 U5061 ( .A1(n6271), .A2(n6081), .ZN(n6234) );
  CLKBUF_X1 U5062 ( .A(n8858), .Z(n4589) );
  NAND2_X1 U5063 ( .A1(n9505), .A2(n9507), .ZN(n9651) );
  NAND2_X1 U5064 ( .A1(n7105), .A2(n7104), .ZN(n9945) );
  NAND2_X1 U5065 ( .A1(n6080), .A2(n6079), .ZN(n6085) );
  NOR2_X1 U5066 ( .A1(n9317), .A2(n9318), .ZN(n6928) );
  AOI21_X1 U5067 ( .B1(n4732), .B2(n4734), .A(n5158), .ZN(n4731) );
  OR2_X1 U5068 ( .A1(n5805), .A2(n8398), .ZN(n6236) );
  AOI21_X1 U5069 ( .B1(n4437), .B2(n4984), .A(n4980), .ZN(n4979) );
  CLKBUF_X1 U5070 ( .A(n7102), .Z(n8335) );
  NAND2_X1 U5071 ( .A1(n7100), .A2(n7099), .ZN(n7119) );
  XNOR2_X1 U5072 ( .A(n6102), .B(n6101), .ZN(n10109) );
  AND2_X1 U5073 ( .A1(n6873), .A2(n6872), .ZN(n9241) );
  NAND2_X1 U5074 ( .A1(n6648), .A2(n9195), .ZN(n9197) );
  XNOR2_X1 U5075 ( .A(n6075), .B(SI_29_), .ZN(n7098) );
  NAND2_X2 U5076 ( .A1(n7054), .A2(n7053), .ZN(n9675) );
  AND2_X1 U5077 ( .A1(n9497), .A2(n9434), .ZN(n9693) );
  NAND2_X1 U5078 ( .A1(n9959), .A2(n9946), .ZN(n9434) );
  NAND2_X1 U5079 ( .A1(n4581), .A2(n5796), .ZN(n6075) );
  NAND2_X1 U5080 ( .A1(n5761), .A2(n5760), .ZN(n8762) );
  NAND2_X1 U5081 ( .A1(n6932), .A2(n6931), .ZN(n9680) );
  NAND2_X2 U5082 ( .A1(n4591), .A2(n6910), .ZN(n9959) );
  OR2_X1 U5083 ( .A1(n9034), .A2(n8578), .ZN(n6213) );
  XNOR2_X1 U5084 ( .A(n6070), .B(n6069), .ZN(n8409) );
  NAND2_X1 U5085 ( .A1(n5722), .A2(n5721), .ZN(n9034) );
  XNOR2_X1 U5087 ( .A(n5740), .B(n5739), .ZN(n9117) );
  AND2_X1 U5088 ( .A1(n4474), .A2(n4442), .ZN(n4812) );
  NAND2_X1 U5089 ( .A1(n5770), .A2(n5769), .ZN(n5785) );
  INV_X1 U5090 ( .A(n5115), .ZN(n4410) );
  AND2_X1 U5091 ( .A1(n9397), .A2(n9838), .ZN(n9868) );
  NAND2_X1 U5092 ( .A1(n9253), .A2(n6576), .ZN(n6595) );
  AOI22_X1 U5093 ( .A1(n8627), .A2(n8628), .B1(n6038), .B2(n8633), .ZN(n8643)
         );
  AND2_X1 U5094 ( .A1(n8825), .A2(n8465), .ZN(n6204) );
  NAND2_X1 U5095 ( .A1(n8119), .A2(n9460), .ZN(n8118) );
  NAND2_X1 U5096 ( .A1(n6852), .A2(n6851), .ZN(n9763) );
  AND2_X1 U5097 ( .A1(n4472), .A2(n8654), .ZN(n8636) );
  CLKBUF_X1 U5098 ( .A(n9054), .Z(n4558) );
  XNOR2_X1 U5099 ( .A(n5696), .B(n5695), .ZN(n8245) );
  XNOR2_X1 U5100 ( .A(n9996), .B(n9792), .ZN(n9783) );
  NAND2_X1 U5101 ( .A1(n5668), .A2(n5667), .ZN(n8825) );
  OR2_X1 U5102 ( .A1(n9866), .A2(n9881), .ZN(n9397) );
  AND2_X1 U5103 ( .A1(n5135), .A2(n5828), .ZN(n5134) );
  NAND2_X1 U5104 ( .A1(n5968), .A2(n7274), .ZN(n8649) );
  NAND2_X2 U5105 ( .A1(n6822), .A2(n6821), .ZN(n9996) );
  NAND2_X1 U5106 ( .A1(n8115), .A2(n9380), .ZN(n9901) );
  NAND2_X1 U5107 ( .A1(n5652), .A2(n5651), .ZN(n9060) );
  XNOR2_X1 U5108 ( .A(n5579), .B(n5578), .ZN(n7547) );
  AND2_X1 U5109 ( .A1(n5997), .A2(n8296), .ZN(n8256) );
  NAND2_X1 U5110 ( .A1(n5537), .A2(n5536), .ZN(n8998) );
  CLKBUF_X1 U5111 ( .A(n9086), .Z(n4626) );
  OAI21_X1 U5112 ( .B1(n7898), .B2(n5366), .A(n5365), .ZN(n10253) );
  NAND2_X1 U5113 ( .A1(n6780), .A2(n6779), .ZN(n10084) );
  NAND2_X1 U5114 ( .A1(n6654), .A2(n6653), .ZN(n10048) );
  XNOR2_X1 U5115 ( .A(n5574), .B(n5533), .ZN(n7489) );
  NAND2_X1 U5116 ( .A1(n6678), .A2(n6677), .ZN(n10042) );
  OAI21_X1 U5117 ( .B1(n10283), .B2(n5290), .A(n5289), .ZN(n10274) );
  NAND2_X1 U5118 ( .A1(n5043), .A2(n5047), .ZN(n5574) );
  AND2_X1 U5119 ( .A1(n7854), .A2(n7853), .ZN(n7856) );
  NAND2_X1 U5120 ( .A1(n6629), .A2(n6628), .ZN(n10095) );
  NAND2_X1 U5121 ( .A1(n6823), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6854) );
  INV_X1 U5122 ( .A(n6824), .ZN(n6823) );
  NAND2_X1 U5123 ( .A1(n7075), .A2(n8151), .ZN(n8002) );
  OR2_X1 U5124 ( .A1(n8548), .A2(n8473), .ZN(n6155) );
  NAND2_X1 U5125 ( .A1(n5498), .A2(n5497), .ZN(n5516) );
  INV_X1 U5126 ( .A(n9157), .ZN(n4411) );
  NAND2_X1 U5127 ( .A1(n6604), .A2(n6603), .ZN(n7027) );
  NAND2_X1 U5128 ( .A1(n5438), .A2(n5437), .ZN(n8444) );
  OR2_X1 U5129 ( .A1(n8226), .A2(n8339), .ZN(n8233) );
  AND2_X1 U5130 ( .A1(n9360), .A2(n9351), .ZN(n7824) );
  NAND2_X1 U5131 ( .A1(n4762), .A2(n5410), .ZN(n8226) );
  AND2_X1 U5132 ( .A1(n5960), .A2(n7966), .ZN(n7758) );
  NAND2_X1 U5133 ( .A1(n6746), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6782) );
  INV_X1 U5134 ( .A(n6748), .ZN(n6746) );
  NAND2_X1 U5135 ( .A1(n8609), .A2(n10297), .ZN(n6116) );
  INV_X1 U5136 ( .A(n7812), .ZN(n9593) );
  AND2_X2 U5137 ( .A1(n6496), .A2(n6495), .ZN(n7811) );
  NOR2_X2 U5138 ( .A1(n6473), .A2(n6472), .ZN(n7812) );
  NAND4_X2 U5139 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n10285)
         );
  AOI21_X1 U5140 ( .B1(n4497), .B2(n4721), .A(n4443), .ZN(n4719) );
  NAND4_X2 U5141 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n9594)
         );
  INV_X1 U5142 ( .A(n10231), .ZN(n7652) );
  NAND4_X2 U5143 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n9592)
         );
  NAND3_X2 U5144 ( .A1(n6431), .A2(n6430), .A3(n4450), .ZN(n9595) );
  INV_X2 U5145 ( .A(n4424), .ZN(n5845) );
  AND2_X2 U5146 ( .A1(n6374), .A2(n6373), .ZN(n6906) );
  INV_X1 U5148 ( .A(n6418), .ZN(n6537) );
  CLKBUF_X3 U5149 ( .A(n6399), .Z(n8316) );
  AND3_X2 U5150 ( .A1(n6417), .A2(n6416), .A3(n6415), .ZN(n10225) );
  AND2_X1 U5151 ( .A1(n7838), .A2(n5854), .ZN(n7384) );
  AND2_X2 U5152 ( .A1(n6326), .A2(n6324), .ZN(n6937) );
  INV_X2 U5153 ( .A(n5286), .ZN(n6106) );
  NAND2_X1 U5154 ( .A1(n6962), .A2(n6343), .ZN(n6358) );
  INV_X1 U5155 ( .A(n7751), .ZN(n5854) );
  AND2_X1 U5156 ( .A1(n6392), .A2(n6391), .ZN(n6396) );
  OR2_X1 U5157 ( .A1(n4406), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5224) );
  AND2_X1 U5158 ( .A1(n5042), .A2(n5555), .ZN(n5041) );
  AND2_X1 U5159 ( .A1(n6336), .A2(n6335), .ZN(n6962) );
  NAND2_X1 U5160 ( .A1(n6367), .A2(n6973), .ZN(n8177) );
  NAND2_X1 U5161 ( .A1(n6321), .A2(n6320), .ZN(n8336) );
  NAND2_X1 U5162 ( .A1(n5811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U5163 ( .A1(n4622), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6609) );
  AOI21_X1 U5164 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n7458), .A(n7450), .ZN(
        n7217) );
  XNOR2_X1 U5165 ( .A(n5351), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7179) );
  MUX2_X1 U5166 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6333), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6336) );
  NAND3_X1 U5167 ( .A1(n4547), .A2(n4590), .A3(n5276), .ZN(n5326) );
  MUX2_X1 U5168 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6338), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6339) );
  AND2_X1 U5169 ( .A1(n5375), .A2(n5357), .ZN(n5358) );
  INV_X1 U5170 ( .A(n6584), .ZN(n4622) );
  XNOR2_X1 U5171 ( .A(n5228), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5229) );
  XNOR2_X1 U5172 ( .A(n6349), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U5173 ( .A1(n6558), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6584) );
  INV_X2 U5174 ( .A(n10108), .ZN(n8337) );
  NAND2_X1 U5175 ( .A1(n5377), .A2(SI_7_), .ZN(n5420) );
  NAND2_X1 U5176 ( .A1(n6361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6349) );
  AND2_X1 U5177 ( .A1(n6539), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U5178 ( .A1(n10102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U5179 ( .A(n6434), .B(n6433), .ZN(n7222) );
  AND2_X1 U5180 ( .A1(n6516), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U5181 ( .A1(n6432), .A2(n4737), .ZN(n7221) );
  NOR2_X1 U5182 ( .A1(n6498), .A2(n6497), .ZN(n6516) );
  OR2_X1 U5183 ( .A1(n5259), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5319) );
  INV_X4 U5184 ( .A(n5302), .ZN(n6393) );
  NAND2_X1 U5185 ( .A1(n6466), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6498) );
  AND2_X1 U5186 ( .A1(n6475), .A2(n6312), .ZN(n4682) );
  AND2_X1 U5187 ( .A1(n6311), .A2(n6345), .ZN(n5039) );
  AND4_X1 U5188 ( .A1(n6718), .A2(n6368), .A3(n6362), .A4(n6365), .ZN(n6313)
         );
  AND2_X1 U5189 ( .A1(n6310), .A2(n6309), .ZN(n6312) );
  AND4_X1 U5190 ( .A1(n6345), .A2(n6718), .A3(n6719), .A4(n6344), .ZN(n6347)
         );
  INV_X1 U5191 ( .A(n6468), .ZN(n6466) );
  NAND2_X1 U5192 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6468) );
  NOR2_X1 U5193 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4792) );
  NOR2_X1 U5194 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4791) );
  NOR2_X1 U5195 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6345) );
  INV_X1 U5196 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5108) );
  INV_X4 U5197 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5198 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5856) );
  INV_X1 U5199 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U5200 ( .A1(n9441), .A2(n4412), .ZN(n9442) );
  AND2_X1 U5201 ( .A1(n7088), .A2(n4618), .ZN(n4414) );
  NAND2_X2 U5202 ( .A1(n5229), .A2(n5233), .ZN(n5292) );
  OAI21_X1 U5203 ( .B1(n9678), .B2(n10211), .A(n7087), .ZN(n4619) );
  CLKBUF_X1 U5204 ( .A(n9193), .Z(n4415) );
  CLKBUF_X1 U5205 ( .A(n7511), .Z(n4416) );
  AND2_X1 U5206 ( .A1(n9128), .A2(n9127), .ZN(n4417) );
  NOR2_X1 U5207 ( .A1(n4417), .A2(n9219), .ZN(n9129) );
  INV_X1 U5208 ( .A(n6944), .ZN(n4418) );
  NOR2_X1 U5209 ( .A1(n9127), .A2(n9128), .ZN(n9219) );
  XNOR2_X2 U5210 ( .A(n4419), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6387) );
  NOR2_X1 U5211 ( .A1(n6334), .A2(n6651), .ZN(n4419) );
  NAND2_X2 U5212 ( .A1(n9197), .A2(n6649), .ZN(n9277) );
  MUX2_X1 U5213 ( .A(n9490), .B(n9483), .S(n9449), .Z(n9424) );
  OAI21_X1 U5214 ( .B1(n5302), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n4632), .ZN(
        n5253) );
  NAND2_X1 U5215 ( .A1(n5067), .A2(n10276), .ZN(n5066) );
  NAND2_X1 U5216 ( .A1(n4720), .A2(n4719), .ZN(n5634) );
  NOR2_X2 U5217 ( .A1(n8002), .A2(n8070), .ZN(n8001) );
  OR2_X2 U5218 ( .A1(n8070), .A2(n9152), .ZN(n9365) );
  NAND2_X2 U5219 ( .A1(n6387), .A2(n4429), .ZN(n4420) );
  NAND2_X2 U5220 ( .A1(n6387), .A2(n4429), .ZN(n4421) );
  INV_X1 U5221 ( .A(n4660), .ZN(n4659) );
  OAI21_X1 U5222 ( .B1(n9425), .B2(n9424), .A(n9493), .ZN(n4660) );
  NAND2_X1 U5223 ( .A1(n9837), .A2(n7067), .ZN(n9839) );
  INV_X1 U5224 ( .A(n5229), .ZN(n9108) );
  NAND3_X4 U5225 ( .A1(n5180), .A2(n5197), .A3(n6385), .ZN(n6400) );
  AND2_X2 U5226 ( .A1(n6383), .A2(n6382), .ZN(n5197) );
  NAND2_X2 U5227 ( .A1(n6384), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6385) );
  INV_X4 U5228 ( .A(n4427), .ZN(n8313) );
  NOR2_X2 U5229 ( .A1(n7797), .A2(n5068), .ZN(n8013) );
  NOR2_X2 U5230 ( .A1(n7690), .A2(n7689), .ZN(n7797) );
  AND2_X1 U5231 ( .A1(n6374), .A2(n6373), .ZN(n4422) );
  AND2_X1 U5232 ( .A1(n6374), .A2(n6373), .ZN(n4423) );
  INV_X2 U5233 ( .A(n4404), .ZN(n4424) );
  NAND2_X2 U5234 ( .A1(n6595), .A2(n6594), .ZN(n9295) );
  NOR2_X2 U5235 ( .A1(n9243), .A2(n6895), .ZN(n9209) );
  NAND2_X1 U5236 ( .A1(n5243), .A2(n7161), .ZN(n4425) );
  XNOR2_X1 U5237 ( .A(n5405), .B(n5404), .ZN(n7190) );
  NAND2_X1 U5238 ( .A1(n6876), .A2(n6875), .ZN(n9735) );
  NAND2_X1 U5239 ( .A1(n9365), .A2(n7995), .ZN(n9350) );
  OAI21_X2 U5240 ( .B1(n9872), .B2(n7037), .A(n7036), .ZN(n9867) );
  XNOR2_X1 U5241 ( .A(n5620), .B(n5808), .ZN(n7751) );
  AND2_X1 U5242 ( .A1(n8336), .A2(n6326), .ZN(n6520) );
  NAND3_X2 U5243 ( .A1(n5167), .A2(n9540), .A3(n9456), .ZN(n7976) );
  OR2_X2 U5244 ( .A1(n9464), .A2(n7061), .ZN(n9540) );
  OAI21_X2 U5245 ( .B1(n5405), .B2(n5404), .A(n5422), .ZN(n5406) );
  XNOR2_X2 U5246 ( .A(n5209), .B(n10387), .ZN(n5841) );
  NOR2_X2 U5247 ( .A1(n9464), .A2(n7060), .ZN(n9535) );
  OR2_X1 U5248 ( .A1(n5302), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5216) );
  OAI21_X2 U5249 ( .B1(n7805), .B2(n7806), .A(n7807), .ZN(n7866) );
  NAND2_X2 U5250 ( .A1(n6487), .A2(n7842), .ZN(n7805) );
  NOR2_X1 U5251 ( .A1(n9959), .A2(n9961), .ZN(n5060) );
  NAND2_X1 U5252 ( .A1(n5531), .A2(SI_14_), .ZN(n5047) );
  NOR2_X1 U5253 ( .A1(n8459), .A2(n5076), .ZN(n5075) );
  INV_X1 U5254 ( .A(n8371), .ZN(n5076) );
  AND2_X1 U5255 ( .A1(n4440), .A2(n5733), .ZN(n4823) );
  OR2_X1 U5256 ( .A1(n9675), .A2(n9947), .ZN(n9504) );
  NAND2_X1 U5257 ( .A1(n9675), .A2(n9947), .ZN(n9427) );
  OR2_X1 U5258 ( .A1(n9959), .A2(n9946), .ZN(n9497) );
  AND2_X1 U5259 ( .A1(n4923), .A2(n7047), .ZN(n4922) );
  NAND2_X1 U5260 ( .A1(n4925), .A2(n4927), .ZN(n4923) );
  NAND2_X1 U5261 ( .A1(n7132), .A2(n5057), .ZN(n5056) );
  INV_X1 U5262 ( .A(n5059), .ZN(n5057) );
  INV_X1 U5263 ( .A(n5595), .ZN(n4725) );
  INV_X1 U5264 ( .A(n5292), .ZN(n5799) );
  INV_X1 U5265 ( .A(n4733), .ZN(n4732) );
  OAI21_X1 U5266 ( .B1(n7070), .B2(n4734), .A(n9693), .ZN(n4733) );
  AND2_X1 U5267 ( .A1(n9521), .A2(n9451), .ZN(n7184) );
  NAND2_X1 U5268 ( .A1(n6186), .A2(n4755), .ZN(n4754) );
  AND2_X1 U5269 ( .A1(n6189), .A2(n6247), .ZN(n4755) );
  NAND2_X1 U5270 ( .A1(n9388), .A2(n4673), .ZN(n4671) );
  AND2_X1 U5271 ( .A1(n4674), .A2(n9840), .ZN(n4673) );
  NAND2_X1 U5272 ( .A1(n6203), .A2(n4465), .ZN(n4563) );
  INV_X1 U5273 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5200) );
  AOI211_X1 U5274 ( .C1(n9428), .C2(n9497), .A(n9449), .B(n9433), .ZN(n9430)
         );
  NAND2_X1 U5275 ( .A1(n9418), .A2(n4656), .ZN(n4655) );
  INV_X1 U5276 ( .A(n8457), .ZN(n8377) );
  NOR2_X1 U5277 ( .A1(n8351), .A2(n5092), .ZN(n5091) );
  INV_X1 U5278 ( .A(n8341), .ZN(n5092) );
  XNOR2_X1 U5279 ( .A(n5232), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U5280 ( .A1(n8204), .A2(n5995), .ZN(n5996) );
  AOI21_X1 U5281 ( .B1(n4855), .B2(n4854), .A(n4850), .ZN(n5968) );
  NAND2_X1 U5282 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  NOR2_X1 U5283 ( .A1(n4859), .A2(n4856), .ZN(n4855) );
  NAND2_X1 U5284 ( .A1(n4531), .A2(n5967), .ZN(n4851) );
  INV_X1 U5285 ( .A(n5653), .ZN(n5641) );
  OR2_X1 U5286 ( .A1(n9028), .A2(n8755), .ZN(n6221) );
  INV_X1 U5287 ( .A(n5694), .ZN(n4806) );
  INV_X1 U5288 ( .A(n6195), .ZN(n5116) );
  OR2_X1 U5289 ( .A1(n9045), .A2(n8817), .ZN(n6246) );
  OR2_X1 U5290 ( .A1(n9054), .A2(n8816), .ZN(n8797) );
  OR2_X1 U5291 ( .A1(n9060), .A2(n8855), .ZN(n6196) );
  OR2_X1 U5292 ( .A1(n8871), .A2(n8883), .ZN(n6247) );
  OR2_X1 U5293 ( .A1(n9071), .A2(n8894), .ZN(n6261) );
  OR2_X1 U5294 ( .A1(n8902), .A2(n8908), .ZN(n6181) );
  INV_X1 U5295 ( .A(n6156), .ZN(n5136) );
  OAI21_X1 U5296 ( .B1(n9102), .B2(n8931), .A(n5824), .ZN(n5825) );
  AND2_X1 U5297 ( .A1(n5211), .A2(n5138), .ZN(n5137) );
  OR2_X1 U5298 ( .A1(n7867), .A2(n7868), .ZN(n5000) );
  NAND2_X1 U5299 ( .A1(n7867), .A2(n7868), .ZN(n4999) );
  INV_X1 U5300 ( .A(n4999), .ZN(n4998) );
  OR2_X1 U5301 ( .A1(n7119), .A2(n9671), .ZN(n9505) );
  AND2_X1 U5302 ( .A1(n4943), .A2(n5156), .ZN(n4941) );
  NAND2_X1 U5303 ( .A1(n9693), .A2(n7052), .ZN(n4947) );
  INV_X1 U5304 ( .A(n4925), .ZN(n4924) );
  NAND2_X1 U5305 ( .A1(n9788), .A2(n9789), .ZN(n9794) );
  NAND2_X1 U5306 ( .A1(n7045), .A2(n7044), .ZN(n9787) );
  NOR2_X1 U5307 ( .A1(n4460), .A2(n4954), .ZN(n4953) );
  OR2_X1 U5308 ( .A1(n10084), .A2(n9233), .ZN(n9410) );
  OR2_X1 U5309 ( .A1(n10034), .A2(n10039), .ZN(n9393) );
  NOR2_X1 U5310 ( .A1(n7007), .A2(n7074), .ZN(n7603) );
  NAND2_X1 U5311 ( .A1(n5785), .A2(n5787), .ZN(n6070) );
  NAND2_X1 U5312 ( .A1(n5735), .A2(n5734), .ZN(n5755) );
  INV_X1 U5313 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6362) );
  AOI21_X1 U5314 ( .B1(n4723), .B2(n5045), .A(n4722), .ZN(n4721) );
  INV_X1 U5315 ( .A(n5594), .ZN(n4722) );
  NAND2_X1 U5316 ( .A1(n5594), .A2(n5559), .ZN(n5595) );
  NAND2_X1 U5317 ( .A1(n5493), .A2(SI_13_), .ZN(n5515) );
  NAND2_X1 U5318 ( .A1(n5463), .A2(SI_12_), .ZN(n5491) );
  INV_X1 U5319 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U5320 ( .A1(n5428), .A2(n5426), .ZN(n4951) );
  XNOR2_X1 U5321 ( .A(n5430), .B(SI_9_), .ZN(n5424) );
  NAND2_X1 U5322 ( .A1(n5302), .A2(n7164), .ZN(n4632) );
  INV_X1 U5323 ( .A(n5083), .ZN(n5082) );
  OAI21_X1 U5324 ( .B1(n8487), .B2(n5084), .A(n8574), .ZN(n5083) );
  XNOR2_X1 U5325 ( .A(n8762), .B(n8394), .ZN(n8392) );
  OR2_X1 U5326 ( .A1(n8360), .A2(n8893), .ZN(n8361) );
  INV_X1 U5327 ( .A(n5066), .ZN(n5064) );
  AOI21_X1 U5328 ( .B1(n5072), .B2(n5074), .A(n5070), .ZN(n5069) );
  INV_X1 U5329 ( .A(n8541), .ZN(n5070) );
  NAND2_X1 U5330 ( .A1(n9021), .A2(n8737), .ZN(n6284) );
  AND2_X1 U5331 ( .A1(n5768), .A2(n5767), .ZN(n8401) );
  NAND2_X1 U5332 ( .A1(n5233), .A2(n9108), .ZN(n5291) );
  NAND2_X1 U5333 ( .A1(n5992), .A2(n7956), .ZN(n7961) );
  NAND2_X1 U5334 ( .A1(n7959), .A2(n7957), .ZN(n5992) );
  OR2_X1 U5335 ( .A1(n5561), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5446) );
  OR2_X1 U5336 ( .A1(n5968), .A2(n7274), .ZN(n5969) );
  INV_X1 U5337 ( .A(n4823), .ZN(n4822) );
  AOI21_X1 U5338 ( .B1(n4823), .B2(n4821), .A(n4820), .ZN(n4819) );
  AND2_X1 U5339 ( .A1(n4440), .A2(n4508), .ZN(n4820) );
  OR2_X1 U5340 ( .A1(n8871), .A2(n8601), .ZN(n5609) );
  OR2_X1 U5341 ( .A1(n5584), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5586) );
  INV_X1 U5342 ( .A(n5125), .ZN(n8395) );
  NAND2_X1 U5343 ( .A1(n6237), .A2(n7404), .ZN(n10254) );
  AOI21_X1 U5344 ( .B1(n4831), .B2(n4829), .A(n4479), .ZN(n4828) );
  INV_X1 U5345 ( .A(n4834), .ZN(n4829) );
  NAND2_X1 U5346 ( .A1(n8271), .A2(n8345), .ZN(n5458) );
  INV_X1 U5347 ( .A(n10254), .ZN(n10284) );
  AND2_X1 U5348 ( .A1(n7402), .A2(n6237), .ZN(n10286) );
  INV_X1 U5349 ( .A(n8853), .ZN(n10289) );
  INV_X1 U5350 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10387) );
  INV_X1 U5351 ( .A(n6715), .ZN(n4991) );
  NAND2_X1 U5352 ( .A1(n4986), .A2(n4989), .ZN(n4985) );
  NAND2_X1 U5353 ( .A1(n6840), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6879) );
  INV_X1 U5354 ( .A(n6854), .ZN(n6840) );
  AND2_X1 U5355 ( .A1(n6972), .A2(n7111), .ZN(n6991) );
  AND3_X1 U5356 ( .A1(n4971), .A2(n9613), .A3(n4970), .ZN(n10178) );
  NAND2_X1 U5357 ( .A1(n9504), .A2(n9427), .ZN(n9475) );
  OR2_X1 U5358 ( .A1(n9667), .A2(n6465), .ZN(n6987) );
  INV_X1 U5359 ( .A(n5060), .ZN(n5058) );
  OR2_X1 U5360 ( .A1(n9711), .A2(n7070), .ZN(n4631) );
  INV_X1 U5361 ( .A(n4840), .ZN(n4839) );
  INV_X1 U5362 ( .A(n4932), .ZN(n4929) );
  OR2_X1 U5363 ( .A1(n10001), .A2(n9992), .ZN(n9403) );
  NAND2_X1 U5364 ( .A1(n7121), .A2(n9643), .ZN(n9652) );
  INV_X1 U5365 ( .A(n7119), .ZN(n9659) );
  AND2_X1 U5366 ( .A1(n9672), .A2(n7086), .ZN(n7087) );
  NAND2_X1 U5367 ( .A1(n9950), .A2(n10241), .ZN(n4596) );
  NOR2_X1 U5368 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6310) );
  NOR2_X1 U5369 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6309) );
  INV_X1 U5370 ( .A(n8779), .ZN(n8755) );
  INV_X1 U5371 ( .A(n8788), .ZN(n8817) );
  NAND2_X1 U5372 ( .A1(n4705), .A2(n5779), .ZN(n8757) );
  NAND2_X1 U5373 ( .A1(n8399), .A2(n5799), .ZN(n4705) );
  INV_X1 U5374 ( .A(n8401), .ZN(n8768) );
  OR2_X1 U5375 ( .A1(n4429), .A2(n5048), .ZN(n7215) );
  NAND2_X1 U5376 ( .A1(n9710), .A2(n9431), .ZN(n9694) );
  NAND2_X1 U5377 ( .A1(n8335), .A2(n7103), .ZN(n7105) );
  NAND2_X1 U5378 ( .A1(n6128), .A2(n6127), .ZN(n6144) );
  INV_X1 U5379 ( .A(n6165), .ZN(n4772) );
  INV_X1 U5380 ( .A(n9353), .ZN(n4644) );
  OR2_X1 U5381 ( .A1(n7060), .A2(n9449), .ZN(n4640) );
  AOI21_X1 U5382 ( .B1(n4646), .B2(n4643), .A(n9342), .ZN(n4642) );
  INV_X1 U5383 ( .A(n9362), .ZN(n4643) );
  AOI21_X1 U5384 ( .B1(n9355), .B2(n9354), .A(n9449), .ZN(n4638) );
  NAND2_X1 U5385 ( .A1(n9355), .A2(n9354), .ZN(n4639) );
  AND2_X1 U5386 ( .A1(n6263), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5387 ( .A1(n8926), .A2(n4773), .ZN(n4768) );
  NAND2_X1 U5388 ( .A1(n4753), .A2(n4752), .ZN(n6193) );
  NAND2_X1 U5389 ( .A1(n6187), .A2(n6241), .ZN(n4752) );
  NAND2_X1 U5390 ( .A1(n4754), .A2(n6237), .ZN(n4753) );
  AOI21_X1 U5391 ( .B1(n4677), .B2(n4676), .A(n4453), .ZN(n4667) );
  NOR2_X1 U5392 ( .A1(n4672), .A2(n9556), .ZN(n4670) );
  NOR2_X1 U5393 ( .A1(n4672), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U5394 ( .A1(n4676), .A2(n4453), .ZN(n4669) );
  NAND2_X1 U5395 ( .A1(n9422), .A2(n9736), .ZN(n4665) );
  NOR2_X1 U5396 ( .A1(n6213), .A2(n6241), .ZN(n4760) );
  AND2_X1 U5397 ( .A1(n6243), .A2(n6246), .ZN(n4567) );
  NAND2_X1 U5398 ( .A1(n6212), .A2(n4821), .ZN(n4761) );
  INV_X1 U5399 ( .A(n9454), .ZN(n4608) );
  NOR2_X1 U5400 ( .A1(n4610), .A2(n10213), .ZN(n4609) );
  INV_X1 U5401 ( .A(n5104), .ZN(n5103) );
  NAND2_X1 U5402 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5099) );
  INV_X1 U5403 ( .A(n5099), .ZN(n5095) );
  NAND2_X1 U5404 ( .A1(n4411), .A2(n9590), .ZN(n9373) );
  INV_X1 U5405 ( .A(n5047), .ZN(n5046) );
  INV_X1 U5406 ( .A(n5982), .ZN(n4891) );
  NOR2_X1 U5407 ( .A1(n4434), .A2(n8231), .ZN(n4874) );
  NOR2_X1 U5408 ( .A1(n8083), .A2(n5962), .ZN(n4873) );
  NAND2_X1 U5409 ( .A1(n5966), .A2(n8288), .ZN(n4854) );
  AND2_X1 U5410 ( .A1(n8654), .A2(n6001), .ZN(n4904) );
  NAND2_X1 U5411 ( .A1(n4866), .A2(n4865), .ZN(n4869) );
  AND2_X1 U5412 ( .A1(n4867), .A2(n4538), .ZN(n4865) );
  NOR2_X1 U5413 ( .A1(n5125), .A2(n5122), .ZN(n5121) );
  AND2_X1 U5414 ( .A1(n4714), .A2(n4713), .ZN(n4712) );
  INV_X1 U5415 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n4713) );
  AND2_X1 U5416 ( .A1(n5566), .A2(n4703), .ZN(n4702) );
  INV_X1 U5417 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4703) );
  INV_X1 U5418 ( .A(n5586), .ZN(n5567) );
  AND2_X1 U5419 ( .A1(n4828), .A2(n4470), .ZN(n4825) );
  INV_X1 U5420 ( .A(n4819), .ZN(n4817) );
  AND2_X1 U5421 ( .A1(n9040), .A2(n8493), .ZN(n6215) );
  AND2_X1 U5422 ( .A1(n4477), .A2(n4809), .ZN(n4808) );
  INV_X1 U5423 ( .A(n4812), .ZN(n4811) );
  OR2_X1 U5424 ( .A1(n9040), .A2(n8493), .ZN(n6243) );
  NOR2_X1 U5425 ( .A1(n5833), .A2(n5119), .ZN(n5118) );
  NOR2_X1 U5426 ( .A1(n6248), .A2(n4832), .ZN(n4831) );
  INV_X1 U5427 ( .A(n5489), .ZN(n4832) );
  INV_X1 U5428 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5203) );
  INV_X1 U5429 ( .A(n4997), .ZN(n4996) );
  OAI21_X1 U5430 ( .B1(n5000), .B2(n4998), .A(n6552), .ZN(n4997) );
  AND2_X1 U5431 ( .A1(n9250), .A2(n6571), .ZN(n6572) );
  NOR4_X1 U5432 ( .A1(n9469), .A2(n9556), .A3(n9878), .A4(n9468), .ZN(n9470)
         );
  AOI21_X1 U5433 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10148), .A(n10140), .ZN(
        n9612) );
  NOR2_X1 U5434 ( .A1(n6935), .A2(n6934), .ZN(n4620) );
  OR2_X1 U5435 ( .A1(n9680), .A2(n9954), .ZN(n9498) );
  INV_X1 U5436 ( .A(n4620), .ZN(n6980) );
  NAND2_X1 U5437 ( .A1(n6911), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6935) );
  INV_X1 U5438 ( .A(n6913), .ZN(n6911) );
  NAND2_X1 U5439 ( .A1(n4624), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6913) );
  OR2_X1 U5440 ( .A1(n9961), .A2(n9953), .ZN(n9486) );
  INV_X1 U5441 ( .A(n9402), .ZN(n4841) );
  NOR2_X1 U5442 ( .A1(n10084), .A2(n10009), .ZN(n5055) );
  OR2_X1 U5443 ( .A1(n10009), .A2(n9822), .ZN(n9411) );
  AND2_X1 U5444 ( .A1(n10048), .A2(n10058), .ZN(n9389) );
  INV_X1 U5445 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5446 ( .B1(n9916), .B2(n4937), .A(n7035), .ZN(n4936) );
  INV_X1 U5447 ( .A(n7034), .ZN(n4937) );
  AND2_X1 U5448 ( .A1(n9373), .A2(n8024), .ZN(n9456) );
  NAND2_X1 U5449 ( .A1(n5161), .A2(n7058), .ZN(n4679) );
  INV_X1 U5450 ( .A(n9526), .ZN(n5162) );
  AND2_X1 U5451 ( .A1(n5022), .A2(n5020), .ZN(n5019) );
  AND2_X1 U5452 ( .A1(n5751), .A2(n5720), .ZN(n5734) );
  AND2_X1 U5453 ( .A1(n5716), .A2(n5701), .ZN(n5715) );
  NAND2_X1 U5454 ( .A1(n5015), .A2(n5012), .ZN(n6361) );
  NOR2_X1 U5455 ( .A1(n4462), .A2(n5013), .ZN(n5012) );
  NAND2_X1 U5456 ( .A1(n6348), .A2(n5014), .ZN(n5013) );
  OR2_X1 U5457 ( .A1(n6553), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U5458 ( .A1(n5354), .A2(SI_6_), .ZN(n5375) );
  NAND2_X1 U5459 ( .A1(n5334), .A2(SI_5_), .ZN(n5352) );
  NAND2_X1 U5460 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  AOI21_X1 U5461 ( .B1(n5091), .B2(n5089), .A(n5088), .ZN(n5087) );
  INV_X1 U5462 ( .A(n8212), .ZN(n5089) );
  INV_X1 U5463 ( .A(n8350), .ZN(n5088) );
  INV_X1 U5464 ( .A(n5091), .ZN(n5090) );
  AOI21_X1 U5465 ( .B1(n5075), .B2(n5073), .A(n4501), .ZN(n5072) );
  INV_X1 U5466 ( .A(n5078), .ZN(n5073) );
  INV_X1 U5467 ( .A(n5075), .ZN(n5074) );
  INV_X1 U5469 ( .A(n10287), .ZN(n7528) );
  OR2_X1 U5470 ( .A1(n7796), .A2(n7795), .ZN(n5068) );
  NOR2_X1 U5471 ( .A1(n6274), .A2(n7838), .ZN(n6275) );
  AND2_X1 U5472 ( .A1(n5631), .A2(n5630), .ZN(n8563) );
  OR2_X1 U5473 ( .A1(n5291), .A2(n4586), .ZN(n5234) );
  AOI21_X1 U5474 ( .B1(n4849), .B2(n5222), .A(n5948), .ZN(n7351) );
  AND2_X1 U5475 ( .A1(n5947), .A2(n5257), .ZN(n4849) );
  XNOR2_X1 U5476 ( .A(n7163), .B(n7624), .ZN(n8616) );
  OR2_X1 U5477 ( .A1(n5842), .A2(n4586), .ZN(n4587) );
  INV_X1 U5478 ( .A(n5946), .ZN(n6014) );
  NAND2_X1 U5479 ( .A1(n4890), .A2(n8614), .ZN(n4893) );
  NOR2_X1 U5480 ( .A1(n7166), .A2(n4891), .ZN(n4890) );
  NAND2_X1 U5481 ( .A1(n5989), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4906) );
  INV_X1 U5482 ( .A(n7562), .ZN(n4864) );
  AOI21_X1 U5483 ( .B1(n7562), .B2(n4863), .A(n4539), .ZN(n4862) );
  OR2_X1 U5484 ( .A1(n5956), .A2(n7168), .ZN(n5957) );
  NAND2_X1 U5485 ( .A1(n7431), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U5486 ( .A1(n5961), .A2(n7967), .ZN(n7970) );
  NOR2_X1 U5487 ( .A1(n7202), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U5488 ( .A1(n4911), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7202), .B2(
        n4910), .ZN(n4909) );
  INV_X1 U5489 ( .A(n8288), .ZN(n4859) );
  INV_X1 U5490 ( .A(n4854), .ZN(n8250) );
  NAND2_X1 U5491 ( .A1(n8250), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U5492 ( .A1(n8256), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U5493 ( .A1(n6000), .A2(n7274), .ZN(n8654) );
  NAND2_X1 U5494 ( .A1(n4848), .A2(n8648), .ZN(n8652) );
  AND2_X1 U5495 ( .A1(n8676), .A2(n4605), .ZN(n4430) );
  NAND2_X1 U5496 ( .A1(n5971), .A2(n7490), .ZN(n4605) );
  OAI21_X1 U5497 ( .B1(n8643), .B2(n8644), .A(n4527), .ZN(n8666) );
  NOR2_X1 U5498 ( .A1(n8716), .A2(n8715), .ZN(n8723) );
  NAND2_X1 U5499 ( .A1(n8738), .A2(n5775), .ZN(n8399) );
  NAND2_X1 U5500 ( .A1(n5706), .A2(n5705), .ZN(n5725) );
  INV_X1 U5501 ( .A(n5707), .ZN(n5706) );
  AOI21_X1 U5502 ( .B1(n8848), .B2(n5799), .A(n5657), .ZN(n8855) );
  AND2_X1 U5503 ( .A1(n5832), .A2(n6176), .ZN(n5110) );
  AND4_X1 U5504 ( .A1(n5456), .A2(n5455), .A3(n5454), .A4(n5453), .ZN(n8473)
         );
  NAND2_X1 U5505 ( .A1(n5368), .A2(n4709), .ZN(n5412) );
  NAND2_X1 U5506 ( .A1(n5368), .A2(n5367), .ZN(n5394) );
  NAND4_X1 U5507 ( .A1(n5293), .A2(n10294), .A3(n4716), .A4(n5312), .ZN(n5369)
         );
  INV_X1 U5508 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4716) );
  AND2_X1 U5509 ( .A1(n6221), .A2(n6222), .ZN(n8766) );
  OAI21_X1 U5510 ( .B1(n8858), .B2(n4498), .A(n5112), .ZN(n5835) );
  AND3_X1 U5511 ( .A1(n4561), .A2(n5113), .A3(n6246), .ZN(n5112) );
  NAND2_X1 U5512 ( .A1(n4813), .A2(n4812), .ZN(n8802) );
  NAND2_X1 U5513 ( .A1(n5639), .A2(n5638), .ZN(n9054) );
  NAND2_X1 U5514 ( .A1(n4589), .A2(n5118), .ZN(n5117) );
  AND2_X1 U5515 ( .A1(n8844), .A2(n8843), .ZN(n8841) );
  AND3_X1 U5516 ( .A1(n5589), .A2(n5588), .A3(n5587), .ZN(n8908) );
  AND3_X1 U5517 ( .A1(n5547), .A2(n5546), .A3(n5545), .ZN(n8893) );
  AOI21_X1 U5518 ( .B1(n5134), .B2(n5130), .A(n4488), .ZN(n5129) );
  NOR2_X1 U5519 ( .A1(n5825), .A2(n5136), .ZN(n5128) );
  INV_X1 U5520 ( .A(n4831), .ZN(n4830) );
  NOR2_X1 U5521 ( .A1(n5490), .A2(n4835), .ZN(n4834) );
  OR2_X1 U5522 ( .A1(n8482), .A2(n8931), .ZN(n5489) );
  AOI21_X1 U5523 ( .B1(n4431), .B2(n5189), .A(n4441), .ZN(n4798) );
  NAND2_X1 U5524 ( .A1(n4503), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U5525 ( .A1(n4464), .A2(n4431), .ZN(n4796) );
  OAI21_X1 U5526 ( .B1(n5401), .B2(n4803), .A(n4801), .ZN(n4800) );
  NAND2_X1 U5527 ( .A1(n8179), .A2(n7385), .ZN(n10330) );
  NAND4_X1 U5528 ( .A1(n5140), .A2(n5139), .A3(n5182), .A4(n5137), .ZN(n5226)
         );
  NAND2_X1 U5529 ( .A1(n4836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5228) );
  CLKBUF_X1 U5530 ( .A(n5258), .Z(n5259) );
  INV_X1 U5531 ( .A(n6594), .ZN(n4593) );
  NAND2_X1 U5532 ( .A1(n4621), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6632) );
  INV_X1 U5533 ( .A(n6609), .ZN(n4621) );
  XNOR2_X1 U5534 ( .A(n6909), .B(n8316), .ZN(n6927) );
  INV_X1 U5535 ( .A(n6741), .ZN(n4990) );
  NAND2_X1 U5536 ( .A1(n4983), .A2(n4987), .ZN(n4982) );
  NAND2_X1 U5537 ( .A1(n7511), .A2(n7510), .ZN(n6445) );
  AOI21_X1 U5538 ( .B1(n6400), .B2(n4422), .A(n6401), .ZN(n6403) );
  XNOR2_X1 U5539 ( .A(n4542), .B(n6399), .ZN(n6402) );
  NAND2_X1 U5540 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  AND2_X1 U5541 ( .A1(n10067), .A2(n9509), .ZN(n9567) );
  NOR2_X1 U5542 ( .A1(n5048), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7447) );
  OAI21_X1 U5543 ( .B1(n7221), .B2(P1_REG2_REG_2__SCAN_IN), .A(n4959), .ZN(
        n7453) );
  NAND2_X1 U5544 ( .A1(n7221), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4959) );
  OAI21_X1 U5545 ( .B1(n7221), .B2(P1_REG1_REG_2__SCAN_IN), .A(n7220), .ZN(
        n7457) );
  NAND2_X1 U5546 ( .A1(n7221), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U5547 ( .A1(n7264), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4965) );
  OR2_X1 U5548 ( .A1(n7246), .A2(n4504), .ZN(n4961) );
  AND2_X1 U5549 ( .A1(n7541), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4974) );
  NOR2_X1 U5550 ( .A1(n8088), .A2(n8087), .ZN(n8089) );
  NAND2_X1 U5551 ( .A1(n8089), .A2(n8090), .ZN(n9610) );
  OR2_X1 U5552 ( .A1(n10132), .A2(n10133), .ZN(n4968) );
  OR2_X1 U5553 ( .A1(n10144), .A2(n4750), .ZN(n4748) );
  OR2_X1 U5554 ( .A1(n10129), .A2(n4749), .ZN(n4747) );
  OR2_X1 U5555 ( .A1(n10144), .A2(n10130), .ZN(n4749) );
  OR2_X1 U5556 ( .A1(n10157), .A2(n4972), .ZN(n4970) );
  OR2_X1 U5557 ( .A1(n10166), .A2(n6701), .ZN(n4972) );
  OR2_X1 U5558 ( .A1(n4452), .A2(n10166), .ZN(n4971) );
  OR2_X1 U5559 ( .A1(n10157), .A2(n6701), .ZN(n4973) );
  NOR2_X1 U5560 ( .A1(n10190), .A2(n9614), .ZN(n4976) );
  NAND2_X1 U5561 ( .A1(n4620), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9653) );
  NOR2_X1 U5562 ( .A1(n7071), .A2(n5158), .ZN(n5157) );
  NAND2_X1 U5563 ( .A1(n5156), .A2(n9426), .ZN(n5155) );
  NOR2_X1 U5564 ( .A1(n4946), .A2(n4945), .ZN(n4944) );
  INV_X1 U5565 ( .A(n7051), .ZN(n4945) );
  INV_X1 U5566 ( .A(n4947), .ZN(n4946) );
  NAND2_X1 U5567 ( .A1(n4947), .A2(n4484), .ZN(n4943) );
  NAND2_X1 U5568 ( .A1(n9712), .A2(n10212), .ZN(n4629) );
  AND2_X1 U5569 ( .A1(n9736), .A2(n9480), .ZN(n5170) );
  INV_X1 U5570 ( .A(n9736), .ZN(n9721) );
  NAND2_X1 U5571 ( .A1(n7069), .A2(n9480), .ZN(n9722) );
  OAI21_X1 U5572 ( .B1(n4580), .B2(n4693), .A(n4691), .ZN(n7069) );
  AND2_X1 U5573 ( .A1(n6885), .A2(n6884), .ZN(n9750) );
  AOI21_X2 U5574 ( .B1(n4839), .B2(n4841), .A(n4838), .ZN(n4837) );
  INV_X1 U5575 ( .A(n9419), .ZN(n4838) );
  AOI21_X1 U5576 ( .B1(n4928), .B2(n4926), .A(n4491), .ZN(n4925) );
  INV_X1 U5577 ( .A(n4458), .ZN(n4926) );
  OR2_X1 U5578 ( .A1(n10001), .A2(n9779), .ZN(n4932) );
  AND2_X1 U5579 ( .A1(n6830), .A2(n6829), .ZN(n9792) );
  OR2_X1 U5580 ( .A1(n9777), .A2(n6465), .ZN(n6830) );
  NAND2_X1 U5582 ( .A1(n4625), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6804) );
  AND2_X1 U5583 ( .A1(n9847), .A2(n9831), .ZN(n9826) );
  OR2_X1 U5584 ( .A1(n10084), .A2(n9842), .ZN(n4956) );
  AND2_X1 U5585 ( .A1(n9411), .A2(n9561), .ZN(n9806) );
  NOR2_X1 U5586 ( .A1(n7043), .A2(n4958), .ZN(n4957) );
  INV_X1 U5587 ( .A(n7041), .ZN(n4958) );
  NOR2_X1 U5588 ( .A1(n9878), .A2(n4686), .ZN(n4685) );
  INV_X1 U5589 ( .A(n7065), .ZN(n4686) );
  NAND2_X1 U5590 ( .A1(n9901), .A2(n9550), .ZN(n7066) );
  NAND2_X1 U5591 ( .A1(n9393), .A2(n9391), .ZN(n9878) );
  NAND2_X1 U5592 ( .A1(n8118), .A2(n7033), .ZN(n9917) );
  AND2_X1 U5593 ( .A1(n6689), .A2(n6688), .ZN(n9912) );
  OR2_X1 U5594 ( .A1(n7027), .A2(n9203), .ZN(n9366) );
  NAND2_X1 U5595 ( .A1(n9157), .A2(n7028), .ZN(n8024) );
  NAND2_X1 U5596 ( .A1(n9366), .A2(n9376), .ZN(n9461) );
  INV_X1 U5597 ( .A(n9456), .ZN(n7987) );
  NAND2_X1 U5598 ( .A1(n7602), .A2(n7056), .ZN(n7743) );
  NAND2_X1 U5599 ( .A1(n9117), .A2(n7103), .ZN(n4591) );
  AND2_X1 U5600 ( .A1(n4469), .A2(n9716), .ZN(n9962) );
  AND2_X1 U5601 ( .A1(n6811), .A2(n6810), .ZN(n9992) );
  AND2_X1 U5602 ( .A1(n7184), .A2(n7448), .ZN(n10053) );
  AND2_X1 U5603 ( .A1(n7594), .A2(n7092), .ZN(n7112) );
  AND2_X1 U5604 ( .A1(n7993), .A2(n8177), .ZN(n5181) );
  AND3_X2 U5605 ( .A1(n6346), .A2(n6313), .A3(n5039), .ZN(n4681) );
  INV_X1 U5606 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6315) );
  XNOR2_X1 U5607 ( .A(n5770), .B(n5769), .ZN(n9113) );
  XNOR2_X1 U5608 ( .A(n5735), .B(n5734), .ZN(n9120) );
  INV_X1 U5609 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6370) );
  OAI21_X1 U5610 ( .B1(n5532), .B2(n4724), .A(n4721), .ZN(n5613) );
  NAND2_X1 U5611 ( .A1(n4726), .A2(n5041), .ZN(n5596) );
  NAND2_X1 U5612 ( .A1(n5532), .A2(n5044), .ZN(n4726) );
  NAND2_X1 U5613 ( .A1(n5471), .A2(n5468), .ZN(n5462) );
  NOR2_X1 U5614 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  XNOR2_X1 U5615 ( .A(n5462), .B(n5461), .ZN(n7231) );
  OAI21_X1 U5616 ( .B1(n5431), .B2(SI_10_), .A(n5468), .ZN(n5433) );
  AND2_X1 U5617 ( .A1(n5420), .A2(n5380), .ZN(n5381) );
  NOR2_X1 U5618 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6308) );
  NAND2_X1 U5619 ( .A1(n6414), .A2(n6413), .ZN(n6432) );
  NAND2_X1 U5620 ( .A1(n6412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U5621 ( .A1(n4575), .A2(n8411), .ZN(n8414) );
  NAND2_X1 U5622 ( .A1(n8572), .A2(n4576), .ZN(n4575) );
  INV_X1 U5623 ( .A(n8412), .ZN(n4576) );
  NAND2_X1 U5624 ( .A1(n5081), .A2(n5080), .ZN(n8413) );
  AOI21_X1 U5625 ( .B1(n5082), .B2(n5084), .A(n4486), .ZN(n5080) );
  INV_X1 U5626 ( .A(n7572), .ZN(n5067) );
  AOI21_X1 U5627 ( .B1(n8837), .B2(n5799), .A(n5645), .ZN(n8816) );
  NAND2_X1 U5628 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  NAND2_X1 U5629 ( .A1(n8489), .A2(n8389), .ZN(n8573) );
  NAND2_X1 U5630 ( .A1(n5692), .A2(n5691), .ZN(n8788) );
  NAND2_X1 U5631 ( .A1(n5675), .A2(n5674), .ZN(n8834) );
  INV_X1 U5632 ( .A(n8473), .ZN(n8603) );
  NAND2_X1 U5633 ( .A1(n8620), .A2(n4782), .ZN(n7331) );
  OR2_X1 U5634 ( .A1(n6016), .A2(n8619), .ZN(n4782) );
  NOR2_X1 U5635 ( .A1(n7331), .A2(n7332), .ZN(n7330) );
  OR2_X1 U5636 ( .A1(n6020), .A2(n6021), .ZN(n4788) );
  AOI21_X1 U5637 ( .B1(n7179), .B2(n6025), .A(n7551), .ZN(n7757) );
  AND2_X1 U5638 ( .A1(n4786), .A2(n4785), .ZN(n8189) );
  NAND2_X1 U5639 ( .A1(n6031), .A2(n8083), .ZN(n4785) );
  OAI22_X1 U5640 ( .A1(n8189), .A2(n8190), .B1(n6032), .B2(n7197), .ZN(n8248)
         );
  OAI21_X1 U5641 ( .B1(n8735), .B2(n8734), .A(n4572), .ZN(n4571) );
  AND2_X1 U5642 ( .A1(n8733), .A2(n4573), .ZN(n4572) );
  INV_X1 U5643 ( .A(n8725), .ZN(n4573) );
  AND2_X1 U5644 ( .A1(n8757), .A2(n10284), .ZN(n8956) );
  NAND2_X1 U5645 ( .A1(n5742), .A2(n5741), .ZN(n9028) );
  NAND2_X1 U5646 ( .A1(n9117), .A2(n6106), .ZN(n5742) );
  NAND2_X1 U5647 ( .A1(n5624), .A2(n5623), .ZN(n8987) );
  INV_X1 U5648 ( .A(n8744), .ZN(n10292) );
  INV_X1 U5649 ( .A(n8912), .ZN(n10293) );
  NAND2_X1 U5650 ( .A1(n8409), .A2(n6106), .ZN(n5773) );
  INV_X1 U5651 ( .A(n5805), .ZN(n8745) );
  NAND2_X1 U5652 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  NAND2_X1 U5653 ( .A1(n8600), .A2(n10284), .ZN(n5920) );
  NAND2_X1 U5654 ( .A1(n8751), .A2(n6226), .ZN(n5923) );
  XNOR2_X1 U5655 ( .A(n8765), .B(n8766), .ZN(n9031) );
  INV_X1 U5656 ( .A(n9101), .ZN(n9093) );
  OR2_X1 U5657 ( .A1(n7400), .A2(n5906), .ZN(n5913) );
  AND3_X1 U5658 ( .A1(n6709), .A2(n6708), .A3(n6707), .ZN(n10039) );
  INV_X1 U5659 ( .A(n7027), .ZN(n9308) );
  AND2_X1 U5660 ( .A1(n6991), .A2(n6989), .ZN(n9326) );
  AND3_X1 U5661 ( .A1(n6730), .A2(n6729), .A3(n6728), .ZN(n9881) );
  INV_X1 U5662 ( .A(n9320), .ZN(n9340) );
  INV_X1 U5663 ( .A(n9946), .ZN(n9712) );
  INV_X1 U5664 ( .A(n9750), .ZN(n9974) );
  INV_X1 U5665 ( .A(n9769), .ZN(n9983) );
  NAND2_X1 U5666 ( .A1(n6860), .A2(n6859), .ZN(n9973) );
  INV_X1 U5667 ( .A(n9233), .ZN(n9842) );
  INV_X1 U5668 ( .A(n9203), .ZN(n10054) );
  AND2_X1 U5669 ( .A1(n4961), .A2(n4960), .ZN(n7292) );
  NOR2_X1 U5670 ( .A1(n4963), .A2(n4964), .ZN(n4960) );
  AND2_X1 U5671 ( .A1(n7290), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4964) );
  NOR2_X1 U5672 ( .A1(n7540), .A2(n4745), .ZN(n7542) );
  AND2_X1 U5673 ( .A1(n7541), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4745) );
  OR2_X1 U5674 ( .A1(n9632), .A2(n10164), .ZN(n9633) );
  INV_X1 U5675 ( .A(n9629), .ZN(n9635) );
  NAND2_X1 U5676 ( .A1(n7135), .A2(n4949), .ZN(n4948) );
  INV_X1 U5677 ( .A(n9649), .ZN(n4949) );
  NAND2_X1 U5678 ( .A1(n5147), .A2(n9651), .ZN(n5146) );
  OAI21_X1 U5679 ( .B1(n9651), .B2(n5149), .A(n5142), .ZN(n5141) );
  NAND2_X1 U5680 ( .A1(n8409), .A2(n7103), .ZN(n7054) );
  NAND2_X1 U5681 ( .A1(n7042), .A2(n7041), .ZN(n9818) );
  AND2_X1 U5682 ( .A1(n9893), .A2(n7650), .ZN(n9928) );
  NAND2_X1 U5683 ( .A1(n5194), .A2(n4409), .ZN(n5165) );
  INV_X1 U5684 ( .A(n9675), .ZN(n7132) );
  NAND2_X1 U5685 ( .A1(n9959), .A2(n10063), .ZN(n4696) );
  NOR2_X1 U5686 ( .A1(n10243), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5035) );
  NOR2_X1 U5687 ( .A1(n9640), .A2(n10002), .ZN(n5030) );
  OAI21_X1 U5688 ( .B1(n9643), .B2(n9945), .A(n10067), .ZN(n5032) );
  NAND2_X1 U5689 ( .A1(n9445), .A2(n5034), .ZN(n5033) );
  NAND2_X1 U5690 ( .A1(n7135), .A2(n7134), .ZN(n7136) );
  NOR2_X1 U5691 ( .A1(n9659), .A2(n10090), .ZN(n7140) );
  INV_X1 U5692 ( .A(n4619), .ZN(n4618) );
  AOI21_X1 U5693 ( .B1(n9988), .B2(n4729), .A(n4595), .ZN(n10071) );
  INV_X1 U5694 ( .A(n9951), .ZN(n4729) );
  NAND2_X1 U5695 ( .A1(n4596), .A2(n4478), .ZN(n4595) );
  NAND2_X1 U5696 ( .A1(n9952), .A2(n9988), .ZN(n4697) );
  NAND2_X1 U5697 ( .A1(n9957), .A2(n9958), .ZN(n4699) );
  OAI21_X1 U5698 ( .B1(n6144), .B2(n6131), .A(n4614), .ZN(n4613) );
  AND2_X1 U5699 ( .A1(n6150), .A2(n8130), .ZN(n4551) );
  MUX2_X1 U5700 ( .A(n6138), .B(n6137), .S(n6241), .Z(n6152) );
  NOR2_X1 U5701 ( .A1(n4772), .A2(n6169), .ZN(n4771) );
  NAND2_X1 U5702 ( .A1(n4645), .A2(n4641), .ZN(n9375) );
  OAI22_X1 U5703 ( .A1(n9349), .A2(n4639), .B1(n4638), .B2(n4485), .ZN(n4641)
         );
  OAI21_X1 U5704 ( .B1(n9363), .B2(n4647), .A(n4642), .ZN(n4645) );
  AOI21_X1 U5705 ( .B1(n6186), .B2(n4604), .A(n4500), .ZN(n4603) );
  AND2_X1 U5706 ( .A1(n9463), .A2(n9342), .ZN(n4675) );
  AND2_X1 U5707 ( .A1(n4471), .A2(n9840), .ZN(n4672) );
  INV_X1 U5708 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U5709 ( .A1(n4658), .A2(n9423), .ZN(n4657) );
  NOR2_X1 U5710 ( .A1(n9425), .A2(n4665), .ZN(n4658) );
  AND2_X1 U5711 ( .A1(n4664), .A2(n4662), .ZN(n4656) );
  NOR2_X1 U5712 ( .A1(n9425), .A2(n4663), .ZN(n4662) );
  INV_X1 U5713 ( .A(n4665), .ZN(n4664) );
  OAI21_X1 U5714 ( .B1(n4667), .B2(n4666), .A(n9412), .ZN(n9414) );
  OAI21_X1 U5715 ( .B1(n4758), .B2(n4761), .A(n4759), .ZN(n4757) );
  AOI21_X1 U5716 ( .B1(n6211), .B2(n4821), .A(n4760), .ZN(n4759) );
  INV_X1 U5717 ( .A(n6218), .ZN(n6219) );
  INV_X1 U5718 ( .A(n5967), .ZN(n4856) );
  AND2_X1 U5719 ( .A1(n5967), .A2(n4858), .ZN(n4853) );
  XNOR2_X1 U5720 ( .A(n4623), .B(n9342), .ZN(n9429) );
  AND2_X1 U5721 ( .A1(n9456), .A2(n4499), .ZN(n4607) );
  INV_X1 U5722 ( .A(n4956), .ZN(n4954) );
  INV_X1 U5723 ( .A(n5016), .ZN(n7074) );
  AOI21_X1 U5724 ( .B1(n5024), .B2(n5027), .A(n5023), .ZN(n5022) );
  INV_X1 U5725 ( .A(n5715), .ZN(n5023) );
  NAND2_X1 U5726 ( .A1(n5024), .A2(n5678), .ZN(n5020) );
  INV_X1 U5727 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U5728 ( .A1(n5615), .A2(n5614), .ZN(n5632) );
  NAND2_X1 U5729 ( .A1(n5557), .A2(n5556), .ZN(n5594) );
  INV_X1 U5730 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4701) );
  INV_X1 U5731 ( .A(n5403), .ZN(n5421) );
  INV_X1 U5732 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5213) );
  INV_X1 U5733 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5211) );
  AND2_X1 U5734 ( .A1(n6238), .A2(n6237), .ZN(n5172) );
  NOR2_X1 U5735 ( .A1(n5257), .A2(n6012), .ZN(n5948) );
  NOR2_X1 U5736 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5202) );
  OR2_X1 U5737 ( .A1(n5991), .A2(n7763), .ZN(n4914) );
  INV_X1 U5738 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5407) );
  INV_X1 U5739 ( .A(n4457), .ZN(n4911) );
  INV_X1 U5740 ( .A(n5993), .ZN(n4910) );
  NAND2_X1 U5741 ( .A1(n4903), .A2(n6001), .ZN(n4902) );
  AOI21_X1 U5742 ( .B1(n6003), .B2(n4886), .A(n4534), .ZN(n4885) );
  NOR2_X1 U5743 ( .A1(n6049), .A2(n6048), .ZN(n8716) );
  INV_X1 U5744 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n4706) );
  AND2_X1 U5745 ( .A1(n5723), .A2(n4708), .ZN(n4707) );
  INV_X1 U5746 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4708) );
  INV_X1 U5747 ( .A(n5725), .ZN(n5724) );
  AND2_X1 U5748 ( .A1(n5640), .A2(n10592), .ZN(n4714) );
  NAND2_X1 U5749 ( .A1(n5567), .A2(n4702), .ZN(n5625) );
  AND2_X1 U5750 ( .A1(n5367), .A2(n4710), .ZN(n4709) );
  INV_X1 U5751 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4710) );
  INV_X1 U5752 ( .A(n5369), .ZN(n5368) );
  INV_X1 U5753 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5312) );
  INV_X1 U5754 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U5755 ( .A1(n10294), .A2(n5293), .ZN(n5313) );
  INV_X1 U5756 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U5757 ( .A1(n9034), .A2(n8578), .ZN(n6218) );
  INV_X1 U5758 ( .A(n5118), .ZN(n5114) );
  AND2_X1 U5759 ( .A1(n4562), .A2(n8799), .ZN(n4561) );
  OR2_X1 U5760 ( .A1(n6204), .A2(n8797), .ZN(n4562) );
  NAND2_X1 U5761 ( .A1(n5117), .A2(n4410), .ZN(n8798) );
  INV_X1 U5762 ( .A(n6172), .ZN(n5132) );
  AND2_X1 U5763 ( .A1(n6156), .A2(n8345), .ZN(n5126) );
  NAND2_X1 U5764 ( .A1(n5105), .A2(n4481), .ZN(n10259) );
  AOI21_X1 U5765 ( .B1(n5858), .B2(P2_IR_REG_31__SCAN_IN), .A(n5098), .ZN(
        n5097) );
  NAND2_X1 U5766 ( .A1(n5099), .A2(n5866), .ZN(n5098) );
  NAND2_X1 U5767 ( .A1(n5096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  NOR3_X1 U5768 ( .A1(n5095), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5094) );
  INV_X1 U5769 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5198) );
  OR2_X1 U5770 ( .A1(n5350), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5384) );
  INV_X1 U5771 ( .A(n6674), .ZN(n4989) );
  AOI21_X1 U5772 ( .B1(n5006), .B2(n5007), .A(n5005), .ZN(n5004) );
  INV_X1 U5773 ( .A(n9187), .ZN(n5005) );
  INV_X1 U5774 ( .A(n5010), .ZN(n5006) );
  NOR2_X1 U5775 ( .A1(n6660), .A2(n6659), .ZN(n6681) );
  NAND2_X1 U5776 ( .A1(n5154), .A2(n5155), .ZN(n5153) );
  INV_X1 U5777 ( .A(n9475), .ZN(n5154) );
  NAND2_X1 U5778 ( .A1(n10072), .A2(n5060), .ZN(n5059) );
  INV_X1 U5779 ( .A(n4624), .ZN(n6899) );
  INV_X1 U5780 ( .A(n4839), .ZN(n4687) );
  INV_X1 U5781 ( .A(n4837), .ZN(n4693) );
  INV_X1 U5782 ( .A(n9389), .ZN(n9543) );
  AND2_X1 U5783 ( .A1(n9592), .A2(n7811), .ZN(n7820) );
  AND2_X1 U5784 ( .A1(n10231), .A2(n7637), .ZN(n5052) );
  NAND2_X1 U5785 ( .A1(n7098), .A2(n7103), .ZN(n7100) );
  NAND2_X1 U5786 ( .A1(n7074), .A2(n7073), .ZN(n7739) );
  INV_X1 U5787 ( .A(n5752), .ZN(n5753) );
  AND2_X1 U5788 ( .A1(n5787), .A2(n5758), .ZN(n5769) );
  INV_X1 U5789 ( .A(n5695), .ZN(n5027) );
  AOI21_X1 U5790 ( .B1(n5695), .B2(n5026), .A(n5025), .ZN(n5024) );
  INV_X1 U5791 ( .A(n5697), .ZN(n5025) );
  INV_X1 U5792 ( .A(n5677), .ZN(n5026) );
  INV_X1 U5793 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U5794 ( .A1(n5532), .A2(n4468), .ZN(n4720) );
  NAND2_X1 U5795 ( .A1(n5044), .A2(n5046), .ZN(n5042) );
  OR2_X1 U5796 ( .A1(n5432), .A2(n5038), .ZN(n5037) );
  NAND2_X1 U5797 ( .A1(n5431), .A2(SI_10_), .ZN(n5468) );
  NAND2_X1 U5798 ( .A1(n5403), .A2(n5402), .ZN(n5422) );
  INV_X1 U5799 ( .A(SI_8_), .ZN(n5402) );
  NAND2_X1 U5800 ( .A1(n5277), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5278) );
  OAI211_X1 U5801 ( .C1(n5277), .C2(P1_DATAO_REG_0__SCAN_IN), .A(n5216), .B(
        SI_0_), .ZN(n5217) );
  INV_X1 U5802 ( .A(n8389), .ZN(n5084) );
  AND2_X1 U5803 ( .A1(n8378), .A2(n8376), .ZN(n8457) );
  OR2_X1 U5804 ( .A1(n8377), .A2(n8456), .ZN(n8460) );
  OR2_X1 U5805 ( .A1(n8524), .A2(n8377), .ZN(n8459) );
  INV_X1 U5806 ( .A(n8834), .ZN(n8465) );
  AND2_X1 U5807 ( .A1(n8389), .A2(n8387), .ZN(n8487) );
  AND2_X1 U5808 ( .A1(n8214), .A2(n8211), .ZN(n8212) );
  NOR2_X1 U5809 ( .A1(n8372), .A2(n5079), .ZN(n5078) );
  INV_X1 U5810 ( .A(n8369), .ZN(n5079) );
  NAND2_X1 U5811 ( .A1(n8342), .A2(n8341), .ZN(n8470) );
  NOR2_X1 U5812 ( .A1(n4778), .A2(n4617), .ZN(n4616) );
  INV_X1 U5813 ( .A(n6231), .ZN(n4617) );
  NAND2_X1 U5814 ( .A1(n4779), .A2(n6233), .ZN(n4778) );
  AND2_X1 U5815 ( .A1(n6239), .A2(n6237), .ZN(n4568) );
  OAI21_X1 U5816 ( .B1(n6010), .B2(P2_REG1_REG_0__SCAN_IN), .A(n4574), .ZN(
        n7298) );
  NAND2_X1 U5817 ( .A1(n6010), .A2(n5109), .ZN(n4574) );
  AOI21_X1 U5818 ( .B1(n6014), .B2(n5979), .A(n5980), .ZN(n7353) );
  NAND2_X1 U5819 ( .A1(n4887), .A2(n7166), .ZN(n7308) );
  NAND2_X1 U5820 ( .A1(n8614), .A2(n5982), .ZN(n4887) );
  AOI21_X1 U5821 ( .B1(n7166), .B2(n4891), .A(n4889), .ZN(n4888) );
  NAND2_X1 U5822 ( .A1(n5954), .A2(n7316), .ZN(n7320) );
  NAND2_X1 U5823 ( .A1(n4905), .A2(n7557), .ZN(n7559) );
  INV_X1 U5824 ( .A(n4906), .ZN(n4905) );
  AND2_X1 U5825 ( .A1(n4914), .A2(n7957), .ZN(n7759) );
  NAND2_X1 U5826 ( .A1(n5991), .A2(n7763), .ZN(n7957) );
  NAND2_X1 U5827 ( .A1(n7970), .A2(n4434), .ZN(n4878) );
  NAND2_X1 U5828 ( .A1(n7961), .A2(n4457), .ZN(n4913) );
  OAI21_X1 U5829 ( .B1(n7970), .B2(n4875), .A(n4872), .ZN(n5963) );
  NOR2_X1 U5830 ( .A1(n7202), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4875) );
  NOR2_X1 U5831 ( .A1(n4874), .A2(n4873), .ZN(n4872) );
  NAND2_X1 U5832 ( .A1(n7970), .A2(n5962), .ZN(n4871) );
  OR2_X1 U5833 ( .A1(n4877), .A2(n4876), .ZN(n8195) );
  NAND2_X1 U5834 ( .A1(n4878), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4877) );
  INV_X1 U5835 ( .A(n8193), .ZN(n4876) );
  NAND2_X1 U5836 ( .A1(n7961), .A2(n5993), .ZN(n4908) );
  INV_X1 U5837 ( .A(n8297), .ZN(n4897) );
  OR2_X1 U5838 ( .A1(n5996), .A2(n8251), .ZN(n5997) );
  AND2_X1 U5839 ( .A1(n8649), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4847) );
  AND2_X1 U5840 ( .A1(n6042), .A2(n7490), .ZN(n4784) );
  NAND2_X1 U5841 ( .A1(n4430), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U5842 ( .A1(n4430), .A2(n4532), .ZN(n4866) );
  OAI211_X1 U5843 ( .C1(n8689), .C2(n8688), .A(n4885), .B(n6047), .ZN(n4881)
         );
  NOR2_X1 U5844 ( .A1(n6047), .A2(n8688), .ZN(n4879) );
  OR2_X1 U5845 ( .A1(n4885), .A2(n6047), .ZN(n4882) );
  AOI21_X1 U5846 ( .B1(n8395), .B2(n5124), .A(n4494), .ZN(n5123) );
  INV_X1 U5847 ( .A(n6226), .ZN(n5124) );
  OR2_X1 U5848 ( .A1(n5774), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U5849 ( .A1(n5641), .A2(n4712), .ZN(n5686) );
  NAND2_X1 U5850 ( .A1(n5641), .A2(n4533), .ZN(n5707) );
  INV_X1 U5851 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U5852 ( .A1(n5641), .A2(n4714), .ZN(n5669) );
  NAND2_X1 U5853 ( .A1(n5567), .A2(n4526), .ZN(n5653) );
  NAND2_X1 U5854 ( .A1(n5593), .A2(n5592), .ZN(n8864) );
  OAI21_X1 U5855 ( .B1(n8881), .B2(n8880), .A(n5590), .ZN(n5591) );
  NAND2_X1 U5856 ( .A1(n5567), .A2(n5566), .ZN(n5602) );
  NAND2_X1 U5857 ( .A1(n5542), .A2(n5541), .ZN(n5584) );
  INV_X1 U5858 ( .A(n5543), .ZN(n5542) );
  AND2_X1 U5859 ( .A1(n4827), .A2(n5530), .ZN(n4826) );
  NAND2_X1 U5860 ( .A1(n5508), .A2(n5507), .ZN(n5524) );
  INV_X1 U5861 ( .A(n5509), .ZN(n5508) );
  OR2_X1 U5862 ( .A1(n5524), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5543) );
  INV_X1 U5863 ( .A(n8920), .ZN(n8477) );
  OAI21_X1 U5864 ( .B1(n8270), .B2(n8345), .A(n6156), .ZN(n7151) );
  OR2_X1 U5865 ( .A1(n5451), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U5866 ( .A1(n5482), .A2(n10485), .ZN(n5509) );
  INV_X1 U5867 ( .A(n5483), .ZN(n5482) );
  OR2_X1 U5868 ( .A1(n5439), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5451) );
  AND2_X1 U5869 ( .A1(n6150), .A2(n7940), .ZN(n10258) );
  AND4_X1 U5870 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n10255)
         );
  AND3_X1 U5871 ( .A1(n7419), .A2(n5840), .A3(n10330), .ZN(n7902) );
  NAND2_X1 U5872 ( .A1(n7407), .A2(n7392), .ZN(n7713) );
  AND2_X1 U5873 ( .A1(n8737), .A2(n8736), .ZN(n9019) );
  NAND2_X1 U5874 ( .A1(n8768), .A2(n10286), .ZN(n5919) );
  AOI21_X1 U5875 ( .B1(n4816), .B2(n4822), .A(n4496), .ZN(n4814) );
  NOR2_X1 U5876 ( .A1(n4817), .A2(n8753), .ZN(n4816) );
  OR2_X1 U5877 ( .A1(n8762), .A2(n8401), .ZN(n6226) );
  NOR2_X1 U5878 ( .A1(n4811), .A2(n4806), .ZN(n4805) );
  AND2_X1 U5879 ( .A1(n6244), .A2(n6243), .ZN(n8786) );
  AND2_X1 U5880 ( .A1(n4813), .A2(n4442), .ZN(n8844) );
  INV_X1 U5881 ( .A(n8878), .ZN(n8881) );
  NAND2_X1 U5882 ( .A1(n5523), .A2(n5522), .ZN(n9086) );
  INV_X1 U5883 ( .A(n7937), .ZN(n10324) );
  AND2_X1 U5884 ( .A1(n8179), .A2(n7384), .ZN(n10317) );
  OAI21_X1 U5885 ( .B1(n5858), .B2(n5857), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5865) );
  MUX2_X1 U5886 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5221), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5222) );
  NOR2_X1 U5887 ( .A1(n10118), .A2(n8310), .ZN(n6343) );
  OR2_X1 U5888 ( .A1(n6867), .A2(n9241), .ZN(n9141) );
  NAND2_X1 U5889 ( .A1(n9595), .A2(n8313), .ZN(n6439) );
  NAND2_X1 U5890 ( .A1(n7866), .A2(n5000), .ZN(n4995) );
  NOR2_X1 U5891 ( .A1(n9265), .A2(n5011), .ZN(n5010) );
  INV_X1 U5892 ( .A(n6800), .ZN(n5011) );
  INV_X1 U5893 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10500) );
  AND2_X1 U5894 ( .A1(n6649), .A2(n6647), .ZN(n9195) );
  OR2_X1 U5895 ( .A1(n6726), .A2(n6725), .ZN(n6748) );
  AND2_X1 U5896 ( .A1(n6572), .A2(n4993), .ZN(n4992) );
  NAND2_X1 U5897 ( .A1(n4996), .A2(n4998), .ZN(n4993) );
  AND2_X1 U5898 ( .A1(n6817), .A2(n6818), .ZN(n9265) );
  NAND2_X1 U5899 ( .A1(n9277), .A2(n9278), .ZN(n9276) );
  AND2_X1 U5900 ( .A1(n6865), .A2(n6864), .ZN(n9286) );
  AND2_X1 U5901 ( .A1(n9194), .A2(n6624), .ZN(n9296) );
  INV_X1 U5902 ( .A(n6798), .ZN(n9161) );
  AND2_X1 U5903 ( .A1(n6508), .A2(n6509), .ZN(n7806) );
  INV_X1 U5904 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U5905 ( .A1(n4546), .A2(n4545), .ZN(n6929) );
  INV_X1 U5906 ( .A(n9210), .ZN(n4545) );
  INV_X1 U5907 ( .A(n9209), .ZN(n4546) );
  NOR2_X1 U5908 ( .A1(n6927), .A2(n6926), .ZN(n9318) );
  NAND2_X1 U5909 ( .A1(n9221), .A2(n9220), .ZN(n9223) );
  NAND2_X1 U5910 ( .A1(n6681), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U5911 ( .A1(n6703), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6726) );
  INV_X1 U5912 ( .A(n6705), .ZN(n6703) );
  INV_X1 U5913 ( .A(n8177), .ZN(n9521) );
  NOR4_X1 U5914 ( .A1(n9651), .A2(n9475), .A3(n5156), .A4(n9474), .ZN(n9477)
         );
  NOR4_X1 U5915 ( .A1(n4692), .A2(n4663), .A3(n9783), .A4(n9472), .ZN(n9473)
         );
  AND2_X1 U5916 ( .A1(n6789), .A2(n6788), .ZN(n9233) );
  AND2_X1 U5917 ( .A1(n7452), .A2(n7453), .ZN(n7450) );
  AND2_X1 U5918 ( .A1(n7456), .A2(n7457), .ZN(n7454) );
  OR2_X1 U5919 ( .A1(n7224), .A2(n7223), .ZN(n4742) );
  NAND2_X1 U5920 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U5921 ( .A1(n7248), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4741) );
  OR2_X1 U5922 ( .A1(n7246), .A2(n7245), .ZN(n4966) );
  NAND2_X1 U5923 ( .A1(n7533), .A2(n7534), .ZN(n7768) );
  NAND2_X1 U5924 ( .A1(n4565), .A2(n4564), .ZN(n7854) );
  INV_X1 U5925 ( .A(n7771), .ZN(n4564) );
  INV_X1 U5926 ( .A(n7770), .ZN(n4565) );
  OR2_X1 U5927 ( .A1(n10129), .A2(n10130), .ZN(n4751) );
  AND2_X1 U5928 ( .A1(n4968), .A2(n4967), .ZN(n10142) );
  NAND2_X1 U5929 ( .A1(n10136), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4967) );
  NOR2_X1 U5930 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  AND2_X1 U5931 ( .A1(n4747), .A2(n4447), .ZN(n9622) );
  INV_X1 U5932 ( .A(n5150), .ZN(n5149) );
  OAI21_X1 U5933 ( .B1(n5151), .B2(n9475), .A(n9427), .ZN(n5150) );
  NAND2_X1 U5934 ( .A1(n5152), .A2(n5155), .ZN(n5151) );
  INV_X1 U5935 ( .A(n5157), .ZN(n5152) );
  NAND2_X1 U5936 ( .A1(n5149), .A2(n5143), .ZN(n5142) );
  NAND2_X1 U5937 ( .A1(n5153), .A2(n5145), .ZN(n5143) );
  INV_X1 U5938 ( .A(n5153), .ZN(n5147) );
  AOI21_X1 U5939 ( .B1(n4941), .B2(n4940), .A(n4490), .ZN(n4939) );
  AND2_X1 U5940 ( .A1(n6980), .A2(n6936), .ZN(n9681) );
  NAND2_X1 U5941 ( .A1(n6839), .A2(n6838), .ZN(n9752) );
  AOI21_X1 U5942 ( .B1(n4922), .B2(n4924), .A(n4492), .ZN(n4919) );
  INV_X1 U5943 ( .A(n9996), .ZN(n5053) );
  NAND2_X1 U5944 ( .A1(n4438), .A2(n9847), .ZN(n5175) );
  INV_X1 U5945 ( .A(n4625), .ZN(n6784) );
  NAND2_X1 U5946 ( .A1(n9847), .A2(n5055), .ZN(n9810) );
  AND2_X1 U5947 ( .A1(n6770), .A2(n6769), .ZN(n9822) );
  AOI21_X1 U5948 ( .B1(n4935), .B2(n4937), .A(n4489), .ZN(n4933) );
  AND2_X1 U5949 ( .A1(n9463), .A2(n9462), .ZN(n9903) );
  NAND2_X1 U5950 ( .A1(n9917), .A2(n9916), .ZN(n9915) );
  NAND2_X1 U5951 ( .A1(n8001), .A2(n4435), .ZN(n8120) );
  AND2_X1 U5952 ( .A1(n8001), .A2(n4411), .ZN(n8033) );
  NAND2_X1 U5953 ( .A1(n9456), .A2(n8028), .ZN(n7029) );
  AND2_X1 U5954 ( .A1(n9893), .A2(n10053), .ZN(n9898) );
  NAND2_X1 U5955 ( .A1(n5052), .A2(n7738), .ZN(n7666) );
  NAND2_X1 U5956 ( .A1(n5162), .A2(n4679), .ZN(n5159) );
  NAND2_X1 U5957 ( .A1(n7738), .A2(n10231), .ZN(n7630) );
  OAI21_X1 U5958 ( .B1(n7743), .B2(n7057), .A(n9528), .ZN(n7641) );
  INV_X1 U5959 ( .A(n9629), .ZN(n6372) );
  OR2_X1 U5960 ( .A1(n6463), .A2(n6325), .ZN(n6331) );
  INV_X1 U5961 ( .A(n7135), .ZN(n9650) );
  NOR2_X1 U5962 ( .A1(n5145), .A2(n7133), .ZN(n7134) );
  OR2_X1 U5963 ( .A1(n9649), .A2(n10211), .ZN(n7133) );
  OAI21_X1 U5964 ( .B1(n9651), .B2(n7128), .A(n7127), .ZN(n7129) );
  NAND2_X1 U5965 ( .A1(n7489), .A2(n7103), .ZN(n6699) );
  OR2_X1 U5966 ( .A1(n7273), .A2(n6650), .ZN(n6654) );
  NAND2_X1 U5967 ( .A1(n5755), .A2(n5751), .ZN(n5740) );
  INV_X1 U5968 ( .A(n6361), .ZN(n6363) );
  INV_X1 U5969 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6368) );
  NAND3_X1 U5970 ( .A1(n6346), .A2(n6347), .A3(n6475), .ZN(n6742) );
  OR2_X1 U5971 ( .A1(n5574), .A2(SI_15_), .ZN(n5575) );
  AND2_X1 U5972 ( .A1(n5515), .A2(n5496), .ZN(n5497) );
  NAND2_X1 U5973 ( .A1(n5460), .A2(n5459), .ZN(n5472) );
  NAND2_X1 U5974 ( .A1(n5491), .A2(n5465), .ZN(n5474) );
  AND2_X1 U5975 ( .A1(n4952), .A2(n5432), .ZN(n4950) );
  NAND2_X1 U5976 ( .A1(n4951), .A2(n4952), .ZN(n5434) );
  OR2_X1 U5977 ( .A1(n6577), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6578) );
  INV_X1 U5978 ( .A(n5334), .ZN(n5062) );
  NAND2_X1 U5979 ( .A1(n4844), .A2(SI_4_), .ZN(n5328) );
  NAND2_X1 U5980 ( .A1(n5279), .A2(SI_3_), .ZN(n5327) );
  NAND2_X1 U5981 ( .A1(n5253), .A2(n5252), .ZN(n5275) );
  AND4_X1 U5982 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n10257)
         );
  NAND2_X1 U5983 ( .A1(n4579), .A2(n8369), .ZN(n8447) );
  OR2_X1 U5984 ( .A1(n8392), .A2(n8401), .ZN(n8393) );
  AND2_X1 U5985 ( .A1(n5713), .A2(n5712), .ZN(n8493) );
  NAND2_X1 U5986 ( .A1(n8586), .A2(n8361), .ZN(n8499) );
  AND2_X1 U5987 ( .A1(n5183), .A2(n8361), .ZN(n5093) );
  NAND2_X1 U5988 ( .A1(n8213), .A2(n8212), .ZN(n8342) );
  NAND2_X1 U5989 ( .A1(n5077), .A2(n8371), .ZN(n8523) );
  NAND2_X1 U5990 ( .A1(n4579), .A2(n5078), .ZN(n5077) );
  AOI21_X1 U5991 ( .B1(n5087), .B2(n5090), .A(n4493), .ZN(n5085) );
  OAI21_X1 U5992 ( .B1(n4579), .B2(n5074), .A(n5072), .ZN(n8540) );
  AND4_X1 U5993 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n8171)
         );
  NAND2_X1 U5994 ( .A1(n7401), .A2(n8912), .ZN(n8568) );
  INV_X1 U5995 ( .A(n8594), .ZN(n8566) );
  INV_X1 U5996 ( .A(n9028), .ZN(n8583) );
  INV_X1 U5997 ( .A(n8592), .ZN(n8580) );
  INV_X1 U5998 ( .A(n8568), .ZN(n8597) );
  NAND2_X1 U5999 ( .A1(n8585), .A2(n8359), .ZN(n8586) );
  AND2_X1 U6000 ( .A1(n8588), .A2(n8584), .ZN(n8359) );
  INV_X1 U6001 ( .A(n8570), .ZN(n8587) );
  AND2_X1 U6002 ( .A1(n6284), .A2(n4428), .ZN(n4601) );
  AOI21_X1 U6003 ( .B1(n6281), .B2(n6280), .A(n6279), .ZN(n6295) );
  NAND2_X1 U6004 ( .A1(n5749), .A2(n5748), .ZN(n8779) );
  INV_X1 U6005 ( .A(n8563), .ZN(n8866) );
  INV_X1 U6006 ( .A(n8171), .ZN(n8607) );
  INV_X1 U6007 ( .A(n10257), .ZN(n8608) );
  NAND4_X1 U6008 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n10287)
         );
  OR2_X2 U6009 ( .A1(n5237), .A2(n5236), .ZN(n8609) );
  OR2_X1 U6010 ( .A1(n4424), .A2(n6012), .ZN(n5241) );
  OR2_X1 U6011 ( .A1(n6013), .A2(n6014), .ZN(n4783) );
  AND2_X1 U6012 ( .A1(n6018), .A2(n4892), .ZN(n4789) );
  NAND2_X1 U6013 ( .A1(n7428), .A2(n4585), .ZN(n7552) );
  OR2_X1 U6014 ( .A1(n6023), .A2(n5986), .ZN(n4585) );
  NOR2_X1 U6015 ( .A1(n7552), .A2(n7553), .ZN(n7551) );
  NAND2_X1 U6016 ( .A1(n4907), .A2(n7556), .ZN(n7561) );
  OAI21_X1 U6017 ( .B1(n7431), .B2(n4864), .A(n4862), .ZN(n7565) );
  AND2_X1 U6018 ( .A1(n6027), .A2(n6028), .ZN(n4787) );
  NAND2_X1 U6019 ( .A1(n8201), .A2(n4913), .ZN(n8073) );
  OAI21_X1 U6020 ( .B1(n8250), .B2(n4859), .A(n4857), .ZN(n8291) );
  NAND2_X1 U6021 ( .A1(n4901), .A2(n8653), .ZN(n8657) );
  NAND2_X1 U6022 ( .A1(n4866), .A2(n4867), .ZN(n8679) );
  AOI21_X1 U6023 ( .B1(n8694), .B2(n8711), .A(n8710), .ZN(n8713) );
  AND2_X1 U6024 ( .A1(n5704), .A2(n5703), .ZN(n8792) );
  AOI21_X1 U6025 ( .B1(n8832), .B2(n4541), .A(n8814), .ZN(n8815) );
  AND2_X1 U6026 ( .A1(n8820), .A2(n8813), .ZN(n4541) );
  NAND2_X1 U6027 ( .A1(n5831), .A2(n6176), .ZN(n8874) );
  CLKBUF_X1 U6028 ( .A(n8872), .Z(n8873) );
  NAND2_X1 U6029 ( .A1(n5601), .A2(n5600), .ZN(n8871) );
  NAND2_X1 U6030 ( .A1(n7201), .A2(n6106), .ZN(n4762) );
  INV_X1 U6031 ( .A(n10331), .ZN(n10268) );
  INV_X1 U6032 ( .A(n7392), .ZN(n7427) );
  INV_X1 U6033 ( .A(n8956), .ZN(n4612) );
  CLKBUF_X1 U6034 ( .A(n8774), .Z(n8775) );
  INV_X1 U6035 ( .A(n8792), .ZN(n9040) );
  NAND2_X1 U6036 ( .A1(n8245), .A2(n6106), .ZN(n5685) );
  NAND2_X1 U6037 ( .A1(n5117), .A2(n6195), .ZN(n8828) );
  NAND2_X1 U6038 ( .A1(n4589), .A2(n6189), .ZN(n8840) );
  NAND2_X1 U6039 ( .A1(n5565), .A2(n5564), .ZN(n9071) );
  NAND2_X1 U6040 ( .A1(n5133), .A2(n5134), .ZN(n8925) );
  OAI21_X1 U6041 ( .B1(n5458), .B2(n4830), .A(n4828), .ZN(n8919) );
  NAND2_X1 U6042 ( .A1(n4833), .A2(n5489), .ZN(n8930) );
  NAND2_X1 U6043 ( .A1(n5458), .A2(n4834), .ZN(n4833) );
  AND2_X1 U6044 ( .A1(n4802), .A2(n4799), .ZN(n8237) );
  INV_X1 U6045 ( .A(n4800), .ZN(n4799) );
  NAND2_X1 U6046 ( .A1(n8307), .A2(n9119), .ZN(n7237) );
  AND2_X1 U6047 ( .A1(n10387), .A2(n5101), .ZN(n5100) );
  INV_X1 U6048 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5101) );
  NOR2_X1 U6049 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4916) );
  AND2_X1 U6050 ( .A1(n6666), .A2(n6665), .ZN(n10058) );
  NAND2_X1 U6051 ( .A1(n6426), .A2(n6425), .ZN(n7511) );
  NAND2_X1 U6052 ( .A1(n5003), .A2(n5007), .ZN(n9186) );
  NAND2_X1 U6053 ( .A1(n4598), .A2(n5010), .ZN(n5003) );
  AND2_X1 U6054 ( .A1(n6920), .A2(n6919), .ZN(n9946) );
  INV_X1 U6055 ( .A(n6929), .ZN(n9208) );
  INV_X1 U6056 ( .A(n9217), .ZN(n4980) );
  NAND2_X1 U6057 ( .A1(n6445), .A2(n6444), .ZN(n7787) );
  OAI21_X1 U6058 ( .B1(n4598), .B2(n6801), .A(n6800), .ZN(n9268) );
  AND2_X1 U6059 ( .A1(n6638), .A2(n6637), .ZN(n9911) );
  AND2_X1 U6060 ( .A1(n6905), .A2(n6904), .ZN(n9953) );
  OR2_X1 U6061 ( .A1(n9714), .A2(n6465), .ZN(n6905) );
  AND2_X1 U6062 ( .A1(n6991), .A2(n6977), .ZN(n9320) );
  INV_X1 U6063 ( .A(n9440), .ZN(n9444) );
  NAND2_X1 U6064 ( .A1(n9445), .A2(n9446), .ZN(n4648) );
  INV_X1 U6065 ( .A(n9567), .ZN(n9516) );
  INV_X1 U6066 ( .A(n9947), .ZN(n9657) );
  INV_X1 U6067 ( .A(n9954), .ZN(n9669) );
  INV_X1 U6068 ( .A(n9953), .ZN(n9701) );
  INV_X1 U6069 ( .A(n9822), .ZN(n9586) );
  INV_X1 U6070 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7229) );
  NAND2_X1 U6071 ( .A1(n5048), .A2(n10383), .ZN(n10122) );
  INV_X1 U6072 ( .A(n4742), .ZN(n7247) );
  AND2_X1 U6073 ( .A1(n4740), .A2(n4739), .ZN(n7479) );
  INV_X1 U6074 ( .A(n7480), .ZN(n4739) );
  INV_X1 U6075 ( .A(n4740), .ZN(n7481) );
  NOR2_X1 U6076 ( .A1(n7479), .A2(n4738), .ZN(n7253) );
  NOR2_X1 U6077 ( .A1(n7249), .A2(n7250), .ZN(n4738) );
  AND2_X1 U6078 ( .A1(n4966), .A2(n4965), .ZN(n7267) );
  NAND2_X1 U6079 ( .A1(n4961), .A2(n4962), .ZN(n7289) );
  AOI21_X1 U6080 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n7264), .A(n7259), .ZN(
        n7262) );
  NOR2_X1 U6081 ( .A1(n7292), .A2(n7291), .ZN(n7467) );
  NOR2_X1 U6082 ( .A1(n7467), .A2(n4975), .ZN(n7470) );
  AND2_X1 U6083 ( .A1(n7468), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4975) );
  NOR2_X1 U6084 ( .A1(n7470), .A2(n7469), .ZN(n7532) );
  NOR2_X1 U6085 ( .A1(n7466), .A2(n7465), .ZN(n7540) );
  NOR2_X1 U6086 ( .A1(n7464), .A2(n4746), .ZN(n7466) );
  AND2_X1 U6087 ( .A1(n7468), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U6088 ( .A1(n7542), .A2(n7543), .ZN(n7772) );
  NAND2_X1 U6089 ( .A1(n7768), .A2(n4566), .ZN(n7770) );
  OR2_X1 U6090 ( .A1(n7773), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4566) );
  NOR2_X1 U6091 ( .A1(n7860), .A2(n7859), .ZN(n8096) );
  NOR2_X1 U6092 ( .A1(n7857), .A2(n4744), .ZN(n7860) );
  AND2_X1 U6093 ( .A1(n7858), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4744) );
  NOR2_X1 U6094 ( .A1(n7856), .A2(n7855), .ZN(n8088) );
  NOR2_X1 U6095 ( .A1(n8096), .A2(n4743), .ZN(n8098) );
  AND2_X1 U6096 ( .A1(n8097), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U6097 ( .A1(n8098), .A2(n8099), .ZN(n9619) );
  OR2_X1 U6098 ( .A1(n9620), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4969) );
  INV_X1 U6099 ( .A(n4968), .ZN(n10131) );
  NAND2_X1 U6100 ( .A1(n4747), .A2(n4748), .ZN(n10143) );
  AND2_X1 U6101 ( .A1(n4751), .A2(n4750), .ZN(n10145) );
  XNOR2_X1 U6102 ( .A(n9622), .B(n9621), .ZN(n10155) );
  NAND2_X1 U6103 ( .A1(n4735), .A2(n4736), .ZN(n10170) );
  AND2_X1 U6104 ( .A1(n4433), .A2(n10171), .ZN(n4735) );
  NAND2_X1 U6105 ( .A1(n4971), .A2(n4970), .ZN(n10165) );
  OR2_X1 U6106 ( .A1(n10194), .A2(n10195), .ZN(n10197) );
  NAND2_X1 U6107 ( .A1(n10176), .A2(n9615), .ZN(n10189) );
  XNOR2_X1 U6108 ( .A(n9643), .B(n5034), .ZN(n4543) );
  AND2_X1 U6109 ( .A1(n7084), .A2(n7083), .ZN(n9671) );
  NAND2_X1 U6110 ( .A1(n9708), .A2(n4944), .ZN(n4942) );
  NAND2_X1 U6111 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U6112 ( .A1(n9710), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U6113 ( .A1(n9974), .A2(n10053), .ZN(n4628) );
  NAND2_X1 U6114 ( .A1(n9120), .A2(n7103), .ZN(n6897) );
  NAND2_X1 U6115 ( .A1(n4839), .A2(n4580), .ZN(n4690) );
  AND2_X1 U6116 ( .A1(n6845), .A2(n6844), .ZN(n9769) );
  NAND2_X1 U6117 ( .A1(n9773), .A2(n9402), .ZN(n9757) );
  NAND2_X1 U6118 ( .A1(n4921), .A2(n4925), .ZN(n9756) );
  NAND2_X1 U6119 ( .A1(n4584), .A2(n4928), .ZN(n4921) );
  NAND2_X1 U6120 ( .A1(n4930), .A2(n4932), .ZN(n9784) );
  NAND2_X1 U6121 ( .A1(n4931), .A2(n4458), .ZN(n4930) );
  INV_X1 U6122 ( .A(n4584), .ZN(n4931) );
  NAND2_X1 U6123 ( .A1(n4580), .A2(n9403), .ZN(n9775) );
  NAND2_X1 U6124 ( .A1(n4955), .A2(n4956), .ZN(n9803) );
  NAND2_X1 U6125 ( .A1(n7066), .A2(n7065), .ZN(n9879) );
  INV_X1 U6126 ( .A(n10048), .ZN(n7076) );
  AND2_X1 U6127 ( .A1(n6615), .A2(n6614), .ZN(n9203) );
  NAND2_X1 U6128 ( .A1(n5167), .A2(n9540), .ZN(n7978) );
  NAND2_X1 U6129 ( .A1(n6937), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5180) );
  OR3_X1 U6130 ( .A1(n10015), .A2(n10014), .A3(n10013), .ZN(n10082) );
  OR2_X1 U6131 ( .A1(n7209), .A2(n6650), .ZN(n6629) );
  NAND2_X2 U6132 ( .A1(n6556), .A2(n6555), .ZN(n8070) );
  AND2_X1 U6133 ( .A1(n10099), .A2(n10098), .ZN(n10208) );
  NOR2_X1 U6134 ( .A1(n5169), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5168) );
  INV_X1 U6135 ( .A(n6962), .ZN(n10115) );
  INV_X1 U6136 ( .A(n9522), .ZN(n7837) );
  INV_X1 U6137 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7204) );
  XNOR2_X1 U6138 ( .A(n6534), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U6139 ( .A1(n5428), .A2(n5383), .ZN(n7189) );
  AND2_X1 U6140 ( .A1(n6494), .A2(n6526), .ZN(n7290) );
  NAND2_X1 U6141 ( .A1(n4436), .A2(n6412), .ZN(n4737) );
  NAND2_X1 U6142 ( .A1(n7571), .A2(n5066), .ZN(n7576) );
  NAND2_X1 U6143 ( .A1(n4570), .A2(n4569), .ZN(P2_U3200) );
  NAND2_X1 U6144 ( .A1(n8726), .A2(n8727), .ZN(n4569) );
  NOR2_X1 U6145 ( .A1(n4571), .A2(n8724), .ZN(n4570) );
  NAND2_X1 U6146 ( .A1(n5943), .A2(n5942), .ZN(P2_U3205) );
  INV_X1 U6147 ( .A(n5941), .ZN(n5942) );
  OAI21_X1 U6148 ( .B1(n8954), .B2(n8941), .A(n5940), .ZN(n5941) );
  OAI22_X1 U6149 ( .A1(n8745), .A2(n9018), .B1(n10672), .B2(n5900), .ZN(n5901)
         );
  NAND2_X1 U6150 ( .A1(n8950), .A2(n8949), .ZN(n8953) );
  NAND2_X1 U6151 ( .A1(n8965), .A2(n4556), .ZN(P2_U3485) );
  INV_X1 U6152 ( .A(n4557), .ZN(n4556) );
  OAI21_X1 U6153 ( .B1(n9031), .B2(n9010), .A(n8964), .ZN(n4557) );
  OAI22_X1 U6154 ( .A1(n8745), .A2(n9101), .B1(n10336), .B2(n5914), .ZN(n5915)
         );
  INV_X1 U6155 ( .A(n5925), .ZN(n5926) );
  OAI21_X1 U6156 ( .B1(n8954), .B2(n9096), .A(n5924), .ZN(n5925) );
  NAND2_X1 U6157 ( .A1(n9030), .A2(n4554), .ZN(P2_U3453) );
  INV_X1 U6158 ( .A(n4555), .ZN(n4554) );
  OAI21_X1 U6159 ( .B1(n9031), .B2(n9096), .A(n9029), .ZN(n4555) );
  XNOR2_X1 U6160 ( .A(n4577), .B(n9225), .ZN(n9230) );
  INV_X1 U6161 ( .A(n4683), .ZN(P1_U3554) );
  AOI21_X1 U6162 ( .B1(n9596), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n4684), .ZN(
        n4683) );
  NOR2_X1 U6163 ( .A1(n9596), .A2(n7364), .ZN(n4684) );
  AOI21_X1 U6164 ( .B1(n10169), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9638), .ZN(
        n4978) );
  NAND2_X1 U6165 ( .A1(n9630), .A2(n9629), .ZN(n9637) );
  NAND2_X1 U6166 ( .A1(n9636), .A2(n9635), .ZN(n4977) );
  AOI21_X1 U6167 ( .B1(n9663), .B2(n9928), .A(n9662), .ZN(n9664) );
  XNOR2_X1 U6168 ( .A(n4948), .B(n5145), .ZN(n9663) );
  AND2_X1 U6169 ( .A1(n9945), .A2(n10063), .ZN(n4544) );
  AOI21_X1 U6170 ( .B1(n7138), .B2(n5194), .A(n5164), .ZN(n5163) );
  NAND2_X1 U6171 ( .A1(n5195), .A2(n5165), .ZN(n5164) );
  INV_X1 U6172 ( .A(n7116), .ZN(n7117) );
  OAI22_X1 U6173 ( .A1(n7132), .A2(n10032), .B1(n10252), .B2(n10514), .ZN(
        n7116) );
  AOI21_X1 U6174 ( .B1(n9680), .B2(n10063), .A(n4728), .ZN(n4727) );
  NOR2_X1 U6175 ( .A1(n10252), .A2(n10460), .ZN(n4728) );
  AOI21_X1 U6176 ( .B1(n10073), .B2(n10252), .A(n4694), .ZN(n9960) );
  NAND2_X1 U6177 ( .A1(n4696), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U6178 ( .A1(n4409), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n4695) );
  OAI21_X1 U6179 ( .B1(n9639), .B2(n5031), .A(n5029), .ZN(n10066) );
  NAND2_X1 U6180 ( .A1(n9941), .A2(n10243), .ZN(n5031) );
  AOI21_X1 U6181 ( .B1(n5030), .B2(n10243), .A(n5035), .ZN(n5029) );
  NOR2_X1 U6182 ( .A1(n7140), .A2(n7142), .ZN(n7143) );
  NOR2_X1 U6183 ( .A1(n10243), .A2(n7141), .ZN(n7142) );
  INV_X1 U6184 ( .A(n4843), .ZN(n4842) );
  OAI22_X1 U6185 ( .A1(n10072), .A2(n10090), .B1(n10243), .B2(n10565), .ZN(
        n4843) );
  INV_X1 U6186 ( .A(n4634), .ZN(n4633) );
  OAI22_X1 U6187 ( .A1(n10074), .A2(n10090), .B1(n10243), .B2(n6915), .ZN(
        n4634) );
  OAI222_X1 U6188 ( .A1(n10116), .A2(n8410), .B1(n8337), .B2(n9112), .C1(n4429), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI21_X1 U6189 ( .B1(n10111), .B2(n8337), .A(n5049), .ZN(P1_U3328) );
  INV_X1 U6190 ( .A(n5050), .ZN(n5049) );
  OAI222_X1 U6191 ( .A1(n10116), .A2(n8178), .B1(n8337), .B2(n8180), .C1(n8177), .C2(P1_U3086), .ZN(P1_U3333) );
  OAI222_X1 U6192 ( .A1(n10116), .A2(n10519), .B1(P1_U3086), .B2(n7993), .C1(
        n8337), .C2(n7994), .ZN(P1_U3334) );
  OAI222_X1 U6193 ( .A1(n10116), .A2(n7754), .B1(n8337), .B2(n7753), .C1(n9629), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U6194 ( .A1(n10116), .A2(n10623), .B1(n8337), .B2(n7612), .C1(
        n10201), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI222_X1 U6195 ( .A1(n10116), .A2(n7548), .B1(n8337), .B2(n7550), .C1(n9618), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U6196 ( .A1(n10116), .A2(n7493), .B1(n8337), .B2(n7492), .C1(
        P1_U3086), .C2(n9621), .ZN(P1_U3340) );
  OAI222_X1 U6197 ( .A1(n10116), .A2(n10549), .B1(n8337), .B2(n7329), .C1(
        P1_U3086), .C2(n7328), .ZN(P1_U3341) );
  OAI222_X1 U6198 ( .A1(n10116), .A2(n7234), .B1(n8337), .B2(n7233), .C1(
        P1_U3086), .C2(n7862), .ZN(P1_U3344) );
  OR2_X1 U6199 ( .A1(n8444), .A2(n8604), .ZN(n4431) );
  AND2_X1 U6200 ( .A1(n4535), .A2(n8201), .ZN(n4432) );
  INV_X1 U6201 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6651) );
  XNOR2_X1 U6202 ( .A(n6355), .B(n6354), .ZN(n6386) );
  OR2_X1 U6203 ( .A1(n9622), .A2(n9621), .ZN(n4433) );
  AND2_X1 U6204 ( .A1(n5962), .A2(n8083), .ZN(n4434) );
  AND2_X1 U6205 ( .A1(n9308), .A2(n4411), .ZN(n4435) );
  AND2_X1 U6206 ( .A1(n4900), .A2(n4448), .ZN(n6003) );
  AND2_X1 U6207 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4436) );
  NOR2_X1 U6208 ( .A1(n5971), .A2(n7490), .ZN(n5972) );
  AND2_X1 U6209 ( .A1(n4990), .A2(n4982), .ZN(n4437) );
  AND2_X1 U6210 ( .A1(n5055), .A2(n5054), .ZN(n4438) );
  AND4_X1 U6211 ( .A1(n6271), .A2(n6284), .A3(n6272), .A4(n8753), .ZN(n4439)
         );
  NAND2_X1 U6212 ( .A1(n8583), .A2(n8755), .ZN(n4440) );
  AND2_X1 U6213 ( .A1(n8444), .A2(n8604), .ZN(n4441) );
  INV_X1 U6214 ( .A(n9434), .ZN(n5158) );
  NAND2_X1 U6215 ( .A1(n8987), .A2(n8866), .ZN(n4442) );
  AND2_X1 U6216 ( .A1(n5612), .A2(SI_18_), .ZN(n4443) );
  NAND2_X1 U6217 ( .A1(n4502), .A2(n6341), .ZN(n5169) );
  NAND2_X1 U6218 ( .A1(n6236), .A2(n6081), .ZN(n6242) );
  INV_X1 U6219 ( .A(n6242), .ZN(n4779) );
  AND2_X1 U6220 ( .A1(n4435), .A2(n5061), .ZN(n4444) );
  XNOR2_X1 U6221 ( .A(n5612), .B(n5597), .ZN(n5611) );
  AND2_X1 U6222 ( .A1(n6837), .A2(n6836), .ZN(n4445) );
  AND2_X1 U6223 ( .A1(n6457), .A2(n6444), .ZN(n4446) );
  INV_X1 U6224 ( .A(n10032), .ZN(n10063) );
  INV_X1 U6225 ( .A(n8296), .ZN(n4898) );
  NAND2_X1 U6226 ( .A1(n4847), .A2(n5969), .ZN(n8634) );
  AND2_X1 U6227 ( .A1(n4748), .A2(n4525), .ZN(n4447) );
  AND2_X1 U6228 ( .A1(n4902), .A2(n4899), .ZN(n4448) );
  INV_X1 U6229 ( .A(n8688), .ZN(n4886) );
  NAND2_X1 U6230 ( .A1(n4908), .A2(n7202), .ZN(n8201) );
  OR2_X1 U6231 ( .A1(n9862), .A2(n9866), .ZN(n4449) );
  AND2_X1 U6232 ( .A1(n6429), .A2(n6428), .ZN(n4450) );
  AND2_X1 U6233 ( .A1(n7068), .A2(n9403), .ZN(n4451) );
  INV_X1 U6234 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4599) );
  OR2_X1 U6235 ( .A1(n9612), .A2(n9621), .ZN(n4452) );
  INV_X1 U6236 ( .A(n9758), .ZN(n4663) );
  OR2_X1 U6237 ( .A1(n10155), .A2(n10154), .ZN(n4736) );
  NAND2_X1 U6238 ( .A1(n9840), .A2(n9449), .ZN(n4453) );
  NAND2_X1 U6239 ( .A1(n6346), .A2(n6475), .ZN(n6626) );
  OR2_X1 U6240 ( .A1(n9731), .A2(n5058), .ZN(n4454) );
  OR2_X1 U6241 ( .A1(n6337), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U6242 ( .A1(n5641), .A2(n5640), .ZN(n4456) );
  AND2_X1 U6243 ( .A1(n5993), .A2(n8083), .ZN(n4457) );
  NAND2_X1 U6244 ( .A1(n10001), .A2(n9779), .ZN(n4458) );
  OR2_X1 U6245 ( .A1(n9643), .A2(n5033), .ZN(n4459) );
  NOR2_X1 U6246 ( .A1(n10009), .A2(n9586), .ZN(n4460) );
  NAND2_X1 U6247 ( .A1(n8167), .A2(n8168), .ZN(n8213) );
  INV_X1 U6248 ( .A(n4724), .ZN(n4723) );
  NAND2_X1 U6249 ( .A1(n5041), .A2(n4725), .ZN(n4724) );
  INV_X1 U6250 ( .A(n9651), .ZN(n5145) );
  AND2_X1 U6251 ( .A1(n4882), .A2(n4883), .ZN(n4461) );
  INV_X1 U6252 ( .A(n7060), .ZN(n9359) );
  NAND2_X1 U6253 ( .A1(n6368), .A2(n6370), .ZN(n4462) );
  NAND2_X1 U6254 ( .A1(n4690), .A2(n4837), .ZN(n9742) );
  OR2_X1 U6255 ( .A1(n5531), .A2(SI_14_), .ZN(n4463) );
  AND2_X1 U6256 ( .A1(n5419), .A2(n5388), .ZN(n4464) );
  XNOR2_X1 U6257 ( .A(n7006), .B(n6400), .ZN(n9457) );
  NAND2_X1 U6258 ( .A1(n5222), .A2(n5257), .ZN(n5946) );
  AND2_X1 U6259 ( .A1(n6202), .A2(n8820), .ZN(n4465) );
  AND4_X1 U6260 ( .A1(n6155), .A2(n6257), .A3(n8233), .A4(n6241), .ZN(n4466)
         );
  OR3_X1 U6261 ( .A1(n6742), .A2(P1_IR_REG_17__SCAN_IN), .A3(n4462), .ZN(n4467) );
  AND2_X1 U6262 ( .A1(n4721), .A2(n5611), .ZN(n4468) );
  OR2_X1 U6263 ( .A1(n9731), .A2(n9961), .ZN(n4469) );
  NAND2_X1 U6264 ( .A1(n4626), .A2(n8932), .ZN(n4470) );
  NAND2_X1 U6265 ( .A1(n4880), .A2(n4879), .ZN(n4883) );
  NAND2_X1 U6266 ( .A1(n6213), .A2(n6218), .ZN(n8777) );
  INV_X1 U6267 ( .A(n8777), .ZN(n4821) );
  AND3_X1 U6268 ( .A1(n9398), .A2(n9342), .A3(n9397), .ZN(n4471) );
  OR2_X1 U6269 ( .A1(n6000), .A2(n7274), .ZN(n4472) );
  AND3_X1 U6270 ( .A1(n8786), .A2(n4821), .A3(n8766), .ZN(n4473) );
  AND2_X1 U6271 ( .A1(n8829), .A2(n8843), .ZN(n4474) );
  AND2_X1 U6272 ( .A1(n9021), .A2(n6287), .ZN(n4475) );
  AND4_X1 U6273 ( .A1(n5202), .A2(n5201), .A3(n5322), .A4(n5320), .ZN(n4476)
         );
  INV_X1 U6274 ( .A(n9945), .ZN(n5034) );
  INV_X1 U6275 ( .A(n8851), .ZN(n4810) );
  NAND4_X1 U6276 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n10276)
         );
  OR2_X1 U6277 ( .A1(n8987), .A2(n8563), .ZN(n6189) );
  INV_X1 U6278 ( .A(n6189), .ZN(n5119) );
  INV_X1 U6279 ( .A(n5045), .ZN(n5044) );
  OAI21_X1 U6280 ( .B1(n4463), .B2(n5046), .A(n5549), .ZN(n5045) );
  AND2_X1 U6281 ( .A1(n8801), .A2(n8803), .ZN(n4477) );
  NOR2_X1 U6282 ( .A1(n9949), .A2(n9948), .ZN(n4478) );
  NAND2_X2 U6283 ( .A1(n5773), .A2(n5772), .ZN(n8951) );
  INV_X1 U6284 ( .A(n8951), .ZN(n4704) );
  INV_X1 U6285 ( .A(n4928), .ZN(n4927) );
  NOR2_X1 U6286 ( .A1(n4929), .A2(n7046), .ZN(n4928) );
  AND2_X1 U6287 ( .A1(n9092), .A2(n8920), .ZN(n4479) );
  AND3_X1 U6288 ( .A1(n4779), .A2(n6230), .A3(n6229), .ZN(n4480) );
  NAND2_X1 U6289 ( .A1(n6762), .A2(n6761), .ZN(n10009) );
  AND2_X1 U6290 ( .A1(n6590), .A2(n6589), .ZN(n7028) );
  INV_X1 U6291 ( .A(n7028), .ZN(n9590) );
  INV_X1 U6292 ( .A(n7006), .ZN(n7073) );
  AND2_X1 U6293 ( .A1(n6226), .A2(n6227), .ZN(n8753) );
  INV_X1 U6294 ( .A(n8753), .ZN(n5122) );
  INV_X1 U6295 ( .A(n5189), .ZN(n4801) );
  AND2_X1 U6296 ( .A1(n5106), .A2(n6147), .ZN(n4481) );
  NOR4_X1 U6297 ( .A1(n9453), .A2(n9452), .A3(n7059), .A4(n9451), .ZN(n4482)
         );
  AND2_X1 U6298 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4483) );
  NAND2_X1 U6299 ( .A1(n9690), .A2(n7052), .ZN(n4484) );
  INV_X1 U6300 ( .A(n4984), .ZN(n4983) );
  NAND2_X1 U6301 ( .A1(n4985), .A2(n4991), .ZN(n4984) );
  INV_X1 U6302 ( .A(n5419), .ZN(n4803) );
  NOR2_X1 U6303 ( .A1(n4644), .A2(n4640), .ZN(n4485) );
  OR2_X1 U6304 ( .A1(n8411), .A2(n8412), .ZN(n4486) );
  NAND2_X1 U6305 ( .A1(n9961), .A2(n9953), .ZN(n9431) );
  INV_X1 U6306 ( .A(n9431), .ZN(n4734) );
  INV_X1 U6307 ( .A(n4963), .ZN(n4962) );
  NOR2_X1 U6308 ( .A1(n7266), .A2(n4965), .ZN(n4963) );
  AND2_X1 U6309 ( .A1(n4444), .A2(n7076), .ZN(n4487) );
  AND2_X1 U6310 ( .A1(n9086), .A2(n8907), .ZN(n4488) );
  NOR2_X1 U6311 ( .A1(n10042), .A2(n9588), .ZN(n4489) );
  NOR2_X1 U6312 ( .A1(n9680), .A2(n9669), .ZN(n4490) );
  INV_X1 U6313 ( .A(n4987), .ZN(n4986) );
  NAND2_X1 U6314 ( .A1(n6716), .A2(n4988), .ZN(n4987) );
  NAND2_X1 U6315 ( .A1(n4580), .A2(n4451), .ZN(n9773) );
  INV_X1 U6316 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5808) );
  AND2_X1 U6317 ( .A1(n9996), .A2(n9982), .ZN(n4491) );
  NAND2_X1 U6318 ( .A1(n5815), .A2(n6116), .ZN(n6250) );
  INV_X1 U6319 ( .A(n10067), .ZN(n9445) );
  INV_X1 U6320 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9104) );
  AND2_X1 U6321 ( .A1(n9763), .A2(n9973), .ZN(n4492) );
  NOR2_X1 U6322 ( .A1(n8353), .A2(n8352), .ZN(n4493) );
  NOR2_X1 U6323 ( .A1(n8951), .A2(n5838), .ZN(n4494) );
  OR2_X1 U6324 ( .A1(n6742), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n4495) );
  INV_X1 U6325 ( .A(n5040), .ZN(n6340) );
  NAND2_X1 U6326 ( .A1(n4681), .A2(n4682), .ZN(n5040) );
  NOR2_X1 U6327 ( .A1(n8768), .A2(n8762), .ZN(n4496) );
  AND2_X1 U6328 ( .A1(n9421), .A2(n9480), .ZN(n9743) );
  INV_X1 U6329 ( .A(n9743), .ZN(n4692) );
  INV_X1 U6330 ( .A(n4647), .ZN(n4646) );
  NAND2_X1 U6331 ( .A1(n9374), .A2(n9364), .ZN(n4647) );
  AND2_X1 U6332 ( .A1(n4724), .A2(n5611), .ZN(n4497) );
  OR2_X1 U6333 ( .A1(n6204), .A2(n5115), .ZN(n4498) );
  AND3_X1 U6334 ( .A1(n9455), .A2(n4609), .A3(n4608), .ZN(n4499) );
  NAND2_X1 U6335 ( .A1(n6247), .A2(n6261), .ZN(n4500) );
  NAND2_X1 U6336 ( .A1(n8378), .A2(n8460), .ZN(n4501) );
  AND2_X1 U6337 ( .A1(n6315), .A2(n6314), .ZN(n4502) );
  AND2_X1 U6338 ( .A1(n4431), .A2(n5419), .ZN(n4503) );
  INV_X1 U6339 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6365) );
  OR2_X1 U6340 ( .A1(n7266), .A2(n7245), .ZN(n4504) );
  AND2_X1 U6341 ( .A1(n6180), .A2(n6237), .ZN(n4505) );
  INV_X1 U6342 ( .A(n7166), .ZN(n4892) );
  AND3_X1 U6343 ( .A1(n4883), .A2(n4882), .A3(n4881), .ZN(n4506) );
  NOR2_X1 U6344 ( .A1(n6956), .A2(n6955), .ZN(n4507) );
  AND2_X1 U6345 ( .A1(n9498), .A2(n9426), .ZN(n9686) );
  INV_X1 U6346 ( .A(n9686), .ZN(n5156) );
  AND2_X1 U6347 ( .A1(n9028), .A2(n8779), .ZN(n4508) );
  AND2_X1 U6348 ( .A1(n5430), .A2(n5429), .ZN(n4509) );
  AND2_X1 U6349 ( .A1(n6180), .A2(n6179), .ZN(n4510) );
  INV_X1 U6350 ( .A(n5008), .ZN(n5007) );
  OAI21_X1 U6351 ( .B1(n9265), .B2(n5009), .A(n9264), .ZN(n5008) );
  INV_X1 U6352 ( .A(n8578), .ZN(n8789) );
  AND2_X1 U6353 ( .A1(n5731), .A2(n5730), .ZN(n8578) );
  AND2_X1 U6354 ( .A1(n5149), .A2(n5145), .ZN(n4511) );
  AND2_X1 U6355 ( .A1(n6134), .A2(n6147), .ZN(n4512) );
  NAND2_X1 U6356 ( .A1(n5693), .A2(n8817), .ZN(n4513) );
  AOI21_X1 U6357 ( .B1(n8689), .B2(n8687), .A(n8688), .ZN(n4884) );
  AND2_X1 U6358 ( .A1(n6181), .A2(n6174), .ZN(n4514) );
  AND2_X1 U6359 ( .A1(n4973), .A2(n4452), .ZN(n4515) );
  AND2_X1 U6360 ( .A1(n5037), .A2(n5475), .ZN(n4516) );
  AND2_X1 U6361 ( .A1(n4709), .A2(n5411), .ZN(n4517) );
  AND2_X1 U6362 ( .A1(n4736), .A2(n4433), .ZN(n4518) );
  AND2_X1 U6363 ( .A1(n4882), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4519) );
  AND2_X1 U6364 ( .A1(n8014), .A2(n8608), .ZN(n4520) );
  AND2_X1 U6365 ( .A1(n5137), .A2(n10387), .ZN(n4521) );
  INV_X1 U6366 ( .A(n5470), .ZN(n5038) );
  INV_X1 U6367 ( .A(n6173), .ZN(n4773) );
  INV_X1 U6368 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5214) );
  AND2_X1 U6369 ( .A1(n8395), .A2(n4473), .ZN(n4522) );
  INV_X1 U6370 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6371 ( .A1(n4871), .A2(n7202), .ZN(n8193) );
  INV_X1 U6372 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4846) );
  OAI21_X1 U6373 ( .B1(n7658), .B2(n7059), .A(n9537), .ZN(n7704) );
  AND2_X1 U6374 ( .A1(n4995), .A2(n4999), .ZN(n4523) );
  NOR2_X1 U6375 ( .A1(n5205), .A2(n5389), .ZN(n5619) );
  INV_X1 U6376 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4863) );
  INV_X1 U6377 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6378 ( .A1(n9915), .A2(n7034), .ZN(n9887) );
  NAND2_X1 U6379 ( .A1(n5818), .A2(n6130), .ZN(n7893) );
  NAND2_X1 U6380 ( .A1(n6803), .A2(n6802), .ZN(n10001) );
  INV_X1 U6381 ( .A(n10001), .ZN(n5054) );
  AOI21_X1 U6382 ( .B1(n8296), .B2(n10488), .A(n4897), .ZN(n4896) );
  NAND2_X1 U6383 ( .A1(n4444), .A2(n8001), .ZN(n4524) );
  NAND2_X1 U6384 ( .A1(n7893), .A2(n6141), .ZN(n7920) );
  INV_X1 U6385 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4586) );
  INV_X1 U6386 ( .A(n8894), .ZN(n8865) );
  AND3_X1 U6387 ( .A1(n5571), .A2(n5570), .A3(n5569), .ZN(n8894) );
  NAND2_X1 U6388 ( .A1(n10148), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4525) );
  AND2_X1 U6389 ( .A1(n4702), .A2(n10589), .ZN(n4526) );
  INV_X1 U6390 ( .A(n7830), .ZN(n7075) );
  INV_X1 U6391 ( .A(n9680), .ZN(n10072) );
  OR2_X1 U6392 ( .A1(n8645), .A2(n6040), .ZN(n4527) );
  OR2_X1 U6393 ( .A1(n6029), .A2(n7198), .ZN(n4528) );
  OR2_X1 U6394 ( .A1(n9051), .A2(n9101), .ZN(n4529) );
  AND2_X1 U6395 ( .A1(n8649), .A2(n5969), .ZN(n4530) );
  INV_X1 U6396 ( .A(n7490), .ZN(n4899) );
  AND2_X1 U6397 ( .A1(n8177), .A2(n9635), .ZN(n9449) );
  AND2_X1 U6398 ( .A1(n5181), .A2(n7837), .ZN(n10002) );
  INV_X1 U6399 ( .A(n8653), .ZN(n4903) );
  AND2_X1 U6400 ( .A1(n7667), .A2(n7811), .ZN(n7705) );
  XOR2_X1 U6401 ( .A(n8294), .B(P2_REG1_REG_12__SCAN_IN), .Z(n4531) );
  INV_X1 U6402 ( .A(n10095), .ZN(n5061) );
  AND2_X1 U6403 ( .A1(n4870), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4532) );
  AND2_X1 U6404 ( .A1(n4712), .A2(n4711), .ZN(n4533) );
  AND2_X1 U6405 ( .A1(n8684), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4534) );
  AND2_X1 U6406 ( .A1(n4913), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4535) );
  INV_X1 U6407 ( .A(n8677), .ZN(n4870) );
  AND2_X1 U6408 ( .A1(n5989), .A2(n7557), .ZN(n4536) );
  AND2_X1 U6409 ( .A1(n4707), .A2(n4706), .ZN(n4537) );
  OR2_X1 U6410 ( .A1(n6043), .A2(n5973), .ZN(n4538) );
  INV_X1 U6411 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10294) );
  INV_X1 U6412 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5138) );
  XOR2_X1 U6413 ( .A(n7179), .B(P2_REG1_REG_6__SCAN_IN), .Z(n4539) );
  AND2_X1 U6414 ( .A1(n4893), .A2(n7308), .ZN(n4540) );
  INV_X1 U6415 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4700) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4918) );
  INV_X1 U6417 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4588) );
  INV_X1 U6418 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n4858) );
  OAI222_X1 U6419 ( .A1(n8338), .A2(n10116), .B1(n8337), .B2(n8407), .C1(
        P1_U3086), .C2(n8336), .ZN(P1_U3325) );
  OAI222_X1 U6420 ( .A1(n10116), .A2(n7176), .B1(n8337), .B2(n7175), .C1(
        P1_U3086), .C2(n7249), .ZN(P1_U3351) );
  OAI222_X1 U6421 ( .A1(n10116), .A2(n7204), .B1(n8337), .B2(n7203), .C1(n7536), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X2 U6422 ( .A1(n7161), .A2(P1_U3086), .ZN(n10116) );
  OAI222_X1 U6423 ( .A1(n10116), .A2(n4918), .B1(n8337), .B2(n7162), .C1(n7218), .C2(P1_U3086), .ZN(P1_U3354) );
  OAI222_X1 U6424 ( .A1(n10116), .A2(n8312), .B1(P1_U3086), .B2(n8311), .C1(
        n8337), .C2(n9109), .ZN(P1_U3326) );
  OAI222_X1 U6425 ( .A1(n10116), .A2(n7210), .B1(n8337), .B2(n7209), .C1(n8092), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI22_X1 U6426 ( .A1(n5048), .A2(P1_U3086), .B1(n10116), .B2(n10112), .ZN(
        n5050) );
  NAND2_X1 U6427 ( .A1(n8864), .A2(n5609), .ZN(n5610) );
  NAND2_X1 U6428 ( .A1(n9050), .A2(n4529), .ZN(P2_U3449) );
  NAND2_X2 U6429 ( .A1(n5244), .A2(n7409), .ZN(n5815) );
  NAND2_X1 U6430 ( .A1(n8852), .A2(n8851), .ZN(n4813) );
  NAND2_X1 U6431 ( .A1(n6397), .A2(n6398), .ZN(n4542) );
  NAND2_X1 U6432 ( .A1(n4578), .A2(n9224), .ZN(n4577) );
  NAND2_X1 U6433 ( .A1(n4482), .A2(n4607), .ZN(n9459) );
  OR2_X1 U6435 ( .A1(n9944), .A2(n4544), .ZN(P1_U3552) );
  NAND2_X4 U6436 ( .A1(n4420), .A2(n6393), .ZN(n6650) );
  NOR2_X4 U6437 ( .A1(n7739), .A2(n7740), .ZN(n7738) );
  NOR2_X2 U6438 ( .A1(n9918), .A2(n10042), .ZN(n9890) );
  NOR2_X4 U6439 ( .A1(n4449), .A2(n10020), .ZN(n9847) );
  AOI21_X1 U6440 ( .B1(n5004), .B2(n5008), .A(n4445), .ZN(n5002) );
  NAND2_X1 U6441 ( .A1(n6800), .A2(n6801), .ZN(n5009) );
  NAND2_X1 U6442 ( .A1(n5036), .A2(n4516), .ZN(n5492) );
  AOI21_X1 U6443 ( .B1(n9639), .B2(n10002), .A(n9640), .ZN(n10065) );
  NAND2_X1 U6444 ( .A1(n5272), .A2(n5275), .ZN(n4547) );
  OAI21_X2 U6445 ( .B1(n6083), .B2(n6082), .A(n6234), .ZN(n6096) );
  OAI21_X1 U6446 ( .B1(n5785), .B2(n5786), .A(n5795), .ZN(n4582) );
  OAI21_X1 U6447 ( .B1(n5131), .B2(n8270), .A(n5129), .ZN(n8916) );
  OAI21_X1 U6448 ( .B1(n6303), .B2(n4548), .A(n6302), .ZN(P2_U3296) );
  NAND4_X1 U6449 ( .A1(n6293), .A2(n6295), .A3(n6292), .A4(n6294), .ZN(n4548)
         );
  NAND2_X1 U6450 ( .A1(n5492), .A2(n5491), .ZN(n5498) );
  OAI21_X1 U6451 ( .B1(n9433), .B2(n9498), .A(n9504), .ZN(n4623) );
  NAND2_X2 U6452 ( .A1(n5516), .A2(n5515), .ZN(n5532) );
  AND3_X1 U6453 ( .A1(n6270), .A2(n4522), .A3(n4779), .ZN(n4606) );
  OR4_X2 U6454 ( .A1(n6266), .A2(n6265), .A3(n8898), .A4(n6264), .ZN(n6267) );
  NAND2_X1 U6455 ( .A1(n5576), .A2(n5575), .ZN(n5579) );
  NAND2_X1 U6456 ( .A1(n4549), .A2(n8881), .ZN(n4756) );
  NAND2_X1 U6457 ( .A1(n6175), .A2(n4505), .ZN(n4549) );
  NAND2_X1 U6458 ( .A1(n4550), .A2(n6152), .ZN(n6154) );
  NAND2_X1 U6459 ( .A1(n6151), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U6460 ( .A1(n4552), .A2(n7131), .ZN(n9437) );
  NAND4_X1 U6461 ( .A1(n9435), .A2(n9499), .A3(n9434), .A4(n9449), .ZN(n4552)
         );
  NAND2_X1 U6462 ( .A1(n4553), .A2(n6126), .ZN(n6128) );
  NAND2_X1 U6463 ( .A1(n6119), .A2(n6118), .ZN(n4553) );
  NAND3_X1 U6464 ( .A1(n6163), .A2(n4763), .A3(n6162), .ZN(n4615) );
  NAND2_X1 U6465 ( .A1(n4563), .A2(n6209), .ZN(n6214) );
  INV_X1 U6466 ( .A(n9439), .ZN(n4650) );
  NAND2_X1 U6467 ( .A1(n5492), .A2(n5476), .ZN(n7209) );
  NAND2_X1 U6468 ( .A1(n5837), .A2(n6221), .ZN(n8752) );
  NAND2_X1 U6469 ( .A1(n4560), .A2(n4559), .ZN(n5499) );
  INV_X1 U6470 ( .A(n5497), .ZN(n4559) );
  INV_X1 U6471 ( .A(n5498), .ZN(n4560) );
  OAI21_X1 U6472 ( .B1(n4808), .B2(n4806), .A(n4513), .ZN(n4804) );
  INV_X1 U6473 ( .A(n7273), .ZN(n4583) );
  NAND2_X1 U6474 ( .A1(n8776), .A2(n5733), .ZN(n8767) );
  AND2_X1 U6475 ( .A1(n9479), .A2(n4648), .ZN(n9584) );
  MUX2_X1 U6476 ( .A(n9441), .B(n9449), .S(n9945), .Z(n9439) );
  NAND2_X1 U6477 ( .A1(n4691), .A2(n4693), .ZN(n4689) );
  INV_X1 U6478 ( .A(n8915), .ZN(n6263) );
  NAND2_X1 U6479 ( .A1(n6232), .A2(n4616), .ZN(n4775) );
  NAND2_X1 U6480 ( .A1(n6486), .A2(n6485), .ZN(n7842) );
  AOI21_X2 U6481 ( .B1(n6893), .B2(n6892), .A(n9239), .ZN(n9243) );
  NAND2_X1 U6482 ( .A1(n7394), .A2(n7393), .ZN(n7496) );
  AND2_X1 U6483 ( .A1(n7277), .A2(n6380), .ZN(n7362) );
  NAND2_X1 U6484 ( .A1(n7278), .A2(n7279), .ZN(n7277) );
  NAND3_X2 U6485 ( .A1(n7523), .A2(n7522), .A3(n7524), .ZN(n7571) );
  OAI21_X2 U6486 ( .B1(n5874), .B2(n5873), .A(n5890), .ZN(n5875) );
  NAND2_X1 U6487 ( .A1(n8419), .A2(n8420), .ZN(n8585) );
  NAND2_X2 U6488 ( .A1(n5877), .A2(n5876), .ZN(n7194) );
  OR2_X2 U6489 ( .A1(n7194), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5894) );
  INV_X1 U6490 ( .A(n5809), .ZN(n5807) );
  NAND2_X1 U6491 ( .A1(n5809), .A2(n5808), .ZN(n5858) );
  AND2_X2 U6492 ( .A1(n5619), .A2(n5618), .ZN(n5809) );
  NAND2_X1 U6493 ( .A1(n8561), .A2(n8560), .ZN(n8370) );
  NAND2_X1 U6494 ( .A1(n4981), .A2(n4979), .ZN(n9232) );
  NAND2_X1 U6495 ( .A1(n6760), .A2(n6759), .ZN(n9160) );
  NAND2_X1 U6496 ( .A1(n4594), .A2(n4593), .ZN(n5018) );
  NAND2_X1 U6497 ( .A1(n8017), .A2(n8016), .ZN(n8166) );
  OAI21_X1 U6498 ( .B1(n4650), .B2(n9444), .A(n4649), .ZN(n9479) );
  OAI211_X1 U6499 ( .C1(n9417), .C2(n9416), .A(n9415), .B(n9414), .ZN(n9418)
         );
  NAND2_X1 U6500 ( .A1(n9610), .A2(n4969), .ZN(n10132) );
  NOR2_X1 U6501 ( .A1(n7532), .A2(n4974), .ZN(n7533) );
  AOI21_X1 U6502 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n7248), .A(n7243), .ZN(
        n7478) );
  NAND2_X1 U6503 ( .A1(n6288), .A2(n4475), .ZN(n6289) );
  NAND2_X1 U6504 ( .A1(n6214), .A2(n4567), .ZN(n6216) );
  NAND3_X1 U6505 ( .A1(n4776), .A2(n4775), .A3(n4568), .ZN(n4777) );
  OAI21_X2 U6506 ( .B1(n7953), .B2(n7954), .A(n4528), .ZN(n8075) );
  NOR2_X1 U6507 ( .A1(n7330), .A2(n4789), .ZN(n7307) );
  NAND2_X1 U6508 ( .A1(n7430), .A2(n7429), .ZN(n7428) );
  NAND2_X1 U6509 ( .A1(n8622), .A2(n8621), .ZN(n8620) );
  AOI22_X2 U6510 ( .A1(n8787), .A2(n5714), .B1(n8807), .B2(n9040), .ZN(n8778)
         );
  NAND2_X1 U6511 ( .A1(n7305), .A2(n4788), .ZN(n7430) );
  NAND2_X1 U6512 ( .A1(n7346), .A2(n4783), .ZN(n8622) );
  NAND2_X1 U6513 ( .A1(n4812), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U6514 ( .A1(n4818), .A2(n4819), .ZN(n8754) );
  NOR2_X1 U6515 ( .A1(n8958), .A2(n8957), .ZN(n9024) );
  OAI21_X2 U6516 ( .B1(n8388), .B2(n5084), .A(n5082), .ZN(n8572) );
  INV_X1 U6517 ( .A(n9329), .ZN(n4578) );
  INV_X1 U6518 ( .A(n6595), .ZN(n4594) );
  NOR2_X1 U6519 ( .A1(n8013), .A2(n4520), .ZN(n8017) );
  INV_X1 U6520 ( .A(n4582), .ZN(n4581) );
  NAND2_X1 U6521 ( .A1(n4410), .A2(n5114), .ZN(n5111) );
  NAND2_X1 U6522 ( .A1(n4439), .A2(n4606), .ZN(n4715) );
  AOI21_X2 U6523 ( .B1(n10109), .B2(n6106), .A(n6105), .ZN(n9021) );
  NAND2_X1 U6524 ( .A1(n4583), .A2(n6106), .ZN(n5506) );
  NAND2_X1 U6525 ( .A1(n5499), .A2(n5516), .ZN(n7273) );
  OAI21_X2 U6526 ( .B1(n8900), .B2(n8898), .A(n6180), .ZN(n8879) );
  NAND2_X1 U6527 ( .A1(n8856), .A2(n4810), .ZN(n8858) );
  INV_X1 U6528 ( .A(n7209), .ZN(n4592) );
  AOI21_X1 U6529 ( .B1(n5426), .B2(n5427), .A(n4509), .ZN(n4952) );
  INV_X1 U6530 ( .A(n4944), .ZN(n4940) );
  NAND2_X1 U6531 ( .A1(n7736), .A2(n7010), .ZN(n7647) );
  NAND2_X1 U6532 ( .A1(n10073), .A2(n10243), .ZN(n4635) );
  NAND2_X4 U6533 ( .A1(n6395), .A2(n6396), .ZN(n7006) );
  NAND2_X1 U6534 ( .A1(n7307), .A2(n7306), .ZN(n7305) );
  OAI22_X1 U6535 ( .A1(n8681), .A2(n8680), .B1(n6044), .B2(n8684), .ZN(n8698)
         );
  NAND2_X1 U6536 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  AOI21_X1 U6537 ( .B1(n8666), .B2(n8665), .A(n4784), .ZN(n8681) );
  NAND2_X1 U6538 ( .A1(n6056), .A2(n8704), .ZN(n6064) );
  NOR2_X1 U6539 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  NAND2_X1 U6540 ( .A1(n7347), .A2(n7348), .ZN(n7346) );
  OAI21_X2 U6541 ( .B1(n6010), .B2(n4588), .A(n4587), .ZN(n6011) );
  NAND2_X1 U6542 ( .A1(n8075), .A2(n8074), .ZN(n4786) );
  NAND2_X1 U6543 ( .A1(n4592), .A2(n6106), .ZN(n5481) );
  AND2_X2 U6544 ( .A1(n9724), .A2(n9483), .ZN(n9711) );
  NAND3_X1 U6545 ( .A1(n4688), .A2(n4689), .A3(n5170), .ZN(n9724) );
  NAND2_X1 U6546 ( .A1(n5148), .A2(n5155), .ZN(n7118) );
  NAND3_X1 U6547 ( .A1(n5273), .A2(n5275), .A3(n5274), .ZN(n4590) );
  NAND2_X1 U6548 ( .A1(n5376), .A2(n5375), .ZN(n5382) );
  OAI21_X1 U6549 ( .B1(n5646), .B2(n5648), .A(n5647), .ZN(n5636) );
  NAND2_X1 U6550 ( .A1(n7088), .A2(n4618), .ZN(n7115) );
  NAND3_X1 U6551 ( .A1(n9967), .A2(n7050), .A3(n4941), .ZN(n4938) );
  NAND2_X1 U6552 ( .A1(n8872), .A2(n6247), .ZN(n8856) );
  NAND2_X1 U6553 ( .A1(n7042), .A2(n4957), .ZN(n4955) );
  NAND3_X1 U6554 ( .A1(n5018), .A2(n9295), .A3(n6598), .ZN(n9148) );
  NAND2_X1 U6555 ( .A1(n7019), .A2(n7018), .ZN(n7700) );
  NAND2_X1 U6556 ( .A1(n4597), .A2(n9528), .ZN(n9453) );
  INV_X1 U6557 ( .A(n7057), .ZN(n4597) );
  OR2_X1 U6558 ( .A1(n10225), .A2(n6537), .ZN(n6419) );
  NAND2_X1 U6559 ( .A1(n7785), .A2(n6462), .ZN(n6483) );
  NAND2_X1 U6560 ( .A1(n4994), .A2(n4992), .ZN(n9253) );
  NAND2_X1 U6561 ( .A1(n7497), .A2(n7498), .ZN(n7523) );
  XNOR2_X2 U6562 ( .A(n5813), .B(n4599), .ZN(n7838) );
  NAND2_X1 U6563 ( .A1(n8367), .A2(n8366), .ZN(n8561) );
  NAND2_X1 U6564 ( .A1(n4600), .A2(n4599), .ZN(n5811) );
  INV_X1 U6565 ( .A(n5858), .ZN(n4600) );
  NAND2_X1 U6566 ( .A1(n5086), .A2(n5085), .ZN(n8533) );
  NAND2_X2 U6567 ( .A1(n8485), .A2(n8486), .ZN(n8388) );
  NAND2_X1 U6568 ( .A1(n6285), .A2(n4601), .ZN(n6293) );
  NAND2_X1 U6569 ( .A1(n4602), .A2(n5230), .ZN(n5237) );
  NAND2_X1 U6570 ( .A1(n4404), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U6571 ( .A1(n6178), .A2(n4514), .ZN(n6175) );
  NAND2_X1 U6572 ( .A1(n4603), .A2(n6183), .ZN(n6184) );
  AND2_X1 U6573 ( .A1(n6178), .A2(n4510), .ZN(n4604) );
  XNOR2_X2 U6574 ( .A(n5232), .B(n5231), .ZN(n8408) );
  OAI21_X1 U6575 ( .B1(n9741), .B2(n7049), .A(n7048), .ZN(n9737) );
  NAND2_X1 U6576 ( .A1(n7700), .A2(n7020), .ZN(n7024) );
  NAND2_X1 U6577 ( .A1(n4635), .A2(n4633), .ZN(P1_U3516) );
  INV_X1 U6578 ( .A(n9457), .ZN(n4610) );
  OR2_X2 U6579 ( .A1(n6650), .A2(n7162), .ZN(n6395) );
  OR2_X1 U6580 ( .A1(n5951), .A2(n7166), .ZN(n5952) );
  NAND2_X1 U6581 ( .A1(n7431), .A2(n4862), .ZN(n4861) );
  OR4_X2 U6582 ( .A1(n8829), .A2(n8843), .A3(n6267), .A4(n8851), .ZN(n6268) );
  NAND3_X2 U6583 ( .A1(n4681), .A2(n4682), .A3(n5168), .ZN(n10102) );
  NAND2_X1 U6584 ( .A1(n5127), .A2(n5126), .ZN(n5135) );
  NOR2_X1 U6585 ( .A1(n6096), .A2(n6095), .ZN(n6281) );
  NAND2_X1 U6586 ( .A1(n4951), .A2(n4950), .ZN(n5471) );
  OAI21_X2 U6587 ( .B1(n5662), .B2(n5661), .A(n5660), .ZN(n5679) );
  NAND2_X1 U6588 ( .A1(n4655), .A2(n4654), .ZN(n9428) );
  NAND2_X1 U6589 ( .A1(n9443), .A2(n9445), .ZN(n4649) );
  NOR2_X1 U6590 ( .A1(n9430), .A2(n9429), .ZN(n9438) );
  NAND2_X1 U6591 ( .A1(n5333), .A2(n5332), .ZN(n5340) );
  INV_X1 U6592 ( .A(n4652), .ZN(n4651) );
  NAND2_X1 U6593 ( .A1(n9024), .A2(n10672), .ZN(n8962) );
  NAND2_X1 U6594 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  INV_X1 U6595 ( .A(n5097), .ZN(n5874) );
  INV_X1 U6596 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U6597 ( .A1(n4715), .A2(n6275), .ZN(n6288) );
  NAND2_X1 U6598 ( .A1(n8334), .A2(n8323), .ZN(n8332) );
  NAND2_X1 U6599 ( .A1(n4613), .A2(n4512), .ZN(n6135) );
  AND2_X1 U6600 ( .A1(n6145), .A2(n6130), .ZN(n4614) );
  NAND2_X1 U6601 ( .A1(n4615), .A2(n7148), .ZN(n6166) );
  NAND2_X1 U6602 ( .A1(n4765), .A2(n6152), .ZN(n4764) );
  INV_X1 U6603 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U6604 ( .A1(n5227), .A2(n5100), .ZN(n5102) );
  NAND2_X1 U6605 ( .A1(n7704), .A2(n9535), .ZN(n5167) );
  NAND2_X1 U6606 ( .A1(n7066), .A2(n4685), .ZN(n9880) );
  OAI21_X2 U6607 ( .B1(n9711), .B2(n4734), .A(n4732), .ZN(n9696) );
  NAND2_X1 U6608 ( .A1(n4942), .A2(n4943), .ZN(n9687) );
  OAI21_X1 U6609 ( .B1(n10071), .B2(n4409), .A(n4727), .ZN(P1_U3549) );
  OAI21_X1 U6610 ( .B1(n10071), .B2(n7144), .A(n4842), .ZN(P1_U3517) );
  OAI21_X1 U6611 ( .B1(n9438), .B2(n9437), .A(n9436), .ZN(n9441) );
  NOR3_X2 U6612 ( .A1(n6879), .A2(n6878), .A3(n6877), .ZN(n4624) );
  NOR2_X2 U6613 ( .A1(n6782), .A2(n6781), .ZN(n4625) );
  OAI21_X2 U6614 ( .B1(n6232), .B2(n6233), .A(n4480), .ZN(n4776) );
  NAND2_X1 U6615 ( .A1(n8060), .A2(n5213), .ZN(n4781) );
  OAI21_X1 U6616 ( .B1(n5302), .B2(n4918), .A(n4917), .ZN(n5215) );
  NAND2_X1 U6617 ( .A1(n4934), .A2(n4933), .ZN(n9872) );
  NAND2_X2 U6618 ( .A1(n9967), .A2(n7050), .ZN(n9708) );
  INV_X1 U6619 ( .A(n5560), .ZN(n4790) );
  NAND4_X1 U6620 ( .A1(n4791), .A2(n4792), .A3(n4793), .A4(n5198), .ZN(n5560)
         );
  NAND2_X1 U6621 ( .A1(n4636), .A2(n5187), .ZN(n6224) );
  NAND2_X1 U6622 ( .A1(n4757), .A2(n6217), .ZN(n4636) );
  AND3_X2 U6623 ( .A1(n4637), .A2(n4777), .A3(n7838), .ZN(n6285) );
  NAND2_X1 U6624 ( .A1(n4774), .A2(n5171), .ZN(n4637) );
  NAND2_X1 U6625 ( .A1(n4764), .A2(n4466), .ZN(n4763) );
  NAND2_X1 U6626 ( .A1(n4769), .A2(n4767), .ZN(n6178) );
  NAND2_X1 U6627 ( .A1(n6139), .A2(n8129), .ZN(n4765) );
  INV_X1 U6628 ( .A(n6214), .ZN(n4758) );
  AOI21_X1 U6629 ( .B1(n9375), .B2(n9365), .A(n9377), .ZN(n9368) );
  INV_X1 U6630 ( .A(n9423), .ZN(n4661) );
  AND2_X1 U6631 ( .A1(n4653), .A2(n4651), .ZN(n9432) );
  OAI21_X1 U6632 ( .B1(n4661), .B2(n4665), .A(n9424), .ZN(n4652) );
  NAND3_X1 U6633 ( .A1(n9418), .A2(n9758), .A3(n4664), .ZN(n4653) );
  AND2_X1 U6634 ( .A1(n4657), .A2(n4659), .ZN(n4654) );
  INV_X2 U6635 ( .A(n6937), .ZN(n6465) );
  NAND2_X1 U6636 ( .A1(n4671), .A2(n4670), .ZN(n4666) );
  OAI211_X1 U6637 ( .C1(n4677), .C2(n4453), .A(n4671), .B(n4668), .ZN(n9413)
         );
  AND2_X1 U6638 ( .A1(n9525), .A2(n4675), .ZN(n4674) );
  INV_X1 U6639 ( .A(n9395), .ZN(n4676) );
  NAND2_X1 U6640 ( .A1(n9396), .A2(n9547), .ZN(n4677) );
  NAND3_X1 U6641 ( .A1(n4680), .A2(n9346), .A3(n4678), .ZN(n7658) );
  NAND4_X1 U6642 ( .A1(n5162), .A2(n9529), .A3(n9528), .A4(n7743), .ZN(n4678)
         );
  NAND3_X1 U6643 ( .A1(n5162), .A2(n4679), .A3(n9529), .ZN(n4680) );
  NAND2_X1 U6644 ( .A1(n7658), .A2(n9449), .ZN(n9345) );
  AND2_X2 U6645 ( .A1(n6411), .A2(n6308), .ZN(n6475) );
  AND4_X2 U6646 ( .A1(n6307), .A2(n6304), .A3(n6306), .A4(n6305), .ZN(n6346)
         );
  NAND2_X1 U6647 ( .A1(n7007), .A2(n5016), .ZN(n7587) );
  AOI21_X1 U6648 ( .B1(n7007), .B2(n9527), .A(n7993), .ZN(n9530) );
  XNOR2_X1 U6649 ( .A(n7007), .B(n9527), .ZN(n10213) );
  AOI22_X1 U6650 ( .A1(n10212), .A2(n7009), .B1(n7007), .B2(n10053), .ZN(n7605) );
  INV_X1 U6651 ( .A(n7007), .ZN(n7364) );
  NAND2_X1 U6652 ( .A1(n9794), .A2(n4691), .ZN(n4688) );
  MUX2_X1 U6653 ( .A(n4701), .B(n4700), .S(n7161), .Z(n5403) );
  AND2_X4 U6654 ( .A1(n4781), .A2(n4717), .ZN(n5302) );
  NAND2_X1 U6655 ( .A1(n5724), .A2(n4707), .ZN(n5762) );
  NAND2_X1 U6656 ( .A1(n5724), .A2(n4537), .ZN(n5774) );
  NAND2_X1 U6657 ( .A1(n5724), .A2(n5723), .ZN(n5743) );
  NAND2_X1 U6658 ( .A1(n5368), .A2(n4517), .ZN(n5439) );
  NAND3_X1 U6659 ( .A1(n5312), .A2(n10294), .A3(n5293), .ZN(n5344) );
  INV_X1 U6660 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4718) );
  NAND2_X1 U6661 ( .A1(n5326), .A2(n5325), .ZN(n5333) );
  INV_X1 U6662 ( .A(n5217), .ZN(n5273) );
  NAND2_X1 U6663 ( .A1(n9711), .A2(n4732), .ZN(n4730) );
  NAND2_X1 U6664 ( .A1(n4730), .A2(n4731), .ZN(n9679) );
  NAND2_X1 U6665 ( .A1(n9711), .A2(n7070), .ZN(n9710) );
  OR2_X2 U6666 ( .A1(n5679), .A2(n5678), .ZN(n5028) );
  NAND2_X1 U6667 ( .A1(n10170), .A2(n9623), .ZN(n10181) );
  INV_X1 U6668 ( .A(n4736), .ZN(n10153) );
  INV_X1 U6669 ( .A(n4751), .ZN(n10128) );
  NAND2_X1 U6670 ( .A1(n10136), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4750) );
  NAND2_X2 U6671 ( .A1(n4756), .A2(n6177), .ZN(n6186) );
  NAND2_X1 U6672 ( .A1(n6166), .A2(n4771), .ZN(n4766) );
  NAND2_X1 U6673 ( .A1(n4766), .A2(n6168), .ZN(n4770) );
  NAND3_X1 U6674 ( .A1(n6171), .A2(n4770), .A3(n4773), .ZN(n4769) );
  NAND2_X1 U6675 ( .A1(n6166), .A2(n6165), .ZN(n6170) );
  NAND3_X1 U6676 ( .A1(n4776), .A2(n6239), .A3(n4775), .ZN(n4774) );
  NAND2_X1 U6677 ( .A1(n5278), .A2(n4780), .ZN(n5279) );
  NAND2_X1 U6678 ( .A1(n5302), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4780) );
  MUX2_X1 U6679 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n6010), .Z(n6015) );
  NAND4_X1 U6680 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5182), .ZN(n5210)
         );
  NAND2_X1 U6681 ( .A1(n4790), .A2(n5178), .ZN(n5205) );
  NAND2_X1 U6682 ( .A1(n10253), .A2(n4464), .ZN(n4802) );
  OAI211_X2 U6683 ( .C1(n4797), .C2(n4796), .A(n4798), .B(n4794), .ZN(n8271)
         );
  INV_X1 U6684 ( .A(n5401), .ZN(n4795) );
  INV_X1 U6685 ( .A(n10253), .ZN(n4797) );
  NAND2_X1 U6686 ( .A1(n7943), .A2(n5401), .ZN(n8136) );
  NAND2_X1 U6687 ( .A1(n10253), .A2(n5388), .ZN(n7943) );
  INV_X1 U6688 ( .A(n8852), .ZN(n4807) );
  AOI21_X2 U6689 ( .B1(n4807), .B2(n4805), .A(n4804), .ZN(n8787) );
  OR2_X1 U6690 ( .A1(n8778), .A2(n4822), .ZN(n4818) );
  NAND2_X1 U6691 ( .A1(n8778), .A2(n8777), .ZN(n8776) );
  NAND2_X1 U6692 ( .A1(n4815), .A2(n4814), .ZN(n5918) );
  NAND2_X1 U6693 ( .A1(n8778), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U6694 ( .A1(n5458), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U6695 ( .A1(n4824), .A2(n4826), .ZN(n8906) );
  NAND3_X1 U6696 ( .A1(n4828), .A2(n4830), .A3(n4470), .ZN(n4827) );
  NAND2_X1 U6697 ( .A1(n5458), .A2(n5457), .ZN(n7146) );
  INV_X1 U6698 ( .A(n5457), .ZN(n4835) );
  NAND4_X1 U6699 ( .A1(n5140), .A2(n5139), .A3(n4521), .A4(n5182), .ZN(n4836)
         );
  AND2_X2 U6700 ( .A1(n9880), .A2(n9393), .ZN(n9856) );
  OAI21_X2 U6701 ( .B1(n7189), .B2(n6650), .A(n6528), .ZN(n7917) );
  INV_X1 U6702 ( .A(n5305), .ZN(n4844) );
  NAND2_X1 U6703 ( .A1(n5303), .A2(n4845), .ZN(n5305) );
  NAND2_X1 U6704 ( .A1(n5302), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U6705 ( .A1(n8634), .A2(n8649), .ZN(n4848) );
  NAND2_X1 U6706 ( .A1(n7351), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7350) );
  AOI21_X1 U6707 ( .B1(n8288), .B2(n4858), .A(n4531), .ZN(n4857) );
  NAND2_X1 U6708 ( .A1(n8288), .A2(n4853), .ZN(n4852) );
  NAND2_X1 U6709 ( .A1(n4864), .A2(n4862), .ZN(n4860) );
  NAND3_X1 U6710 ( .A1(n4861), .A2(n5958), .A3(n4860), .ZN(n5959) );
  OR2_X2 U6711 ( .A1(n8676), .A2(n8677), .ZN(n4867) );
  NOR2_X2 U6712 ( .A1(n5974), .A2(n4868), .ZN(n8695) );
  NOR2_X1 U6713 ( .A1(n4869), .A2(n8702), .ZN(n4868) );
  NAND2_X1 U6714 ( .A1(n8193), .A2(n4878), .ZN(n8079) );
  INV_X1 U6715 ( .A(n8689), .ZN(n4880) );
  NAND3_X1 U6716 ( .A1(n4883), .A2(n4519), .A3(n4881), .ZN(n8729) );
  OAI211_X1 U6717 ( .C1(n8614), .C2(n4892), .A(n4893), .B(n4888), .ZN(n7311)
         );
  OAI21_X1 U6718 ( .B1(n8256), .B2(n4898), .A(n4896), .ZN(n8299) );
  NAND3_X1 U6719 ( .A1(n4895), .A2(n5999), .A3(n4894), .ZN(n6000) );
  NAND2_X1 U6720 ( .A1(n4896), .A2(n4898), .ZN(n4894) );
  NAND2_X1 U6721 ( .A1(n8256), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U6722 ( .A1(n4900), .A2(n4902), .ZN(n6002) );
  NAND2_X1 U6723 ( .A1(n8635), .A2(n4904), .ZN(n4900) );
  NAND2_X1 U6724 ( .A1(n8635), .A2(n8654), .ZN(n4901) );
  NAND2_X1 U6725 ( .A1(n4906), .A2(n7557), .ZN(n4907) );
  OAI21_X1 U6726 ( .B1(n7961), .B2(n4912), .A(n4909), .ZN(n5994) );
  NAND3_X1 U6727 ( .A1(n4914), .A2(P2_REG2_REG_7__SCAN_IN), .A3(n7957), .ZN(
        n7959) );
  NAND2_X2 U6728 ( .A1(n4915), .A2(n5259), .ZN(n7163) );
  AOI21_X2 U6729 ( .B1(n5257), .B2(n4483), .A(n4916), .ZN(n4915) );
  NAND2_X1 U6730 ( .A1(n5988), .A2(n7168), .ZN(n7557) );
  NAND2_X1 U6731 ( .A1(n7312), .A2(n5985), .ZN(n5988) );
  NAND2_X1 U6732 ( .A1(n5987), .A2(n5986), .ZN(n5989) );
  AND2_X2 U6733 ( .A1(n5957), .A2(n7562), .ZN(n7431) );
  OR2_X1 U6734 ( .A1(n5215), .A2(SI_1_), .ZN(n5274) );
  NAND2_X1 U6735 ( .A1(n5302), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U6736 ( .A1(n9787), .A2(n4922), .ZN(n4920) );
  NAND2_X1 U6737 ( .A1(n9917), .A2(n4935), .ZN(n4934) );
  NAND2_X1 U6738 ( .A1(n9708), .A2(n7051), .ZN(n9691) );
  NAND2_X1 U6739 ( .A1(n4955), .A2(n4953), .ZN(n7045) );
  INV_X1 U6740 ( .A(n4966), .ZN(n7263) );
  INV_X1 U6741 ( .A(n4973), .ZN(n10156) );
  NAND2_X1 U6742 ( .A1(n10176), .A2(n4976), .ZN(n10192) );
  NAND2_X1 U6743 ( .A1(n10192), .A2(n9616), .ZN(n9617) );
  NAND3_X1 U6744 ( .A1(n9637), .A2(n4978), .A3(n4977), .ZN(P1_U3262) );
  NAND2_X1 U6745 ( .A1(n9277), .A2(n4437), .ZN(n4981) );
  OR2_X1 U6746 ( .A1(n9278), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U6747 ( .A1(n7866), .A2(n4996), .ZN(n4994) );
  NAND2_X1 U6748 ( .A1(n9160), .A2(n5004), .ZN(n5001) );
  NAND2_X1 U6749 ( .A1(n5001), .A2(n5002), .ZN(n9136) );
  NAND2_X1 U6750 ( .A1(n6445), .A2(n4446), .ZN(n7785) );
  INV_X1 U6751 ( .A(n6742), .ZN(n5015) );
  AND2_X1 U6752 ( .A1(n6418), .A2(n5016), .ZN(n6357) );
  INV_X1 U6753 ( .A(n6356), .ZN(n5017) );
  NAND2_X1 U6754 ( .A1(n5018), .A2(n9295), .ZN(n9149) );
  AND2_X2 U6755 ( .A1(n9321), .A2(n4507), .ZN(n8334) );
  NAND2_X1 U6756 ( .A1(n6340), .A2(n6341), .ZN(n6337) );
  NOR2_X2 U6757 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8060) );
  NAND2_X1 U6758 ( .A1(n5021), .A2(n5019), .ZN(n5717) );
  NAND2_X1 U6759 ( .A1(n5679), .A2(n5024), .ZN(n5021) );
  NAND2_X1 U6760 ( .A1(n5028), .A2(n5677), .ZN(n5696) );
  NAND2_X1 U6761 ( .A1(n5434), .A2(n5470), .ZN(n5036) );
  NOR2_X2 U6762 ( .A1(n5040), .A2(n5169), .ZN(n6334) );
  NAND2_X1 U6763 ( .A1(n5532), .A2(n4463), .ZN(n5043) );
  INV_X1 U6764 ( .A(n6387), .ZN(n9518) );
  CLKBUF_X1 U6765 ( .A(n6387), .Z(n5048) );
  MUX2_X1 U6766 ( .A(n9598), .B(n7446), .S(n5048), .Z(n7449) );
  AND3_X2 U6767 ( .A1(n5052), .A2(n5051), .A3(n7738), .ZN(n7667) );
  AND3_X2 U6768 ( .A1(n4438), .A2(n9847), .A3(n5053), .ZN(n9760) );
  NOR2_X4 U6769 ( .A1(n5056), .A2(n9731), .ZN(n7101) );
  NAND2_X1 U6770 ( .A1(n5062), .A2(n5335), .ZN(n5336) );
  MUX2_X1 U6771 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n5302), .Z(n5334) );
  NAND2_X1 U6772 ( .A1(n7571), .A2(n5063), .ZN(n5065) );
  NOR2_X1 U6773 ( .A1(n5064), .A2(n7575), .ZN(n5063) );
  INV_X1 U6774 ( .A(n5065), .ZN(n7688) );
  AND2_X2 U6775 ( .A1(n5065), .A2(n7687), .ZN(n7690) );
  NAND2_X1 U6776 ( .A1(n8370), .A2(n5072), .ZN(n5071) );
  NAND2_X1 U6777 ( .A1(n8388), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U6778 ( .A1(n8388), .A2(n5082), .ZN(n5081) );
  NAND2_X1 U6779 ( .A1(n8213), .A2(n5087), .ZN(n5086) );
  NAND2_X1 U6780 ( .A1(n8586), .A2(n5093), .ZN(n8363) );
  NAND2_X1 U6781 ( .A1(n5809), .A2(n5094), .ZN(n5096) );
  NAND2_X2 U6782 ( .A1(n5102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6783 ( .A1(n5818), .A2(n5103), .ZN(n5105) );
  OAI21_X1 U6784 ( .B1(n6130), .B2(n6133), .A(n6145), .ZN(n5104) );
  NAND2_X1 U6785 ( .A1(n6145), .A2(n6133), .ZN(n5106) );
  NAND3_X1 U6786 ( .A1(n5107), .A2(n5108), .A3(n5203), .ZN(n5258) );
  INV_X2 U6787 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5107) );
  NOR2_X1 U6788 ( .A1(n5257), .A2(n5109), .ZN(n5980) );
  NAND2_X1 U6789 ( .A1(n5831), .A2(n5110), .ZN(n8872) );
  OR2_X1 U6790 ( .A1(n6204), .A2(n5111), .ZN(n5113) );
  NAND2_X1 U6791 ( .A1(n8752), .A2(n8753), .ZN(n8751) );
  NAND2_X1 U6792 ( .A1(n8752), .A2(n5121), .ZN(n5120) );
  NOR2_X1 U6793 ( .A1(n5128), .A2(n6172), .ZN(n5130) );
  INV_X1 U6794 ( .A(n5825), .ZN(n5127) );
  NAND2_X1 U6795 ( .A1(n8270), .A2(n5128), .ZN(n5133) );
  NAND2_X1 U6796 ( .A1(n5134), .A2(n5132), .ZN(n5131) );
  NAND3_X1 U6797 ( .A1(n5140), .A2(n5139), .A3(n5182), .ZN(n5862) );
  INV_X2 U6798 ( .A(n5389), .ZN(n5139) );
  INV_X2 U6799 ( .A(n5205), .ZN(n5140) );
  NAND2_X1 U6800 ( .A1(n9696), .A2(n4511), .ZN(n5144) );
  NAND2_X1 U6801 ( .A1(n9696), .A2(n5157), .ZN(n5148) );
  OAI211_X1 U6802 ( .C1(n9696), .C2(n5146), .A(n5144), .B(n5141), .ZN(n9648)
         );
  NAND3_X1 U6803 ( .A1(n5162), .A2(n9528), .A3(n7743), .ZN(n5160) );
  NAND2_X1 U6804 ( .A1(n7057), .A2(n9528), .ZN(n5161) );
  NAND2_X1 U6805 ( .A1(n7626), .A2(n9529), .ZN(n9343) );
  NAND2_X1 U6806 ( .A1(n5160), .A2(n5159), .ZN(n7626) );
  NAND2_X1 U6807 ( .A1(n7139), .A2(n5194), .ZN(n5166) );
  NAND2_X1 U6808 ( .A1(n5166), .A2(n5163), .ZN(P1_U3551) );
  NOR2_X1 U6809 ( .A1(n7139), .A2(n7138), .ZN(n7145) );
  NAND2_X2 U6810 ( .A1(n9537), .A2(n9533), .ZN(n7059) );
  NAND2_X1 U6811 ( .A1(n7115), .A2(n10243), .ZN(n7095) );
  NAND2_X1 U6812 ( .A1(n8948), .A2(n10672), .ZN(n8950) );
  NAND2_X1 U6813 ( .A1(n9942), .A2(n9941), .ZN(n10068) );
  NAND2_X1 U6814 ( .A1(n10068), .A2(n10252), .ZN(n9943) );
  INV_X1 U6815 ( .A(n6427), .ZN(n6512) );
  INV_X1 U6816 ( .A(n6483), .ZN(n6486) );
  AND2_X1 U6817 ( .A1(n7390), .A2(n8609), .ZN(n7391) );
  INV_X1 U6818 ( .A(n8609), .ZN(n5244) );
  NAND2_X1 U6819 ( .A1(n9761), .A2(n9977), .ZN(n9744) );
  AND2_X2 U6820 ( .A1(n9760), .A2(n9985), .ZN(n9761) );
  AOI21_X1 U6821 ( .B1(n9321), .B2(n6958), .A(n6957), .ZN(n6978) );
  XNOR2_X1 U6822 ( .A(n5923), .B(n8395), .ZN(n8954) );
  OAI21_X2 U6823 ( .B1(n5634), .B2(n5633), .A(n5632), .ZN(n5646) );
  NAND2_X1 U6824 ( .A1(n6947), .A2(n6379), .ZN(n6380) );
  AND2_X1 U6825 ( .A1(n8742), .A2(n10317), .ZN(n5855) );
  NAND2_X1 U6826 ( .A1(n6319), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n6320) );
  INV_X2 U6827 ( .A(n10337), .ZN(n10336) );
  INV_X1 U6828 ( .A(n10672), .ZN(n8960) );
  NAND2_X1 U6829 ( .A1(n6271), .A2(n6240), .ZN(n5171) );
  OR2_X1 U6830 ( .A1(n10067), .A2(n10032), .ZN(n5173) );
  AND2_X1 U6831 ( .A1(n7094), .A2(n5196), .ZN(n5174) );
  OR2_X1 U6832 ( .A1(n8992), .A2(n8883), .ZN(n5176) );
  AND2_X1 U6833 ( .A1(n9652), .A2(n7130), .ZN(n5177) );
  AND3_X1 U6834 ( .A1(n5407), .A2(n5200), .A3(n5199), .ZN(n5178) );
  OR2_X1 U6835 ( .A1(n10072), .A2(n9335), .ZN(n5179) );
  INV_X1 U6836 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6341) );
  AND4_X1 U6837 ( .A1(n5856), .A2(n5208), .A3(n5207), .A4(n5206), .ZN(n5182)
         );
  OR2_X1 U6838 ( .A1(n8497), .A2(n8908), .ZN(n5183) );
  OR2_X1 U6839 ( .A1(n9079), .A2(n9078), .ZN(P2_U3438) );
  OR2_X1 U6840 ( .A1(n8997), .A2(n8996), .ZN(P2_U3475) );
  OR2_X1 U6841 ( .A1(n8905), .A2(n8904), .ZN(P2_U3217) );
  AND2_X1 U6842 ( .A1(n8766), .A2(n6220), .ZN(n5187) );
  NAND2_X1 U6843 ( .A1(n9486), .A2(n9431), .ZN(n9709) );
  AND2_X1 U6844 ( .A1(n8226), .A2(n8605), .ZN(n5189) );
  AND3_X1 U6845 ( .A1(n6137), .A2(n6256), .A3(n10258), .ZN(n5190) );
  INV_X1 U6846 ( .A(n9140), .ZN(n6867) );
  NOR2_X1 U6847 ( .A1(n8523), .A2(n8524), .ZN(n5191) );
  AND2_X1 U6848 ( .A1(n6235), .A2(n6241), .ZN(n5192) );
  OR2_X1 U6849 ( .A1(n10252), .A2(n10534), .ZN(n5193) );
  OR2_X1 U6850 ( .A1(n10252), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5194) );
  AND2_X1 U6851 ( .A1(n7649), .A2(n10215), .ZN(n10211) );
  INV_X1 U6852 ( .A(n10211), .ZN(n10241) );
  INV_X1 U6853 ( .A(n9933), .ZN(n9854) );
  AND2_X1 U6854 ( .A1(n7595), .A2(n9891), .ZN(n9933) );
  OR2_X1 U6855 ( .A1(n9659), .A2(n10032), .ZN(n5195) );
  OR2_X1 U6856 ( .A1(n10243), .A2(n10393), .ZN(n5196) );
  AND2_X2 U6857 ( .A1(n7112), .A2(n7111), .ZN(n10252) );
  INV_X1 U6858 ( .A(n10090), .ZN(n7093) );
  AND2_X1 U6859 ( .A1(n6123), .A2(n6237), .ZN(n6124) );
  AOI21_X1 U6860 ( .B1(n6125), .B2(n6241), .A(n6124), .ZN(n6126) );
  AND2_X1 U6861 ( .A1(n10258), .A2(n6147), .ZN(n6148) );
  INV_X1 U6862 ( .A(n9449), .ZN(n9342) );
  NAND2_X1 U6863 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  OAI21_X1 U6864 ( .B1(n9358), .B2(n9357), .A(n9356), .ZN(n9361) );
  NAND2_X1 U6865 ( .A1(n9386), .A2(n9385), .ZN(n9390) );
  NAND2_X1 U6866 ( .A1(n6219), .A2(n6241), .ZN(n6220) );
  INV_X1 U6867 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5201) );
  NOR2_X1 U6868 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n6311) );
  INV_X1 U6869 ( .A(n7788), .ZN(n6457) );
  INV_X1 U6870 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6314) );
  INV_X1 U6871 ( .A(n9034), .ZN(n5732) );
  INV_X1 U6872 ( .A(n9614), .ZN(n9615) );
  INV_X1 U6873 ( .A(n9783), .ZN(n7068) );
  INV_X1 U6874 ( .A(n8532), .ZN(n8355) );
  XNOR2_X1 U6875 ( .A(n7520), .B(n7409), .ZN(n7390) );
  NAND2_X1 U6876 ( .A1(n5226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5209) );
  AND2_X1 U6877 ( .A1(n5676), .A2(n8813), .ZN(n8801) );
  INV_X1 U6878 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6879 ( .A1(n5894), .A2(n7237), .ZN(n7383) );
  NAND2_X1 U6880 ( .A1(n5732), .A2(n8578), .ZN(n5733) );
  INV_X1 U6881 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6583) );
  INV_X1 U6882 ( .A(n9709), .ZN(n7070) );
  NAND2_X1 U6883 ( .A1(n7914), .A2(n9591), .ZN(n9351) );
  INV_X1 U6884 ( .A(n5552), .ZN(n5572) );
  AND2_X1 U6885 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  AND2_X1 U6886 ( .A1(n5324), .A2(n5330), .ZN(n5325) );
  OR2_X1 U6887 ( .A1(n5302), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5303) );
  OR2_X1 U6888 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  INV_X1 U6889 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10485) );
  INV_X1 U6890 ( .A(n7713), .ZN(n5814) );
  OR2_X1 U6891 ( .A1(n6241), .A2(n5839), .ZN(n7419) );
  NOR2_X1 U6892 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  AND2_X1 U6893 ( .A1(n8097), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8087) );
  OR2_X1 U6894 ( .A1(n10172), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9623) );
  OAI21_X2 U6895 ( .B1(n6075), .B2(n10613), .A(n6074), .ZN(n6099) );
  AND2_X1 U6896 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U6897 ( .A1(n8365), .A2(n8894), .ZN(n8366) );
  INV_X1 U6898 ( .A(n8601), .ZN(n8883) );
  INV_X1 U6899 ( .A(n10286), .ZN(n10256) );
  OR2_X1 U6900 ( .A1(n5930), .A2(n7383), .ZN(n5904) );
  AND2_X1 U6901 ( .A1(n5905), .A2(n7386), .ZN(n8853) );
  OR2_X1 U6902 ( .A1(n7151), .A2(n7150), .ZN(n9014) );
  AND2_X1 U6903 ( .A1(n6136), .A2(n8130), .ZN(n7944) );
  NAND2_X1 U6904 ( .A1(n7373), .A2(n7241), .ZN(n6297) );
  OR2_X1 U6905 ( .A1(n9699), .A2(n6465), .ZN(n6920) );
  OR2_X1 U6906 ( .A1(n6512), .A2(n6328), .ZN(n6329) );
  AND2_X1 U6907 ( .A1(n9410), .A2(n9409), .ZN(n9820) );
  AND2_X1 U6908 ( .A1(n5697), .A2(n5683), .ZN(n5695) );
  INV_X1 U6909 ( .A(n5340), .ZN(n5337) );
  INV_X1 U6910 ( .A(n5326), .ZN(n5282) );
  NAND2_X1 U6911 ( .A1(n7382), .A2(n7381), .ZN(n8594) );
  AND2_X1 U6912 ( .A1(n6094), .A2(n5804), .ZN(n8398) );
  NAND2_X1 U6913 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  INV_X1 U6914 ( .A(n8717), .ZN(n8632) );
  INV_X1 U6915 ( .A(n8655), .ZN(n8730) );
  OR2_X1 U6916 ( .A1(n8133), .A2(n8137), .ZN(n8234) );
  OR2_X1 U6917 ( .A1(n6297), .A2(n5935), .ZN(n8912) );
  INV_X1 U6918 ( .A(n9018), .ZN(n9007) );
  AND2_X1 U6919 ( .A1(n5895), .A2(n5904), .ZN(n5933) );
  NAND2_X1 U6920 ( .A1(n6196), .A2(n6195), .ZN(n8843) );
  INV_X1 U6921 ( .A(n10330), .ZN(n10316) );
  OR2_X1 U6922 ( .A1(n7902), .A2(n10317), .ZN(n10327) );
  INV_X1 U6923 ( .A(n5619), .ZN(n5598) );
  AND2_X1 U6924 ( .A1(n8322), .A2(n9320), .ZN(n8323) );
  INV_X1 U6925 ( .A(n9335), .ZN(n9272) );
  OR2_X1 U6926 ( .A1(n6994), .A2(n6993), .ZN(n9338) );
  INV_X1 U6927 ( .A(n7854), .ZN(n7769) );
  OR2_X1 U6928 ( .A1(n10127), .A2(n7215), .ZN(n10164) );
  INV_X1 U6929 ( .A(n10202), .ZN(n10183) );
  AND2_X1 U6930 ( .A1(n9403), .A2(n9401), .ZN(n9789) );
  NAND2_X1 U6931 ( .A1(n6999), .A2(n10099), .ZN(n9891) );
  NAND2_X1 U6932 ( .A1(n9943), .A2(n5193), .ZN(n9944) );
  INV_X1 U6933 ( .A(n7637), .ZN(n7781) );
  AND2_X1 U6934 ( .A1(n7072), .A2(n9447), .ZN(n10210) );
  AND2_X1 U6935 ( .A1(n5181), .A2(n7003), .ZN(n10049) );
  INV_X1 U6936 ( .A(n10210), .ZN(n9988) );
  INV_X1 U6937 ( .A(n10057), .ZN(n10212) );
  AND2_X1 U6938 ( .A1(n7185), .A2(n6976), .ZN(n10099) );
  INV_X1 U6939 ( .A(n9451), .ZN(n7993) );
  INV_X1 U6940 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6719) );
  INV_X1 U6941 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6474) );
  AND2_X1 U6942 ( .A1(n7398), .A2(n7397), .ZN(n8570) );
  INV_X1 U6943 ( .A(n8493), .ZN(n8807) );
  INV_X1 U6944 ( .A(n8893), .ZN(n8921) );
  INV_X1 U6945 ( .A(n10255), .ZN(n8606) );
  INV_X1 U6946 ( .A(n8704), .ZN(n8722) );
  NAND2_X1 U6947 ( .A1(n10282), .A2(n5937), .ZN(n8941) );
  INV_X1 U6948 ( .A(n5901), .ZN(n5902) );
  XNOR2_X1 U6949 ( .A(n8775), .B(n4821), .ZN(n9037) );
  NAND2_X1 U6950 ( .A1(n10336), .A2(n10327), .ZN(n9096) );
  AND2_X1 U6951 ( .A1(n5913), .A2(n5912), .ZN(n10337) );
  AND2_X1 U6952 ( .A1(n7372), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7241) );
  INV_X1 U6953 ( .A(n6301), .ZN(n8179) );
  INV_X1 U6954 ( .A(n6028), .ZN(n7763) );
  AND2_X1 U6955 ( .A1(n7212), .A2(n7187), .ZN(n10169) );
  INV_X1 U6956 ( .A(n4611), .ZN(n9977) );
  INV_X1 U6957 ( .A(n9338), .ZN(n9303) );
  INV_X1 U6958 ( .A(n9763), .ZN(n9985) );
  AND2_X1 U6959 ( .A1(n7000), .A2(n9891), .ZN(n9335) );
  INV_X1 U6960 ( .A(n9792), .ZN(n9982) );
  INV_X1 U6961 ( .A(n9912), .ZN(n9588) );
  INV_X1 U6962 ( .A(n10169), .ZN(n10207) );
  INV_X1 U6963 ( .A(n9928), .ZN(n9909) );
  INV_X1 U6964 ( .A(n10243), .ZN(n7144) );
  INV_X1 U6965 ( .A(n10208), .ZN(n10209) );
  INV_X1 U6966 ( .A(n8718), .ZN(P2_U3893) );
  NAND2_X1 U6967 ( .A1(n5927), .A2(n5926), .ZN(P2_U3455) );
  AND2_X1 U6968 ( .A1(n7185), .A2(n7157), .ZN(P1_U3973) );
  OAI21_X1 U6969 ( .B1(n4414), .B2(n4409), .A(n7117), .ZN(P1_U3550) );
  NAND2_X1 U6970 ( .A1(n7095), .A2(n5174), .ZN(P1_U3518) );
  INV_X2 U6971 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5320) );
  INV_X1 U6972 ( .A(n5258), .ZN(n5204) );
  NAND2_X1 U6973 ( .A1(n4476), .A2(n5204), .ZN(n5389) );
  NOR2_X1 U6974 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5208) );
  NOR2_X1 U6975 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5207) );
  NOR2_X1 U6976 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5206) );
  NAND2_X1 U6977 ( .A1(n5210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5212) );
  XNOR2_X2 U6978 ( .A(n5212), .B(n5211), .ZN(n5842) );
  NAND2_X1 U6979 ( .A1(n5243), .A2(n7161), .ZN(n5286) );
  NAND2_X1 U6980 ( .A1(n5215), .A2(SI_1_), .ZN(n5271) );
  AND2_X1 U6981 ( .A1(n5271), .A2(n5274), .ZN(n5218) );
  NAND2_X1 U6982 ( .A1(n5218), .A2(n5273), .ZN(n5251) );
  INV_X1 U6983 ( .A(n5218), .ZN(n5219) );
  NAND2_X1 U6984 ( .A1(n5219), .A2(n5217), .ZN(n5220) );
  AND2_X1 U6985 ( .A1(n5251), .A2(n5220), .ZN(n6394) );
  OR2_X1 U6986 ( .A1(n4425), .A2(n6394), .ZN(n5225) );
  NAND2_X1 U6987 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5221) );
  NAND2_X1 U6988 ( .A1(n5621), .A2(n5946), .ZN(n5223) );
  INV_X1 U6989 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5231) );
  AND2_X4 U6990 ( .A1(n8408), .A2(n9108), .ZN(n6086) );
  NAND2_X1 U6991 ( .A1(n6086), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5230) );
  INV_X1 U6992 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7716) );
  OR2_X1 U6993 ( .A1(n5292), .A2(n7716), .ZN(n5235) );
  INV_X1 U6994 ( .A(n7409), .ZN(n10297) );
  INV_X1 U6995 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U6996 ( .A1(n6086), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5240) );
  INV_X1 U6997 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7415) );
  OR2_X1 U6998 ( .A1(n5292), .A2(n7415), .ZN(n5239) );
  OR2_X1 U6999 ( .A1(n5291), .A2(n5109), .ZN(n5238) );
  NAND4_X2 U7000 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n6109)
         );
  NAND2_X1 U7001 ( .A1(n7161), .A2(SI_0_), .ZN(n5242) );
  XNOR2_X1 U7002 ( .A(n5242), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9125) );
  MUX2_X1 U7003 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9125), .S(n5243), .Z(n7392) );
  NAND2_X1 U7004 ( .A1(n6109), .A2(n7392), .ZN(n7717) );
  NAND2_X1 U7005 ( .A1(n6250), .A2(n7717), .ZN(n5246) );
  NAND2_X1 U7006 ( .A1(n5244), .A2(n10297), .ZN(n5245) );
  NAND2_X1 U7007 ( .A1(n5246), .A2(n5245), .ZN(n7616) );
  OR2_X1 U7008 ( .A1(n4424), .A2(n10338), .ZN(n5250) );
  INV_X1 U7009 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7621) );
  OR2_X1 U7010 ( .A1(n5292), .A2(n7621), .ZN(n5249) );
  INV_X1 U7011 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7624) );
  OR2_X1 U7012 ( .A1(n5291), .A2(n7624), .ZN(n5248) );
  NAND2_X1 U7013 ( .A1(n6086), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U7014 ( .A1(n5251), .A2(n5271), .ZN(n5256) );
  INV_X1 U7015 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7173) );
  INV_X1 U7016 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7164) );
  INV_X1 U7017 ( .A(SI_2_), .ZN(n5252) );
  INV_X1 U7018 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U7019 ( .A1(n5254), .A2(SI_2_), .ZN(n5276) );
  AND2_X1 U7020 ( .A1(n5275), .A2(n5276), .ZN(n5255) );
  XNOR2_X1 U7021 ( .A(n5256), .B(n5255), .ZN(n7174) );
  OR2_X1 U7022 ( .A1(n5286), .A2(n7174), .ZN(n5262) );
  OR2_X1 U7023 ( .A1(n6104), .A2(n7164), .ZN(n5261) );
  INV_X1 U7024 ( .A(n7163), .ZN(n8619) );
  NAND2_X1 U7025 ( .A1(n4407), .A2(n8619), .ZN(n5260) );
  XNOR2_X1 U7026 ( .A(n10287), .B(n10302), .ZN(n7615) );
  NAND2_X1 U7027 ( .A1(n7616), .A2(n7615), .ZN(n5264) );
  NAND2_X1 U7028 ( .A1(n7528), .A2(n10302), .ZN(n5263) );
  NAND2_X1 U7029 ( .A1(n5264), .A2(n5263), .ZN(n10283) );
  OR2_X1 U7030 ( .A1(n5292), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U7031 ( .A1(n6086), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5267) );
  OR2_X1 U7032 ( .A1(n5291), .A2(n4889), .ZN(n5266) );
  INV_X1 U7033 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10340) );
  OR2_X1 U7034 ( .A1(n4424), .A2(n10340), .ZN(n5265) );
  NAND2_X1 U7035 ( .A1(n5259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5269) );
  MUX2_X1 U7036 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5269), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5270) );
  INV_X1 U7037 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7165) );
  OR2_X1 U7038 ( .A1(n4405), .A2(n7165), .ZN(n5288) );
  INV_X1 U7039 ( .A(n5271), .ZN(n5272) );
  INV_X1 U7040 ( .A(n5279), .ZN(n5281) );
  INV_X1 U7041 ( .A(SI_3_), .ZN(n5280) );
  NAND2_X1 U7042 ( .A1(n5281), .A2(n5280), .ZN(n5324) );
  NAND2_X1 U7043 ( .A1(n5327), .A2(n5324), .ZN(n5283) );
  NAND2_X1 U7044 ( .A1(n5282), .A2(n5283), .ZN(n5285) );
  INV_X1 U7045 ( .A(n5283), .ZN(n5284) );
  NAND2_X1 U7046 ( .A1(n5326), .A2(n5284), .ZN(n5301) );
  NAND2_X1 U7047 ( .A1(n5285), .A2(n5301), .ZN(n7170) );
  OR2_X1 U7048 ( .A1(n4425), .A2(n7170), .ZN(n5287) );
  OAI211_X1 U7049 ( .C1(n5243), .C2(n7166), .A(n5288), .B(n5287), .ZN(n6121)
         );
  NOR2_X1 U7050 ( .A1(n10276), .A2(n6121), .ZN(n5290) );
  NAND2_X1 U7051 ( .A1(n10276), .A2(n6121), .ZN(n5289) );
  NAND2_X1 U7052 ( .A1(n5845), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U7053 ( .A1(n5844), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U7054 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5294) );
  AND2_X1 U7055 ( .A1(n5313), .A2(n5294), .ZN(n7577) );
  OR2_X1 U7056 ( .A1(n5292), .A2(n7577), .ZN(n5297) );
  INV_X1 U7057 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5295) );
  OR2_X1 U7058 ( .A1(n5848), .A2(n5295), .ZN(n5296) );
  NAND2_X1 U7059 ( .A1(n5319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5300) );
  XNOR2_X2 U7060 ( .A(n5300), .B(n5320), .ZN(n7325) );
  OR2_X1 U7061 ( .A1(n6104), .A2(n4846), .ZN(n5309) );
  NAND2_X1 U7062 ( .A1(n5301), .A2(n5327), .ZN(n5307) );
  INV_X1 U7063 ( .A(SI_4_), .ZN(n5304) );
  NAND2_X1 U7064 ( .A1(n5305), .A2(n5304), .ZN(n5330) );
  AND2_X1 U7065 ( .A1(n5330), .A2(n5328), .ZN(n5306) );
  XNOR2_X1 U7066 ( .A(n5307), .B(n5306), .ZN(n7175) );
  OR2_X1 U7067 ( .A1(n5286), .A2(n7175), .ZN(n5308) );
  OAI211_X1 U7068 ( .C1(n5243), .C2(n7325), .A(n5309), .B(n5308), .ZN(n10311)
         );
  AND2_X1 U7069 ( .A1(n10285), .A2(n10311), .ZN(n5311) );
  NAND2_X1 U7070 ( .A1(n7894), .A2(n7573), .ZN(n5310) );
  OAI21_X1 U7071 ( .B1(n10274), .B2(n5311), .A(n5310), .ZN(n7898) );
  NAND2_X1 U7072 ( .A1(n5844), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U7073 ( .A1(n6086), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5317) );
  OR2_X1 U7074 ( .A1(n4424), .A2(n4863), .ZN(n5316) );
  NAND2_X1 U7075 ( .A1(n5313), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5314) );
  AND2_X1 U7076 ( .A1(n5344), .A2(n5314), .ZN(n7691) );
  OR2_X1 U7077 ( .A1(n5292), .A2(n7691), .ZN(n5315) );
  NAND4_X1 U7078 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n10275)
         );
  INV_X1 U7079 ( .A(n5319), .ZN(n5321) );
  NAND2_X1 U7080 ( .A1(n5321), .A2(n5320), .ZN(n5350) );
  NAND2_X1 U7081 ( .A1(n5350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5323) );
  XNOR2_X1 U7082 ( .A(n5323), .B(n5322), .ZN(n7168) );
  INV_X1 U7083 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7167) );
  OR2_X1 U7084 ( .A1(n4405), .A2(n7167), .ZN(n5343) );
  INV_X1 U7085 ( .A(n5327), .ZN(n5331) );
  INV_X1 U7086 ( .A(n5328), .ZN(n5329) );
  AOI21_X1 U7087 ( .B1(n5331), .B2(n5330), .A(n5329), .ZN(n5332) );
  INV_X1 U7088 ( .A(SI_5_), .ZN(n5335) );
  NAND2_X1 U7089 ( .A1(n5352), .A2(n5336), .ZN(n5338) );
  NAND2_X1 U7090 ( .A1(n5337), .A2(n5338), .ZN(n5341) );
  INV_X1 U7091 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U7092 ( .A1(n5340), .A2(n5339), .ZN(n5353) );
  NAND2_X1 U7093 ( .A1(n5341), .A2(n5353), .ZN(n7172) );
  OR2_X1 U7094 ( .A1(n5286), .A2(n7172), .ZN(n5342) );
  OAI211_X1 U7095 ( .C1(n5243), .C2(n7168), .A(n5343), .B(n5342), .ZN(n10315)
         );
  INV_X1 U7096 ( .A(n10315), .ZN(n5819) );
  NAND2_X1 U7097 ( .A1(n7930), .A2(n5819), .ZN(n7895) );
  NAND2_X1 U7098 ( .A1(n6086), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5349) );
  INV_X1 U7099 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10546) );
  OR2_X1 U7100 ( .A1(n4424), .A2(n10546), .ZN(n5348) );
  NAND2_X1 U7101 ( .A1(n5344), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5345) );
  AND2_X1 U7102 ( .A1(n5369), .A2(n5345), .ZN(n7935) );
  OR2_X1 U7103 ( .A1(n5292), .A2(n7935), .ZN(n5347) );
  INV_X1 U7104 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7934) );
  OR2_X1 U7105 ( .A1(n6091), .A2(n7934), .ZN(n5346) );
  NAND2_X1 U7106 ( .A1(n5384), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5351) );
  AOI22_X1 U7107 ( .A1(n5622), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4407), .B2(
        n7179), .ZN(n5362) );
  NAND2_X1 U7108 ( .A1(n5353), .A2(n5352), .ZN(n5359) );
  MUX2_X1 U7109 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6393), .Z(n5354) );
  INV_X1 U7110 ( .A(n5354), .ZN(n5356) );
  INV_X1 U7111 ( .A(SI_6_), .ZN(n5355) );
  NAND2_X1 U7112 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U7113 ( .A1(n5359), .A2(n5358), .ZN(n5376) );
  OR2_X1 U7114 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  AND2_X1 U7115 ( .A1(n5376), .A2(n5360), .ZN(n7177) );
  NAND2_X1 U7116 ( .A1(n7177), .A2(n6106), .ZN(n5361) );
  NAND2_X1 U7117 ( .A1(n5362), .A2(n5361), .ZN(n7937) );
  NAND2_X1 U7118 ( .A1(n10257), .A2(n10324), .ZN(n7928) );
  NAND2_X1 U7119 ( .A1(n7895), .A2(n7928), .ZN(n5366) );
  NAND2_X1 U7120 ( .A1(n10275), .A2(n10315), .ZN(n7923) );
  NAND2_X1 U7121 ( .A1(n7923), .A2(n10257), .ZN(n5364) );
  AND2_X1 U7122 ( .A1(n8608), .A2(n10315), .ZN(n5363) );
  AOI22_X1 U7123 ( .A1(n5364), .A2(n7937), .B1(n5363), .B2(n10275), .ZN(n5365)
         );
  NAND2_X1 U7124 ( .A1(n6086), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5374) );
  INV_X1 U7125 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10273) );
  OR2_X1 U7126 ( .A1(n6091), .A2(n10273), .ZN(n5373) );
  INV_X1 U7127 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10345) );
  OR2_X1 U7128 ( .A1(n4424), .A2(n10345), .ZN(n5372) );
  NAND2_X1 U7129 ( .A1(n5369), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5370) );
  AND2_X1 U7130 ( .A1(n5394), .A2(n5370), .ZN(n10266) );
  OR2_X1 U7131 ( .A1(n5292), .A2(n10266), .ZN(n5371) );
  MUX2_X1 U7132 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6393), .Z(n5377) );
  INV_X1 U7133 ( .A(n5377), .ZN(n5379) );
  INV_X1 U7134 ( .A(SI_7_), .ZN(n5378) );
  NAND2_X1 U7135 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND2_X2 U7136 ( .A1(n5382), .A2(n5381), .ZN(n5428) );
  OR2_X1 U7137 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  OR2_X1 U7138 ( .A1(n7189), .A2(n4425), .ZN(n5387) );
  OAI21_X1 U7139 ( .B1(n5384), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5385) );
  XNOR2_X1 U7140 ( .A(n5385), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6028) );
  AOI22_X1 U7141 ( .A1(n5622), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4407), .B2(
        n6028), .ZN(n5386) );
  AND2_X2 U7142 ( .A1(n5387), .A2(n5386), .ZN(n10331) );
  NAND2_X1 U7143 ( .A1(n8171), .A2(n10331), .ZN(n5388) );
  NAND2_X1 U7144 ( .A1(n10268), .A2(n8607), .ZN(n7942) );
  INV_X1 U7145 ( .A(n7942), .ZN(n5400) );
  XNOR2_X1 U7146 ( .A(n5421), .B(SI_8_), .ZN(n5404) );
  NAND2_X1 U7147 ( .A1(n7190), .A2(n6106), .ZN(n5392) );
  NAND2_X1 U7148 ( .A1(n5389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U7149 ( .A(n5390), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7964) );
  AOI22_X1 U7150 ( .A1(n5622), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4407), .B2(
        n7964), .ZN(n5391) );
  NAND2_X1 U7151 ( .A1(n5392), .A2(n5391), .ZN(n8163) );
  NAND2_X1 U7152 ( .A1(n5844), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5399) );
  INV_X1 U7153 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5393) );
  OR2_X1 U7154 ( .A1(n4424), .A2(n5393), .ZN(n5398) );
  NAND2_X1 U7155 ( .A1(n5394), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5395) );
  AND2_X1 U7156 ( .A1(n5412), .A2(n5395), .ZN(n8182) );
  OR2_X1 U7157 ( .A1(n5292), .A2(n8182), .ZN(n5397) );
  INV_X1 U7158 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7950) );
  OR2_X1 U7159 ( .A1(n5848), .A2(n7950), .ZN(n5396) );
  OR2_X1 U7160 ( .A1(n8163), .A2(n10255), .ZN(n6136) );
  NAND2_X1 U7161 ( .A1(n8163), .A2(n10255), .ZN(n8130) );
  NOR2_X1 U7162 ( .A1(n5400), .A2(n7944), .ZN(n5401) );
  OR2_X1 U7163 ( .A1(n8163), .A2(n8606), .ZN(n8135) );
  MUX2_X1 U7164 ( .A(n7229), .B(n7204), .S(n6393), .Z(n5430) );
  NAND2_X1 U7165 ( .A1(n5139), .A2(n5407), .ZN(n5561) );
  NAND2_X1 U7166 ( .A1(n5561), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5408) );
  MUX2_X1 U7167 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5408), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5409) );
  AND2_X1 U7168 ( .A1(n5409), .A2(n5446), .ZN(n8083) );
  AOI22_X1 U7169 ( .A1(n5622), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4407), .B2(
        n8083), .ZN(n5410) );
  NAND2_X1 U7170 ( .A1(n5845), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7171 ( .A1(n6086), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5416) );
  INV_X1 U7172 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10577) );
  OR2_X1 U7173 ( .A1(n6091), .A2(n10577), .ZN(n5415) );
  NAND2_X1 U7174 ( .A1(n5412), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5413) );
  AND2_X1 U7175 ( .A1(n5439), .A2(n5413), .ZN(n8216) );
  OR2_X1 U7176 ( .A1(n5292), .A2(n8216), .ZN(n5414) );
  NAND4_X1 U7177 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n8605)
         );
  OR2_X1 U7178 ( .A1(n8226), .A2(n8605), .ZN(n5418) );
  AND2_X1 U7179 ( .A1(n8135), .A2(n5418), .ZN(n5419) );
  INV_X1 U7180 ( .A(n5422), .ZN(n5427) );
  INV_X1 U7181 ( .A(n5420), .ZN(n5423) );
  AOI22_X1 U7182 ( .A1(n5423), .A2(n5422), .B1(SI_8_), .B2(n5421), .ZN(n5425)
         );
  INV_X1 U7183 ( .A(SI_9_), .ZN(n5429) );
  MUX2_X1 U7184 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6393), .Z(n5431) );
  INV_X1 U7185 ( .A(n5433), .ZN(n5432) );
  NAND2_X1 U7186 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  NAND2_X1 U7187 ( .A1(n5471), .A2(n5435), .ZN(n7196) );
  OR2_X1 U7188 ( .A1(n7196), .A2(n5286), .ZN(n5438) );
  NAND2_X1 U7189 ( .A1(n5446), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U7190 ( .A(n5436), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8200) );
  AOI22_X1 U7191 ( .A1(n5622), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4407), .B2(
        n8200), .ZN(n5437) );
  NAND2_X1 U7192 ( .A1(n5844), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U7193 ( .A1(n5845), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7194 ( .A1(n5439), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5440) );
  AND2_X1 U7195 ( .A1(n5451), .A2(n5440), .ZN(n8442) );
  OR2_X1 U7196 ( .A1(n5292), .A2(n8442), .ZN(n5443) );
  INV_X1 U7197 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5441) );
  OR2_X1 U7198 ( .A1(n5848), .A2(n5441), .ZN(n5442) );
  NAND4_X1 U7199 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n8604)
         );
  MUX2_X1 U7200 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6393), .Z(n5467) );
  XNOR2_X1 U7201 ( .A(n5467), .B(SI_11_), .ZN(n5461) );
  NAND2_X1 U7202 ( .A1(n7231), .A2(n6106), .ZN(n5450) );
  INV_X1 U7203 ( .A(n5446), .ZN(n5448) );
  INV_X1 U7204 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7205 ( .A1(n5448), .A2(n5447), .ZN(n5503) );
  NAND2_X1 U7206 ( .A1(n5503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5477) );
  XNOR2_X1 U7207 ( .A(n5477), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6035) );
  AOI22_X1 U7208 ( .A1(n5622), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4407), .B2(
        n6035), .ZN(n5449) );
  NAND2_X2 U7209 ( .A1(n5450), .A2(n5449), .ZN(n8548) );
  NAND2_X1 U7210 ( .A1(n5845), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5456) );
  INV_X1 U7211 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10488) );
  OR2_X1 U7212 ( .A1(n6091), .A2(n10488), .ZN(n5455) );
  NAND2_X1 U7213 ( .A1(n5451), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5452) );
  AND2_X1 U7214 ( .A1(n5483), .A2(n5452), .ZN(n8281) );
  OR2_X1 U7215 ( .A1(n5292), .A2(n8281), .ZN(n5454) );
  INV_X1 U7216 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8275) );
  OR2_X1 U7217 ( .A1(n5848), .A2(n8275), .ZN(n5453) );
  NAND2_X1 U7218 ( .A1(n8548), .A2(n8473), .ZN(n6156) );
  NAND2_X1 U7219 ( .A1(n8548), .A2(n8603), .ZN(n5457) );
  INV_X1 U7220 ( .A(n5467), .ZN(n5460) );
  INV_X1 U7221 ( .A(SI_11_), .ZN(n5459) );
  OAI21_X1 U7222 ( .B1(n5462), .B2(n5461), .A(n5472), .ZN(n5466) );
  MUX2_X1 U7223 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6393), .Z(n5463) );
  INV_X1 U7224 ( .A(n5463), .ZN(n5464) );
  INV_X1 U7225 ( .A(SI_12_), .ZN(n10492) );
  NAND2_X1 U7226 ( .A1(n5464), .A2(n10492), .ZN(n5465) );
  NAND2_X1 U7227 ( .A1(n5466), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U7228 ( .A1(n5467), .A2(SI_11_), .ZN(n5469) );
  INV_X1 U7229 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7230 ( .A1(n5477), .A2(n5501), .ZN(n5478) );
  NAND2_X1 U7231 ( .A1(n5478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U7232 ( .A(n5479), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8294) );
  AOI22_X1 U7233 ( .A1(n5622), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4407), .B2(
        n8294), .ZN(n5480) );
  NAND2_X1 U7234 ( .A1(n5845), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7235 ( .A1(n6086), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7236 ( .A1(n5483), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5484) );
  AND2_X1 U7237 ( .A1(n5509), .A2(n5484), .ZN(n8480) );
  OR2_X1 U7238 ( .A1(n5292), .A2(n8480), .ZN(n5486) );
  INV_X1 U7239 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7240 ( .A1(n6091), .A2(n5998), .ZN(n5485) );
  NAND4_X1 U7241 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n8931)
         );
  AND2_X1 U7242 ( .A1(n8482), .A2(n8931), .ZN(n5490) );
  MUX2_X1 U7243 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6393), .Z(n5493) );
  INV_X1 U7244 ( .A(n5493), .ZN(n5495) );
  INV_X1 U7245 ( .A(SI_13_), .ZN(n5494) );
  NAND2_X1 U7246 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  INV_X1 U7247 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7248 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  OR2_X1 U7249 ( .A1(n5503), .A2(n5502), .ZN(n5518) );
  NAND2_X1 U7250 ( .A1(n5518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5504) );
  XNOR2_X1 U7251 ( .A(n5504), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8633) );
  AOI22_X1 U7252 ( .A1(n5622), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4407), .B2(
        n8633), .ZN(n5505) );
  NAND2_X2 U7253 ( .A1(n5506), .A2(n5505), .ZN(n9092) );
  NAND2_X1 U7254 ( .A1(n5845), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7255 ( .A1(n6086), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5513) );
  INV_X1 U7256 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7257 ( .A1(n5509), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5510) );
  AND2_X1 U7258 ( .A1(n5524), .A2(n5510), .ZN(n8934) );
  OR2_X1 U7259 ( .A1(n5292), .A2(n8934), .ZN(n5512) );
  INV_X1 U7260 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10520) );
  OR2_X1 U7261 ( .A1(n6091), .A2(n10520), .ZN(n5511) );
  NAND4_X1 U7262 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n8920)
         );
  NOR2_X1 U7263 ( .A1(n9092), .A2(n8920), .ZN(n6248) );
  MUX2_X1 U7264 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6393), .Z(n5531) );
  XNOR2_X1 U7265 ( .A(n5531), .B(SI_14_), .ZN(n5517) );
  XNOR2_X1 U7266 ( .A(n5532), .B(n5517), .ZN(n7326) );
  NAND2_X1 U7267 ( .A1(n7326), .A2(n6106), .ZN(n5523) );
  OAI21_X1 U7268 ( .B1(n5518), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5520) );
  INV_X1 U7269 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7270 ( .A1(n5520), .A2(n5519), .ZN(n5534) );
  OR2_X1 U7271 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  AND2_X1 U7272 ( .A1(n5534), .A2(n5521), .ZN(n6039) );
  AOI22_X1 U7273 ( .A1(n5622), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4407), .B2(
        n6039), .ZN(n5522) );
  NAND2_X1 U7274 ( .A1(n5845), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7275 ( .A1(n5524), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7276 ( .A1(n5543), .A2(n5525), .ZN(n8923) );
  NAND2_X1 U7277 ( .A1(n5799), .A2(n8923), .ZN(n5528) );
  INV_X1 U7278 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9085) );
  OR2_X1 U7279 ( .A1(n5848), .A2(n9085), .ZN(n5527) );
  INV_X1 U7280 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8927) );
  OR2_X1 U7281 ( .A1(n6091), .A2(n8927), .ZN(n5526) );
  NAND4_X1 U7282 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n8932)
         );
  OR2_X1 U7283 ( .A1(n4626), .A2(n8932), .ZN(n5530) );
  MUX2_X1 U7284 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6393), .Z(n5552) );
  XNOR2_X1 U7285 ( .A(n5552), .B(SI_15_), .ZN(n5533) );
  NAND2_X1 U7286 ( .A1(n7489), .A2(n6106), .ZN(n5537) );
  NAND2_X1 U7287 ( .A1(n5534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5535) );
  XNOR2_X1 U7288 ( .A(n5535), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7490) );
  AOI22_X1 U7289 ( .A1(n7490), .A2(n4407), .B1(n5622), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5536) );
  INV_X1 U7290 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10652) );
  OR2_X1 U7291 ( .A1(n6091), .A2(n10652), .ZN(n5540) );
  INV_X1 U7292 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5538) );
  OR2_X1 U7293 ( .A1(n4424), .A2(n5538), .ZN(n5539) );
  AND2_X1 U7294 ( .A1(n5540), .A2(n5539), .ZN(n5547) );
  INV_X1 U7295 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7296 ( .A1(n5543), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7297 ( .A1(n5584), .A2(n5544), .ZN(n8911) );
  NAND2_X1 U7298 ( .A1(n8911), .A2(n5799), .ZN(n5546) );
  NAND2_X1 U7299 ( .A1(n6086), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7300 ( .A1(n8998), .A2(n8893), .ZN(n6179) );
  NOR2_X1 U7301 ( .A1(n8998), .A2(n8921), .ZN(n5548) );
  AOI21_X2 U7302 ( .B1(n8906), .B2(n8915), .A(n5548), .ZN(n8890) );
  INV_X1 U7303 ( .A(SI_15_), .ZN(n10621) );
  INV_X1 U7304 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7549) );
  INV_X1 U7305 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7548) );
  MUX2_X1 U7306 ( .A(n7549), .B(n7548), .S(n6393), .Z(n5577) );
  INV_X1 U7307 ( .A(SI_16_), .ZN(n5550) );
  AOI22_X1 U7308 ( .A1(n10621), .A2(n5572), .B1(n5577), .B2(n5550), .ZN(n5549)
         );
  OAI21_X1 U7309 ( .B1(n5572), .B2(n10621), .A(n5550), .ZN(n5554) );
  INV_X1 U7310 ( .A(n5577), .ZN(n5553) );
  AND2_X1 U7311 ( .A1(SI_16_), .A2(SI_15_), .ZN(n5551) );
  AOI22_X1 U7312 ( .A1(n5554), .A2(n5553), .B1(n5552), .B2(n5551), .ZN(n5555)
         );
  INV_X1 U7313 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7509) );
  INV_X1 U7314 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7275) );
  MUX2_X1 U7315 ( .A(n7509), .B(n7275), .S(n6393), .Z(n5557) );
  INV_X1 U7316 ( .A(SI_17_), .ZN(n5556) );
  INV_X1 U7317 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U7318 ( .A1(n5558), .A2(SI_17_), .ZN(n5559) );
  XNOR2_X1 U7319 ( .A(n5596), .B(n5595), .ZN(n7505) );
  NAND2_X1 U7320 ( .A1(n7505), .A2(n6106), .ZN(n5565) );
  OR2_X1 U7321 ( .A1(n5561), .A2(n5560), .ZN(n5580) );
  OAI21_X1 U7322 ( .B1(n5580), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5562) );
  MUX2_X1 U7323 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5562), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5563) );
  NAND2_X1 U7324 ( .A1(n5563), .A2(n5598), .ZN(n8702) );
  INV_X1 U7325 ( .A(n8702), .ZN(n6047) );
  AOI22_X1 U7326 ( .A1(n5622), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4407), .B2(
        n6047), .ZN(n5564) );
  INV_X1 U7327 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7328 ( .A1(n5586), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7329 ( .A1(n5602), .A2(n5568), .ZN(n8887) );
  NAND2_X1 U7330 ( .A1(n8887), .A2(n5799), .ZN(n5571) );
  AOI22_X1 U7331 ( .A1(n5844), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n5845), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7332 ( .A1(n6086), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7333 ( .A1(n9071), .A2(n8894), .ZN(n6176) );
  NAND2_X1 U7334 ( .A1(n6261), .A2(n6176), .ZN(n8878) );
  NAND2_X1 U7335 ( .A1(n5574), .A2(SI_15_), .ZN(n5573) );
  NAND2_X1 U7336 ( .A1(n5573), .A2(n5572), .ZN(n5576) );
  XNOR2_X1 U7337 ( .A(n5577), .B(SI_16_), .ZN(n5578) );
  NAND2_X1 U7338 ( .A1(n7547), .A2(n6106), .ZN(n5583) );
  NAND2_X1 U7339 ( .A1(n5580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5581) );
  XNOR2_X1 U7340 ( .A(n5581), .B(P2_IR_REG_16__SCAN_IN), .ZN(n6043) );
  AOI22_X1 U7341 ( .A1(n5622), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4407), .B2(
        n6043), .ZN(n5582) );
  NAND2_X2 U7342 ( .A1(n5583), .A2(n5582), .ZN(n8902) );
  NAND2_X1 U7343 ( .A1(n5584), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7344 ( .A1(n5586), .A2(n5585), .ZN(n8901) );
  NAND2_X1 U7345 ( .A1(n8901), .A2(n5799), .ZN(n5589) );
  AOI22_X1 U7346 ( .A1(n5844), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n5845), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7347 ( .A1(n6086), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7348 ( .A1(n8902), .A2(n8908), .ZN(n6180) );
  NAND3_X1 U7349 ( .A1(n8890), .A2(n8878), .A3(n8898), .ZN(n5593) );
  INV_X1 U7350 ( .A(n8908), .ZN(n8602) );
  NAND2_X1 U7351 ( .A1(n8902), .A2(n8602), .ZN(n8880) );
  NAND2_X1 U7352 ( .A1(n9071), .A2(n8865), .ZN(n5590) );
  INV_X1 U7353 ( .A(n5591), .ZN(n5592) );
  MUX2_X1 U7354 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6393), .Z(n5612) );
  INV_X1 U7355 ( .A(SI_18_), .ZN(n5597) );
  XNOR2_X1 U7356 ( .A(n5613), .B(n5611), .ZN(n7585) );
  NAND2_X1 U7357 ( .A1(n7585), .A2(n6106), .ZN(n5601) );
  NAND2_X1 U7358 ( .A1(n5598), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5599) );
  XNOR2_X1 U7359 ( .A(n5599), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8727) );
  AOI22_X1 U7360 ( .A1(n5622), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4407), .B2(
        n8727), .ZN(n5600) );
  NAND2_X1 U7361 ( .A1(n5602), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7362 ( .A1(n5625), .A2(n5603), .ZN(n8562) );
  NAND2_X1 U7363 ( .A1(n8562), .A2(n5799), .ZN(n5608) );
  INV_X1 U7364 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U7365 ( .A1(n5844), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7366 ( .A1(n6086), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U7367 ( .C1(n4424), .C2(n10517), .A(n5605), .B(n5604), .ZN(n5606)
         );
  INV_X1 U7368 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U7369 ( .A1(n5608), .A2(n5607), .ZN(n8601) );
  INV_X1 U7370 ( .A(n8871), .ZN(n8992) );
  NAND2_X1 U7371 ( .A1(n5610), .A2(n5176), .ZN(n8852) );
  INV_X1 U7372 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7752) );
  INV_X1 U7373 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7754) );
  MUX2_X1 U7374 ( .A(n7752), .B(n7754), .S(n6393), .Z(n5615) );
  INV_X1 U7375 ( .A(SI_19_), .ZN(n5614) );
  INV_X1 U7376 ( .A(n5615), .ZN(n5616) );
  NAND2_X1 U7377 ( .A1(n5616), .A2(SI_19_), .ZN(n5617) );
  NAND2_X1 U7378 ( .A1(n5632), .A2(n5617), .ZN(n5633) );
  XNOR2_X1 U7379 ( .A(n5634), .B(n5633), .ZN(n7750) );
  NAND2_X1 U7380 ( .A1(n7750), .A2(n6106), .ZN(n5624) );
  INV_X1 U7381 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7382 ( .A1(n5807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5620) );
  AOI22_X1 U7383 ( .A1(n5622), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5854), .B2(
        n4407), .ZN(n5623) );
  INV_X1 U7384 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U7385 ( .A1(n5625), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7386 ( .A1(n5653), .A2(n5626), .ZN(n8859) );
  NAND2_X1 U7387 ( .A1(n8859), .A2(n5799), .ZN(n5631) );
  INV_X1 U7388 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U7389 ( .A1(n5844), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7390 ( .A1(n6086), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U7391 ( .C1(n4424), .C2(n10545), .A(n5628), .B(n5627), .ZN(n5629)
         );
  INV_X1 U7392 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7393 ( .A1(n8987), .A2(n8563), .ZN(n6188) );
  NAND2_X1 U7394 ( .A1(n6189), .A2(n6188), .ZN(n8851) );
  INV_X1 U7395 ( .A(SI_20_), .ZN(n5648) );
  INV_X1 U7396 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7840) );
  INV_X1 U7397 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7836) );
  MUX2_X1 U7398 ( .A(n7840), .B(n7836), .S(n5277), .Z(n5647) );
  NAND2_X1 U7399 ( .A1(n5646), .A2(n5648), .ZN(n5635) );
  INV_X1 U7400 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7992) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10519) );
  MUX2_X1 U7402 ( .A(n7992), .B(n10519), .S(n6393), .Z(n5658) );
  XNOR2_X1 U7403 ( .A(n5658), .B(SI_21_), .ZN(n5637) );
  NAND2_X1 U7404 ( .A1(n7991), .A2(n6106), .ZN(n5639) );
  OR2_X1 U7405 ( .A1(n4405), .A2(n7992), .ZN(n5638) );
  INV_X1 U7406 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5640) );
  INV_X1 U7407 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U7408 ( .A1(n4456), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7409 ( .A1(n5669), .A2(n5642), .ZN(n8837) );
  INV_X1 U7410 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U7411 ( .A1(n5844), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7412 ( .A1(n5845), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U7413 ( .C1(n9053), .C2(n5848), .A(n5644), .B(n5643), .ZN(n5645)
         );
  INV_X1 U7414 ( .A(n5647), .ZN(n5649) );
  XNOR2_X1 U7415 ( .A(n5649), .B(n5648), .ZN(n5650) );
  XNOR2_X1 U7416 ( .A(n5646), .B(n5650), .ZN(n7835) );
  NAND2_X1 U7417 ( .A1(n7835), .A2(n6106), .ZN(n5652) );
  OR2_X1 U7418 ( .A1(n6104), .A2(n7840), .ZN(n5651) );
  NAND2_X1 U7419 ( .A1(n5653), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7420 ( .A1(n4456), .A2(n5654), .ZN(n8848) );
  INV_X1 U7421 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U7422 ( .A1(n6086), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7423 ( .A1(n5845), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5655) );
  OAI211_X1 U7424 ( .C1(n6091), .C2(n8847), .A(n5656), .B(n5655), .ZN(n5657)
         );
  NAND2_X1 U7425 ( .A1(n9060), .A2(n8855), .ZN(n6195) );
  NOR2_X1 U7426 ( .A1(n5659), .A2(SI_21_), .ZN(n5661) );
  NAND2_X1 U7427 ( .A1(n5659), .A2(SI_21_), .ZN(n5660) );
  INV_X1 U7428 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8181) );
  INV_X1 U7429 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8178) );
  MUX2_X1 U7430 ( .A(n8181), .B(n8178), .S(n6393), .Z(n5664) );
  INV_X1 U7431 ( .A(SI_22_), .ZN(n5663) );
  NAND2_X1 U7432 ( .A1(n5664), .A2(n5663), .ZN(n5677) );
  INV_X1 U7433 ( .A(n5664), .ZN(n5665) );
  NAND2_X1 U7434 ( .A1(n5665), .A2(SI_22_), .ZN(n5666) );
  NAND2_X1 U7435 ( .A1(n5677), .A2(n5666), .ZN(n5678) );
  XNOR2_X1 U7436 ( .A(n5679), .B(n5678), .ZN(n8176) );
  NAND2_X1 U7437 ( .A1(n8176), .A2(n6106), .ZN(n5668) );
  OR2_X1 U7438 ( .A1(n6104), .A2(n8181), .ZN(n5667) );
  NAND2_X1 U7439 ( .A1(n5669), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7440 ( .A1(n5686), .A2(n5670), .ZN(n8543) );
  NAND2_X1 U7441 ( .A1(n8543), .A2(n5799), .ZN(n5675) );
  INV_X1 U7442 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U7443 ( .A1(n5845), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5672) );
  INV_X1 U7444 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8818) );
  OR2_X1 U7445 ( .A1(n6091), .A2(n8818), .ZN(n5671) );
  OAI211_X1 U7446 ( .C1(n10655), .C2(n5848), .A(n5672), .B(n5671), .ZN(n5673)
         );
  INV_X1 U7447 ( .A(n5673), .ZN(n5674) );
  OR2_X1 U7448 ( .A1(n8825), .A2(n8834), .ZN(n8803) );
  INV_X1 U7449 ( .A(n8855), .ZN(n8833) );
  NOR2_X1 U7450 ( .A1(n9060), .A2(n8833), .ZN(n8830) );
  NAND2_X1 U7451 ( .A1(n8829), .A2(n8830), .ZN(n5676) );
  INV_X1 U7452 ( .A(n8816), .ZN(n8845) );
  OR2_X1 U7453 ( .A1(n9054), .A2(n8845), .ZN(n8813) );
  INV_X1 U7454 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10501) );
  INV_X1 U7455 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8243) );
  MUX2_X1 U7456 ( .A(n10501), .B(n8243), .S(n6393), .Z(n5681) );
  INV_X1 U7457 ( .A(SI_23_), .ZN(n5680) );
  NAND2_X1 U7458 ( .A1(n5681), .A2(n5680), .ZN(n5697) );
  INV_X1 U7459 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U7460 ( .A1(n5682), .A2(SI_23_), .ZN(n5683) );
  OR2_X1 U7461 ( .A1(n4405), .A2(n10501), .ZN(n5684) );
  NAND2_X2 U7462 ( .A1(n5685), .A2(n5684), .ZN(n9045) );
  NAND2_X1 U7463 ( .A1(n5686), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7464 ( .A1(n5707), .A2(n5687), .ZN(n8810) );
  NAND2_X1 U7465 ( .A1(n8810), .A2(n5799), .ZN(n5692) );
  INV_X1 U7466 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10574) );
  NAND2_X1 U7467 ( .A1(n5844), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7468 ( .A1(n5845), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5688) );
  OAI211_X1 U7469 ( .C1(n10574), .C2(n5848), .A(n5689), .B(n5688), .ZN(n5690)
         );
  INV_X1 U7470 ( .A(n5690), .ZN(n5691) );
  AOI22_X1 U7471 ( .A1(n9045), .A2(n8788), .B1(n8834), .B2(n8825), .ZN(n5694)
         );
  INV_X1 U7472 ( .A(n9045), .ZN(n5693) );
  INV_X1 U7473 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8306) );
  INV_X1 U7474 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8308) );
  MUX2_X1 U7475 ( .A(n8306), .B(n8308), .S(n6393), .Z(n5699) );
  INV_X1 U7476 ( .A(SI_24_), .ZN(n5698) );
  NAND2_X1 U7477 ( .A1(n5699), .A2(n5698), .ZN(n5716) );
  INV_X1 U7478 ( .A(n5699), .ZN(n5700) );
  NAND2_X1 U7479 ( .A1(n5700), .A2(SI_24_), .ZN(n5701) );
  NAND2_X1 U7480 ( .A1(n8305), .A2(n6106), .ZN(n5704) );
  OR2_X1 U7481 ( .A1(n4405), .A2(n8306), .ZN(n5703) );
  INV_X1 U7482 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7483 ( .A1(n5707), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7484 ( .A1(n5725), .A2(n5708), .ZN(n8794) );
  NAND2_X1 U7485 ( .A1(n8794), .A2(n5799), .ZN(n5713) );
  INV_X1 U7486 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U7487 ( .A1(n5844), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7488 ( .A1(n5845), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5709) );
  OAI211_X1 U7489 ( .C1(n9039), .C2(n5848), .A(n5710), .B(n5709), .ZN(n5711)
         );
  INV_X1 U7490 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7491 ( .A1(n8792), .A2(n8493), .ZN(n5714) );
  NAND2_X1 U7492 ( .A1(n5717), .A2(n5716), .ZN(n5735) );
  INV_X1 U7493 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9122) );
  INV_X1 U7494 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10563) );
  MUX2_X1 U7495 ( .A(n9122), .B(n10563), .S(n6393), .Z(n5718) );
  INV_X1 U7496 ( .A(SI_25_), .ZN(n10595) );
  NAND2_X1 U7497 ( .A1(n5718), .A2(n10595), .ZN(n5751) );
  INV_X1 U7498 ( .A(n5718), .ZN(n5719) );
  NAND2_X1 U7499 ( .A1(n5719), .A2(SI_25_), .ZN(n5720) );
  NAND2_X1 U7500 ( .A1(n9120), .A2(n6106), .ZN(n5722) );
  OR2_X1 U7501 ( .A1(n6104), .A2(n9122), .ZN(n5721) );
  INV_X1 U7502 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7503 ( .A1(n5725), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7504 ( .A1(n5743), .A2(n5726), .ZN(n8782) );
  NAND2_X1 U7505 ( .A1(n8782), .A2(n5799), .ZN(n5731) );
  INV_X1 U7506 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U7507 ( .A1(n5844), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7508 ( .A1(n6086), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5727) );
  OAI211_X1 U7509 ( .C1(n4424), .C2(n10609), .A(n5728), .B(n5727), .ZN(n5729)
         );
  INV_X1 U7510 ( .A(n5729), .ZN(n5730) );
  INV_X1 U7511 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9118) );
  INV_X1 U7512 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10113) );
  MUX2_X1 U7513 ( .A(n9118), .B(n10113), .S(n6393), .Z(n5737) );
  INV_X1 U7514 ( .A(SI_26_), .ZN(n5736) );
  NAND2_X1 U7515 ( .A1(n5737), .A2(n5736), .ZN(n5750) );
  INV_X1 U7516 ( .A(n5737), .ZN(n5738) );
  NAND2_X1 U7517 ( .A1(n5738), .A2(SI_26_), .ZN(n5752) );
  AND2_X1 U7518 ( .A1(n5750), .A2(n5752), .ZN(n5739) );
  OR2_X1 U7519 ( .A1(n6104), .A2(n9118), .ZN(n5741) );
  NAND2_X1 U7520 ( .A1(n5743), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7521 ( .A1(n5762), .A2(n5744), .ZN(n8771) );
  NAND2_X1 U7522 ( .A1(n8771), .A2(n5799), .ZN(n5749) );
  INV_X1 U7523 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U7524 ( .A1(n5844), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5746) );
  INV_X1 U7525 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10505) );
  OR2_X1 U7526 ( .A1(n4424), .A2(n10505), .ZN(n5745) );
  OAI211_X1 U7527 ( .C1(n10590), .C2(n5848), .A(n5746), .B(n5745), .ZN(n5747)
         );
  INV_X1 U7528 ( .A(n5747), .ZN(n5748) );
  AND2_X1 U7529 ( .A1(n5751), .A2(n5750), .ZN(n5754) );
  INV_X1 U7530 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5759) );
  INV_X1 U7531 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10112) );
  MUX2_X1 U7532 ( .A(n5759), .B(n10112), .S(n5277), .Z(n5756) );
  INV_X1 U7533 ( .A(SI_27_), .ZN(n10554) );
  NAND2_X1 U7534 ( .A1(n5756), .A2(n10554), .ZN(n5787) );
  INV_X1 U7535 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7536 ( .A1(n5757), .A2(SI_27_), .ZN(n5758) );
  NAND2_X1 U7537 ( .A1(n9113), .A2(n6106), .ZN(n5761) );
  OR2_X1 U7538 ( .A1(n4405), .A2(n5759), .ZN(n5760) );
  NAND2_X1 U7539 ( .A1(n5762), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7540 ( .A1(n5774), .A2(n5763), .ZN(n8758) );
  NAND2_X1 U7541 ( .A1(n8758), .A2(n5799), .ZN(n5768) );
  INV_X1 U7542 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U7543 ( .A1(n5844), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7544 ( .A1(n5845), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U7545 ( .C1(n10449), .C2(n5848), .A(n5765), .B(n5764), .ZN(n5766)
         );
  INV_X1 U7546 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7547 ( .A1(n8762), .A2(n8401), .ZN(n6227) );
  INV_X1 U7548 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5771) );
  INV_X1 U7549 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8410) );
  MUX2_X1 U7550 ( .A(n5771), .B(n8410), .S(n5277), .Z(n5788) );
  XNOR2_X1 U7551 ( .A(n5788), .B(SI_28_), .ZN(n6069) );
  OR2_X1 U7552 ( .A1(n6104), .A2(n5771), .ZN(n5772) );
  NAND2_X1 U7553 ( .A1(n5774), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5775) );
  INV_X1 U7554 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10612) );
  INV_X1 U7555 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5936) );
  OR2_X1 U7556 ( .A1(n6091), .A2(n5936), .ZN(n5777) );
  INV_X1 U7557 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10506) );
  OR2_X1 U7558 ( .A1(n4424), .A2(n10506), .ZN(n5776) );
  OAI211_X1 U7559 ( .C1(n5848), .C2(n10612), .A(n5777), .B(n5776), .ZN(n5778)
         );
  INV_X1 U7560 ( .A(n5778), .ZN(n5779) );
  NOR2_X1 U7561 ( .A1(n8951), .A2(n8757), .ZN(n5780) );
  INV_X1 U7562 ( .A(n8757), .ZN(n5838) );
  OAI22_X1 U7563 ( .A1(n5918), .A2(n5780), .B1(n5838), .B2(n4704), .ZN(n5806)
         );
  INV_X1 U7564 ( .A(n5788), .ZN(n5789) );
  NAND2_X1 U7565 ( .A1(n5789), .A2(SI_28_), .ZN(n5781) );
  INV_X1 U7566 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10636) );
  INV_X1 U7567 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8312) );
  MUX2_X1 U7568 ( .A(n10636), .B(n8312), .S(n6393), .Z(n5783) );
  NAND2_X1 U7569 ( .A1(n5781), .A2(n5783), .ZN(n5786) );
  INV_X1 U7570 ( .A(SI_28_), .ZN(n5782) );
  NAND2_X1 U7571 ( .A1(n5788), .A2(n5782), .ZN(n6071) );
  INV_X1 U7572 ( .A(n5783), .ZN(n6072) );
  AND3_X1 U7573 ( .A1(n6071), .A2(n5787), .A3(n6072), .ZN(n5784) );
  NAND2_X1 U7574 ( .A1(n5785), .A2(n5784), .ZN(n5796) );
  INV_X1 U7575 ( .A(n5786), .ZN(n5794) );
  INV_X1 U7576 ( .A(n5787), .ZN(n5793) );
  OAI21_X1 U7577 ( .B1(n6072), .B2(SI_28_), .A(n5788), .ZN(n5792) );
  NAND2_X1 U7578 ( .A1(n6072), .A2(SI_28_), .ZN(n5790) );
  NAND2_X1 U7579 ( .A1(n5790), .A2(n5789), .ZN(n5791) );
  AOI22_X1 U7580 ( .A1(n5794), .A2(n5793), .B1(n5792), .B2(n5791), .ZN(n5795)
         );
  NAND2_X1 U7581 ( .A1(n7098), .A2(n6106), .ZN(n5798) );
  OR2_X1 U7582 ( .A1(n6104), .A2(n10636), .ZN(n5797) );
  NAND2_X1 U7583 ( .A1(n5798), .A2(n5797), .ZN(n5805) );
  INV_X1 U7584 ( .A(n8738), .ZN(n5800) );
  NAND2_X1 U7585 ( .A1(n5800), .A2(n5799), .ZN(n6094) );
  INV_X1 U7586 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7587 ( .A1(n6086), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7588 ( .A1(n5844), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5801) );
  OAI211_X1 U7589 ( .C1(n4424), .C2(n5900), .A(n5802), .B(n5801), .ZN(n5803)
         );
  INV_X1 U7590 ( .A(n5803), .ZN(n5804) );
  NAND2_X1 U7591 ( .A1(n5805), .A2(n8398), .ZN(n6081) );
  XNOR2_X1 U7592 ( .A(n5806), .B(n6242), .ZN(n5853) );
  XNOR2_X2 U7593 ( .A(n5810), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7594 ( .A1(n6301), .A2(n5854), .ZN(n5905) );
  XNOR2_X2 U7595 ( .A(n5812), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7596 ( .A1(n5858), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5813) );
  INV_X1 U7597 ( .A(n7838), .ZN(n6273) );
  NAND2_X1 U7598 ( .A1(n6114), .A2(n6273), .ZN(n7386) );
  INV_X1 U7599 ( .A(n6109), .ZN(n7407) );
  NAND2_X1 U7600 ( .A1(n7715), .A2(n5814), .ZN(n7714) );
  NAND2_X1 U7601 ( .A1(n7714), .A2(n5815), .ZN(n7613) );
  INV_X1 U7602 ( .A(n7615), .ZN(n6252) );
  NAND2_X1 U7603 ( .A1(n7613), .A2(n6252), .ZN(n5816) );
  INV_X1 U7604 ( .A(n10302), .ZN(n7501) );
  NAND2_X1 U7605 ( .A1(n7528), .A2(n7501), .ZN(n6120) );
  NAND2_X1 U7606 ( .A1(n5816), .A2(n6120), .ZN(n10290) );
  XNOR2_X1 U7607 ( .A(n10276), .B(n6121), .ZN(n10291) );
  NAND2_X1 U7608 ( .A1(n10290), .A2(n10291), .ZN(n5817) );
  NAND2_X1 U7609 ( .A1(n7617), .A2(n6121), .ZN(n6140) );
  NAND2_X1 U7610 ( .A1(n5817), .A2(n6140), .ZN(n10278) );
  XNOR2_X1 U7611 ( .A(n10285), .B(n10311), .ZN(n10279) );
  NAND2_X1 U7612 ( .A1(n10278), .A2(n10279), .ZN(n5818) );
  NAND2_X1 U7613 ( .A1(n7894), .A2(n10311), .ZN(n6130) );
  NAND2_X1 U7614 ( .A1(n10275), .A2(n5819), .ZN(n6141) );
  NAND2_X1 U7615 ( .A1(n10257), .A2(n7937), .ZN(n6132) );
  NAND2_X1 U7616 ( .A1(n7930), .A2(n10315), .ZN(n7921) );
  AND2_X1 U7617 ( .A1(n6132), .A2(n7921), .ZN(n6145) );
  NAND2_X1 U7618 ( .A1(n8608), .A2(n10324), .ZN(n6147) );
  INV_X1 U7619 ( .A(n8605), .ZN(n8339) );
  NAND2_X1 U7620 ( .A1(n8226), .A2(n8339), .ZN(n6249) );
  AND2_X1 U7621 ( .A1(n6249), .A2(n8130), .ZN(n6137) );
  NAND2_X1 U7622 ( .A1(n8444), .A2(n8554), .ZN(n6256) );
  NAND2_X1 U7623 ( .A1(n8171), .A2(n10268), .ZN(n6150) );
  NAND2_X1 U7624 ( .A1(n10331), .A2(n8607), .ZN(n7940) );
  NAND2_X1 U7625 ( .A1(n10259), .A2(n5190), .ZN(n5823) );
  INV_X1 U7626 ( .A(n6137), .ZN(n5820) );
  AND2_X1 U7627 ( .A1(n6136), .A2(n7940), .ZN(n8129) );
  OR2_X1 U7628 ( .A1(n8444), .A2(n8554), .ZN(n6257) );
  OAI211_X1 U7629 ( .C1(n5820), .C2(n8129), .A(n8233), .B(n6257), .ZN(n5821)
         );
  NAND2_X1 U7630 ( .A1(n5821), .A2(n6256), .ZN(n5822) );
  NAND2_X1 U7631 ( .A1(n5823), .A2(n5822), .ZN(n8270) );
  NAND2_X1 U7632 ( .A1(n9092), .A2(n8477), .ZN(n5824) );
  INV_X1 U7633 ( .A(n8931), .ZN(n8352) );
  OR2_X1 U7634 ( .A1(n8482), .A2(n8352), .ZN(n8938) );
  NAND2_X1 U7635 ( .A1(n8938), .A2(n8477), .ZN(n5827) );
  INV_X1 U7636 ( .A(n9092), .ZN(n6167) );
  AND2_X1 U7637 ( .A1(n8920), .A2(n8931), .ZN(n5826) );
  AOI22_X1 U7638 ( .A1(n5827), .A2(n6167), .B1(n9102), .B2(n5826), .ZN(n5828)
         );
  INV_X1 U7639 ( .A(n8932), .ZN(n8907) );
  NOR2_X1 U7640 ( .A1(n9086), .A2(n8907), .ZN(n6172) );
  INV_X1 U7641 ( .A(n8916), .ZN(n5829) );
  NAND2_X1 U7642 ( .A1(n5829), .A2(n6179), .ZN(n5830) );
  NAND2_X1 U7643 ( .A1(n5830), .A2(n6174), .ZN(n8900) );
  NAND2_X1 U7644 ( .A1(n8879), .A2(n6261), .ZN(n5831) );
  NAND2_X1 U7645 ( .A1(n8871), .A2(n8883), .ZN(n6185) );
  NAND2_X1 U7646 ( .A1(n6247), .A2(n6185), .ZN(n8875) );
  INV_X1 U7647 ( .A(n8875), .ZN(n5832) );
  INV_X1 U7648 ( .A(n6196), .ZN(n5833) );
  INV_X1 U7649 ( .A(n6201), .ZN(n5834) );
  OR2_X1 U7650 ( .A1(n8825), .A2(n8465), .ZN(n8799) );
  NAND2_X1 U7651 ( .A1(n9045), .A2(n8817), .ZN(n6245) );
  NAND2_X1 U7652 ( .A1(n8774), .A2(n6218), .ZN(n5836) );
  NAND2_X1 U7653 ( .A1(n5836), .A2(n6213), .ZN(n8765) );
  NAND2_X1 U7654 ( .A1(n9028), .A2(n8755), .ZN(n6222) );
  NAND2_X1 U7655 ( .A1(n8765), .A2(n8766), .ZN(n5837) );
  NAND2_X2 U7656 ( .A1(n6301), .A2(n6114), .ZN(n6241) );
  AND2_X1 U7657 ( .A1(n7838), .A2(n4428), .ZN(n5867) );
  INV_X1 U7658 ( .A(n5867), .ZN(n5839) );
  AOI21_X1 U7659 ( .B1(n8179), .B2(n6273), .A(n5854), .ZN(n5840) );
  NAND2_X1 U7660 ( .A1(n8742), .A2(n7902), .ZN(n5852) );
  INV_X1 U7661 ( .A(n5841), .ZN(n6299) );
  INV_X4 U7662 ( .A(n6010), .ZN(n6298) );
  NAND2_X1 U7663 ( .A1(n6299), .A2(n6010), .ZN(n5843) );
  NAND2_X1 U7664 ( .A1(n5243), .A2(n5843), .ZN(n7404) );
  INV_X1 U7665 ( .A(n7404), .ZN(n7402) );
  INV_X1 U7666 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10446) );
  NAND2_X1 U7667 ( .A1(n5844), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7668 ( .A1(n5845), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5846) );
  OAI211_X1 U7669 ( .C1(n10446), .C2(n5848), .A(n5847), .B(n5846), .ZN(n5849)
         );
  INV_X1 U7670 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U7671 ( .A1(n6094), .A2(n5850), .ZN(n8599) );
  AOI21_X1 U7672 ( .B1(P2_B_REG_SCAN_IN), .B2(n5243), .A(n10254), .ZN(n8736)
         );
  AOI22_X1 U7673 ( .A1(n10286), .A2(n8757), .B1(n8599), .B2(n8736), .ZN(n5851)
         );
  OAI211_X1 U7674 ( .C1(n5853), .C2(n8853), .A(n5852), .B(n5851), .ZN(n8743)
         );
  NOR2_X1 U7675 ( .A1(n8743), .A2(n5855), .ZN(n5917) );
  NAND2_X1 U7676 ( .A1(n5856), .A2(n4599), .ZN(n5857) );
  INV_X1 U7677 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5866) );
  INV_X1 U7678 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7679 ( .A1(n5861), .A2(n5868), .ZN(n5859) );
  NAND2_X1 U7680 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U7681 ( .A(n5860), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7682 ( .A(n5861), .B(P2_IR_REG_24__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7683 ( .A1(n5862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5863) );
  XNOR2_X1 U7684 ( .A(n5863), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5890) );
  AND2_X1 U7685 ( .A1(n5893), .A2(n5890), .ZN(n5864) );
  NAND2_X1 U7686 ( .A1(n5889), .A2(n5864), .ZN(n7373) );
  XNOR2_X1 U7687 ( .A(n5865), .B(n5866), .ZN(n7372) );
  OR2_X1 U7688 ( .A1(n6241), .A2(n5867), .ZN(n7371) );
  NAND2_X1 U7689 ( .A1(n5868), .A2(P2_B_REG_SCAN_IN), .ZN(n5871) );
  INV_X1 U7690 ( .A(P2_B_REG_SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7691 ( .A1(n5869), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5870) );
  NAND4_X1 U7692 ( .A1(n5874), .A2(P2_IR_REG_25__SCAN_IN), .A3(n5871), .A4(
        n5870), .ZN(n5877) );
  OAI21_X1 U7693 ( .B1(n5871), .B2(P2_IR_REG_25__SCAN_IN), .A(n5870), .ZN(
        n5872) );
  INV_X1 U7694 ( .A(n5872), .ZN(n5873) );
  INV_X1 U7695 ( .A(n5875), .ZN(n5876) );
  NOR4_X1 U7696 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n10410) );
  NOR2_X1 U7697 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n5880) );
  NOR4_X1 U7698 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5879) );
  NOR4_X1 U7699 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5878) );
  NAND4_X1 U7700 ( .A1(n10410), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n5886)
         );
  NOR4_X1 U7701 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5884) );
  NOR4_X1 U7702 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5883) );
  NOR4_X1 U7703 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5882) );
  NOR4_X1 U7704 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5881) );
  NAND4_X1 U7705 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n5885)
         );
  NOR2_X1 U7706 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  OR2_X1 U7707 ( .A1(n7194), .A2(n5887), .ZN(n5907) );
  NAND2_X1 U7708 ( .A1(n7371), .A2(n5907), .ZN(n5888) );
  NOR2_X1 U7709 ( .A1(n6297), .A2(n5888), .ZN(n5895) );
  INV_X1 U7710 ( .A(n5889), .ZN(n9124) );
  INV_X1 U7711 ( .A(n5890), .ZN(n9119) );
  NAND2_X1 U7712 ( .A1(n9124), .A2(n9119), .ZN(n7240) );
  INV_X1 U7713 ( .A(n7194), .ZN(n5891) );
  INV_X1 U7714 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10637) );
  NAND2_X1 U7715 ( .A1(n5891), .A2(n10637), .ZN(n5892) );
  NAND2_X1 U7716 ( .A1(n7240), .A2(n5892), .ZN(n5930) );
  INV_X1 U7717 ( .A(n5893), .ZN(n8307) );
  AND2_X1 U7718 ( .A1(n10317), .A2(n7385), .ZN(n5934) );
  NOR2_X1 U7719 ( .A1(n5934), .A2(n7383), .ZN(n5898) );
  INV_X1 U7720 ( .A(n5930), .ZN(n5897) );
  NAND3_X1 U7721 ( .A1(n6301), .A2(n6273), .A3(n4428), .ZN(n5896) );
  NAND2_X1 U7722 ( .A1(n6241), .A2(n5896), .ZN(n5928) );
  MUX2_X1 U7723 ( .A(n5898), .B(n5897), .S(n5928), .Z(n5899) );
  AND2_X2 U7724 ( .A1(n5933), .A2(n5899), .ZN(n10672) );
  NAND2_X1 U7725 ( .A1(n10672), .A2(n10316), .ZN(n9018) );
  OAI21_X1 U7726 ( .B1(n5917), .B2(n8960), .A(n5902), .ZN(P2_U3488) );
  INV_X1 U7727 ( .A(n5907), .ZN(n5903) );
  NOR2_X1 U7728 ( .A1(n5904), .A2(n5903), .ZN(n7377) );
  INV_X1 U7729 ( .A(n6297), .ZN(n7193) );
  NAND2_X1 U7730 ( .A1(n7377), .A2(n7193), .ZN(n7400) );
  NOR2_X1 U7731 ( .A1(n5905), .A2(n7838), .ZN(n5909) );
  NAND2_X1 U7732 ( .A1(n5909), .A2(n7385), .ZN(n7370) );
  AND2_X1 U7733 ( .A1(n7370), .A2(n7419), .ZN(n5906) );
  AND2_X1 U7734 ( .A1(n7383), .A2(n5907), .ZN(n5908) );
  NAND2_X1 U7735 ( .A1(n5930), .A2(n5908), .ZN(n7379) );
  NOR2_X1 U7736 ( .A1(n7379), .A2(n6297), .ZN(n7406) );
  AND2_X1 U7737 ( .A1(n6241), .A2(n10330), .ZN(n5911) );
  INV_X1 U7738 ( .A(n5909), .ZN(n5910) );
  NAND2_X1 U7739 ( .A1(n5911), .A2(n5910), .ZN(n7395) );
  OR2_X1 U7740 ( .A1(n10330), .A2(n7384), .ZN(n8791) );
  NAND2_X1 U7741 ( .A1(n7395), .A2(n8791), .ZN(n7369) );
  NAND2_X1 U7742 ( .A1(n7406), .A2(n7369), .ZN(n5912) );
  NAND2_X1 U7743 ( .A1(n10336), .A2(n10316), .ZN(n9101) );
  INV_X1 U7744 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5914) );
  INV_X1 U7745 ( .A(n5915), .ZN(n5916) );
  OAI21_X1 U7746 ( .B1(n5917), .B2(n10337), .A(n5916), .ZN(P2_U3456) );
  XNOR2_X1 U7747 ( .A(n5918), .B(n5125), .ZN(n5922) );
  INV_X1 U7748 ( .A(n8398), .ZN(n8600) );
  AOI21_X1 U7749 ( .B1(n5922), .B2(n10289), .A(n5921), .ZN(n8948) );
  MUX2_X1 U7750 ( .A(n10612), .B(n8948), .S(n10336), .Z(n5927) );
  NAND2_X1 U7751 ( .A1(n8951), .A2(n9093), .ZN(n5924) );
  INV_X1 U7752 ( .A(n5928), .ZN(n5931) );
  AND2_X1 U7753 ( .A1(n7383), .A2(n5928), .ZN(n5929) );
  AOI21_X1 U7754 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(n5932) );
  NAND2_X1 U7755 ( .A1(n5933), .A2(n5932), .ZN(n5938) );
  INV_X1 U7756 ( .A(n5934), .ZN(n5935) );
  NAND2_X2 U7757 ( .A1(n5938), .A2(n8912), .ZN(n10282) );
  MUX2_X1 U7758 ( .A(n5936), .B(n8948), .S(n10282), .Z(n5943) );
  AND2_X1 U7759 ( .A1(n7384), .A2(n6114), .ZN(n7614) );
  OR2_X1 U7760 ( .A1(n7902), .A2(n7614), .ZN(n5937) );
  INV_X1 U7761 ( .A(n5938), .ZN(n5939) );
  INV_X1 U7762 ( .A(n8791), .ZN(n8936) );
  NAND2_X1 U7763 ( .A1(n5939), .A2(n8936), .ZN(n8744) );
  AOI22_X1 U7764 ( .A1(n8951), .A2(n10292), .B1(n10293), .B2(n8399), .ZN(n5940) );
  NAND2_X1 U7765 ( .A1(n7373), .A2(n6241), .ZN(n5944) );
  NAND2_X1 U7766 ( .A1(n5944), .A2(n7372), .ZN(n6057) );
  NAND2_X1 U7767 ( .A1(n6057), .A2(n5243), .ZN(n5945) );
  NAND2_X1 U7768 ( .A1(n5945), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U7769 ( .A(n4428), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6051) );
  INV_X1 U7770 ( .A(n6043), .ZN(n8684) );
  NAND2_X1 U7771 ( .A1(n5107), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5947) );
  INV_X1 U7772 ( .A(n5948), .ZN(n5949) );
  NAND2_X1 U7773 ( .A1(n7350), .A2(n5949), .ZN(n8611) );
  XNOR2_X1 U7774 ( .A(n7163), .B(n10338), .ZN(n8612) );
  NAND2_X1 U7775 ( .A1(n8611), .A2(n8612), .ZN(n8610) );
  NAND2_X1 U7776 ( .A1(n7163), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7777 ( .A1(n8610), .A2(n5950), .ZN(n5951) );
  NAND2_X1 U7778 ( .A1(n5951), .A2(n7166), .ZN(n7317) );
  AND2_X1 U7779 ( .A1(n7317), .A2(n5952), .ZN(n7334) );
  NAND2_X1 U7780 ( .A1(n7334), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U7781 ( .A1(n7333), .A2(n7317), .ZN(n5954) );
  INV_X1 U7782 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5953) );
  XNOR2_X1 U7783 ( .A(n7325), .B(n5953), .ZN(n7316) );
  NAND2_X1 U7784 ( .A1(n7325), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7785 ( .A1(n7320), .A2(n5955), .ZN(n5956) );
  NAND2_X1 U7786 ( .A1(n5956), .A2(n7168), .ZN(n7562) );
  OR2_X1 U7787 ( .A1(n7179), .A2(n10546), .ZN(n5958) );
  OR2_X1 U7788 ( .A1(n5959), .A2(n7763), .ZN(n5960) );
  NAND2_X1 U7789 ( .A1(n5959), .A2(n7763), .ZN(n7966) );
  NAND2_X1 U7790 ( .A1(n7965), .A2(n7966), .ZN(n5961) );
  XNOR2_X1 U7791 ( .A(n7964), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7967) );
  INV_X1 U7792 ( .A(n7964), .ZN(n7198) );
  NAND2_X1 U7793 ( .A1(n7198), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5962) );
  INV_X1 U7794 ( .A(n8083), .ZN(n7202) );
  INV_X1 U7795 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8231) );
  XNOR2_X1 U7796 ( .A(n8200), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U7797 ( .A1(n5963), .A2(n8192), .ZN(n8197) );
  INV_X1 U7798 ( .A(n8200), .ZN(n7197) );
  NAND2_X1 U7799 ( .A1(n7197), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7800 ( .A1(n8197), .A2(n5964), .ZN(n5965) );
  INV_X1 U7801 ( .A(n6035), .ZN(n8251) );
  OR2_X1 U7802 ( .A1(n5965), .A2(n8251), .ZN(n5966) );
  NAND2_X1 U7803 ( .A1(n5965), .A2(n8251), .ZN(n8288) );
  INV_X1 U7804 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9016) );
  OR2_X1 U7805 ( .A1(n8294), .A2(n9016), .ZN(n5967) );
  INV_X1 U7806 ( .A(n8633), .ZN(n7274) );
  XNOR2_X1 U7807 ( .A(n6039), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8648) );
  INV_X1 U7808 ( .A(n6039), .ZN(n8645) );
  NAND2_X1 U7809 ( .A1(n8645), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5970) );
  INV_X1 U7810 ( .A(n5972), .ZN(n8676) );
  INV_X1 U7811 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7812 ( .A(n6043), .B(n5973), .ZN(n8677) );
  NAND2_X1 U7813 ( .A1(n8695), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8694) );
  INV_X1 U7814 ( .A(n5974), .ZN(n8711) );
  OR2_X1 U7815 ( .A1(n8727), .A2(n10517), .ZN(n5976) );
  NAND2_X1 U7816 ( .A1(n8727), .A2(n10517), .ZN(n5975) );
  NAND2_X1 U7817 ( .A1(n5976), .A2(n5975), .ZN(n8710) );
  INV_X1 U7818 ( .A(n5976), .ZN(n5977) );
  NOR2_X1 U7819 ( .A1(n8713), .A2(n5977), .ZN(n5978) );
  XOR2_X1 U7820 ( .A(n6051), .B(n5978), .Z(n6068) );
  NOR2_X1 U7821 ( .A1(n5841), .A2(P2_U3151), .ZN(n9110) );
  NAND2_X1 U7822 ( .A1(n6057), .A2(n9110), .ZN(n7300) );
  OR2_X1 U7823 ( .A1(n7300), .A2(n6010), .ZN(n8734) );
  NAND2_X1 U7824 ( .A1(n5107), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7825 ( .A1(n7353), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7352) );
  INV_X1 U7826 ( .A(n5980), .ZN(n5981) );
  NAND2_X1 U7827 ( .A1(n7352), .A2(n5981), .ZN(n8615) );
  NAND2_X1 U7828 ( .A1(n8615), .A2(n8616), .ZN(n8614) );
  NAND2_X1 U7829 ( .A1(n7163), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7830 ( .A1(n7311), .A2(n7308), .ZN(n5984) );
  INV_X1 U7831 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7832 ( .A(n7325), .B(n5983), .ZN(n7309) );
  NAND2_X1 U7833 ( .A1(n5984), .A2(n7309), .ZN(n7312) );
  NAND2_X1 U7834 ( .A1(n7325), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5985) );
  INV_X1 U7835 ( .A(n5988), .ZN(n5987) );
  INV_X1 U7836 ( .A(n7168), .ZN(n5986) );
  XNOR2_X1 U7837 ( .A(n7179), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7556) );
  OR2_X1 U7838 ( .A1(n7179), .A2(n7934), .ZN(n5990) );
  NAND2_X1 U7839 ( .A1(n7561), .A2(n5990), .ZN(n5991) );
  XNOR2_X1 U7840 ( .A(n7964), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U7841 ( .A1(n7198), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5993) );
  XNOR2_X1 U7842 ( .A(n8200), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U7843 ( .A1(n5994), .A2(n8202), .ZN(n8204) );
  NAND2_X1 U7844 ( .A1(n7197), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7845 ( .A1(n5996), .A2(n8251), .ZN(n8296) );
  XNOR2_X1 U7846 ( .A(n8294), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8297) );
  OR2_X1 U7847 ( .A1(n8294), .A2(n5998), .ZN(n5999) );
  NAND2_X1 U7848 ( .A1(n8636), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8635) );
  XNOR2_X1 U7849 ( .A(n6039), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U7850 ( .A1(n8645), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6001) );
  AOI21_X1 U7851 ( .B1(n6002), .B2(n7490), .A(n6003), .ZN(n8671) );
  NAND2_X1 U7852 ( .A1(n8671), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8689) );
  INV_X1 U7853 ( .A(n6003), .ZN(n8687) );
  INV_X1 U7854 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7855 ( .A(n6043), .B(n6004), .ZN(n8688) );
  INV_X1 U7856 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8869) );
  OR2_X1 U7857 ( .A1(n8727), .A2(n8869), .ZN(n6006) );
  NAND2_X1 U7858 ( .A1(n8727), .A2(n8869), .ZN(n6005) );
  NAND2_X1 U7859 ( .A1(n6006), .A2(n6005), .ZN(n8728) );
  AOI21_X1 U7860 ( .B1(n8729), .B2(n4461), .A(n8728), .ZN(n8732) );
  INV_X1 U7861 ( .A(n6006), .ZN(n6007) );
  NOR2_X1 U7862 ( .A1(n8732), .A2(n6007), .ZN(n6008) );
  XNOR2_X1 U7863 ( .A(n5854), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6050) );
  XNOR2_X1 U7864 ( .A(n6008), .B(n6050), .ZN(n6009) );
  OR2_X1 U7865 ( .A1(n7300), .A2(n6298), .ZN(n8655) );
  NOR2_X1 U7866 ( .A1(n6009), .A2(n8655), .ZN(n6066) );
  MUX2_X1 U7867 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6298), .Z(n6026) );
  INV_X1 U7868 ( .A(n6026), .ZN(n6027) );
  MUX2_X1 U7869 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6298), .Z(n6024) );
  INV_X1 U7870 ( .A(n6024), .ZN(n6025) );
  MUX2_X1 U7871 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6298), .Z(n6022) );
  INV_X1 U7872 ( .A(n6022), .ZN(n6023) );
  INV_X1 U7873 ( .A(n7325), .ZN(n6021) );
  MUX2_X1 U7874 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6298), .Z(n6019) );
  INV_X1 U7875 ( .A(n6019), .ZN(n6020) );
  MUX2_X1 U7876 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5842), .Z(n6017) );
  INV_X1 U7877 ( .A(n6017), .ZN(n6018) );
  INV_X1 U7878 ( .A(n6015), .ZN(n6016) );
  INV_X1 U7879 ( .A(n6011), .ZN(n6013) );
  XNOR2_X1 U7880 ( .A(n6014), .B(n6011), .ZN(n7347) );
  NAND2_X1 U7881 ( .A1(n7298), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7348) );
  XNOR2_X1 U7882 ( .A(n6015), .B(n8619), .ZN(n8621) );
  XNOR2_X1 U7883 ( .A(n6017), .B(n7166), .ZN(n7332) );
  XOR2_X1 U7884 ( .A(n7325), .B(n6019), .Z(n7306) );
  XOR2_X1 U7885 ( .A(n7168), .B(n6022), .Z(n7429) );
  XOR2_X1 U7886 ( .A(n7179), .B(n6024), .Z(n7553) );
  XOR2_X1 U7887 ( .A(n6028), .B(n6026), .Z(n7756) );
  MUX2_X1 U7888 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6298), .Z(n6029) );
  XOR2_X1 U7889 ( .A(n7964), .B(n6029), .Z(n7954) );
  MUX2_X1 U7890 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6298), .Z(n6030) );
  XNOR2_X1 U7891 ( .A(n6030), .B(n8083), .ZN(n8074) );
  INV_X1 U7892 ( .A(n6030), .ZN(n6031) );
  MUX2_X1 U7893 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6298), .Z(n6032) );
  XOR2_X1 U7894 ( .A(n8200), .B(n6032), .Z(n8190) );
  MUX2_X1 U7895 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6298), .Z(n6033) );
  XNOR2_X1 U7896 ( .A(n6033), .B(n6035), .ZN(n8249) );
  INV_X1 U7897 ( .A(n6033), .ZN(n6034) );
  MUX2_X1 U7898 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6298), .Z(n6036) );
  XOR2_X1 U7899 ( .A(n8294), .B(n6036), .Z(n8286) );
  INV_X1 U7900 ( .A(n8294), .ZN(n7208) );
  MUX2_X1 U7901 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6298), .Z(n6037) );
  XNOR2_X1 U7902 ( .A(n6037), .B(n8633), .ZN(n8628) );
  INV_X1 U7903 ( .A(n6037), .ZN(n6038) );
  MUX2_X1 U7904 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6298), .Z(n6040) );
  XOR2_X1 U7905 ( .A(n6039), .B(n6040), .Z(n8644) );
  MUX2_X1 U7906 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6298), .Z(n6041) );
  XNOR2_X1 U7907 ( .A(n7490), .B(n6041), .ZN(n8665) );
  INV_X1 U7908 ( .A(n6041), .ZN(n6042) );
  MUX2_X1 U7909 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6298), .Z(n6044) );
  XOR2_X1 U7910 ( .A(n6043), .B(n6044), .Z(n8680) );
  MUX2_X1 U7911 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n6298), .Z(n6045) );
  XNOR2_X1 U7912 ( .A(n6045), .B(n6047), .ZN(n8697) );
  INV_X1 U7913 ( .A(n6045), .ZN(n6046) );
  MUX2_X1 U7914 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6298), .Z(n6048) );
  NAND2_X1 U7915 ( .A1(n6049), .A2(n6048), .ZN(n8714) );
  OAI21_X1 U7916 ( .B1(n8716), .B2(n8727), .A(n8714), .ZN(n6054) );
  INV_X1 U7917 ( .A(n6050), .ZN(n6052) );
  MUX2_X1 U7918 ( .A(n6052), .B(n6051), .S(n6298), .Z(n6053) );
  XNOR2_X1 U7919 ( .A(n6054), .B(n6053), .ZN(n6056) );
  INV_X1 U7920 ( .A(n7241), .ZN(n6055) );
  OR2_X2 U7921 ( .A1(n7373), .A2(n6055), .ZN(n8718) );
  NOR2_X1 U7922 ( .A1(n8718), .A2(n6299), .ZN(n8704) );
  NOR2_X1 U7923 ( .A1(n6298), .A2(P2_U3151), .ZN(n9114) );
  NAND2_X1 U7924 ( .A1(n6057), .A2(n9114), .ZN(n6058) );
  MUX2_X1 U7925 ( .A(n8718), .B(n6058), .S(n5841), .Z(n8717) );
  INV_X1 U7926 ( .A(n7372), .ZN(n6059) );
  NOR2_X1 U7927 ( .A1(n7373), .A2(n6059), .ZN(n6060) );
  OR2_X1 U7928 ( .A1(P2_U3150), .A2(n6060), .ZN(n8721) );
  INV_X1 U7929 ( .A(n8721), .ZN(n8699) );
  NOR2_X1 U7930 ( .A1(n10589), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8450) );
  AOI21_X1 U7931 ( .B1(n8699), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8450), .ZN(
        n6061) );
  OAI21_X1 U7932 ( .B1(n4428), .B2(n8717), .A(n6061), .ZN(n6062) );
  INV_X1 U7933 ( .A(n6062), .ZN(n6063) );
  OAI21_X1 U7934 ( .B1(n6068), .B2(n8734), .A(n6067), .ZN(P2_U3201) );
  INV_X1 U7935 ( .A(n6236), .ZN(n6082) );
  INV_X1 U7936 ( .A(SI_29_), .ZN(n10613) );
  NAND2_X1 U7937 ( .A1(n6070), .A2(n6069), .ZN(n6073) );
  NAND3_X1 U7938 ( .A1(n6073), .A2(n6072), .A3(n6071), .ZN(n6074) );
  INV_X1 U7939 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8338) );
  INV_X1 U7940 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8406) );
  MUX2_X1 U7941 ( .A(n8338), .B(n8406), .S(n7161), .Z(n6076) );
  INV_X1 U7942 ( .A(SI_30_), .ZN(n10587) );
  NAND2_X1 U7943 ( .A1(n6076), .A2(n10587), .ZN(n6097) );
  INV_X1 U7944 ( .A(n6076), .ZN(n6077) );
  NAND2_X1 U7945 ( .A1(n6077), .A2(SI_30_), .ZN(n6078) );
  NAND2_X1 U7946 ( .A1(n6097), .A2(n6078), .ZN(n6098) );
  XNOR2_X1 U7947 ( .A(n6099), .B(n6098), .ZN(n7102) );
  NAND2_X1 U7948 ( .A1(n7102), .A2(n6106), .ZN(n6080) );
  OR2_X1 U7949 ( .A1(n4405), .A2(n8406), .ZN(n6079) );
  INV_X1 U7950 ( .A(n8599), .ZN(n6084) );
  NAND2_X1 U7951 ( .A1(n6085), .A2(n6084), .ZN(n6271) );
  AOI21_X1 U7952 ( .B1(n6096), .B2(n6272), .A(n7386), .ZN(n6283) );
  INV_X1 U7953 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7954 ( .A1(n6086), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6089) );
  INV_X1 U7955 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6087) );
  OR2_X1 U7956 ( .A1(n4424), .A2(n6087), .ZN(n6088) );
  OAI211_X1 U7957 ( .C1(n6091), .C2(n6090), .A(n6089), .B(n6088), .ZN(n6092)
         );
  INV_X1 U7958 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7959 ( .A1(n6094), .A2(n6093), .ZN(n8737) );
  NAND2_X1 U7960 ( .A1(n8737), .A2(n5854), .ZN(n6286) );
  OR2_X1 U7961 ( .A1(n6085), .A2(n7386), .ZN(n6095) );
  INV_X1 U7962 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10105) );
  INV_X1 U7963 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6103) );
  MUX2_X1 U7964 ( .A(n10105), .B(n6103), .S(n7161), .Z(n6100) );
  XNOR2_X1 U7965 ( .A(n6100), .B(SI_31_), .ZN(n6101) );
  NOR2_X1 U7966 ( .A1(n4406), .A2(n6103), .ZN(n6105) );
  NAND2_X1 U7967 ( .A1(n9021), .A2(n5854), .ZN(n6107) );
  OAI22_X1 U7968 ( .A1(n6283), .A2(n6286), .B1(n6281), .B2(n6107), .ZN(n6108)
         );
  INV_X1 U7969 ( .A(n6108), .ZN(n6277) );
  NAND2_X1 U7970 ( .A1(n6109), .A2(n7427), .ZN(n6251) );
  NAND2_X1 U7971 ( .A1(n6251), .A2(n6274), .ZN(n6110) );
  NAND2_X1 U7972 ( .A1(n6110), .A2(n6241), .ZN(n6112) );
  NAND3_X1 U7973 ( .A1(n6116), .A2(n6251), .A3(n6301), .ZN(n6111) );
  NAND2_X1 U7974 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  OAI21_X1 U7975 ( .B1(n6274), .B2(n7713), .A(n6113), .ZN(n6115) );
  MUX2_X2 U7976 ( .A(n6241), .B(n6115), .S(n5815), .Z(n6119) );
  NOR2_X1 U7977 ( .A1(n6116), .A2(n6237), .ZN(n6117) );
  NOR2_X1 U7978 ( .A1(n7615), .A2(n6117), .ZN(n6118) );
  NAND2_X1 U7979 ( .A1(n6140), .A2(n6120), .ZN(n6125) );
  NAND2_X1 U7980 ( .A1(n10276), .A2(n7521), .ZN(n6129) );
  NAND2_X1 U7981 ( .A1(n10287), .A2(n10302), .ZN(n6122) );
  NAND2_X1 U7982 ( .A1(n6129), .A2(n6122), .ZN(n6123) );
  NAND2_X1 U7983 ( .A1(n10285), .A2(n7573), .ZN(n6142) );
  MUX2_X1 U7984 ( .A(n6142), .B(n6130), .S(n6237), .Z(n6127) );
  INV_X1 U7985 ( .A(n6129), .ZN(n6131) );
  INV_X1 U7986 ( .A(n6141), .ZN(n6133) );
  NAND2_X1 U7987 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  NAND2_X1 U7988 ( .A1(n6135), .A2(n10258), .ZN(n6139) );
  AND2_X1 U7989 ( .A1(n8233), .A2(n6136), .ZN(n6138) );
  INV_X1 U7990 ( .A(n6140), .ZN(n6143) );
  OAI211_X1 U7991 ( .C1(n6144), .C2(n6143), .A(n6142), .B(n6141), .ZN(n6146)
         );
  NAND2_X1 U7992 ( .A1(n6146), .A2(n6145), .ZN(n6149) );
  NAND2_X1 U7993 ( .A1(n6149), .A2(n6148), .ZN(n6151) );
  AND4_X1 U7994 ( .A1(n6156), .A2(n6237), .A3(n6256), .A4(n6249), .ZN(n6153)
         );
  NAND2_X1 U7995 ( .A1(n6154), .A2(n6153), .ZN(n6163) );
  NAND4_X1 U7996 ( .A1(n6155), .A2(n8554), .A3(n8444), .A4(n6241), .ZN(n6161)
         );
  INV_X1 U7997 ( .A(n8444), .ZN(n8343) );
  NAND4_X1 U7998 ( .A1(n6156), .A2(n8343), .A3(n6237), .A4(n8604), .ZN(n6160)
         );
  NOR2_X1 U7999 ( .A1(n8473), .A2(n6241), .ZN(n6158) );
  OAI21_X1 U8000 ( .B1(n6237), .B2(n8603), .A(n8548), .ZN(n6157) );
  OAI21_X1 U8001 ( .B1(n6158), .B2(n8548), .A(n6157), .ZN(n6159) );
  AND3_X1 U8002 ( .A1(n6161), .A2(n6160), .A3(n6159), .ZN(n6162) );
  XNOR2_X1 U8003 ( .A(n8482), .B(n8931), .ZN(n7148) );
  MUX2_X1 U8004 ( .A(n6237), .B(n8352), .S(n8482), .Z(n6164) );
  OAI21_X1 U8005 ( .B1(n6241), .B2(n8931), .A(n6164), .ZN(n6165) );
  INV_X1 U8006 ( .A(n6248), .ZN(n6169) );
  MUX2_X1 U8007 ( .A(n6167), .B(n8477), .S(n6241), .Z(n6168) );
  NAND2_X1 U8008 ( .A1(n6170), .A2(n4479), .ZN(n6171) );
  OR2_X1 U8009 ( .A1(n6172), .A2(n4488), .ZN(n8926) );
  MUX2_X1 U8010 ( .A(n4488), .B(n6172), .S(n6237), .Z(n6173) );
  NAND2_X1 U8011 ( .A1(n6185), .A2(n6176), .ZN(n6264) );
  NAND2_X1 U8012 ( .A1(n6264), .A2(n6237), .ZN(n6177) );
  NAND2_X1 U8013 ( .A1(n6181), .A2(n6241), .ZN(n6182) );
  NAND2_X1 U8014 ( .A1(n6186), .A2(n6182), .ZN(n6183) );
  NAND2_X1 U8015 ( .A1(n6184), .A2(n6188), .ZN(n6194) );
  INV_X1 U8016 ( .A(n6185), .ZN(n6187) );
  AND2_X1 U8017 ( .A1(n6195), .A2(n6188), .ZN(n6191) );
  NOR2_X1 U8018 ( .A1(n8843), .A2(n5119), .ZN(n6190) );
  MUX2_X1 U8019 ( .A(n6191), .B(n6190), .S(n6241), .Z(n6192) );
  AND2_X1 U8020 ( .A1(n6201), .A2(n6195), .ZN(n6198) );
  AND2_X1 U8021 ( .A1(n8797), .A2(n6196), .ZN(n6197) );
  MUX2_X1 U8022 ( .A(n6198), .B(n6197), .S(n6237), .Z(n6199) );
  NAND2_X1 U8023 ( .A1(n6200), .A2(n6199), .ZN(n6203) );
  XNOR2_X1 U8024 ( .A(n8825), .B(n8834), .ZN(n8820) );
  MUX2_X1 U8025 ( .A(n6201), .B(n8797), .S(n6241), .Z(n6202) );
  INV_X1 U8026 ( .A(n6204), .ZN(n6205) );
  NAND2_X1 U8027 ( .A1(n6245), .A2(n6205), .ZN(n6207) );
  NAND2_X1 U8028 ( .A1(n6246), .A2(n8799), .ZN(n6206) );
  MUX2_X1 U8029 ( .A(n6207), .B(n6206), .S(n6237), .Z(n6208) );
  INV_X1 U8030 ( .A(n6208), .ZN(n6209) );
  INV_X1 U8031 ( .A(n6245), .ZN(n6210) );
  NOR2_X1 U8032 ( .A1(n6215), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U8033 ( .A1(n6243), .A2(n6237), .ZN(n6211) );
  INV_X1 U8034 ( .A(n6215), .ZN(n6244) );
  NAND3_X1 U8035 ( .A1(n6216), .A2(n6244), .A3(n6241), .ZN(n6217) );
  MUX2_X1 U8036 ( .A(n6222), .B(n6221), .S(n6241), .Z(n6223) );
  NAND2_X1 U8037 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U8038 ( .A1(n6225), .A2(n8753), .ZN(n6232) );
  MUX2_X1 U8039 ( .A(n8757), .B(n8951), .S(n6241), .Z(n6233) );
  MUX2_X1 U8040 ( .A(n6227), .B(n6226), .S(n6241), .Z(n6231) );
  OR2_X1 U8041 ( .A1(n6233), .A2(n6231), .ZN(n6230) );
  AND2_X1 U8042 ( .A1(n8757), .A2(n6241), .ZN(n6228) );
  AOI21_X1 U8043 ( .B1(n8951), .B2(n6237), .A(n6228), .ZN(n6229) );
  INV_X1 U8044 ( .A(n6234), .ZN(n6235) );
  NAND2_X1 U8045 ( .A1(n6272), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U8046 ( .A1(n6272), .A2(n6241), .ZN(n6240) );
  NAND2_X1 U8047 ( .A1(n6246), .A2(n6245), .ZN(n8805) );
  INV_X1 U8048 ( .A(n8820), .ZN(n6269) );
  INV_X1 U8049 ( .A(n6247), .ZN(n6266) );
  OR2_X1 U8050 ( .A1(n6248), .A2(n4479), .ZN(n8939) );
  INV_X1 U8051 ( .A(n8345), .ZN(n8347) );
  AND2_X1 U8052 ( .A1(n8233), .A2(n6249), .ZN(n8132) );
  INV_X1 U8053 ( .A(n6250), .ZN(n7715) );
  AND2_X1 U8054 ( .A1(n7713), .A2(n6251), .ZN(n7421) );
  NAND2_X1 U8055 ( .A1(n7895), .A2(n7923), .ZN(n7897) );
  NAND4_X1 U8056 ( .A1(n7715), .A2(n10258), .A3(n7421), .A4(n7897), .ZN(n6255)
         );
  XNOR2_X1 U8057 ( .A(n10257), .B(n10324), .ZN(n7926) );
  NAND2_X1 U8058 ( .A1(n6252), .A2(n7926), .ZN(n6254) );
  NAND2_X1 U8059 ( .A1(n10291), .A2(n10279), .ZN(n6253) );
  NOR3_X1 U8060 ( .A1(n6255), .A2(n6254), .A3(n6253), .ZN(n6258) );
  AND2_X1 U8061 ( .A1(n6257), .A2(n6256), .ZN(n8236) );
  AND4_X1 U8062 ( .A1(n8132), .A2(n6258), .A3(n8236), .A4(n7944), .ZN(n6259)
         );
  NAND4_X1 U8063 ( .A1(n8939), .A2(n8347), .A3(n6259), .A4(n7148), .ZN(n6260)
         );
  NOR2_X1 U8064 ( .A1(n8926), .A2(n6260), .ZN(n6262) );
  NAND3_X1 U8065 ( .A1(n6263), .A2(n6262), .A3(n6261), .ZN(n6265) );
  NOR3_X1 U8066 ( .A1(n8805), .A2(n6269), .A3(n6268), .ZN(n6270) );
  INV_X1 U8067 ( .A(n9021), .ZN(n6282) );
  INV_X1 U8068 ( .A(n8737), .ZN(n6278) );
  INV_X1 U8069 ( .A(n7385), .ZN(n6274) );
  INV_X1 U8070 ( .A(n6288), .ZN(n6276) );
  NOR3_X1 U8071 ( .A1(n6277), .A2(n6285), .A3(n6276), .ZN(n6303) );
  NAND2_X1 U8072 ( .A1(n6278), .A2(n4428), .ZN(n6290) );
  INV_X1 U8073 ( .A(n6290), .ZN(n6280) );
  NOR2_X1 U8074 ( .A1(n6288), .A2(n5854), .ZN(n6279) );
  NAND3_X1 U8075 ( .A1(n6283), .A2(n4428), .A3(n6282), .ZN(n6294) );
  INV_X1 U8076 ( .A(n6286), .ZN(n6287) );
  NOR2_X1 U8077 ( .A1(n7372), .A2(P2_U3151), .ZN(n6296) );
  OAI211_X1 U8078 ( .C1(n9021), .C2(n6290), .A(n6289), .B(n6296), .ZN(n6291)
         );
  INV_X1 U8079 ( .A(n6296), .ZN(n8246) );
  NOR2_X1 U8080 ( .A1(n6297), .A2(n7419), .ZN(n7380) );
  NAND3_X1 U8081 ( .A1(n7380), .A2(n6299), .A3(n6298), .ZN(n6300) );
  OAI211_X1 U8082 ( .C1(n6301), .C2(n8246), .A(n6300), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6302) );
  NOR2_X1 U8083 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6307) );
  NOR2_X2 U8084 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6306) );
  NOR2_X2 U8085 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6305) );
  NOR2_X2 U8086 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6304) );
  NOR2_X2 U8087 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6411) );
  INV_X1 U8088 ( .A(n10102), .ZN(n6317) );
  NOR2_X1 U8089 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6316) );
  AOI21_X1 U8090 ( .B1(n6317), .B2(n6316), .A(n6651), .ZN(n6319) );
  INV_X1 U8091 ( .A(n6319), .ZN(n6318) );
  INV_X1 U8092 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U8093 ( .A1(n6318), .A2(n10391), .ZN(n6321) );
  INV_X1 U8094 ( .A(n8336), .ZN(n6324) );
  NAND2_X1 U8095 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6322) );
  NAND2_X1 U8096 ( .A1(n6355), .A2(n6322), .ZN(n6323) );
  INV_X1 U8097 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10103) );
  XNOR2_X2 U8098 ( .A(n6323), .B(n10103), .ZN(n6326) );
  INV_X1 U8099 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U8100 ( .A1(n6937), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6332) );
  INV_X1 U8101 ( .A(n6326), .ZN(n8311) );
  INV_X1 U8102 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U8103 ( .A1(n6520), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6330) );
  INV_X1 U8104 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6328) );
  NAND4_X2 U8105 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n7007)
         );
  NAND2_X1 U8106 ( .A1(n4455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6333) );
  INV_X1 U8107 ( .A(n6334), .ZN(n6335) );
  NAND2_X1 U8108 ( .A1(n6337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8109 ( .A1(n6339), .A2(n4455), .ZN(n10118) );
  NAND2_X1 U8110 ( .A1(n5040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6342) );
  XNOR2_X1 U8111 ( .A(n6342), .B(n6341), .ZN(n8310) );
  INV_X1 U8112 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6344) );
  INV_X1 U8113 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8114 ( .A1(n4467), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6350) );
  MUX2_X1 U8115 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6350), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6351) );
  INV_X1 U8116 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7159) );
  INV_X1 U8117 ( .A(SI_0_), .ZN(n6352) );
  NOR2_X1 U8118 ( .A1(n7161), .A2(n6352), .ZN(n6353) );
  XNOR2_X1 U8119 ( .A(n6353), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n7158) );
  INV_X1 U8120 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6354) );
  MUX2_X2 U8121 ( .A(n7159), .B(n7158), .S(n4421), .Z(n9527) );
  INV_X1 U8122 ( .A(n7156), .ZN(n6359) );
  NAND2_X1 U8123 ( .A1(n6359), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8124 ( .A1(n6379), .A2(n6360), .ZN(n7279) );
  NAND2_X1 U8125 ( .A1(n6363), .A2(n6362), .ZN(n6364) );
  NAND2_X1 U8126 ( .A1(n6364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6366) );
  OR2_X1 U8127 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  NAND2_X1 U8128 ( .A1(n6366), .A2(n6365), .ZN(n6973) );
  NAND2_X1 U8129 ( .A1(n4495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8130 ( .A1(n6776), .A2(n6368), .ZN(n6369) );
  NAND2_X1 U8131 ( .A1(n6369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6371) );
  XNOR2_X2 U8132 ( .A(n6371), .B(n6370), .ZN(n9629) );
  NAND2_X1 U8133 ( .A1(n7837), .A2(n9629), .ZN(n7003) );
  INV_X1 U8134 ( .A(n7003), .ZN(n9524) );
  NAND2_X1 U8135 ( .A1(n8177), .A2(n9524), .ZN(n6374) );
  NAND3_X1 U8136 ( .A1(n9451), .A2(n6372), .A3(n7837), .ZN(n7648) );
  NAND2_X1 U8137 ( .A1(n7007), .A2(n4423), .ZN(n6377) );
  OAI22_X1 U8138 ( .A1(n9527), .A2(n4427), .B1(n7159), .B2(n7156), .ZN(n6375)
         );
  INV_X1 U8139 ( .A(n6375), .ZN(n6376) );
  NAND2_X1 U8140 ( .A1(n6377), .A2(n6376), .ZN(n7278) );
  NAND2_X1 U8141 ( .A1(n9451), .A2(n9522), .ZN(n9447) );
  OAI21_X1 U8142 ( .B1(n9451), .B2(n9629), .A(n9447), .ZN(n6378) );
  NOR2_X2 U8143 ( .A1(n5181), .A2(n6378), .ZN(n6399) );
  INV_X1 U8144 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U8145 ( .A1(n6427), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8146 ( .A1(n6520), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8147 ( .A1(n6400), .A2(n4418), .ZN(n6398) );
  INV_X1 U8148 ( .A(n4429), .ZN(n7448) );
  AND2_X1 U8149 ( .A1(n7161), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6388) );
  OAI21_X1 U8150 ( .B1(n7448), .B2(n9518), .A(n6388), .ZN(n6392) );
  INV_X1 U8151 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8152 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6389) );
  OR2_X1 U8153 ( .A1(n4420), .A2(n7218), .ZN(n6391) );
  INV_X1 U8154 ( .A(n6394), .ZN(n7162) );
  NAND2_X1 U8155 ( .A1(n7006), .A2(n6418), .ZN(n6397) );
  AND2_X1 U8156 ( .A1(n7006), .A2(n4418), .ZN(n6401) );
  XNOR2_X1 U8157 ( .A(n6402), .B(n6403), .ZN(n7361) );
  NAND2_X1 U8158 ( .A1(n7362), .A2(n7361), .ZN(n7360) );
  INV_X1 U8159 ( .A(n6402), .ZN(n6404) );
  NAND2_X1 U8160 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  NAND2_X1 U8161 ( .A1(n7360), .A2(n6405), .ZN(n7439) );
  NAND2_X1 U8162 ( .A1(n6937), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6410) );
  INV_X1 U8163 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6406) );
  OR2_X1 U8164 ( .A1(n6463), .A2(n6406), .ZN(n6409) );
  NAND2_X1 U8165 ( .A1(n6520), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8166 ( .A1(n6427), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8167 ( .A1(n7009), .A2(n4418), .ZN(n6420) );
  NAND2_X1 U8168 ( .A1(n4420), .A2(n7161), .ZN(n6488) );
  OR2_X1 U8169 ( .A1(n6488), .A2(n7173), .ZN(n6417) );
  OR2_X1 U8170 ( .A1(n6650), .A2(n7174), .ZN(n6416) );
  INV_X1 U8171 ( .A(n6411), .ZN(n6412) );
  INV_X1 U8172 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6413) );
  OR2_X1 U8173 ( .A1(n4421), .A2(n7221), .ZN(n6415) );
  XNOR2_X1 U8174 ( .A(n6421), .B(n8316), .ZN(n6422) );
  INV_X1 U8175 ( .A(n10225), .ZN(n7740) );
  AOI22_X1 U8176 ( .A1(n7009), .A2(n6906), .B1(n7740), .B2(n8313), .ZN(n6423)
         );
  XNOR2_X1 U8177 ( .A(n6422), .B(n6423), .ZN(n7440) );
  NAND2_X1 U8178 ( .A1(n7439), .A2(n7440), .ZN(n6426) );
  INV_X1 U8179 ( .A(n6422), .ZN(n6424) );
  NAND2_X1 U8180 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  INV_X2 U8181 ( .A(n6512), .ZN(n7106) );
  NAND2_X1 U8182 ( .A1(n7106), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8183 ( .A1(n6384), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U8184 ( .A1(n4408), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6429) );
  INV_X1 U8185 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U8186 ( .A1(n6937), .A2(n7651), .ZN(n6428) );
  INV_X1 U8187 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7169) );
  OR2_X1 U8188 ( .A1(n6930), .A2(n7169), .ZN(n6437) );
  OR2_X1 U8189 ( .A1(n6650), .A2(n7170), .ZN(n6436) );
  NAND2_X1 U8190 ( .A1(n6432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6434) );
  INV_X1 U8191 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6433) );
  OR2_X1 U8192 ( .A1(n4420), .A2(n7222), .ZN(n6435) );
  AND3_X2 U8193 ( .A1(n6437), .A2(n6436), .A3(n6435), .ZN(n10231) );
  OR2_X1 U8194 ( .A1(n10231), .A2(n6537), .ZN(n6438) );
  NAND2_X1 U8195 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  XNOR2_X1 U8196 ( .A(n6440), .B(n8316), .ZN(n6441) );
  AOI22_X1 U8197 ( .A1(n9595), .A2(n6906), .B1(n7652), .B2(n8313), .ZN(n6442)
         );
  XNOR2_X1 U8198 ( .A(n6441), .B(n6442), .ZN(n7510) );
  INV_X1 U8199 ( .A(n6441), .ZN(n6443) );
  NAND2_X1 U8200 ( .A1(n6443), .A2(n6442), .ZN(n6444) );
  NAND2_X1 U8201 ( .A1(n6384), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6449) );
  OAI21_X1 U8202 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n6468), .ZN(n7678) );
  INV_X1 U8203 ( .A(n7678), .ZN(n7791) );
  NAND2_X1 U8204 ( .A1(n6937), .A2(n7791), .ZN(n6448) );
  NAND2_X1 U8205 ( .A1(n7106), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8206 ( .A1(n4408), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8207 ( .A1(n9594), .A2(n8313), .ZN(n6455) );
  OR2_X1 U8208 ( .A1(n6650), .A2(n7175), .ZN(n6453) );
  INV_X1 U8209 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7176) );
  OR2_X1 U8210 ( .A1(n6930), .A2(n7176), .ZN(n6452) );
  OR2_X1 U8211 ( .A1(n6475), .A2(n6651), .ZN(n6450) );
  XNOR2_X1 U8212 ( .A(n6450), .B(n6474), .ZN(n7249) );
  OR2_X1 U8213 ( .A1(n4421), .A2(n7249), .ZN(n6451) );
  OR2_X1 U8214 ( .A1(n7637), .A2(n6537), .ZN(n6454) );
  NAND2_X1 U8215 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  XNOR2_X1 U8216 ( .A(n6456), .B(n6947), .ZN(n6458) );
  AOI22_X1 U8217 ( .A1(n9594), .A2(n6906), .B1(n7781), .B2(n8313), .ZN(n6459)
         );
  XNOR2_X1 U8218 ( .A(n6458), .B(n6459), .ZN(n7788) );
  INV_X1 U8219 ( .A(n6458), .ZN(n6461) );
  INV_X1 U8220 ( .A(n6459), .ZN(n6460) );
  NAND2_X1 U8221 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  CLKBUF_X3 U8222 ( .A(n6463), .Z(n7125) );
  INV_X1 U8223 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U8224 ( .A1(n7106), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6464) );
  OAI21_X1 U8225 ( .B1(n7125), .B2(n7670), .A(n6464), .ZN(n6473) );
  INV_X1 U8226 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U8227 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U8228 ( .A1(n6498), .A2(n6469), .ZN(n7852) );
  INV_X1 U8229 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6470) );
  OR2_X1 U8230 ( .A1(n6982), .A2(n6470), .ZN(n6471) );
  OAI21_X1 U8231 ( .B1(n6465), .B2(n7852), .A(n6471), .ZN(n6472) );
  NAND2_X1 U8232 ( .A1(n6475), .A2(n6474), .ZN(n6489) );
  NAND2_X1 U8233 ( .A1(n6489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6477) );
  INV_X1 U8234 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6476) );
  XNOR2_X1 U8235 ( .A(n6477), .B(n6476), .ZN(n7251) );
  INV_X1 U8236 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7171) );
  OR2_X1 U8237 ( .A1(n6488), .A2(n7171), .ZN(n6479) );
  OR2_X1 U8238 ( .A1(n6650), .A2(n7172), .ZN(n6478) );
  OAI211_X1 U8239 ( .C1(n4420), .C2(n7251), .A(n6479), .B(n6478), .ZN(n7672)
         );
  OAI22_X1 U8240 ( .A1(n7812), .A2(n4427), .B1(n5051), .B2(n6537), .ZN(n6480)
         );
  XNOR2_X1 U8241 ( .A(n6480), .B(n8316), .ZN(n6484) );
  NAND2_X1 U8242 ( .A1(n6483), .A2(n6484), .ZN(n7841) );
  OR2_X1 U8243 ( .A1(n7812), .A2(n8318), .ZN(n6482) );
  NAND2_X1 U8244 ( .A1(n7672), .A2(n8313), .ZN(n6481) );
  AND2_X1 U8245 ( .A1(n6482), .A2(n6481), .ZN(n7844) );
  NAND2_X1 U8246 ( .A1(n7841), .A2(n7844), .ZN(n6487) );
  INV_X1 U8247 ( .A(n6484), .ZN(n6485) );
  NOR2_X1 U8248 ( .A1(n6489), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6533) );
  INV_X1 U8249 ( .A(n6533), .ZN(n6490) );
  NAND2_X1 U8250 ( .A1(n6490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6493) );
  INV_X1 U8251 ( .A(n6493), .ZN(n6491) );
  NAND2_X1 U8252 ( .A1(n6491), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6494) );
  INV_X1 U8253 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U8254 ( .A1(n6493), .A2(n6492), .ZN(n6526) );
  AOI22_X1 U8255 ( .A1(n6778), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6777), .B2(
        n7290), .ZN(n6496) );
  NAND2_X1 U8256 ( .A1(n7177), .A2(n7103), .ZN(n6495) );
  NAND2_X1 U8257 ( .A1(n6384), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6503) );
  INV_X1 U8258 ( .A(n6516), .ZN(n6518) );
  NAND2_X1 U8259 ( .A1(n6498), .A2(n6497), .ZN(n6499) );
  AND2_X1 U8260 ( .A1(n6518), .A2(n6499), .ZN(n7815) );
  NAND2_X1 U8261 ( .A1(n6937), .A2(n7815), .ZN(n6502) );
  NAND2_X1 U8262 ( .A1(n7106), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U8263 ( .A1(n4408), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8264 ( .A1(n9592), .A2(n8313), .ZN(n6504) );
  OAI21_X1 U8265 ( .B1(n7811), .B2(n6537), .A(n6504), .ZN(n6505) );
  XNOR2_X1 U8266 ( .A(n6505), .B(n6947), .ZN(n6508) );
  INV_X1 U8267 ( .A(n7811), .ZN(n7730) );
  NAND2_X1 U8268 ( .A1(n7730), .A2(n8313), .ZN(n6507) );
  NAND2_X1 U8269 ( .A1(n9592), .A2(n6906), .ZN(n6506) );
  AND2_X1 U8270 ( .A1(n6507), .A2(n6506), .ZN(n6509) );
  INV_X1 U8271 ( .A(n6508), .ZN(n6511) );
  INV_X1 U8272 ( .A(n6509), .ZN(n6510) );
  NAND2_X1 U8273 ( .A1(n6511), .A2(n6510), .ZN(n7807) );
  INV_X1 U8274 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6514) );
  INV_X1 U8275 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7913) );
  OR2_X1 U8276 ( .A1(n7122), .A2(n7913), .ZN(n6513) );
  OAI21_X1 U8277 ( .B1(n7125), .B2(n6514), .A(n6513), .ZN(n6515) );
  INV_X1 U8278 ( .A(n6515), .ZN(n6525) );
  INV_X1 U8279 ( .A(n6539), .ZN(n6541) );
  INV_X1 U8280 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8281 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  NAND2_X1 U8282 ( .A1(n6541), .A2(n6519), .ZN(n7827) );
  INV_X2 U8283 ( .A(n6520), .ZN(n6982) );
  INV_X1 U8284 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6521) );
  OR2_X1 U8285 ( .A1(n6982), .A2(n6521), .ZN(n6522) );
  OAI21_X1 U8286 ( .B1(n6465), .B2(n7827), .A(n6522), .ZN(n6523) );
  INV_X1 U8287 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U8288 ( .A1(n6526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6527) );
  XNOR2_X1 U8289 ( .A(n6527), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7468) );
  AOI22_X1 U8290 ( .A1(n6778), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6777), .B2(
        n7468), .ZN(n6528) );
  NAND2_X1 U8291 ( .A1(n7917), .A2(n8313), .ZN(n6529) );
  OAI21_X1 U8292 ( .B1(n7021), .B2(n8318), .A(n6529), .ZN(n7868) );
  NAND2_X1 U8293 ( .A1(n7917), .A2(n6933), .ZN(n6530) );
  OAI21_X1 U8294 ( .B1(n7021), .B2(n4427), .A(n6530), .ZN(n6531) );
  XNOR2_X1 U8295 ( .A(n6531), .B(n8316), .ZN(n7867) );
  NAND2_X1 U8296 ( .A1(n7190), .A2(n7103), .ZN(n6536) );
  NOR2_X1 U8297 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6532) );
  NAND2_X1 U8298 ( .A1(n6533), .A2(n6532), .ZN(n6553) );
  NAND2_X1 U8299 ( .A1(n6553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6534) );
  AOI22_X1 U8300 ( .A1(n6778), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6777), .B2(
        n7541), .ZN(n6535) );
  NAND2_X2 U8301 ( .A1(n6536), .A2(n6535), .ZN(n9183) );
  NAND2_X1 U8302 ( .A1(n9183), .A2(n6933), .ZN(n6548) );
  INV_X1 U8303 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U8304 ( .A1(n7106), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6538) );
  OAI21_X1 U8305 ( .B1(n7125), .B2(n7885), .A(n6538), .ZN(n6546) );
  INV_X1 U8306 ( .A(n6558), .ZN(n6560) );
  INV_X1 U8307 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U8308 ( .A1(n6541), .A2(n6540), .ZN(n6542) );
  NAND2_X1 U8309 ( .A1(n6560), .A2(n6542), .ZN(n9176) );
  INV_X1 U8310 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6543) );
  OR2_X1 U8311 ( .A1(n6982), .A2(n6543), .ZN(n6544) );
  OAI21_X1 U8312 ( .B1(n6465), .B2(n9176), .A(n6544), .ZN(n6545) );
  OR2_X1 U8313 ( .A1(n9257), .A2(n4427), .ZN(n6547) );
  NAND2_X1 U8314 ( .A1(n6548), .A2(n6547), .ZN(n6549) );
  XNOR2_X1 U8315 ( .A(n6549), .B(n6947), .ZN(n9171) );
  NAND2_X1 U8316 ( .A1(n9183), .A2(n8313), .ZN(n6551) );
  OR2_X1 U8317 ( .A1(n9257), .A2(n8318), .ZN(n6550) );
  AND2_X1 U8318 ( .A1(n6551), .A2(n6550), .ZN(n6569) );
  NAND2_X1 U8319 ( .A1(n9171), .A2(n6569), .ZN(n6552) );
  NAND2_X1 U8320 ( .A1(n7201), .A2(n7103), .ZN(n6556) );
  NAND2_X1 U8321 ( .A1(n6577), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U8322 ( .A(n6554), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7773) );
  AOI22_X1 U8323 ( .A1(n6778), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6777), .B2(
        n7773), .ZN(n6555) );
  NAND2_X1 U8324 ( .A1(n8070), .A2(n6933), .ZN(n6566) );
  INV_X1 U8325 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U8326 ( .A1(n7106), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6557) );
  OAI21_X1 U8327 ( .B1(n7125), .B2(n8004), .A(n6557), .ZN(n6564) );
  INV_X1 U8328 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8329 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  NAND2_X1 U8330 ( .A1(n6584), .A2(n6561), .ZN(n9258) );
  INV_X1 U8331 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7539) );
  OR2_X1 U8332 ( .A1(n6982), .A2(n7539), .ZN(n6562) );
  OAI21_X1 U8333 ( .B1(n6465), .B2(n9258), .A(n6562), .ZN(n6563) );
  OR2_X1 U8334 ( .A1(n9152), .A2(n4427), .ZN(n6565) );
  NAND2_X1 U8335 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  XNOR2_X1 U8336 ( .A(n6567), .B(n8316), .ZN(n6573) );
  NOR2_X1 U8337 ( .A1(n9152), .A2(n8318), .ZN(n6568) );
  AOI21_X1 U8338 ( .B1(n8070), .B2(n8313), .A(n6568), .ZN(n6574) );
  XNOR2_X1 U8339 ( .A(n6573), .B(n6574), .ZN(n9250) );
  INV_X1 U8340 ( .A(n9171), .ZN(n6570) );
  INV_X1 U8341 ( .A(n6569), .ZN(n9173) );
  NAND2_X1 U8342 ( .A1(n6570), .A2(n9173), .ZN(n6571) );
  INV_X1 U8343 ( .A(n6573), .ZN(n6575) );
  NAND2_X1 U8344 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  OR2_X1 U8345 ( .A1(n7196), .A2(n6650), .ZN(n6580) );
  NAND2_X1 U8346 ( .A1(n6578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6600) );
  XNOR2_X1 U8347 ( .A(n6600), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7858) );
  AOI22_X1 U8348 ( .A1(n6778), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6777), .B2(
        n7858), .ZN(n6579) );
  NAND2_X2 U8349 ( .A1(n6580), .A2(n6579), .ZN(n9157) );
  NAND2_X1 U8350 ( .A1(n9157), .A2(n6933), .ZN(n6592) );
  INV_X1 U8351 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7979) );
  INV_X1 U8352 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10634) );
  OR2_X1 U8353 ( .A1(n7122), .A2(n10634), .ZN(n6581) );
  OAI21_X1 U8354 ( .B1(n7125), .B2(n7979), .A(n6581), .ZN(n6582) );
  INV_X1 U8355 ( .A(n6582), .ZN(n6590) );
  NAND2_X1 U8356 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U8357 ( .A1(n6609), .A2(n6585), .ZN(n9155) );
  INV_X1 U8358 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6586) );
  OR2_X1 U8359 ( .A1(n6982), .A2(n6586), .ZN(n6587) );
  OAI21_X1 U8360 ( .B1(n6465), .B2(n9155), .A(n6587), .ZN(n6588) );
  INV_X1 U8361 ( .A(n6588), .ZN(n6589) );
  NAND2_X1 U8362 ( .A1(n9590), .A2(n8313), .ZN(n6591) );
  NAND2_X1 U8363 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  XNOR2_X1 U8364 ( .A(n6593), .B(n6947), .ZN(n6594) );
  NAND2_X1 U8365 ( .A1(n9157), .A2(n8313), .ZN(n6597) );
  NAND2_X1 U8366 ( .A1(n9590), .A2(n6906), .ZN(n6596) );
  NAND2_X1 U8367 ( .A1(n6597), .A2(n6596), .ZN(n9150) );
  INV_X1 U8368 ( .A(n9150), .ZN(n6598) );
  NAND2_X1 U8369 ( .A1(n9148), .A2(n9295), .ZN(n6625) );
  NAND2_X1 U8370 ( .A1(n7231), .A2(n7103), .ZN(n6604) );
  INV_X1 U8371 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8372 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  NAND2_X1 U8373 ( .A1(n6601), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6602) );
  XNOR2_X1 U8374 ( .A(n6602), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8097) );
  AOI22_X1 U8375 ( .A1(n6778), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6777), .B2(
        n8097), .ZN(n6603) );
  NAND2_X1 U8376 ( .A1(n7027), .A2(n6933), .ZN(n6617) );
  INV_X1 U8377 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8034) );
  INV_X1 U8378 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6605) );
  OR2_X1 U8379 ( .A1(n7122), .A2(n6605), .ZN(n6606) );
  OAI21_X1 U8380 ( .B1(n7125), .B2(n8034), .A(n6606), .ZN(n6607) );
  INV_X1 U8381 ( .A(n6607), .ZN(n6615) );
  INV_X1 U8382 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8383 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  NAND2_X1 U8384 ( .A1(n6632), .A2(n6610), .ZN(n9302) );
  INV_X1 U8385 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6611) );
  OR2_X1 U8386 ( .A1(n6982), .A2(n6611), .ZN(n6612) );
  OAI21_X1 U8387 ( .B1(n6465), .B2(n9302), .A(n6612), .ZN(n6613) );
  INV_X1 U8388 ( .A(n6613), .ZN(n6614) );
  NAND2_X1 U8389 ( .A1(n10054), .A2(n8313), .ZN(n6616) );
  NAND2_X1 U8390 ( .A1(n6617), .A2(n6616), .ZN(n6618) );
  XNOR2_X1 U8391 ( .A(n6618), .B(n6947), .ZN(n6620) );
  NOR2_X1 U8392 ( .A1(n9203), .A2(n8318), .ZN(n6619) );
  AOI21_X1 U8393 ( .B1(n7027), .B2(n8313), .A(n6619), .ZN(n6621) );
  NAND2_X1 U8394 ( .A1(n6620), .A2(n6621), .ZN(n9194) );
  INV_X1 U8395 ( .A(n6620), .ZN(n6623) );
  INV_X1 U8396 ( .A(n6621), .ZN(n6622) );
  NAND2_X1 U8397 ( .A1(n6623), .A2(n6622), .ZN(n6624) );
  NAND2_X1 U8398 ( .A1(n6625), .A2(n9296), .ZN(n9193) );
  NAND2_X1 U8399 ( .A1(n9193), .A2(n9194), .ZN(n6648) );
  NAND2_X1 U8400 ( .A1(n6626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6627) );
  XNOR2_X1 U8401 ( .A(n6627), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U8402 ( .A1(n6778), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6777), .B2(
        n9620), .ZN(n6628) );
  NAND2_X1 U8403 ( .A1(n10095), .A2(n6933), .ZN(n6640) );
  INV_X1 U8404 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8122) );
  INV_X1 U8405 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8095) );
  OR2_X1 U8406 ( .A1(n6982), .A2(n8095), .ZN(n6630) );
  OAI21_X1 U8407 ( .B1(n7125), .B2(n8122), .A(n6630), .ZN(n6631) );
  INV_X1 U8408 ( .A(n6631), .ZN(n6638) );
  NAND2_X1 U8409 ( .A1(n6632), .A2(n10500), .ZN(n6633) );
  NAND2_X1 U8410 ( .A1(n6660), .A2(n6633), .ZN(n9200) );
  INV_X1 U8411 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6634) );
  OR2_X1 U8412 ( .A1(n7122), .A2(n6634), .ZN(n6635) );
  OAI21_X1 U8413 ( .B1(n6465), .B2(n9200), .A(n6635), .ZN(n6636) );
  INV_X1 U8414 ( .A(n6636), .ZN(n6637) );
  INV_X1 U8415 ( .A(n9911), .ZN(n9589) );
  NAND2_X1 U8416 ( .A1(n9589), .A2(n8313), .ZN(n6639) );
  NAND2_X1 U8417 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  XNOR2_X1 U8418 ( .A(n6641), .B(n6947), .ZN(n6643) );
  NOR2_X1 U8419 ( .A1(n9911), .A2(n8318), .ZN(n6642) );
  AOI21_X1 U8420 ( .B1(n10095), .B2(n8313), .A(n6642), .ZN(n6644) );
  NAND2_X1 U8421 ( .A1(n6643), .A2(n6644), .ZN(n6649) );
  INV_X1 U8422 ( .A(n6643), .ZN(n6646) );
  INV_X1 U8423 ( .A(n6644), .ZN(n6645) );
  NAND2_X1 U8424 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  NOR2_X1 U8425 ( .A1(n6626), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6676) );
  OR2_X1 U8426 ( .A1(n6676), .A2(n6651), .ZN(n6652) );
  XNOR2_X1 U8427 ( .A(n6652), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U8428 ( .A1(n6778), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6777), .B2(
        n10136), .ZN(n6653) );
  NAND2_X1 U8429 ( .A1(n10048), .A2(n6933), .ZN(n6668) );
  INV_X1 U8430 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6657) );
  INV_X1 U8431 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6655) );
  OR2_X1 U8432 ( .A1(n7122), .A2(n6655), .ZN(n6656) );
  OAI21_X1 U8433 ( .B1(n7125), .B2(n6657), .A(n6656), .ZN(n6658) );
  INV_X1 U8434 ( .A(n6658), .ZN(n6666) );
  INV_X1 U8435 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6659) );
  INV_X1 U8436 ( .A(n6681), .ZN(n6683) );
  NAND2_X1 U8437 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  NAND2_X1 U8438 ( .A1(n6683), .A2(n6661), .ZN(n9922) );
  INV_X1 U8439 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6662) );
  OR2_X1 U8440 ( .A1(n6982), .A2(n6662), .ZN(n6663) );
  OAI21_X1 U8441 ( .B1(n6465), .B2(n9922), .A(n6663), .ZN(n6664) );
  INV_X1 U8442 ( .A(n6664), .ZN(n6665) );
  INV_X1 U8443 ( .A(n10058), .ZN(n9897) );
  NAND2_X1 U8444 ( .A1(n9897), .A2(n8313), .ZN(n6667) );
  NAND2_X1 U8445 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  XNOR2_X1 U8446 ( .A(n6669), .B(n8316), .ZN(n6671) );
  NOR2_X1 U8447 ( .A1(n10058), .A2(n8318), .ZN(n6670) );
  AOI21_X1 U8448 ( .B1(n10048), .B2(n8313), .A(n6670), .ZN(n6672) );
  XNOR2_X1 U8449 ( .A(n6671), .B(n6672), .ZN(n9278) );
  INV_X1 U8450 ( .A(n6671), .ZN(n6673) );
  NAND2_X1 U8451 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NAND2_X1 U8452 ( .A1(n7326), .A2(n7103), .ZN(n6678) );
  INV_X1 U8453 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8454 ( .A1(n6676), .A2(n6675), .ZN(n6721) );
  NAND2_X1 U8455 ( .A1(n6721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6695) );
  XNOR2_X1 U8456 ( .A(n6695), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U8457 ( .A1(n6778), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6777), .B2(
        n10148), .ZN(n6677) );
  NAND2_X1 U8458 ( .A1(n10042), .A2(n6933), .ZN(n6691) );
  INV_X1 U8459 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10461) );
  INV_X1 U8460 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10548) );
  OR2_X1 U8461 ( .A1(n6982), .A2(n10548), .ZN(n6679) );
  OAI21_X1 U8462 ( .B1(n7125), .B2(n10461), .A(n6679), .ZN(n6680) );
  INV_X1 U8463 ( .A(n6680), .ZN(n6689) );
  INV_X1 U8464 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U8465 ( .A1(n6683), .A2(n6682), .ZN(n6684) );
  NAND2_X1 U8466 ( .A1(n6705), .A2(n6684), .ZN(n9892) );
  INV_X1 U8467 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6685) );
  OR2_X1 U8468 ( .A1(n7122), .A2(n6685), .ZN(n6686) );
  OAI21_X1 U8469 ( .B1(n6465), .B2(n9892), .A(n6686), .ZN(n6687) );
  INV_X1 U8470 ( .A(n6687), .ZN(n6688) );
  NAND2_X1 U8471 ( .A1(n9588), .A2(n8313), .ZN(n6690) );
  NAND2_X1 U8472 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  XNOR2_X1 U8473 ( .A(n6692), .B(n8316), .ZN(n9128) );
  NAND2_X1 U8474 ( .A1(n10042), .A2(n8313), .ZN(n6694) );
  NAND2_X1 U8475 ( .A1(n9588), .A2(n6906), .ZN(n6693) );
  NAND2_X1 U8476 ( .A1(n6694), .A2(n6693), .ZN(n9126) );
  NAND2_X1 U8477 ( .A1(n9128), .A2(n9126), .ZN(n6716) );
  NAND2_X1 U8478 ( .A1(n6695), .A2(n6718), .ZN(n6696) );
  NAND2_X1 U8479 ( .A1(n6696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6697) );
  XNOR2_X1 U8480 ( .A(n6697), .B(n6719), .ZN(n9621) );
  INV_X1 U8481 ( .A(n9621), .ZN(n10160) );
  AOI22_X1 U8482 ( .A1(n6778), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6777), .B2(
        n10160), .ZN(n6698) );
  NAND2_X2 U8483 ( .A1(n6699), .A2(n6698), .ZN(n10034) );
  NAND2_X1 U8484 ( .A1(n10034), .A2(n6933), .ZN(n6711) );
  INV_X1 U8485 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6701) );
  INV_X1 U8486 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10624) );
  OR2_X1 U8487 ( .A1(n7122), .A2(n10624), .ZN(n6700) );
  OAI21_X1 U8488 ( .B1(n7125), .B2(n6701), .A(n6700), .ZN(n6702) );
  INV_X1 U8489 ( .A(n6702), .ZN(n6709) );
  INV_X1 U8490 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U8491 ( .A1(n6705), .A2(n6704), .ZN(n6706) );
  AND2_X1 U8492 ( .A1(n6726), .A2(n6706), .ZN(n9875) );
  NAND2_X1 U8493 ( .A1(n9875), .A2(n6937), .ZN(n6708) );
  INV_X1 U8494 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10154) );
  OR2_X1 U8495 ( .A1(n6982), .A2(n10154), .ZN(n6707) );
  OR2_X1 U8496 ( .A1(n10039), .A2(n4427), .ZN(n6710) );
  NAND2_X1 U8497 ( .A1(n6711), .A2(n6710), .ZN(n6712) );
  XNOR2_X1 U8498 ( .A(n6712), .B(n8316), .ZN(n6717) );
  NAND2_X1 U8499 ( .A1(n10034), .A2(n8313), .ZN(n6714) );
  OR2_X1 U8500 ( .A1(n10039), .A2(n8318), .ZN(n6713) );
  NAND2_X1 U8501 ( .A1(n6714), .A2(n6713), .ZN(n9331) );
  OAI22_X1 U8502 ( .A1(n6717), .A2(n9331), .B1(n9128), .B2(n9126), .ZN(n6715)
         );
  INV_X1 U8503 ( .A(n9331), .ZN(n6736) );
  INV_X1 U8504 ( .A(n6717), .ZN(n9222) );
  NAND2_X1 U8505 ( .A1(n7547), .A2(n7103), .ZN(n6724) );
  NAND2_X1 U8506 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  OAI21_X1 U8507 ( .B1(n6721), .B2(n6720), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6722) );
  XNOR2_X1 U8508 ( .A(n6722), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U8509 ( .A1(n6778), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6777), .B2(
        n10172), .ZN(n6723) );
  NAND2_X2 U8510 ( .A1(n6724), .A2(n6723), .ZN(n9866) );
  NAND2_X1 U8511 ( .A1(n9866), .A2(n6933), .ZN(n6732) );
  INV_X1 U8512 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8513 ( .A1(n6726), .A2(n6725), .ZN(n6727) );
  AND2_X1 U8514 ( .A1(n6748), .A2(n6727), .ZN(n9858) );
  NAND2_X1 U8515 ( .A1(n9858), .A2(n6937), .ZN(n6730) );
  AOI22_X1 U8516 ( .A1(n6384), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7106), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6729) );
  INV_X1 U8517 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10030) );
  OR2_X1 U8518 ( .A1(n6982), .A2(n10030), .ZN(n6728) );
  INV_X1 U8519 ( .A(n9881), .ZN(n9587) );
  NAND2_X1 U8520 ( .A1(n9587), .A2(n8313), .ZN(n6731) );
  NAND2_X1 U8521 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  XNOR2_X1 U8522 ( .A(n6733), .B(n8316), .ZN(n6737) );
  NAND2_X1 U8523 ( .A1(n9866), .A2(n8313), .ZN(n6735) );
  OR2_X1 U8524 ( .A1(n9881), .A2(n8318), .ZN(n6734) );
  NAND2_X1 U8525 ( .A1(n6735), .A2(n6734), .ZN(n6738) );
  NAND2_X1 U8526 ( .A1(n6737), .A2(n6738), .ZN(n9218) );
  OAI21_X1 U8527 ( .B1(n6736), .B2(n9222), .A(n9218), .ZN(n6741) );
  INV_X1 U8528 ( .A(n6737), .ZN(n6740) );
  INV_X1 U8529 ( .A(n6738), .ZN(n6739) );
  NAND2_X1 U8530 ( .A1(n6740), .A2(n6739), .ZN(n9217) );
  NAND2_X1 U8531 ( .A1(n7505), .A2(n7103), .ZN(n6745) );
  NAND2_X1 U8532 ( .A1(n6742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6743) );
  XNOR2_X1 U8533 ( .A(n6743), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U8534 ( .A1(n6778), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6777), .B2(
        n10184), .ZN(n6744) );
  NAND2_X1 U8535 ( .A1(n10020), .A2(n6933), .ZN(n6753) );
  INV_X1 U8536 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10653) );
  INV_X1 U8537 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U8538 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  NAND2_X1 U8539 ( .A1(n6782), .A2(n6749), .ZN(n9848) );
  OR2_X1 U8540 ( .A1(n9848), .A2(n6465), .ZN(n6751) );
  AOI22_X1 U8541 ( .A1(n6384), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n4408), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n6750) );
  OAI211_X1 U8542 ( .C1(n7122), .C2(n10653), .A(n6751), .B(n6750), .ZN(n10024)
         );
  NAND2_X1 U8543 ( .A1(n10024), .A2(n8313), .ZN(n6752) );
  NAND2_X1 U8544 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  XNOR2_X1 U8545 ( .A(n6754), .B(n8316), .ZN(n6756) );
  AND2_X1 U8546 ( .A1(n10024), .A2(n6906), .ZN(n6755) );
  AOI21_X1 U8547 ( .B1(n10020), .B2(n8313), .A(n6755), .ZN(n6757) );
  XNOR2_X1 U8548 ( .A(n6756), .B(n6757), .ZN(n9231) );
  NAND2_X1 U8549 ( .A1(n9232), .A2(n9231), .ZN(n6760) );
  INV_X1 U8550 ( .A(n6756), .ZN(n6758) );
  NAND2_X1 U8551 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NAND2_X1 U8552 ( .A1(n7750), .A2(n7103), .ZN(n6762) );
  AOI22_X1 U8553 ( .A1(n6778), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9635), .B2(
        n6777), .ZN(n6761) );
  NAND2_X1 U8554 ( .A1(n10009), .A2(n6933), .ZN(n6772) );
  INV_X1 U8555 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6781) );
  INV_X1 U8556 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U8557 ( .A1(n6784), .A2(n6763), .ZN(n6764) );
  NAND2_X1 U8558 ( .A1(n6804), .A2(n6764), .ZN(n9813) );
  OR2_X1 U8559 ( .A1(n9813), .A2(n6465), .ZN(n6770) );
  INV_X1 U8560 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9812) );
  INV_X1 U8561 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10392) );
  OR2_X1 U8562 ( .A1(n7122), .A2(n10392), .ZN(n6767) );
  INV_X1 U8563 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6765) );
  OR2_X1 U8564 ( .A1(n6982), .A2(n6765), .ZN(n6766) );
  OAI211_X1 U8565 ( .C1(n7125), .C2(n9812), .A(n6767), .B(n6766), .ZN(n6768)
         );
  INV_X1 U8566 ( .A(n6768), .ZN(n6769) );
  NAND2_X1 U8567 ( .A1(n9586), .A2(n4418), .ZN(n6771) );
  NAND2_X1 U8568 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  XNOR2_X1 U8569 ( .A(n6773), .B(n8316), .ZN(n9163) );
  NAND2_X1 U8570 ( .A1(n10009), .A2(n8313), .ZN(n6775) );
  NAND2_X1 U8571 ( .A1(n9586), .A2(n6906), .ZN(n6774) );
  NAND2_X1 U8572 ( .A1(n6775), .A2(n6774), .ZN(n6796) );
  NAND2_X1 U8573 ( .A1(n7585), .A2(n7103), .ZN(n6780) );
  XNOR2_X1 U8574 ( .A(n6776), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9625) );
  AOI22_X1 U8575 ( .A1(n6778), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6777), .B2(
        n9625), .ZN(n6779) );
  NAND2_X1 U8576 ( .A1(n10084), .A2(n6933), .ZN(n6791) );
  NAND2_X1 U8577 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  AND2_X1 U8578 ( .A1(n6784), .A2(n6783), .ZN(n9828) );
  NAND2_X1 U8579 ( .A1(n9828), .A2(n6937), .ZN(n6789) );
  NAND2_X1 U8580 ( .A1(n7106), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8581 ( .A1(n4408), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6785) );
  OAI211_X1 U8582 ( .C1(n7125), .C2(n10503), .A(n6786), .B(n6785), .ZN(n6787)
         );
  INV_X1 U8583 ( .A(n6787), .ZN(n6788) );
  NAND2_X1 U8584 ( .A1(n9842), .A2(n4418), .ZN(n6790) );
  NAND2_X1 U8585 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  XNOR2_X1 U8586 ( .A(n6792), .B(n8316), .ZN(n6798) );
  NAND2_X1 U8587 ( .A1(n10084), .A2(n8313), .ZN(n6794) );
  NAND2_X1 U8588 ( .A1(n9842), .A2(n6906), .ZN(n6793) );
  NAND2_X1 U8589 ( .A1(n6794), .A2(n6793), .ZN(n9311) );
  OAI22_X1 U8590 ( .A1(n9163), .A2(n6796), .B1(n6798), .B2(n9311), .ZN(n6801)
         );
  INV_X1 U8591 ( .A(n9311), .ZN(n6795) );
  INV_X1 U8592 ( .A(n6796), .ZN(n9162) );
  OAI21_X1 U8593 ( .B1(n9161), .B2(n6795), .A(n9162), .ZN(n6799) );
  AND2_X1 U8594 ( .A1(n6796), .A2(n9311), .ZN(n6797) );
  AOI22_X1 U8595 ( .A1(n9163), .A2(n6799), .B1(n6798), .B2(n6797), .ZN(n6800)
         );
  NAND2_X1 U8596 ( .A1(n7835), .A2(n7103), .ZN(n6803) );
  OR2_X1 U8597 ( .A1(n6930), .A2(n7836), .ZN(n6802) );
  NAND2_X1 U8598 ( .A1(n10001), .A2(n6933), .ZN(n6813) );
  INV_X1 U8599 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U8600 ( .A1(n6804), .A2(n9269), .ZN(n6805) );
  AND2_X1 U8601 ( .A1(n6824), .A2(n6805), .ZN(n9797) );
  NAND2_X1 U8602 ( .A1(n9797), .A2(n6937), .ZN(n6811) );
  INV_X1 U8603 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8604 ( .A1(n4408), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6807) );
  INV_X1 U8605 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10560) );
  OR2_X1 U8606 ( .A1(n6512), .A2(n10560), .ZN(n6806) );
  OAI211_X1 U8607 ( .C1(n7125), .C2(n6808), .A(n6807), .B(n6806), .ZN(n6809)
         );
  INV_X1 U8608 ( .A(n6809), .ZN(n6810) );
  OR2_X1 U8609 ( .A1(n9992), .A2(n4427), .ZN(n6812) );
  NAND2_X1 U8610 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  XNOR2_X1 U8611 ( .A(n6814), .B(n8316), .ZN(n6817) );
  NAND2_X1 U8612 ( .A1(n10001), .A2(n8313), .ZN(n6816) );
  OR2_X1 U8613 ( .A1(n9992), .A2(n8318), .ZN(n6815) );
  NAND2_X1 U8614 ( .A1(n6816), .A2(n6815), .ZN(n6818) );
  INV_X1 U8615 ( .A(n6817), .ZN(n6820) );
  INV_X1 U8616 ( .A(n6818), .ZN(n6819) );
  NAND2_X1 U8617 ( .A1(n6820), .A2(n6819), .ZN(n9264) );
  NAND2_X1 U8618 ( .A1(n7991), .A2(n7103), .ZN(n6822) );
  OR2_X1 U8619 ( .A1(n6930), .A2(n10519), .ZN(n6821) );
  NAND2_X1 U8620 ( .A1(n9996), .A2(n6933), .ZN(n6832) );
  INV_X1 U8621 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U8622 ( .A1(n6824), .A2(n10647), .ZN(n6825) );
  NAND2_X1 U8623 ( .A1(n6854), .A2(n6825), .ZN(n9777) );
  INV_X1 U8624 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U8625 ( .A1(n7106), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8626 ( .A1(n4408), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6826) );
  OAI211_X1 U8627 ( .C1(n7125), .C2(n9776), .A(n6827), .B(n6826), .ZN(n6828)
         );
  INV_X1 U8628 ( .A(n6828), .ZN(n6829) );
  NAND2_X1 U8629 ( .A1(n9982), .A2(n8313), .ZN(n6831) );
  NAND2_X1 U8630 ( .A1(n6832), .A2(n6831), .ZN(n6833) );
  XNOR2_X1 U8631 ( .A(n6833), .B(n8316), .ZN(n6835) );
  NOR2_X1 U8632 ( .A1(n9792), .A2(n8318), .ZN(n6834) );
  AOI21_X1 U8633 ( .B1(n9996), .B2(n8313), .A(n6834), .ZN(n6836) );
  XNOR2_X1 U8634 ( .A(n6835), .B(n6836), .ZN(n9187) );
  INV_X1 U8635 ( .A(n6835), .ZN(n6837) );
  NAND2_X1 U8636 ( .A1(n8245), .A2(n7103), .ZN(n6839) );
  OR2_X1 U8637 ( .A1(n6930), .A2(n8243), .ZN(n6838) );
  NAND2_X1 U8638 ( .A1(n4611), .A2(n6933), .ZN(n6847) );
  XNOR2_X1 U8639 ( .A(n6879), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U8640 ( .A1(n9747), .A2(n6937), .ZN(n6845) );
  INV_X1 U8641 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U8642 ( .A1(n4408), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6842) );
  INV_X1 U8643 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10535) );
  OR2_X1 U8644 ( .A1(n7122), .A2(n10535), .ZN(n6841) );
  OAI211_X1 U8645 ( .C1(n7125), .C2(n9745), .A(n6842), .B(n6841), .ZN(n6843)
         );
  INV_X1 U8646 ( .A(n6843), .ZN(n6844) );
  OR2_X1 U8647 ( .A1(n9769), .A2(n4427), .ZN(n6846) );
  NAND2_X1 U8648 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  XNOR2_X1 U8649 ( .A(n6848), .B(n8316), .ZN(n6870) );
  NAND2_X1 U8650 ( .A1(n4611), .A2(n8313), .ZN(n6850) );
  OR2_X1 U8651 ( .A1(n9769), .A2(n8318), .ZN(n6849) );
  NAND2_X1 U8652 ( .A1(n6850), .A2(n6849), .ZN(n6871) );
  NAND2_X1 U8653 ( .A1(n6870), .A2(n6871), .ZN(n9140) );
  NAND2_X1 U8654 ( .A1(n8176), .A2(n7103), .ZN(n6852) );
  OR2_X1 U8655 ( .A1(n6930), .A2(n8178), .ZN(n6851) );
  NAND2_X1 U8656 ( .A1(n9763), .A2(n6933), .ZN(n6862) );
  INV_X1 U8657 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8658 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  NAND2_X1 U8659 ( .A1(n6879), .A2(n6855), .ZN(n9765) );
  OR2_X1 U8660 ( .A1(n9765), .A2(n6465), .ZN(n6860) );
  INV_X1 U8661 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9764) );
  NAND2_X1 U8662 ( .A1(n4408), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6857) );
  INV_X1 U8663 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10593) );
  OR2_X1 U8664 ( .A1(n7122), .A2(n10593), .ZN(n6856) );
  OAI211_X1 U8665 ( .C1(n7125), .C2(n9764), .A(n6857), .B(n6856), .ZN(n6858)
         );
  INV_X1 U8666 ( .A(n6858), .ZN(n6859) );
  NAND2_X1 U8667 ( .A1(n9973), .A2(n8313), .ZN(n6861) );
  NAND2_X1 U8668 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  XNOR2_X1 U8669 ( .A(n6863), .B(n6947), .ZN(n9139) );
  NAND2_X1 U8670 ( .A1(n9763), .A2(n4418), .ZN(n6865) );
  NAND2_X1 U8671 ( .A1(n9973), .A2(n6906), .ZN(n6864) );
  NOR2_X1 U8672 ( .A1(n9139), .A2(n9286), .ZN(n6866) );
  NAND2_X1 U8673 ( .A1(n9136), .A2(n6868), .ZN(n6893) );
  INV_X1 U8674 ( .A(n9139), .ZN(n9137) );
  INV_X1 U8675 ( .A(n9286), .ZN(n6869) );
  NOR2_X1 U8676 ( .A1(n9137), .A2(n6869), .ZN(n6874) );
  INV_X1 U8677 ( .A(n6870), .ZN(n6873) );
  INV_X1 U8678 ( .A(n6871), .ZN(n6872) );
  AOI21_X1 U8679 ( .B1(n6874), .B2(n9140), .A(n9241), .ZN(n6892) );
  NAND2_X1 U8680 ( .A1(n8305), .A2(n7103), .ZN(n6876) );
  OR2_X1 U8681 ( .A1(n6930), .A2(n8308), .ZN(n6875) );
  NAND2_X1 U8682 ( .A1(n4426), .A2(n6933), .ZN(n6887) );
  INV_X1 U8683 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6877) );
  INV_X1 U8684 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6878) );
  OAI21_X1 U8685 ( .B1(n6879), .B2(n6877), .A(n6878), .ZN(n6880) );
  AND2_X1 U8686 ( .A1(n6880), .A2(n6899), .ZN(n9728) );
  NAND2_X1 U8687 ( .A1(n9728), .A2(n6937), .ZN(n6885) );
  INV_X1 U8688 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U8689 ( .A1(n7106), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U8690 ( .A1(n4408), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6881) );
  OAI211_X1 U8691 ( .C1(n7125), .C2(n9729), .A(n6882), .B(n6881), .ZN(n6883)
         );
  INV_X1 U8692 ( .A(n6883), .ZN(n6884) );
  NAND2_X1 U8693 ( .A1(n9974), .A2(n8313), .ZN(n6886) );
  NAND2_X1 U8694 ( .A1(n6887), .A2(n6886), .ZN(n6888) );
  XNOR2_X1 U8695 ( .A(n6888), .B(n6947), .ZN(n6891) );
  NOR2_X1 U8696 ( .A1(n9750), .A2(n8318), .ZN(n6889) );
  AOI21_X1 U8697 ( .B1(n4426), .B2(n8313), .A(n6889), .ZN(n6890) );
  NAND2_X1 U8698 ( .A1(n6891), .A2(n6890), .ZN(n6894) );
  OAI21_X1 U8699 ( .B1(n6891), .B2(n6890), .A(n6894), .ZN(n9239) );
  INV_X1 U8700 ( .A(n6894), .ZN(n6895) );
  OR2_X1 U8701 ( .A1(n6930), .A2(n10563), .ZN(n6896) );
  INV_X1 U8702 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U8703 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  NAND2_X1 U8704 ( .A1(n6913), .A2(n6900), .ZN(n9714) );
  INV_X1 U8705 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U8706 ( .A1(n4408), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6902) );
  INV_X1 U8707 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10656) );
  OR2_X1 U8708 ( .A1(n6512), .A2(n10656), .ZN(n6901) );
  OAI211_X1 U8709 ( .C1(n7125), .C2(n9713), .A(n6902), .B(n6901), .ZN(n6903)
         );
  INV_X1 U8710 ( .A(n6903), .ZN(n6904) );
  AOI22_X1 U8711 ( .A1(n9961), .A2(n8313), .B1(n6906), .B2(n9701), .ZN(n6925)
         );
  NAND2_X1 U8712 ( .A1(n9961), .A2(n6933), .ZN(n6908) );
  NAND2_X1 U8713 ( .A1(n9701), .A2(n8313), .ZN(n6907) );
  NAND2_X1 U8714 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  XOR2_X1 U8715 ( .A(n6925), .B(n6927), .Z(n9210) );
  OR2_X1 U8716 ( .A1(n6930), .A2(n10113), .ZN(n6910) );
  INV_X1 U8717 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8718 ( .A1(n6913), .A2(n6912), .ZN(n6914) );
  NAND2_X1 U8719 ( .A1(n6935), .A2(n6914), .ZN(n9699) );
  INV_X1 U8720 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U8721 ( .A1(n4408), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6917) );
  INV_X1 U8722 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6915) );
  OR2_X1 U8723 ( .A1(n7122), .A2(n6915), .ZN(n6916) );
  OAI211_X1 U8724 ( .C1(n7125), .C2(n9698), .A(n6917), .B(n6916), .ZN(n6918)
         );
  INV_X1 U8725 ( .A(n6918), .ZN(n6919) );
  NOR2_X1 U8726 ( .A1(n9946), .A2(n8318), .ZN(n6921) );
  AOI21_X1 U8727 ( .B1(n9959), .B2(n8313), .A(n6921), .ZN(n6952) );
  NAND2_X1 U8728 ( .A1(n9959), .A2(n6933), .ZN(n6923) );
  NAND2_X1 U8729 ( .A1(n9712), .A2(n8313), .ZN(n6922) );
  NAND2_X1 U8730 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  XNOR2_X1 U8731 ( .A(n6924), .B(n8316), .ZN(n6954) );
  XOR2_X1 U8732 ( .A(n6952), .B(n6954), .Z(n9317) );
  INV_X1 U8733 ( .A(n6925), .ZN(n6926) );
  NAND2_X1 U8734 ( .A1(n9113), .A2(n7103), .ZN(n6932) );
  OR2_X1 U8735 ( .A1(n6930), .A2(n10112), .ZN(n6931) );
  NAND2_X1 U8736 ( .A1(n9680), .A2(n6933), .ZN(n6946) );
  INV_X1 U8737 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8738 ( .A1(n6935), .A2(n6934), .ZN(n6936) );
  NAND2_X1 U8739 ( .A1(n9681), .A2(n6937), .ZN(n6943) );
  INV_X1 U8740 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6940) );
  INV_X1 U8741 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10460) );
  OR2_X1 U8742 ( .A1(n6982), .A2(n10460), .ZN(n6939) );
  INV_X1 U8743 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10565) );
  OR2_X1 U8744 ( .A1(n7122), .A2(n10565), .ZN(n6938) );
  OAI211_X1 U8745 ( .C1(n7125), .C2(n6940), .A(n6939), .B(n6938), .ZN(n6941)
         );
  INV_X1 U8746 ( .A(n6941), .ZN(n6942) );
  AND2_X2 U8747 ( .A1(n6943), .A2(n6942), .ZN(n9954) );
  OR2_X1 U8748 ( .A1(n9954), .A2(n4427), .ZN(n6945) );
  NAND2_X1 U8749 ( .A1(n6946), .A2(n6945), .ZN(n6948) );
  XNOR2_X1 U8750 ( .A(n6948), .B(n6947), .ZN(n6951) );
  NOR2_X1 U8751 ( .A1(n9954), .A2(n8318), .ZN(n6949) );
  AOI21_X1 U8752 ( .B1(n9680), .B2(n4418), .A(n6949), .ZN(n6950) );
  NAND2_X1 U8753 ( .A1(n6951), .A2(n6950), .ZN(n8327) );
  OAI21_X1 U8754 ( .B1(n6951), .B2(n6950), .A(n8327), .ZN(n6956) );
  INV_X1 U8755 ( .A(n6952), .ZN(n6953) );
  AND2_X1 U8756 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  INV_X1 U8757 ( .A(n6955), .ZN(n6958) );
  INV_X1 U8758 ( .A(n6956), .ZN(n6957) );
  NAND2_X1 U8759 ( .A1(n10118), .A2(P1_B_REG_SCAN_IN), .ZN(n6960) );
  INV_X1 U8760 ( .A(n8310), .ZN(n6959) );
  MUX2_X1 U8761 ( .A(n6960), .B(P1_B_REG_SCAN_IN), .S(n6959), .Z(n6961) );
  NAND2_X1 U8762 ( .A1(n6961), .A2(n6962), .ZN(n10098) );
  NAND2_X1 U8763 ( .A1(n10115), .A2(n10118), .ZN(n10100) );
  OAI21_X1 U8764 ( .B1(n10098), .B2(P1_D_REG_1__SCAN_IN), .A(n10100), .ZN(
        n7591) );
  NOR4_X1 U8765 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6970) );
  NOR4_X1 U8766 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6969) );
  INV_X1 U8767 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10650) );
  INV_X1 U8768 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10552) );
  INV_X1 U8769 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10576) );
  INV_X1 U8770 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10445) );
  NAND4_X1 U8771 ( .A1(n10650), .A2(n10552), .A3(n10576), .A4(n10445), .ZN(
        n10431) );
  NOR4_X1 U8772 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6966) );
  NOR4_X1 U8773 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6965) );
  NOR4_X1 U8774 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6964) );
  NOR4_X1 U8775 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6963) );
  NAND4_X1 U8776 ( .A1(n6966), .A2(n6965), .A3(n6964), .A4(n6963), .ZN(n6967)
         );
  NOR4_X1 U8777 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10431), .A4(n6967), .ZN(n6968) );
  AND3_X1 U8778 ( .A1(n6970), .A2(n6969), .A3(n6968), .ZN(n6971) );
  NOR2_X1 U8779 ( .A1(n10098), .A2(n6971), .ZN(n7090) );
  NOR2_X1 U8780 ( .A1(n7591), .A2(n7090), .ZN(n6972) );
  NAND2_X1 U8781 ( .A1(n10115), .A2(n8310), .ZN(n10101) );
  OAI21_X1 U8782 ( .B1(n10098), .B2(P1_D_REG_0__SCAN_IN), .A(n10101), .ZN(
        n7592) );
  INV_X1 U8783 ( .A(n7592), .ZN(n7111) );
  INV_X1 U8784 ( .A(n10049), .ZN(n10237) );
  NAND2_X1 U8785 ( .A1(n6973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6975) );
  INV_X1 U8786 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6974) );
  XNOR2_X1 U8787 ( .A(n6975), .B(n6974), .ZN(n7185) );
  AND2_X1 U8788 ( .A1(n7156), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6976) );
  INV_X1 U8789 ( .A(n7184), .ZN(n9515) );
  AND3_X1 U8790 ( .A1(n10237), .A2(n10099), .A3(n9515), .ZN(n6977) );
  OAI21_X1 U8791 ( .B1(n8334), .B2(n6978), .A(n9320), .ZN(n7002) );
  INV_X1 U8792 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6979) );
  NAND2_X1 U8793 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  NAND2_X1 U8794 ( .A1(n9653), .A2(n6981), .ZN(n9667) );
  INV_X1 U8795 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9666) );
  INV_X1 U8796 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10514) );
  OR2_X1 U8797 ( .A1(n6982), .A2(n10514), .ZN(n6984) );
  INV_X1 U8798 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10393) );
  OR2_X1 U8799 ( .A1(n6512), .A2(n10393), .ZN(n6983) );
  OAI211_X1 U8800 ( .C1(n7125), .C2(n9666), .A(n6984), .B(n6983), .ZN(n6985)
         );
  INV_X1 U8801 ( .A(n6985), .ZN(n6986) );
  AND2_X2 U8802 ( .A1(n6987), .A2(n6986), .ZN(n9947) );
  AND2_X1 U8803 ( .A1(n10099), .A2(n9524), .ZN(n6990) );
  INV_X1 U8804 ( .A(n6990), .ZN(n6988) );
  NAND2_X1 U8805 ( .A1(n7184), .A2(n4429), .ZN(n10057) );
  NOR2_X1 U8806 ( .A1(n6988), .A2(n10057), .ZN(n6989) );
  AND2_X1 U8807 ( .A1(n6990), .A2(n10053), .ZN(n9519) );
  NAND2_X1 U8808 ( .A1(n9519), .A2(n6991), .ZN(n9324) );
  INV_X1 U8809 ( .A(n6991), .ZN(n6998) );
  NAND2_X1 U8810 ( .A1(n10002), .A2(n9635), .ZN(n7091) );
  NAND2_X1 U8811 ( .A1(n6998), .A2(n7091), .ZN(n7282) );
  NAND2_X1 U8812 ( .A1(n7184), .A2(n7003), .ZN(n7089) );
  AND2_X1 U8813 ( .A1(n7089), .A2(n7156), .ZN(n6992) );
  AOI21_X1 U8814 ( .B1(n7282), .B2(n6992), .A(P1_U3086), .ZN(n6994) );
  OR2_X1 U8815 ( .A1(n7185), .A2(P1_U3086), .ZN(n9575) );
  INV_X1 U8816 ( .A(n9575), .ZN(n6993) );
  AOI22_X1 U8817 ( .A1(n9681), .A2(n9338), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6995) );
  OAI21_X1 U8818 ( .B1(n9946), .B2(n9324), .A(n6995), .ZN(n6996) );
  AOI21_X1 U8819 ( .B1(n9657), .B2(n9326), .A(n6996), .ZN(n7001) );
  AND2_X1 U8820 ( .A1(n5181), .A2(n9522), .ZN(n7597) );
  NAND2_X1 U8821 ( .A1(n10099), .A2(n7597), .ZN(n6997) );
  OR2_X1 U8822 ( .A1(n6998), .A2(n6997), .ZN(n7000) );
  INV_X1 U8823 ( .A(n7091), .ZN(n6999) );
  NAND3_X1 U8824 ( .A1(n7002), .A2(n7001), .A3(n5179), .ZN(P1_U3214) );
  NAND2_X1 U8825 ( .A1(n7184), .A2(n9524), .ZN(n9935) );
  OAI21_X1 U8826 ( .B1(n8177), .B2(n9635), .A(n7003), .ZN(n7004) );
  INV_X1 U8827 ( .A(n5181), .ZN(n9934) );
  AND2_X1 U8828 ( .A1(n7004), .A2(n9934), .ZN(n7005) );
  NAND2_X1 U8829 ( .A1(n9935), .A2(n7005), .ZN(n7649) );
  NAND2_X1 U8830 ( .A1(n9449), .A2(n7837), .ZN(n10215) );
  NAND2_X1 U8831 ( .A1(n4610), .A2(n7587), .ZN(n7590) );
  INV_X1 U8832 ( .A(n6400), .ZN(n7283) );
  NAND2_X1 U8833 ( .A1(n7283), .A2(n7073), .ZN(n7008) );
  NAND2_X1 U8834 ( .A1(n7590), .A2(n7008), .ZN(n7737) );
  NAND2_X1 U8835 ( .A1(n7009), .A2(n10225), .ZN(n9528) );
  NAND2_X1 U8836 ( .A1(n7737), .A2(n9453), .ZN(n7736) );
  INV_X1 U8837 ( .A(n7009), .ZN(n7514) );
  NAND2_X1 U8838 ( .A1(n7514), .A2(n10225), .ZN(n7010) );
  XNOR2_X2 U8839 ( .A(n9594), .B(n7637), .ZN(n9454) );
  NAND2_X1 U8840 ( .A1(n9595), .A2(n7652), .ZN(n7011) );
  AND2_X1 U8841 ( .A1(n9454), .A2(n7011), .ZN(n7012) );
  NAND2_X1 U8842 ( .A1(n7647), .A2(n7012), .ZN(n7015) );
  NOR2_X1 U8843 ( .A1(n9595), .A2(n7652), .ZN(n7627) );
  NAND2_X1 U8844 ( .A1(n7812), .A2(n5051), .ZN(n7016) );
  INV_X1 U8845 ( .A(n9594), .ZN(n7847) );
  NAND2_X1 U8846 ( .A1(n7847), .A2(n7637), .ZN(n7663) );
  NAND2_X1 U8847 ( .A1(n7016), .A2(n7663), .ZN(n7013) );
  AOI21_X1 U8848 ( .B1(n9454), .B2(n7627), .A(n7013), .ZN(n7014) );
  NAND2_X1 U8849 ( .A1(n7015), .A2(n7014), .ZN(n7019) );
  NAND2_X2 U8850 ( .A1(n9593), .A2(n5051), .ZN(n9537) );
  NAND2_X1 U8851 ( .A1(n7812), .A2(n7672), .ZN(n9533) );
  INV_X1 U8852 ( .A(n7016), .ZN(n7699) );
  INV_X1 U8853 ( .A(n7820), .ZN(n9347) );
  OAI21_X1 U8854 ( .B1(n7059), .B2(n7699), .A(n9452), .ZN(n7017) );
  INV_X1 U8855 ( .A(n7017), .ZN(n7018) );
  INV_X1 U8856 ( .A(n9592), .ZN(n7872) );
  NAND2_X1 U8857 ( .A1(n7872), .A2(n7811), .ZN(n7823) );
  NAND2_X1 U8858 ( .A1(n7021), .A2(n7914), .ZN(n7880) );
  AND2_X1 U8859 ( .A1(n7823), .A2(n7880), .ZN(n7020) );
  NAND2_X1 U8860 ( .A1(n9183), .A2(n9257), .ZN(n9364) );
  NAND2_X1 U8861 ( .A1(n7995), .A2(n9364), .ZN(n7879) );
  NAND2_X1 U8862 ( .A1(n7021), .A2(n7917), .ZN(n9360) );
  NAND2_X1 U8863 ( .A1(n7824), .A2(n7880), .ZN(n7022) );
  AND2_X1 U8864 ( .A1(n7879), .A2(n7022), .ZN(n7023) );
  NAND2_X1 U8865 ( .A1(n7024), .A2(n7023), .ZN(n7883) );
  INV_X1 U8866 ( .A(n9257), .ZN(n8007) );
  OR2_X1 U8867 ( .A1(n9183), .A2(n8007), .ZN(n7025) );
  NAND2_X1 U8868 ( .A1(n7883), .A2(n7025), .ZN(n8000) );
  NAND2_X1 U8869 ( .A1(n8070), .A2(n9152), .ZN(n9374) );
  NAND2_X1 U8870 ( .A1(n9365), .A2(n9374), .ZN(n7999) );
  NAND2_X1 U8871 ( .A1(n8000), .A2(n7999), .ZN(n7985) );
  INV_X1 U8872 ( .A(n9152), .ZN(n9178) );
  OR2_X1 U8873 ( .A1(n8070), .A2(n9178), .ZN(n7986) );
  OR2_X1 U8874 ( .A1(n9157), .A2(n9590), .ZN(n8028) );
  AND2_X1 U8875 ( .A1(n7986), .A2(n8028), .ZN(n7026) );
  NAND2_X1 U8876 ( .A1(n7985), .A2(n7026), .ZN(n7031) );
  NAND2_X1 U8877 ( .A1(n7027), .A2(n9203), .ZN(n9376) );
  AND2_X1 U8878 ( .A1(n9461), .A2(n7029), .ZN(n7030) );
  NAND2_X1 U8879 ( .A1(n7031), .A2(n7030), .ZN(n8031) );
  OR2_X1 U8880 ( .A1(n7027), .A2(n10054), .ZN(n7032) );
  NAND2_X1 U8881 ( .A1(n8031), .A2(n7032), .ZN(n8119) );
  OR2_X1 U8882 ( .A1(n10095), .A2(n9911), .ZN(n9370) );
  NAND2_X1 U8883 ( .A1(n10095), .A2(n9911), .ZN(n9380) );
  OR2_X1 U8884 ( .A1(n10095), .A2(n9589), .ZN(n7033) );
  OR2_X1 U8885 ( .A1(n10048), .A2(n10058), .ZN(n9387) );
  NAND2_X1 U8886 ( .A1(n9387), .A2(n9543), .ZN(n9916) );
  NAND2_X1 U8887 ( .A1(n7076), .A2(n10058), .ZN(n7034) );
  NAND2_X1 U8888 ( .A1(n10042), .A2(n9588), .ZN(n7035) );
  INV_X1 U8889 ( .A(n10039), .ZN(n10023) );
  NOR2_X1 U8890 ( .A1(n10034), .A2(n10023), .ZN(n7037) );
  NAND2_X1 U8891 ( .A1(n10034), .A2(n10023), .ZN(n7036) );
  NAND2_X1 U8892 ( .A1(n9866), .A2(n9881), .ZN(n9838) );
  INV_X1 U8893 ( .A(n9868), .ZN(n9469) );
  NAND2_X1 U8894 ( .A1(n9867), .A2(n9469), .ZN(n7039) );
  NAND2_X1 U8895 ( .A1(n9866), .A2(n9587), .ZN(n7038) );
  NAND2_X1 U8896 ( .A1(n7039), .A2(n7038), .ZN(n9835) );
  OR2_X1 U8897 ( .A1(n10020), .A2(n10024), .ZN(n7040) );
  NAND2_X1 U8898 ( .A1(n9835), .A2(n7040), .ZN(n7042) );
  NAND2_X1 U8899 ( .A1(n10020), .A2(n10024), .ZN(n7041) );
  AND2_X1 U8900 ( .A1(n10084), .A2(n9842), .ZN(n7043) );
  NAND2_X1 U8901 ( .A1(n10009), .A2(n9586), .ZN(n7044) );
  INV_X1 U8902 ( .A(n9992), .ZN(n9779) );
  NOR2_X1 U8903 ( .A1(n9996), .A2(n9982), .ZN(n7046) );
  OR2_X1 U8904 ( .A1(n9763), .A2(n9973), .ZN(n7047) );
  AND2_X1 U8905 ( .A1(n4611), .A2(n9983), .ZN(n7049) );
  OR2_X1 U8906 ( .A1(n4611), .A2(n9983), .ZN(n7048) );
  NAND2_X1 U8907 ( .A1(n9735), .A2(n9750), .ZN(n9490) );
  OR2_X2 U8908 ( .A1(n9737), .A2(n9736), .ZN(n9967) );
  NAND2_X1 U8909 ( .A1(n4426), .A2(n9974), .ZN(n7050) );
  OR2_X1 U8910 ( .A1(n9701), .A2(n9961), .ZN(n7051) );
  NAND2_X1 U8911 ( .A1(n9961), .A2(n9701), .ZN(n9690) );
  NAND2_X1 U8912 ( .A1(n9959), .A2(n9712), .ZN(n7052) );
  NAND2_X1 U8913 ( .A1(n9680), .A2(n9954), .ZN(n9426) );
  OR2_X1 U8914 ( .A1(n6930), .A2(n8410), .ZN(n7053) );
  NAND2_X1 U8915 ( .A1(n5188), .A2(n7135), .ZN(n9678) );
  NAND2_X1 U8916 ( .A1(n7603), .A2(n9457), .ZN(n7602) );
  NAND2_X1 U8917 ( .A1(n7283), .A2(n7006), .ZN(n7056) );
  INV_X1 U8918 ( .A(n9595), .ZN(n7784) );
  NAND2_X1 U8919 ( .A1(n7784), .A2(n7652), .ZN(n7058) );
  AND2_X1 U8920 ( .A1(n9595), .A2(n10231), .ZN(n9526) );
  NAND2_X1 U8921 ( .A1(n9594), .A2(n7637), .ZN(n9529) );
  NAND2_X1 U8922 ( .A1(n7847), .A2(n7781), .ZN(n9346) );
  AND2_X1 U8923 ( .A1(n9364), .A2(n9360), .ZN(n9353) );
  OAI21_X2 U8924 ( .B1(n9350), .B2(n9353), .A(n9374), .ZN(n9464) );
  AND2_X1 U8925 ( .A1(n7995), .A2(n9351), .ZN(n9362) );
  NAND2_X1 U8926 ( .A1(n9365), .A2(n9362), .ZN(n9458) );
  NOR2_X1 U8927 ( .A1(n9458), .A2(n7820), .ZN(n7061) );
  INV_X1 U8928 ( .A(n8024), .ZN(n9377) );
  NOR2_X1 U8929 ( .A1(n9461), .A2(n9377), .ZN(n7062) );
  INV_X1 U8930 ( .A(n9366), .ZN(n9371) );
  NOR2_X1 U8931 ( .A1(n9460), .A2(n9371), .ZN(n7063) );
  OR2_X1 U8932 ( .A1(n10042), .A2(n9912), .ZN(n9463) );
  AND2_X1 U8933 ( .A1(n9463), .A2(n9387), .ZN(n9550) );
  NAND2_X1 U8934 ( .A1(n9463), .A2(n9389), .ZN(n7064) );
  NAND2_X1 U8935 ( .A1(n10042), .A2(n9912), .ZN(n9462) );
  AND2_X1 U8936 ( .A1(n7064), .A2(n9462), .ZN(n7065) );
  NAND2_X1 U8937 ( .A1(n10034), .A2(n10039), .ZN(n9391) );
  XNOR2_X1 U8938 ( .A(n10020), .B(n10024), .ZN(n9840) );
  AND2_X1 U8939 ( .A1(n9840), .A2(n9838), .ZN(n7067) );
  INV_X1 U8940 ( .A(n10024), .ZN(n9861) );
  OR2_X1 U8941 ( .A1(n10020), .A2(n9861), .ZN(n9399) );
  NAND2_X1 U8942 ( .A1(n9839), .A2(n9399), .ZN(n9821) );
  NAND2_X1 U8943 ( .A1(n10084), .A2(n9233), .ZN(n9409) );
  NAND2_X1 U8944 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  NAND2_X1 U8945 ( .A1(n9819), .A2(n9410), .ZN(n9805) );
  NAND2_X1 U8946 ( .A1(n10009), .A2(n9822), .ZN(n9561) );
  NAND2_X1 U8947 ( .A1(n9805), .A2(n9806), .ZN(n9804) );
  NAND2_X1 U8948 ( .A1(n10001), .A2(n9992), .ZN(n9401) );
  NAND2_X1 U8949 ( .A1(n9996), .A2(n9792), .ZN(n9402) );
  XNOR2_X1 U8950 ( .A(n9763), .B(n9973), .ZN(n9758) );
  INV_X1 U8951 ( .A(n9973), .ZN(n9993) );
  NAND2_X1 U8952 ( .A1(n9763), .A2(n9993), .ZN(n9419) );
  OR2_X1 U8953 ( .A1(n9752), .A2(n9769), .ZN(n9421) );
  NAND2_X1 U8954 ( .A1(n9752), .A2(n9769), .ZN(n9480) );
  INV_X1 U8955 ( .A(n9426), .ZN(n7071) );
  NAND2_X1 U8956 ( .A1(n9521), .A2(n9635), .ZN(n7072) );
  NAND2_X1 U8957 ( .A1(n9665), .A2(n9988), .ZN(n7088) );
  NAND2_X1 U8958 ( .A1(n7705), .A2(n7914), .ZN(n7830) );
  INV_X1 U8959 ( .A(n10034), .ZN(n9877) );
  NAND2_X1 U8960 ( .A1(n9890), .A2(n9877), .ZN(n9862) );
  INV_X1 U8961 ( .A(n10084), .ZN(n9831) );
  INV_X1 U8962 ( .A(n10009), .ZN(n9811) );
  OAI21_X1 U8963 ( .B1(n7077), .B2(n7132), .A(n10002), .ZN(n7078) );
  OR2_X1 U8964 ( .A1(n9653), .A2(n6465), .ZN(n7084) );
  INV_X1 U8965 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8966 ( .A1(n4408), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7080) );
  NAND2_X1 U8967 ( .A1(n7106), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7079) );
  OAI211_X1 U8968 ( .C1(n7125), .C2(n7081), .A(n7080), .B(n7079), .ZN(n7082)
         );
  INV_X1 U8969 ( .A(n7082), .ZN(n7083) );
  INV_X1 U8970 ( .A(n10053), .ZN(n10038) );
  OAI22_X1 U8971 ( .A1(n9671), .A2(n10057), .B1(n9954), .B2(n10038), .ZN(n7085) );
  INV_X1 U8972 ( .A(n7085), .ZN(n7086) );
  NAND2_X1 U8973 ( .A1(n10099), .A2(n7089), .ZN(n7280) );
  NOR2_X1 U8974 ( .A1(n7280), .A2(n7090), .ZN(n7594) );
  AND2_X1 U8975 ( .A1(n7091), .A2(n7591), .ZN(n7092) );
  AND2_X2 U8976 ( .A1(n7112), .A2(n7592), .ZN(n10243) );
  NAND2_X1 U8977 ( .A1(n10243), .A2(n10049), .ZN(n10090) );
  NAND2_X1 U8978 ( .A1(n9675), .A2(n7093), .ZN(n7094) );
  INV_X1 U8979 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7113) );
  NAND2_X1 U8980 ( .A1(n10109), .A2(n7103), .ZN(n7097) );
  OR2_X1 U8981 ( .A1(n6930), .A2(n10105), .ZN(n7096) );
  OR2_X1 U8982 ( .A1(n6930), .A2(n8312), .ZN(n7099) );
  OR2_X1 U8983 ( .A1(n6930), .A2(n8338), .ZN(n7104) );
  INV_X1 U8984 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8985 ( .A1(n4408), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8986 ( .A1(n7106), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7107) );
  OAI211_X1 U8987 ( .C1(n7125), .C2(n7109), .A(n7108), .B(n7107), .ZN(n9509)
         );
  AND2_X1 U8988 ( .A1(n9518), .A2(P1_B_REG_SCAN_IN), .ZN(n7110) );
  NOR2_X1 U8989 ( .A1(n10057), .A2(n7110), .ZN(n7126) );
  AND2_X1 U8990 ( .A1(n9509), .A2(n7126), .ZN(n9640) );
  MUX2_X1 U8991 ( .A(n7113), .B(n10065), .S(n10252), .Z(n7114) );
  NAND2_X1 U8992 ( .A1(n10252), .A2(n10049), .ZN(n10032) );
  NAND2_X1 U8993 ( .A1(n7114), .A2(n5173), .ZN(P1_U3553) );
  NAND2_X1 U8994 ( .A1(n7119), .A2(n9671), .ZN(n9507) );
  NOR2_X1 U8995 ( .A1(n9648), .A2(n10210), .ZN(n7139) );
  INV_X1 U8996 ( .A(n7101), .ZN(n7120) );
  INV_X1 U8997 ( .A(n10002), .ZN(n9920) );
  AOI21_X1 U8998 ( .B1(n7120), .B2(n7119), .A(n9920), .ZN(n7121) );
  NAND3_X1 U8999 ( .A1(n9675), .A2(n9657), .A3(n10241), .ZN(n7128) );
  INV_X1 U9000 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9644) );
  INV_X1 U9001 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10534) );
  OR2_X1 U9002 ( .A1(n6982), .A2(n10534), .ZN(n7124) );
  INV_X1 U9003 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10491) );
  OR2_X1 U9004 ( .A1(n7122), .A2(n10491), .ZN(n7123) );
  OAI211_X1 U9005 ( .C1(n7125), .C2(n9644), .A(n7124), .B(n7123), .ZN(n9585)
         );
  AND2_X1 U9006 ( .A1(n9585), .A2(n7126), .ZN(n9654) );
  AOI21_X1 U9007 ( .B1(n9657), .B2(n10053), .A(n9654), .ZN(n7127) );
  INV_X1 U9008 ( .A(n7129), .ZN(n7130) );
  INV_X1 U9009 ( .A(n9651), .ZN(n7131) );
  NAND3_X1 U9010 ( .A1(n9650), .A2(n7131), .A3(n10241), .ZN(n7137) );
  NOR2_X1 U9011 ( .A1(n7132), .A2(n9947), .ZN(n9649) );
  NAND3_X1 U9012 ( .A1(n5177), .A2(n7137), .A3(n7136), .ZN(n7138) );
  INV_X1 U9013 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U9014 ( .B1(n7145), .B2(n7144), .A(n7143), .ZN(P1_U3519) );
  INV_X1 U9015 ( .A(n7148), .ZN(n7150) );
  XNOR2_X1 U9016 ( .A(n7146), .B(n7150), .ZN(n7147) );
  OAI222_X1 U9017 ( .A1(n10256), .A2(n8473), .B1(n10254), .B2(n8477), .C1(
        n8853), .C2(n7147), .ZN(n9013) );
  MUX2_X1 U9018 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n9013), .S(n10282), .Z(n7155) );
  INV_X1 U9019 ( .A(n7151), .ZN(n7149) );
  NOR2_X1 U9020 ( .A1(n7149), .A2(n7148), .ZN(n9012) );
  INV_X1 U9021 ( .A(n9014), .ZN(n7152) );
  NOR3_X1 U9022 ( .A1(n9012), .A2(n7152), .A3(n8941), .ZN(n7154) );
  OAI22_X1 U9023 ( .A1(n9102), .A2(n8744), .B1(n8480), .B2(n8912), .ZN(n7153)
         );
  OR3_X1 U9024 ( .A1(n7155), .A2(n7154), .A3(n7153), .ZN(P2_U3221) );
  NOR2_X1 U9025 ( .A1(n7156), .A2(P1_U3086), .ZN(n7157) );
  XNOR2_X1 U9026 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U9027 ( .A(n7159), .B(n7158), .S(P1_U3086), .Z(n7160) );
  INV_X1 U9028 ( .A(n7160), .ZN(P1_U3355) );
  NOR2_X1 U9029 ( .A1(n7161), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10108) );
  NOR2_X1 U9030 ( .A1(n7161), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9115) );
  INV_X2 U9031 ( .A(n9115), .ZN(n9121) );
  AND2_X1 U9032 ( .A1(n7161), .A2(P2_U3151), .ZN(n8244) );
  INV_X2 U9033 ( .A(n8244), .ZN(n9123) );
  OAI222_X1 U9034 ( .A1(P2_U3151), .A2(n5946), .B1(n9121), .B2(n5214), .C1(
        n7162), .C2(n9123), .ZN(P2_U3294) );
  OAI222_X1 U9035 ( .A1(n9121), .A2(n7164), .B1(n9123), .B2(n7174), .C1(
        P2_U3151), .C2(n7163), .ZN(P2_U3293) );
  OAI222_X1 U9036 ( .A1(P2_U3151), .A2(n7166), .B1(n9123), .B2(n7170), .C1(
        n7165), .C2(n9121), .ZN(P2_U3292) );
  OAI222_X1 U9037 ( .A1(n9121), .A2(n4846), .B1(n9123), .B2(n7175), .C1(
        P2_U3151), .C2(n7325), .ZN(P2_U3291) );
  OAI222_X1 U9038 ( .A1(P2_U3151), .A2(n7168), .B1(n9123), .B2(n7172), .C1(
        n7167), .C2(n9121), .ZN(P2_U3290) );
  OAI222_X1 U9039 ( .A1(n8337), .A2(n7170), .B1(n10116), .B2(n7169), .C1(
        P1_U3086), .C2(n7222), .ZN(P1_U3352) );
  OAI222_X1 U9040 ( .A1(n8337), .A2(n7172), .B1(n10116), .B2(n7171), .C1(
        P1_U3086), .C2(n7251), .ZN(P1_U3350) );
  OAI222_X1 U9041 ( .A1(P1_U3086), .A2(n7221), .B1(n8337), .B2(n7174), .C1(
        n7173), .C2(n10116), .ZN(P1_U3353) );
  INV_X1 U9042 ( .A(n7177), .ZN(n7181) );
  INV_X1 U9043 ( .A(n10116), .ZN(n7506) );
  AOI22_X1 U9044 ( .A1(n7290), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7506), .ZN(n7178) );
  OAI21_X1 U9045 ( .B1(n7181), .B2(n8337), .A(n7178), .ZN(P1_U3349) );
  INV_X1 U9046 ( .A(n7179), .ZN(n7555) );
  INV_X1 U9047 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7180) );
  OAI222_X1 U9048 ( .A1(P2_U3151), .A2(n7555), .B1(n9123), .B2(n7181), .C1(
        n7180), .C2(n9121), .ZN(P2_U3289) );
  AOI22_X1 U9049 ( .A1(n7468), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7506), .ZN(n7182) );
  OAI21_X1 U9050 ( .B1(n7189), .B2(n8337), .A(n7182), .ZN(P1_U3348) );
  INV_X1 U9051 ( .A(n10099), .ZN(n7183) );
  NAND2_X1 U9052 ( .A1(n7183), .A2(n9575), .ZN(n7212) );
  NAND2_X1 U9053 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  AND2_X1 U9054 ( .A1(n7186), .A2(n4421), .ZN(n7211) );
  INV_X1 U9055 ( .A(n7211), .ZN(n7187) );
  NOR2_X1 U9056 ( .A1(n10169), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U9057 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7188) );
  OAI222_X1 U9058 ( .A1(P2_U3151), .A2(n7763), .B1(n9123), .B2(n7189), .C1(
        n7188), .C2(n9121), .ZN(P2_U3288) );
  INV_X1 U9059 ( .A(n7190), .ZN(n7199) );
  AOI22_X1 U9060 ( .A1(n7541), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7506), .ZN(n7191) );
  OAI21_X1 U9061 ( .B1(n7199), .B2(n8337), .A(n7191), .ZN(P1_U3347) );
  AOI22_X1 U9062 ( .A1(n7858), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7506), .ZN(n7192) );
  OAI21_X1 U9063 ( .B1(n7196), .B2(n8337), .A(n7192), .ZN(P1_U3345) );
  AND2_X1 U9064 ( .A1(n7194), .A2(n7193), .ZN(n7236) );
  INV_X1 U9065 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10475) );
  NOR2_X1 U9066 ( .A1(n7236), .A2(n10475), .ZN(P2_U3262) );
  INV_X1 U9067 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U9068 ( .A1(n7236), .A2(n10515), .ZN(P2_U3260) );
  INV_X1 U9069 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10486) );
  NOR2_X1 U9070 ( .A1(n7236), .A2(n10486), .ZN(P2_U3238) );
  INV_X1 U9071 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10646) );
  NOR2_X1 U9072 ( .A1(n7236), .A2(n10646), .ZN(P2_U3246) );
  INV_X1 U9073 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10489) );
  NOR2_X1 U9074 ( .A1(n7236), .A2(n10489), .ZN(P2_U3236) );
  INV_X1 U9075 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U9076 ( .A1(n7236), .A2(n10562), .ZN(P2_U3249) );
  INV_X1 U9077 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10606) );
  NOR2_X1 U9078 ( .A1(n7236), .A2(n10606), .ZN(P2_U3247) );
  INV_X1 U9079 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10573) );
  NOR2_X1 U9080 ( .A1(n7236), .A2(n10573), .ZN(P2_U3256) );
  INV_X1 U9081 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7195) );
  OAI222_X1 U9082 ( .A1(P2_U3151), .A2(n7197), .B1(n9123), .B2(n7196), .C1(
        n7195), .C2(n9121), .ZN(P2_U3285) );
  OAI222_X1 U9083 ( .A1(n9121), .A2(n4700), .B1(n9123), .B2(n7199), .C1(
        P2_U3151), .C2(n7198), .ZN(P2_U3287) );
  NAND2_X1 U9084 ( .A1(n6400), .A2(P1_U3973), .ZN(n7200) );
  OAI21_X1 U9085 ( .B1(P1_U3973), .B2(n5214), .A(n7200), .ZN(P1_U3555) );
  INV_X1 U9086 ( .A(n7201), .ZN(n7203) );
  OAI222_X1 U9087 ( .A1(P2_U3151), .A2(n7202), .B1(n9123), .B2(n7203), .C1(
        n7229), .C2(n9121), .ZN(P2_U3286) );
  INV_X1 U9088 ( .A(n7773), .ZN(n7536) );
  NAND2_X1 U9089 ( .A1(n9509), .A2(P1_U3973), .ZN(n7205) );
  OAI21_X1 U9090 ( .B1(P1_U3973), .B2(n6103), .A(n7205), .ZN(P1_U3585) );
  INV_X1 U9091 ( .A(n7236), .ZN(n7206) );
  AND2_X1 U9092 ( .A1(n7206), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U9093 ( .A1(n7206), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U9094 ( .A1(n7206), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U9095 ( .A1(n7206), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U9096 ( .A1(n7206), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U9097 ( .A1(n7206), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U9098 ( .A1(n7206), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  INV_X1 U9099 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7207) );
  OAI222_X1 U9100 ( .A1(P2_U3151), .A2(n7208), .B1(n9123), .B2(n7209), .C1(
        n7207), .C2(n9121), .ZN(P2_U3283) );
  INV_X1 U9101 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7210) );
  INV_X1 U9102 ( .A(n9620), .ZN(n8092) );
  INV_X1 U9103 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U9104 ( .A1(n7212), .A2(n7211), .ZN(n10127) );
  OR2_X1 U9105 ( .A1(n10127), .A2(n7448), .ZN(n10202) );
  INV_X1 U9106 ( .A(n7222), .ZN(n7248) );
  NAND2_X1 U9107 ( .A1(n10183), .A2(n7248), .ZN(n7213) );
  NAND2_X1 U9108 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n7512) );
  OAI211_X1 U9109 ( .C1(n10607), .C2(n10207), .A(n7213), .B(n7512), .ZN(n7227)
         );
  INV_X1 U9110 ( .A(n7221), .ZN(n7458) );
  XNOR2_X1 U9111 ( .A(n7218), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9599) );
  AND2_X1 U9112 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9598) );
  NAND2_X1 U9113 ( .A1(n9599), .A2(n9598), .ZN(n9597) );
  INV_X1 U9114 ( .A(n7218), .ZN(n9604) );
  NAND2_X1 U9115 ( .A1(n9604), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U9116 ( .A1(n9597), .A2(n7214), .ZN(n7452) );
  XNOR2_X1 U9117 ( .A(n7248), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7216) );
  NOR2_X1 U9118 ( .A1(n7217), .A2(n7216), .ZN(n7243) );
  AOI211_X1 U9119 ( .C1(n7217), .C2(n7216), .A(n7243), .B(n10164), .ZN(n7226)
         );
  XNOR2_X1 U9120 ( .A(n7218), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9602) );
  AND2_X1 U9121 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9601) );
  NAND2_X1 U9122 ( .A1(n9602), .A2(n9601), .ZN(n9600) );
  NAND2_X1 U9123 ( .A1(n9604), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U9124 ( .A1(n9600), .A2(n7219), .ZN(n7456) );
  INV_X1 U9125 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10247) );
  AOI21_X1 U9126 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n7458), .A(n7454), .ZN(
        n7224) );
  XOR2_X1 U9127 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7222), .Z(n7223) );
  OR2_X1 U9128 ( .A1(n10127), .A2(n9518), .ZN(n10152) );
  AOI211_X1 U9129 ( .C1(n7224), .C2(n7223), .A(n7247), .B(n10152), .ZN(n7225)
         );
  OR3_X1 U9130 ( .A1(n7227), .A2(n7226), .A3(n7225), .ZN(P1_U3246) );
  MUX2_X1 U9131 ( .A(n4700), .B(n9257), .S(P1_U3973), .Z(n7228) );
  INV_X1 U9132 ( .A(n7228), .ZN(P1_U3562) );
  MUX2_X1 U9133 ( .A(n7229), .B(n9152), .S(P1_U3973), .Z(n7230) );
  INV_X1 U9134 ( .A(n7230), .ZN(P1_U3563) );
  INV_X1 U9135 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7232) );
  INV_X1 U9136 ( .A(n7231), .ZN(n7233) );
  OAI222_X1 U9137 ( .A1(n9121), .A2(n7232), .B1(n9123), .B2(n7233), .C1(
        P2_U3151), .C2(n8251), .ZN(P2_U3284) );
  INV_X1 U9138 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7234) );
  INV_X1 U9139 ( .A(n8097), .ZN(n7862) );
  AOI22_X1 U9140 ( .A1(n10136), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7506), .ZN(n7235) );
  OAI21_X1 U9141 ( .B1(n7273), .B2(n8337), .A(n7235), .ZN(P1_U3342) );
  INV_X1 U9142 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7239) );
  INV_X1 U9143 ( .A(n7237), .ZN(n7238) );
  AOI22_X1 U9144 ( .A1(n7206), .A2(n7239), .B1(n7238), .B2(n7241), .ZN(
        P2_U3376) );
  INV_X1 U9145 ( .A(n7240), .ZN(n7242) );
  AOI22_X1 U9146 ( .A1(n7206), .A2(n10637), .B1(n7242), .B2(n7241), .ZN(
        P2_U3377) );
  AND2_X1 U9147 ( .A1(n7206), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U9148 ( .A1(n7206), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U9149 ( .A1(n7206), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9150 ( .A1(n7206), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U9151 ( .A1(n7206), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U9152 ( .A1(n7206), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U9153 ( .A1(n7206), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U9154 ( .A1(n7206), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U9155 ( .A1(n7206), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U9156 ( .A1(n7206), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9157 ( .A1(n7206), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U9158 ( .A1(n7206), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U9159 ( .A1(n7206), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U9160 ( .A1(n7206), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U9161 ( .A1(n7206), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  INV_X1 U9162 ( .A(n7249), .ZN(n7482) );
  INV_X1 U9163 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7244) );
  MUX2_X1 U9164 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7244), .S(n7249), .Z(n7477)
         );
  NOR2_X1 U9165 ( .A1(n7478), .A2(n7477), .ZN(n7476) );
  AOI21_X1 U9166 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n7482), .A(n7476), .ZN(
        n7246) );
  INV_X1 U9167 ( .A(n7251), .ZN(n7264) );
  XNOR2_X1 U9168 ( .A(n7264), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n7245) );
  AOI211_X1 U9169 ( .C1(n7246), .C2(n7245), .A(n10164), .B(n7263), .ZN(n7258)
         );
  INV_X1 U9170 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7250) );
  MUX2_X1 U9171 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7250), .S(n7249), .Z(n7480)
         );
  XOR2_X1 U9172 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7251), .Z(n7252) );
  NOR2_X1 U9173 ( .A1(n7253), .A2(n7252), .ZN(n7259) );
  AOI211_X1 U9174 ( .C1(n7253), .C2(n7252), .A(n10152), .B(n7259), .ZN(n7257)
         );
  INV_X1 U9175 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U9176 ( .A1(n10183), .A2(n7264), .ZN(n7254) );
  NAND2_X1 U9177 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7846) );
  OAI211_X1 U9178 ( .C1(n7255), .C2(n10207), .A(n7254), .B(n7846), .ZN(n7256)
         );
  OR3_X1 U9179 ( .A1(n7258), .A2(n7257), .A3(n7256), .ZN(P1_U3248) );
  INV_X1 U9180 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7260) );
  MUX2_X1 U9181 ( .A(n7260), .B(P1_REG1_REG_6__SCAN_IN), .S(n7290), .Z(n7261)
         );
  NOR2_X1 U9182 ( .A1(n7262), .A2(n7261), .ZN(n7286) );
  AOI211_X1 U9183 ( .C1(n7262), .C2(n7261), .A(n10152), .B(n7286), .ZN(n7271)
         );
  INV_X1 U9184 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7265) );
  MUX2_X1 U9185 ( .A(n7265), .B(P1_REG2_REG_6__SCAN_IN), .S(n7290), .Z(n7266)
         );
  AOI211_X1 U9186 ( .C1(n7267), .C2(n7266), .A(n10164), .B(n7289), .ZN(n7270)
         );
  INV_X1 U9187 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U9188 ( .A1(n10183), .A2(n7290), .ZN(n7268) );
  NAND2_X1 U9189 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7810) );
  OAI211_X1 U9190 ( .C1(n10470), .C2(n10207), .A(n7268), .B(n7810), .ZN(n7269)
         );
  OR3_X1 U9191 ( .A1(n7271), .A2(n7270), .A3(n7269), .ZN(P1_U3249) );
  INV_X1 U9192 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7272) );
  OAI222_X1 U9193 ( .A1(P2_U3151), .A2(n7274), .B1(n9123), .B2(n7273), .C1(
        n7272), .C2(n9121), .ZN(P2_U3282) );
  MUX2_X1 U9194 ( .A(n7275), .B(n8894), .S(P2_U3893), .Z(n7276) );
  INV_X1 U9195 ( .A(n7276), .ZN(P2_U3508) );
  OAI21_X1 U9196 ( .B1(n7279), .B2(n7278), .A(n7277), .ZN(n7446) );
  INV_X1 U9197 ( .A(n7280), .ZN(n7281) );
  NAND2_X1 U9198 ( .A1(n7282), .A2(n7281), .ZN(n7443) );
  INV_X1 U9199 ( .A(n9326), .ZN(n9334) );
  OAI22_X1 U9200 ( .A1(n9334), .A2(n7283), .B1(n9335), .B2(n9527), .ZN(n7284)
         );
  AOI21_X1 U9201 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7443), .A(n7284), .ZN(
        n7285) );
  OAI21_X1 U9202 ( .B1(n7446), .B2(n9340), .A(n7285), .ZN(P1_U3232) );
  AOI21_X1 U9203 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n7290), .A(n7286), .ZN(
        n7288) );
  XNOR2_X1 U9204 ( .A(n7468), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n7287) );
  NOR2_X1 U9205 ( .A1(n7288), .A2(n7287), .ZN(n7464) );
  AOI211_X1 U9206 ( .C1(n7288), .C2(n7287), .A(n10152), .B(n7464), .ZN(n7297)
         );
  XNOR2_X1 U9207 ( .A(n7468), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7291) );
  AOI211_X1 U9208 ( .C1(n7292), .C2(n7291), .A(n10164), .B(n7467), .ZN(n7296)
         );
  INV_X1 U9209 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U9210 ( .A1(n10183), .A2(n7468), .ZN(n7293) );
  NAND2_X1 U9211 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7870) );
  OAI211_X1 U9212 ( .C1(n7294), .C2(n10207), .A(n7293), .B(n7870), .ZN(n7295)
         );
  OR3_X1 U9213 ( .A1(n7297), .A2(n7296), .A3(n7295), .ZN(P1_U3250) );
  INV_X1 U9214 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7304) );
  XNOR2_X1 U9215 ( .A(n7298), .B(n5107), .ZN(n7299) );
  AOI21_X1 U9216 ( .B1(n8722), .B2(n7300), .A(n7299), .ZN(n7301) );
  AOI21_X1 U9217 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7301), .ZN(
        n7303) );
  NAND2_X1 U9218 ( .A1(n8632), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7302) );
  OAI211_X1 U9219 ( .C1(n8721), .C2(n7304), .A(n7303), .B(n7302), .ZN(P2_U3182) );
  OAI211_X1 U9220 ( .C1(n7307), .C2(n7306), .A(n7305), .B(n8704), .ZN(n7324)
         );
  INV_X1 U9221 ( .A(n7308), .ZN(n7310) );
  NOR2_X1 U9222 ( .A1(n7310), .A2(n7309), .ZN(n7314) );
  INV_X1 U9223 ( .A(n7312), .ZN(n7313) );
  AOI21_X1 U9224 ( .B1(n7314), .B2(n7311), .A(n7313), .ZN(n7315) );
  NAND2_X1 U9225 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7578) );
  OAI21_X1 U9226 ( .B1(n8655), .B2(n7315), .A(n7578), .ZN(n7322) );
  INV_X1 U9227 ( .A(n7316), .ZN(n7318) );
  NAND3_X1 U9228 ( .A1(n7333), .A2(n7318), .A3(n7317), .ZN(n7319) );
  AOI21_X1 U9229 ( .B1(n7320), .B2(n7319), .A(n8734), .ZN(n7321) );
  AOI211_X1 U9230 ( .C1(n8699), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7322), .B(
        n7321), .ZN(n7323) );
  OAI211_X1 U9231 ( .C1(n8717), .C2(n7325), .A(n7324), .B(n7323), .ZN(P2_U3186) );
  INV_X1 U9232 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7327) );
  INV_X1 U9233 ( .A(n7326), .ZN(n7329) );
  OAI222_X1 U9234 ( .A1(n9121), .A2(n7327), .B1(n9123), .B2(n7329), .C1(
        P2_U3151), .C2(n8645), .ZN(P2_U3281) );
  INV_X1 U9235 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10549) );
  INV_X1 U9236 ( .A(n10148), .ZN(n7328) );
  AOI21_X1 U9237 ( .B1(n7332), .B2(n7331), .A(n7330), .ZN(n7342) );
  INV_X1 U9238 ( .A(n8734), .ZN(n8639) );
  OAI21_X1 U9239 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n7334), .A(n7333), .ZN(
        n7335) );
  AOI22_X1 U9240 ( .A1(n8699), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n8639), .B2(
        n7335), .ZN(n7339) );
  NOR2_X1 U9241 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10294), .ZN(n7526) );
  INV_X1 U9242 ( .A(n7526), .ZN(n7338) );
  OAI21_X1 U9243 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n4540), .A(n7311), .ZN(
        n7336) );
  NAND2_X1 U9244 ( .A1(n8730), .A2(n7336), .ZN(n7337) );
  NAND3_X1 U9245 ( .A1(n7339), .A2(n7338), .A3(n7337), .ZN(n7340) );
  AOI21_X1 U9246 ( .B1(n4892), .B2(n8632), .A(n7340), .ZN(n7341) );
  OAI21_X1 U9247 ( .B1(n7342), .B2(n8722), .A(n7341), .ZN(P2_U3185) );
  INV_X1 U9248 ( .A(n7421), .ZN(n7413) );
  OAI21_X1 U9249 ( .B1(n10289), .B2(n10327), .A(n7413), .ZN(n7344) );
  NOR2_X1 U9250 ( .A1(n5244), .A2(n10254), .ZN(n7422) );
  INV_X1 U9251 ( .A(n7422), .ZN(n7343) );
  OAI211_X1 U9252 ( .C1(n10330), .C2(n7427), .A(n7344), .B(n7343), .ZN(n7416)
         );
  NAND2_X1 U9253 ( .A1(n7416), .A2(n10672), .ZN(n7345) );
  OAI21_X1 U9254 ( .B1(n10672), .B2(n6012), .A(n7345), .ZN(P2_U3459) );
  OAI211_X1 U9255 ( .C1(n7348), .C2(n7347), .A(n8704), .B(n7346), .ZN(n7349)
         );
  OAI21_X1 U9256 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7716), .A(n7349), .ZN(n7358) );
  OAI21_X1 U9257 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n7351), .A(n7350), .ZN(
        n7355) );
  OAI21_X1 U9258 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n7353), .A(n7352), .ZN(
        n7354) );
  AOI22_X1 U9259 ( .A1(n8639), .A2(n7355), .B1(n8730), .B2(n7354), .ZN(n7356)
         );
  INV_X1 U9260 ( .A(n7356), .ZN(n7357) );
  AOI211_X1 U9261 ( .C1(n8699), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7358), .B(
        n7357), .ZN(n7359) );
  OAI21_X1 U9262 ( .B1(n5946), .B2(n8717), .A(n7359), .ZN(P2_U3183) );
  INV_X1 U9263 ( .A(n7443), .ZN(n7368) );
  OAI21_X1 U9264 ( .B1(n7362), .B2(n7361), .A(n7360), .ZN(n7363) );
  NAND2_X1 U9265 ( .A1(n7363), .A2(n9320), .ZN(n7367) );
  OAI22_X1 U9266 ( .A1(n9334), .A2(n7514), .B1(n7364), .B2(n9324), .ZN(n7365)
         );
  AOI21_X1 U9267 ( .B1(n7006), .B2(n9272), .A(n7365), .ZN(n7366) );
  OAI211_X1 U9268 ( .C1(n7368), .C2(n6381), .A(n7367), .B(n7366), .ZN(P1_U3222) );
  INV_X1 U9269 ( .A(n7369), .ZN(n7376) );
  INV_X1 U9270 ( .A(n7370), .ZN(n7396) );
  NAND3_X1 U9271 ( .A1(n7373), .A2(n7372), .A3(n7371), .ZN(n7374) );
  AOI21_X1 U9272 ( .B1(n7379), .B2(n7396), .A(n7374), .ZN(n7375) );
  OAI21_X1 U9273 ( .B1(n7377), .B2(n7376), .A(n7375), .ZN(n7378) );
  NAND2_X1 U9274 ( .A1(n7378), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7382) );
  NAND2_X1 U9275 ( .A1(n7380), .A2(n7379), .ZN(n7381) );
  NOR2_X1 U9276 ( .A1(n8594), .A2(P2_U3151), .ZN(n7504) );
  INV_X1 U9277 ( .A(n7383), .ZN(n7389) );
  NAND2_X1 U9278 ( .A1(n7385), .A2(n7384), .ZN(n7387) );
  AND2_X2 U9279 ( .A1(n7387), .A2(n7386), .ZN(n7388) );
  NAND2_X2 U9280 ( .A1(n7389), .A2(n7388), .ZN(n7520) );
  NOR2_X1 U9281 ( .A1(n8609), .A2(n7390), .ZN(n7494) );
  NOR2_X2 U9282 ( .A1(n7494), .A2(n7391), .ZN(n7394) );
  INV_X4 U9283 ( .A(n7520), .ZN(n8364) );
  OAI21_X1 U9284 ( .B1(n7392), .B2(n8364), .A(n7713), .ZN(n7393) );
  OAI21_X1 U9285 ( .B1(n7394), .B2(n7393), .A(n7496), .ZN(n7399) );
  OR2_X1 U9286 ( .A1(n7400), .A2(n7395), .ZN(n7398) );
  NAND2_X1 U9287 ( .A1(n7406), .A2(n7396), .ZN(n7397) );
  NAND2_X1 U9288 ( .A1(n7399), .A2(n8587), .ZN(n7411) );
  OR2_X1 U9289 ( .A1(n7400), .A2(n8791), .ZN(n7401) );
  NOR2_X1 U9290 ( .A1(n7419), .A2(n7402), .ZN(n7403) );
  NAND2_X1 U9291 ( .A1(n7406), .A2(n7403), .ZN(n8592) );
  NOR2_X1 U9292 ( .A1(n7419), .A2(n7404), .ZN(n7405) );
  NAND2_X1 U9293 ( .A1(n7406), .A2(n7405), .ZN(n8577) );
  OAI22_X1 U9294 ( .A1(n7528), .A2(n8592), .B1(n8577), .B2(n7407), .ZN(n7408)
         );
  AOI21_X1 U9295 ( .B1(n7409), .B2(n8568), .A(n7408), .ZN(n7410) );
  OAI211_X1 U9296 ( .C1(n7504), .C2(n7716), .A(n7411), .B(n7410), .ZN(P2_U3162) );
  OAI22_X1 U9297 ( .A1(n8597), .A2(n7427), .B1(n5244), .B2(n8592), .ZN(n7412)
         );
  AOI21_X1 U9298 ( .B1(n7413), .B2(n8587), .A(n7412), .ZN(n7414) );
  OAI21_X1 U9299 ( .B1(n7504), .B2(n7415), .A(n7414), .ZN(P2_U3172) );
  INV_X1 U9300 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9301 ( .A1(n7416), .A2(n10336), .ZN(n7417) );
  OAI21_X1 U9302 ( .B1(n7418), .B2(n10336), .A(n7417), .ZN(P2_U3390) );
  INV_X1 U9303 ( .A(n7419), .ZN(n7420) );
  NOR3_X1 U9304 ( .A1(n7421), .A2(n7420), .A3(n10316), .ZN(n7424) );
  NOR2_X1 U9305 ( .A1(n8912), .A2(n7415), .ZN(n7423) );
  NOR3_X1 U9306 ( .A1(n7424), .A2(n7423), .A3(n7422), .ZN(n7425) );
  MUX2_X1 U9307 ( .A(n5109), .B(n7425), .S(n10282), .Z(n7426) );
  OAI21_X1 U9308 ( .B1(n8744), .B2(n7427), .A(n7426), .ZN(P2_U3233) );
  OAI211_X1 U9309 ( .C1(n7430), .C2(n7429), .A(n7428), .B(n8704), .ZN(n7438)
         );
  INV_X1 U9310 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7435) );
  OAI21_X1 U9311 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n7431), .A(n7563), .ZN(
        n7433) );
  OAI21_X1 U9312 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n4536), .A(n7559), .ZN(
        n7432) );
  AOI22_X1 U9313 ( .A1(n8639), .A2(n7433), .B1(n8730), .B2(n7432), .ZN(n7434)
         );
  NAND2_X1 U9314 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7692) );
  OAI211_X1 U9315 ( .C1(n8721), .C2(n7435), .A(n7434), .B(n7692), .ZN(n7436)
         );
  AOI21_X1 U9316 ( .B1(n5986), .B2(n8632), .A(n7436), .ZN(n7437) );
  NAND2_X1 U9317 ( .A1(n7438), .A2(n7437), .ZN(P2_U3187) );
  XOR2_X1 U9318 ( .A(n7440), .B(n7439), .Z(n7445) );
  INV_X1 U9319 ( .A(n9324), .ZN(n9332) );
  AOI22_X1 U9320 ( .A1(n9332), .A2(n6400), .B1(n9326), .B2(n9595), .ZN(n7441)
         );
  OAI21_X1 U9321 ( .B1(n10225), .B2(n9335), .A(n7441), .ZN(n7442) );
  AOI21_X1 U9322 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7443), .A(n7442), .ZN(
        n7444) );
  OAI21_X1 U9323 ( .B1(n7445), .B2(n9340), .A(n7444), .ZN(P1_U3237) );
  NOR2_X1 U9324 ( .A1(n4429), .A2(n7447), .ZN(n10120) );
  NOR2_X1 U9325 ( .A1(n10120), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10119) );
  INV_X2 U9326 ( .A(P1_U3973), .ZN(n9596) );
  AOI211_X1 U9327 ( .C1(n7449), .C2(n7448), .A(n10119), .B(n9596), .ZN(n7488)
         );
  INV_X1 U9328 ( .A(n10164), .ZN(n10193) );
  INV_X1 U9329 ( .A(n7450), .ZN(n7451) );
  OAI211_X1 U9330 ( .C1(n7453), .C2(n7452), .A(n10193), .B(n7451), .ZN(n7462)
         );
  AOI22_X1 U9331 ( .A1(n10169), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7461) );
  INV_X1 U9332 ( .A(n10152), .ZN(n10198) );
  INV_X1 U9333 ( .A(n7454), .ZN(n7455) );
  OAI211_X1 U9334 ( .C1(n7457), .C2(n7456), .A(n10198), .B(n7455), .ZN(n7460)
         );
  NAND2_X1 U9335 ( .A1(n10183), .A2(n7458), .ZN(n7459) );
  NAND4_X1 U9336 ( .A1(n7462), .A2(n7461), .A3(n7460), .A4(n7459), .ZN(n7463)
         );
  OR2_X1 U9337 ( .A1(n7488), .A2(n7463), .ZN(P1_U3245) );
  XNOR2_X1 U9338 ( .A(n7541), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7465) );
  AOI211_X1 U9339 ( .C1(n7466), .C2(n7465), .A(n10152), .B(n7540), .ZN(n7475)
         );
  XNOR2_X1 U9340 ( .A(n7541), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7469) );
  AOI211_X1 U9341 ( .C1(n7470), .C2(n7469), .A(n10164), .B(n7532), .ZN(n7474)
         );
  INV_X1 U9342 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7472) );
  NAND2_X1 U9343 ( .A1(n10183), .A2(n7541), .ZN(n7471) );
  NAND2_X1 U9344 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9174) );
  OAI211_X1 U9345 ( .C1(n7472), .C2(n10207), .A(n7471), .B(n9174), .ZN(n7473)
         );
  OR3_X1 U9346 ( .A1(n7475), .A2(n7474), .A3(n7473), .ZN(P1_U3251) );
  AOI211_X1 U9347 ( .C1(n7478), .C2(n7477), .A(n7476), .B(n10164), .ZN(n7487)
         );
  AOI211_X1 U9348 ( .C1(n7481), .C2(n7480), .A(n7479), .B(n10152), .ZN(n7486)
         );
  INV_X1 U9349 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9350 ( .A1(n10183), .A2(n7482), .ZN(n7483) );
  NAND2_X1 U9351 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7782) );
  OAI211_X1 U9352 ( .C1(n7484), .C2(n10207), .A(n7483), .B(n7782), .ZN(n7485)
         );
  OR4_X1 U9353 ( .A1(n7488), .A2(n7487), .A3(n7486), .A4(n7485), .ZN(P1_U3247)
         );
  INV_X1 U9354 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7491) );
  INV_X1 U9355 ( .A(n7489), .ZN(n7492) );
  OAI222_X1 U9356 ( .A1(n9121), .A2(n7491), .B1(n9123), .B2(n7492), .C1(
        P2_U3151), .C2(n4899), .ZN(P2_U3280) );
  INV_X1 U9357 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7493) );
  XNOR2_X1 U9358 ( .A(n8364), .B(n10302), .ZN(n7518) );
  XNOR2_X1 U9359 ( .A(n7518), .B(n7528), .ZN(n7498) );
  INV_X1 U9360 ( .A(n7494), .ZN(n7495) );
  OAI21_X1 U9361 ( .B1(n7498), .B2(n7497), .A(n7523), .ZN(n7499) );
  NAND2_X1 U9362 ( .A1(n7499), .A2(n8587), .ZN(n7503) );
  OAI22_X1 U9363 ( .A1(n7617), .A2(n8592), .B1(n8577), .B2(n5244), .ZN(n7500)
         );
  AOI21_X1 U9364 ( .B1(n7501), .B2(n8568), .A(n7500), .ZN(n7502) );
  OAI211_X1 U9365 ( .C1(n7504), .C2(n7621), .A(n7503), .B(n7502), .ZN(P2_U3177) );
  INV_X1 U9366 ( .A(n7505), .ZN(n7508) );
  AOI22_X1 U9367 ( .A1(n10184), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7506), .ZN(n7507) );
  OAI21_X1 U9368 ( .B1(n7508), .B2(n8337), .A(n7507), .ZN(P1_U3338) );
  OAI222_X1 U9369 ( .A1(n9121), .A2(n7509), .B1(n9123), .B2(n7508), .C1(
        P2_U3151), .C2(n8702), .ZN(P2_U3278) );
  XOR2_X1 U9370 ( .A(n4416), .B(n7510), .Z(n7517) );
  AOI22_X1 U9371 ( .A1(n9272), .A2(n7652), .B1(n9326), .B2(n9594), .ZN(n7513)
         );
  OAI211_X1 U9372 ( .C1(n7514), .C2(n9324), .A(n7513), .B(n7512), .ZN(n7515)
         );
  AOI21_X1 U9373 ( .B1(n7651), .B2(n9338), .A(n7515), .ZN(n7516) );
  OAI21_X1 U9374 ( .B1(n7517), .B2(n9340), .A(n7516), .ZN(P1_U3218) );
  INV_X1 U9375 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U9376 ( .A1(n7519), .A2(n7528), .ZN(n7522) );
  AND2_X1 U9377 ( .A1(n7523), .A2(n7522), .ZN(n7525) );
  XNOR2_X1 U9378 ( .A(n8381), .B(n7521), .ZN(n7572) );
  XNOR2_X1 U9379 ( .A(n7572), .B(n10276), .ZN(n7524) );
  OAI211_X1 U9380 ( .C1(n7525), .C2(n7524), .A(n8587), .B(n7571), .ZN(n7531)
         );
  AOI21_X1 U9381 ( .B1(n8580), .B2(n10285), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9382 ( .B1(n7528), .B2(n8577), .A(n7527), .ZN(n7529) );
  AOI21_X1 U9383 ( .B1(n6121), .B2(n8568), .A(n7529), .ZN(n7530) );
  OAI211_X1 U9384 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8566), .A(n7531), .B(
        n7530), .ZN(P2_U3158) );
  XOR2_X1 U9385 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7773), .Z(n7534) );
  OAI21_X1 U9386 ( .B1(n7534), .B2(n7533), .A(n7768), .ZN(n7538) );
  NAND2_X1 U9387 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U9388 ( .A1(n10169), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n7535) );
  OAI211_X1 U9389 ( .C1(n10202), .C2(n7536), .A(n9256), .B(n7535), .ZN(n7537)
         );
  AOI21_X1 U9390 ( .B1(n7538), .B2(n10193), .A(n7537), .ZN(n7546) );
  XNOR2_X1 U9391 ( .A(n7773), .B(n7539), .ZN(n7543) );
  OAI21_X1 U9392 ( .B1(n7543), .B2(n7542), .A(n7772), .ZN(n7544) );
  NAND2_X1 U9393 ( .A1(n7544), .A2(n10198), .ZN(n7545) );
  NAND2_X1 U9394 ( .A1(n7546), .A2(n7545), .ZN(P1_U3252) );
  INV_X1 U9395 ( .A(n7547), .ZN(n7550) );
  INV_X1 U9396 ( .A(n10172), .ZN(n9618) );
  OAI222_X1 U9397 ( .A1(P2_U3151), .A2(n8684), .B1(n9123), .B2(n7550), .C1(
        n7549), .C2(n9121), .ZN(P2_U3279) );
  AOI21_X1 U9398 ( .B1(n7553), .B2(n7552), .A(n7551), .ZN(n7570) );
  NAND2_X1 U9399 ( .A1(n8699), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9400 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7800) );
  OAI211_X1 U9401 ( .C1(n8717), .C2(n7555), .A(n7554), .B(n7800), .ZN(n7568)
         );
  INV_X1 U9402 ( .A(n7556), .ZN(n7558) );
  NAND3_X1 U9403 ( .A1(n7559), .A2(n7558), .A3(n7557), .ZN(n7560) );
  AOI21_X1 U9404 ( .B1(n7561), .B2(n7560), .A(n8655), .ZN(n7567) );
  NAND3_X1 U9405 ( .A1(n7563), .A2(n4539), .A3(n7562), .ZN(n7564) );
  AOI21_X1 U9406 ( .B1(n7565), .B2(n7564), .A(n8734), .ZN(n7566) );
  NOR3_X1 U9407 ( .A1(n7568), .A2(n7567), .A3(n7566), .ZN(n7569) );
  OAI21_X1 U9408 ( .B1(n7570), .B2(n8722), .A(n7569), .ZN(P2_U3188) );
  XNOR2_X1 U9409 ( .A(n8381), .B(n7573), .ZN(n7574) );
  NAND2_X1 U9410 ( .A1(n7574), .A2(n7894), .ZN(n7687) );
  OAI21_X1 U9411 ( .B1(n7574), .B2(n7894), .A(n7687), .ZN(n7575) );
  AOI21_X1 U9412 ( .B1(n7576), .B2(n7575), .A(n7688), .ZN(n7584) );
  INV_X1 U9413 ( .A(n7577), .ZN(n10280) );
  NAND2_X1 U9414 ( .A1(n8568), .A2(n10311), .ZN(n7581) );
  INV_X1 U9415 ( .A(n7578), .ZN(n7579) );
  AOI21_X1 U9416 ( .B1(n8580), .B2(n10275), .A(n7579), .ZN(n7580) );
  OAI211_X1 U9417 ( .C1(n7617), .C2(n8577), .A(n7581), .B(n7580), .ZN(n7582)
         );
  AOI21_X1 U9418 ( .B1(n10280), .B2(n8594), .A(n7582), .ZN(n7583) );
  OAI21_X1 U9419 ( .B1(n7584), .B2(n8570), .A(n7583), .ZN(P2_U3170) );
  INV_X1 U9420 ( .A(n7585), .ZN(n7612) );
  AOI22_X1 U9421 ( .A1(n8727), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9115), .ZN(n7586) );
  OAI21_X1 U9422 ( .B1(n7612), .B2(n9123), .A(n7586), .ZN(P2_U3277) );
  INV_X1 U9423 ( .A(n7587), .ZN(n7588) );
  NAND2_X1 U9424 ( .A1(n9457), .A2(n7588), .ZN(n7589) );
  NAND2_X1 U9425 ( .A1(n7590), .A2(n7589), .ZN(n10217) );
  INV_X1 U9426 ( .A(n10217), .ZN(n7611) );
  INV_X1 U9427 ( .A(n7591), .ZN(n7593) );
  NAND3_X1 U9428 ( .A1(n7594), .A2(n7593), .A3(n7592), .ZN(n7595) );
  INV_X1 U9429 ( .A(n7648), .ZN(n7596) );
  NAND2_X1 U9430 ( .A1(n9854), .A2(n7596), .ZN(n7610) );
  NAND2_X1 U9431 ( .A1(n9854), .A2(n7597), .ZN(n9926) );
  INV_X1 U9432 ( .A(n9933), .ZN(n9893) );
  INV_X1 U9433 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7598) );
  OAI22_X1 U9434 ( .A1(n9893), .A2(n7598), .B1(n6381), .B2(n9891), .ZN(n7600)
         );
  NAND2_X1 U9435 ( .A1(n9854), .A2(n9629), .ZN(n9863) );
  OAI211_X1 U9436 ( .C1(n7073), .C2(n9527), .A(n10002), .B(n7739), .ZN(n10218)
         );
  NOR2_X1 U9437 ( .A1(n9863), .A2(n10218), .ZN(n7599) );
  AOI211_X1 U9438 ( .C1(n9930), .C2(n7006), .A(n7600), .B(n7599), .ZN(n7609)
         );
  INV_X1 U9439 ( .A(n7649), .ZN(n7601) );
  NAND2_X1 U9440 ( .A1(n10217), .A2(n7601), .ZN(n7607) );
  OAI21_X1 U9441 ( .B1(n7603), .B2(n9457), .A(n7602), .ZN(n7604) );
  NAND2_X1 U9442 ( .A1(n7604), .A2(n9988), .ZN(n7606) );
  NAND3_X1 U9443 ( .A1(n7607), .A2(n7606), .A3(n7605), .ZN(n10221) );
  NAND2_X1 U9444 ( .A1(n10221), .A2(n9893), .ZN(n7608) );
  OAI211_X1 U9445 ( .C1(n7611), .C2(n7610), .A(n7609), .B(n7608), .ZN(P1_U3292) );
  INV_X1 U9446 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10623) );
  INV_X1 U9447 ( .A(n9625), .ZN(n10201) );
  XNOR2_X1 U9448 ( .A(n7613), .B(n7615), .ZN(n10303) );
  NAND2_X1 U9449 ( .A1(n10282), .A2(n7614), .ZN(n10267) );
  INV_X1 U9450 ( .A(n7902), .ZN(n10262) );
  XNOR2_X1 U9451 ( .A(n7616), .B(n7615), .ZN(n7619) );
  OAI22_X1 U9452 ( .A1(n7617), .A2(n10254), .B1(n5244), .B2(n10256), .ZN(n7618) );
  AOI21_X1 U9453 ( .B1(n7619), .B2(n10289), .A(n7618), .ZN(n7620) );
  OAI21_X1 U9454 ( .B1(n10303), .B2(n10262), .A(n7620), .ZN(n10305) );
  OAI22_X1 U9455 ( .A1(n8912), .A2(n7621), .B1(n10302), .B2(n8791), .ZN(n7622)
         );
  NOR2_X1 U9456 ( .A1(n10305), .A2(n7622), .ZN(n7623) );
  MUX2_X1 U9457 ( .A(n7624), .B(n7623), .S(n10282), .Z(n7625) );
  OAI21_X1 U9458 ( .B1(n10303), .B2(n10267), .A(n7625), .ZN(P2_U3231) );
  XOR2_X1 U9459 ( .A(n7626), .B(n9454), .Z(n7677) );
  XNOR2_X1 U9460 ( .A(n9595), .B(n7652), .ZN(n9455) );
  INV_X1 U9461 ( .A(n9455), .ZN(n7646) );
  NAND2_X1 U9462 ( .A1(n7647), .A2(n7646), .ZN(n7645) );
  INV_X1 U9463 ( .A(n7627), .ZN(n7628) );
  NAND2_X1 U9464 ( .A1(n7645), .A2(n7628), .ZN(n7629) );
  NAND2_X1 U9465 ( .A1(n7629), .A2(n9454), .ZN(n7664) );
  OAI21_X1 U9466 ( .B1(n7629), .B2(n9454), .A(n7664), .ZN(n7684) );
  INV_X1 U9467 ( .A(n7684), .ZN(n7633) );
  AOI22_X1 U9468 ( .A1(n9593), .A2(n10212), .B1(n10053), .B2(n9595), .ZN(n7632) );
  AOI21_X1 U9469 ( .B1(n7630), .B2(n7781), .A(n9920), .ZN(n7631) );
  NAND2_X1 U9470 ( .A1(n7631), .A2(n7666), .ZN(n7682) );
  OAI211_X1 U9471 ( .C1(n7633), .C2(n10211), .A(n7632), .B(n7682), .ZN(n7634)
         );
  AOI21_X1 U9472 ( .B1(n7677), .B2(n9988), .A(n7634), .ZN(n7640) );
  AOI22_X1 U9473 ( .A1(n10063), .A2(n7781), .B1(n4409), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7635) );
  OAI21_X1 U9474 ( .B1(n7640), .B2(n4409), .A(n7635), .ZN(P1_U3526) );
  INV_X1 U9475 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7636) );
  OAI22_X1 U9476 ( .A1(n10090), .A2(n7637), .B1(n10243), .B2(n7636), .ZN(n7638) );
  INV_X1 U9477 ( .A(n7638), .ZN(n7639) );
  OAI21_X1 U9478 ( .B1(n7640), .B2(n7144), .A(n7639), .ZN(P1_U3465) );
  XNOR2_X1 U9479 ( .A(n7641), .B(n7646), .ZN(n7642) );
  NAND2_X1 U9480 ( .A1(n7642), .A2(n9988), .ZN(n7644) );
  AOI22_X1 U9481 ( .A1(n10053), .A2(n7009), .B1(n9594), .B2(n10212), .ZN(n7643) );
  NAND2_X1 U9482 ( .A1(n7644), .A2(n7643), .ZN(n10232) );
  INV_X1 U9483 ( .A(n10232), .ZN(n7657) );
  OAI21_X1 U9484 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n10234) );
  NAND2_X1 U9485 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  OAI211_X1 U9486 ( .C1(n7738), .C2(n10231), .A(n7630), .B(n10002), .ZN(n10230) );
  INV_X1 U9487 ( .A(n9891), .ZN(n9932) );
  AOI22_X1 U9488 ( .A1(n9933), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9932), .B2(
        n7651), .ZN(n7654) );
  NAND2_X1 U9489 ( .A1(n9930), .A2(n7652), .ZN(n7653) );
  OAI211_X1 U9490 ( .C1(n10230), .C2(n9863), .A(n7654), .B(n7653), .ZN(n7655)
         );
  AOI21_X1 U9491 ( .B1(n10234), .B2(n9928), .A(n7655), .ZN(n7656) );
  OAI21_X1 U9492 ( .B1(n7657), .B2(n9933), .A(n7656), .ZN(P1_U3290) );
  INV_X1 U9493 ( .A(n7059), .ZN(n7659) );
  XNOR2_X1 U9494 ( .A(n7658), .B(n7659), .ZN(n7660) );
  NAND2_X1 U9495 ( .A1(n7660), .A2(n9988), .ZN(n7662) );
  AOI22_X1 U9496 ( .A1(n10212), .A2(n9592), .B1(n9594), .B2(n10053), .ZN(n7661) );
  NAND2_X1 U9497 ( .A1(n7662), .A2(n7661), .ZN(n10238) );
  INV_X1 U9498 ( .A(n10238), .ZN(n7676) );
  NAND2_X1 U9499 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  NAND2_X1 U9500 ( .A1(n7665), .A2(n7059), .ZN(n7703) );
  OAI21_X1 U9501 ( .B1(n7665), .B2(n7059), .A(n7703), .ZN(n10240) );
  INV_X1 U9502 ( .A(n7666), .ZN(n7669) );
  INV_X1 U9503 ( .A(n7667), .ZN(n7668) );
  OAI211_X1 U9504 ( .C1(n5051), .C2(n7669), .A(n7668), .B(n10002), .ZN(n10236)
         );
  OAI22_X1 U9505 ( .A1(n9893), .A2(n7670), .B1(n7852), .B2(n9891), .ZN(n7671)
         );
  AOI21_X1 U9506 ( .B1(n9930), .B2(n7672), .A(n7671), .ZN(n7673) );
  OAI21_X1 U9507 ( .B1(n10236), .B2(n9863), .A(n7673), .ZN(n7674) );
  AOI21_X1 U9508 ( .B1(n10240), .B2(n9928), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9509 ( .B1(n7676), .B2(n9933), .A(n7675), .ZN(P1_U3288) );
  INV_X1 U9510 ( .A(n7677), .ZN(n7686) );
  NAND2_X1 U9511 ( .A1(n9854), .A2(n9988), .ZN(n9871) );
  NAND2_X1 U9512 ( .A1(n9854), .A2(n10212), .ZN(n9894) );
  INV_X1 U9513 ( .A(n9894), .ZN(n9936) );
  AOI22_X1 U9514 ( .A1(n9936), .A2(n9593), .B1(n9898), .B2(n9595), .ZN(n7681)
         );
  OAI22_X1 U9515 ( .A1(n9893), .A2(n7244), .B1(n7678), .B2(n9891), .ZN(n7679)
         );
  AOI21_X1 U9516 ( .B1(n9930), .B2(n7781), .A(n7679), .ZN(n7680) );
  OAI211_X1 U9517 ( .C1(n9863), .C2(n7682), .A(n7681), .B(n7680), .ZN(n7683)
         );
  AOI21_X1 U9518 ( .B1(n7684), .B2(n9928), .A(n7683), .ZN(n7685) );
  OAI21_X1 U9519 ( .B1(n7686), .B2(n9871), .A(n7685), .ZN(P1_U3289) );
  XNOR2_X1 U9520 ( .A(n8364), .B(n10315), .ZN(n7793) );
  XNOR2_X1 U9521 ( .A(n7793), .B(n7930), .ZN(n7689) );
  AOI21_X1 U9522 ( .B1(n7690), .B2(n7689), .A(n7797), .ZN(n7698) );
  INV_X1 U9523 ( .A(n7691), .ZN(n7904) );
  NAND2_X1 U9524 ( .A1(n8568), .A2(n10315), .ZN(n7695) );
  INV_X1 U9525 ( .A(n7692), .ZN(n7693) );
  AOI21_X1 U9526 ( .B1(n8580), .B2(n8608), .A(n7693), .ZN(n7694) );
  OAI211_X1 U9527 ( .C1(n7894), .C2(n8577), .A(n7695), .B(n7694), .ZN(n7696)
         );
  AOI21_X1 U9528 ( .B1(n7904), .B2(n8594), .A(n7696), .ZN(n7697) );
  OAI21_X1 U9529 ( .B1(n7698), .B2(n8570), .A(n7697), .ZN(P2_U3167) );
  NOR2_X1 U9530 ( .A1(n9452), .A2(n7699), .ZN(n7702) );
  INV_X1 U9531 ( .A(n7700), .ZN(n7701) );
  AOI21_X1 U9532 ( .B1(n7703), .B2(n7702), .A(n7701), .ZN(n7727) );
  XNOR2_X1 U9533 ( .A(n9452), .B(n7704), .ZN(n7729) );
  INV_X1 U9534 ( .A(n9871), .ZN(n9759) );
  NAND2_X1 U9535 ( .A1(n7729), .A2(n9759), .ZN(n7712) );
  INV_X1 U9536 ( .A(n7705), .ZN(n7706) );
  OAI211_X1 U9537 ( .C1(n7811), .C2(n7667), .A(n7706), .B(n10002), .ZN(n7725)
         );
  INV_X1 U9538 ( .A(n7725), .ZN(n7710) );
  AOI22_X1 U9539 ( .A1(n9936), .A2(n9591), .B1(n9898), .B2(n9593), .ZN(n7708)
         );
  AOI22_X1 U9540 ( .A1(n9933), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7815), .B2(
        n9932), .ZN(n7707) );
  OAI211_X1 U9541 ( .C1(n7811), .C2(n9926), .A(n7708), .B(n7707), .ZN(n7709)
         );
  AOI21_X1 U9542 ( .B1(n7710), .B2(n9921), .A(n7709), .ZN(n7711) );
  OAI211_X1 U9543 ( .C1(n7727), .C2(n9909), .A(n7712), .B(n7711), .ZN(P1_U3287) );
  OAI21_X1 U9544 ( .B1(n7715), .B2(n5814), .A(n7714), .ZN(n10300) );
  INV_X1 U9545 ( .A(n8941), .ZN(n7723) );
  OAI22_X1 U9546 ( .A1(n8744), .A2(n10297), .B1(n7716), .B2(n8912), .ZN(n7722)
         );
  XNOR2_X1 U9547 ( .A(n6250), .B(n7717), .ZN(n7718) );
  NAND2_X1 U9548 ( .A1(n7718), .A2(n10289), .ZN(n7720) );
  AOI22_X1 U9549 ( .A1(n10284), .A2(n10287), .B1(n6109), .B2(n10286), .ZN(
        n7719) );
  NAND2_X1 U9550 ( .A1(n7720), .A2(n7719), .ZN(n10298) );
  MUX2_X1 U9551 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10298), .S(n10282), .Z(n7721) );
  AOI211_X1 U9552 ( .C1(n10300), .C2(n7723), .A(n7722), .B(n7721), .ZN(n7724)
         );
  INV_X1 U9553 ( .A(n7724), .ZN(P2_U3232) );
  AOI22_X1 U9554 ( .A1(n10053), .A2(n9593), .B1(n9591), .B2(n10212), .ZN(n7726) );
  OAI211_X1 U9555 ( .C1(n7727), .C2(n10211), .A(n7726), .B(n7725), .ZN(n7728)
         );
  AOI21_X1 U9556 ( .B1(n9988), .B2(n7729), .A(n7728), .ZN(n7735) );
  AOI22_X1 U9557 ( .A1(n10063), .A2(n7730), .B1(n4409), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7731) );
  OAI21_X1 U9558 ( .B1(n7735), .B2(n4409), .A(n7731), .ZN(P1_U3528) );
  INV_X1 U9559 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7732) );
  OAI22_X1 U9560 ( .A1(n10090), .A2(n7811), .B1(n10243), .B2(n7732), .ZN(n7733) );
  INV_X1 U9561 ( .A(n7733), .ZN(n7734) );
  OAI21_X1 U9562 ( .B1(n7735), .B2(n7144), .A(n7734), .ZN(P1_U3471) );
  OAI21_X1 U9563 ( .B1(n9453), .B2(n7737), .A(n7736), .ZN(n10228) );
  AOI211_X1 U9564 ( .C1(n7740), .C2(n7739), .A(n9920), .B(n7738), .ZN(n10223)
         );
  AOI22_X1 U9565 ( .A1(n10223), .A2(n9921), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9932), .ZN(n7741) );
  OAI21_X1 U9566 ( .B1(n10225), .B2(n9926), .A(n7741), .ZN(n7748) );
  INV_X1 U9567 ( .A(n9453), .ZN(n7742) );
  XNOR2_X1 U9568 ( .A(n7743), .B(n7742), .ZN(n7744) );
  NAND2_X1 U9569 ( .A1(n7744), .A2(n9988), .ZN(n7746) );
  AOI22_X1 U9570 ( .A1(n10212), .A2(n9595), .B1(n6400), .B2(n10053), .ZN(n7745) );
  NAND2_X1 U9571 ( .A1(n7746), .A2(n7745), .ZN(n10227) );
  MUX2_X1 U9572 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10227), .S(n9893), .Z(n7747)
         );
  AOI211_X1 U9573 ( .C1(n9928), .C2(n10228), .A(n7748), .B(n7747), .ZN(n7749)
         );
  INV_X1 U9574 ( .A(n7749), .ZN(P1_U3291) );
  INV_X1 U9575 ( .A(n7750), .ZN(n7753) );
  OAI222_X1 U9576 ( .A1(n9121), .A2(n7752), .B1(n9123), .B2(n7753), .C1(
        P2_U3151), .C2(n4428), .ZN(P2_U3276) );
  AOI21_X1 U9577 ( .B1(n7757), .B2(n7756), .A(n7755), .ZN(n7767) );
  OAI21_X1 U9578 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7758), .A(n7965), .ZN(
        n7765) );
  OAI21_X1 U9579 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7759), .A(n7959), .ZN(
        n7760) );
  NAND2_X1 U9580 ( .A1(n7760), .A2(n8730), .ZN(n7762) );
  NOR2_X1 U9581 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5367), .ZN(n8019) );
  AOI21_X1 U9582 ( .B1(n8699), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8019), .ZN(
        n7761) );
  OAI211_X1 U9583 ( .C1(n8717), .C2(n7763), .A(n7762), .B(n7761), .ZN(n7764)
         );
  AOI21_X1 U9584 ( .B1(n8639), .B2(n7765), .A(n7764), .ZN(n7766) );
  OAI21_X1 U9585 ( .B1(n7767), .B2(n8722), .A(n7766), .ZN(P2_U3189) );
  XNOR2_X1 U9586 ( .A(n7858), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7771) );
  AOI211_X1 U9587 ( .C1(n7771), .C2(n7770), .A(n10164), .B(n7769), .ZN(n7780)
         );
  XNOR2_X1 U9588 ( .A(n7858), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7775) );
  OAI21_X1 U9589 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n7773), .A(n7772), .ZN(
        n7774) );
  NOR2_X1 U9590 ( .A1(n7774), .A2(n7775), .ZN(n7857) );
  AOI211_X1 U9591 ( .C1(n7775), .C2(n7774), .A(n10152), .B(n7857), .ZN(n7779)
         );
  INV_X1 U9592 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U9593 ( .A1(n10183), .A2(n7858), .ZN(n7776) );
  NAND2_X1 U9594 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9151) );
  OAI211_X1 U9595 ( .C1(n7777), .C2(n10207), .A(n7776), .B(n9151), .ZN(n7778)
         );
  OR3_X1 U9596 ( .A1(n7780), .A2(n7779), .A3(n7778), .ZN(P1_U3253) );
  AOI22_X1 U9597 ( .A1(n7781), .A2(n9272), .B1(n9593), .B2(n9326), .ZN(n7783)
         );
  OAI211_X1 U9598 ( .C1(n7784), .C2(n9324), .A(n7783), .B(n7782), .ZN(n7790)
         );
  INV_X1 U9599 ( .A(n7785), .ZN(n7786) );
  AOI211_X1 U9600 ( .C1(n7791), .C2(n9338), .A(n7790), .B(n7789), .ZN(n7792)
         );
  INV_X1 U9601 ( .A(n7792), .ZN(P1_U3230) );
  INV_X1 U9602 ( .A(n7793), .ZN(n7794) );
  NOR2_X1 U9603 ( .A1(n7794), .A2(n10275), .ZN(n7796) );
  XNOR2_X1 U9604 ( .A(n8364), .B(n7937), .ZN(n8012) );
  XNOR2_X1 U9605 ( .A(n8012), .B(n10257), .ZN(n7795) );
  INV_X1 U9606 ( .A(n8013), .ZN(n7799) );
  OAI21_X1 U9607 ( .B1(n7797), .B2(n7796), .A(n7795), .ZN(n7798) );
  NAND3_X1 U9608 ( .A1(n7799), .A2(n8587), .A3(n7798), .ZN(n7804) );
  INV_X1 U9609 ( .A(n8577), .ZN(n8590) );
  NAND2_X1 U9610 ( .A1(n8590), .A2(n10275), .ZN(n7801) );
  OAI211_X1 U9611 ( .C1(n8171), .C2(n8592), .A(n7801), .B(n7800), .ZN(n7802)
         );
  AOI21_X1 U9612 ( .B1(n7937), .B2(n8568), .A(n7802), .ZN(n7803) );
  OAI211_X1 U9613 ( .C1(n7935), .C2(n8566), .A(n7804), .B(n7803), .ZN(P2_U3179) );
  INV_X1 U9614 ( .A(n7806), .ZN(n7808) );
  NAND2_X1 U9615 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  XNOR2_X1 U9616 ( .A(n7805), .B(n7809), .ZN(n7818) );
  INV_X1 U9617 ( .A(n7810), .ZN(n7814) );
  OAI22_X1 U9618 ( .A1(n7812), .A2(n9324), .B1(n9335), .B2(n7811), .ZN(n7813)
         );
  AOI211_X1 U9619 ( .C1(n9326), .C2(n9591), .A(n7814), .B(n7813), .ZN(n7817)
         );
  NAND2_X1 U9620 ( .A1(n9338), .A2(n7815), .ZN(n7816) );
  OAI211_X1 U9621 ( .C1(n7818), .C2(n9340), .A(n7817), .B(n7816), .ZN(P1_U3239) );
  NAND2_X1 U9622 ( .A1(n9596), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7819) );
  OAI21_X1 U9623 ( .B1(n9671), .B2(n9596), .A(n7819), .ZN(P1_U3583) );
  OAI21_X1 U9624 ( .B1(n7704), .B2(n7820), .A(n9359), .ZN(n7821) );
  NAND2_X1 U9625 ( .A1(n7821), .A2(n7824), .ZN(n7997) );
  OAI21_X1 U9626 ( .B1(n7824), .B2(n7821), .A(n7997), .ZN(n7822) );
  AND2_X1 U9627 ( .A1(n7822), .A2(n9988), .ZN(n7910) );
  INV_X1 U9628 ( .A(n7910), .ZN(n7834) );
  NAND2_X1 U9629 ( .A1(n7700), .A2(n7823), .ZN(n7826) );
  INV_X1 U9630 ( .A(n7824), .ZN(n7825) );
  NAND2_X1 U9631 ( .A1(n7826), .A2(n7825), .ZN(n7882) );
  OAI21_X1 U9632 ( .B1(n7826), .B2(n7825), .A(n7882), .ZN(n7912) );
  AOI22_X1 U9633 ( .A1(n9936), .A2(n8007), .B1(n9898), .B2(n9592), .ZN(n7829)
         );
  INV_X1 U9634 ( .A(n7827), .ZN(n7874) );
  AOI22_X1 U9635 ( .A1(n9933), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7874), .B2(
        n9932), .ZN(n7828) );
  OAI211_X1 U9636 ( .C1(n7914), .C2(n9926), .A(n7829), .B(n7828), .ZN(n7832)
         );
  OAI211_X1 U9637 ( .C1(n7705), .C2(n7914), .A(n10002), .B(n7830), .ZN(n7909)
         );
  NOR2_X1 U9638 ( .A1(n7909), .A2(n9863), .ZN(n7831) );
  AOI211_X1 U9639 ( .C1(n7912), .C2(n9928), .A(n7832), .B(n7831), .ZN(n7833)
         );
  OAI21_X1 U9640 ( .B1(n7834), .B2(n9933), .A(n7833), .ZN(P1_U3286) );
  INV_X1 U9641 ( .A(n7835), .ZN(n7839) );
  OAI222_X1 U9642 ( .A1(n7837), .A2(P1_U3086), .B1(n8337), .B2(n7839), .C1(
        n7836), .C2(n10116), .ZN(P1_U3335) );
  OAI222_X1 U9643 ( .A1(n9121), .A2(n7840), .B1(n9123), .B2(n7839), .C1(n7838), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  NAND2_X1 U9644 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  XOR2_X1 U9645 ( .A(n7844), .B(n7843), .Z(n7845) );
  NAND2_X1 U9646 ( .A1(n7845), .A2(n9320), .ZN(n7851) );
  INV_X1 U9647 ( .A(n7846), .ZN(n7849) );
  OAI22_X1 U9648 ( .A1(n7847), .A2(n9324), .B1(n9335), .B2(n5051), .ZN(n7848)
         );
  AOI211_X1 U9649 ( .C1(n9326), .C2(n9592), .A(n7849), .B(n7848), .ZN(n7850)
         );
  OAI211_X1 U9650 ( .C1(n9303), .C2(n7852), .A(n7851), .B(n7850), .ZN(P1_U3227) );
  NAND2_X1 U9651 ( .A1(n7858), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7853) );
  XNOR2_X1 U9652 ( .A(n8097), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n7855) );
  AOI211_X1 U9653 ( .C1(n7856), .C2(n7855), .A(n10164), .B(n8088), .ZN(n7865)
         );
  XNOR2_X1 U9654 ( .A(n8097), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7859) );
  AOI211_X1 U9655 ( .C1(n7860), .C2(n7859), .A(n10152), .B(n8096), .ZN(n7864)
         );
  NAND2_X1 U9656 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9301) );
  NAND2_X1 U9657 ( .A1(n10169), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n7861) );
  OAI211_X1 U9658 ( .C1(n10202), .C2(n7862), .A(n9301), .B(n7861), .ZN(n7863)
         );
  OR3_X1 U9659 ( .A1(n7865), .A2(n7864), .A3(n7863), .ZN(P1_U3254) );
  XOR2_X1 U9660 ( .A(n7868), .B(n7867), .Z(n7869) );
  XNOR2_X1 U9661 ( .A(n7866), .B(n7869), .ZN(n7876) );
  AOI22_X1 U9662 ( .A1(n7917), .A2(n9272), .B1(n8007), .B2(n9326), .ZN(n7871)
         );
  OAI211_X1 U9663 ( .C1(n7872), .C2(n9324), .A(n7871), .B(n7870), .ZN(n7873)
         );
  AOI21_X1 U9664 ( .B1(n7874), .B2(n9338), .A(n7873), .ZN(n7875) );
  OAI21_X1 U9665 ( .B1(n7876), .B2(n9340), .A(n7875), .ZN(P1_U3213) );
  NAND2_X1 U9666 ( .A1(n7997), .A2(n9360), .ZN(n7877) );
  XNOR2_X1 U9667 ( .A(n7877), .B(n7879), .ZN(n7878) );
  NOR2_X1 U9668 ( .A1(n7878), .A2(n10210), .ZN(n8146) );
  INV_X1 U9669 ( .A(n8146), .ZN(n7892) );
  INV_X1 U9670 ( .A(n7879), .ZN(n7881) );
  NAND3_X1 U9671 ( .A1(n7882), .A2(n7881), .A3(n7880), .ZN(n7884) );
  NAND2_X1 U9672 ( .A1(n7884), .A2(n7883), .ZN(n8148) );
  OAI22_X1 U9673 ( .A1(n9893), .A2(n7885), .B1(n9176), .B2(n9891), .ZN(n7886)
         );
  AOI21_X1 U9674 ( .B1(n9898), .B2(n9591), .A(n7886), .ZN(n7888) );
  NAND2_X1 U9675 ( .A1(n9930), .A2(n9183), .ZN(n7887) );
  OAI211_X1 U9676 ( .C1(n9152), .C2(n9894), .A(n7888), .B(n7887), .ZN(n7890)
         );
  INV_X1 U9677 ( .A(n9183), .ZN(n8151) );
  OAI211_X1 U9678 ( .C1(n7075), .C2(n8151), .A(n10002), .B(n8002), .ZN(n8145)
         );
  NOR2_X1 U9679 ( .A1(n8145), .A2(n9863), .ZN(n7889) );
  AOI211_X1 U9680 ( .C1(n8148), .C2(n9928), .A(n7890), .B(n7889), .ZN(n7891)
         );
  OAI21_X1 U9681 ( .B1(n7892), .B2(n9933), .A(n7891), .ZN(P1_U3285) );
  XNOR2_X1 U9682 ( .A(n7893), .B(n7897), .ZN(n10318) );
  INV_X1 U9683 ( .A(n10318), .ZN(n7907) );
  INV_X1 U9684 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7903) );
  OAI22_X1 U9685 ( .A1(n7894), .A2(n10256), .B1(n10257), .B2(n10254), .ZN(
        n7901) );
  INV_X1 U9686 ( .A(n7895), .ZN(n7896) );
  NOR2_X1 U9687 ( .A1(n7898), .A2(n7896), .ZN(n7925) );
  AND2_X1 U9688 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  AOI211_X1 U9689 ( .C1(n7925), .C2(n7923), .A(n8853), .B(n7899), .ZN(n7900)
         );
  AOI211_X1 U9690 ( .C1(n7902), .C2(n10318), .A(n7901), .B(n7900), .ZN(n10320)
         );
  MUX2_X1 U9691 ( .A(n7903), .B(n10320), .S(n10282), .Z(n7906) );
  AOI22_X1 U9692 ( .A1(n10292), .A2(n10315), .B1(n10293), .B2(n7904), .ZN(
        n7905) );
  OAI211_X1 U9693 ( .C1(n7907), .C2(n10267), .A(n7906), .B(n7905), .ZN(
        P2_U3228) );
  AOI22_X1 U9694 ( .A1(n8007), .A2(n10212), .B1(n10053), .B2(n9592), .ZN(n7908) );
  NAND2_X1 U9695 ( .A1(n7909), .A2(n7908), .ZN(n7911) );
  AOI211_X1 U9696 ( .C1(n10241), .C2(n7912), .A(n7911), .B(n7910), .ZN(n7919)
         );
  OAI22_X1 U9697 ( .A1(n10090), .A2(n7914), .B1(n10243), .B2(n7913), .ZN(n7915) );
  INV_X1 U9698 ( .A(n7915), .ZN(n7916) );
  OAI21_X1 U9699 ( .B1(n7919), .B2(n7144), .A(n7916), .ZN(P1_U3474) );
  AOI22_X1 U9700 ( .A1(n10063), .A2(n7917), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n4409), .ZN(n7918) );
  OAI21_X1 U9701 ( .B1(n7919), .B2(n4409), .A(n7918), .ZN(P1_U3529) );
  NAND2_X1 U9702 ( .A1(n7920), .A2(n7921), .ZN(n7922) );
  XOR2_X1 U9703 ( .A(n7926), .B(n7922), .Z(n10322) );
  INV_X1 U9704 ( .A(n7923), .ZN(n7924) );
  NOR2_X1 U9705 ( .A1(n7925), .A2(n7924), .ZN(n7927) );
  AOI21_X1 U9706 ( .B1(n7927), .B2(n7926), .A(n8853), .ZN(n7933) );
  INV_X1 U9707 ( .A(n7927), .ZN(n7929) );
  OAI211_X1 U9708 ( .C1(n10257), .C2(n10324), .A(n7929), .B(n7928), .ZN(n7932)
         );
  OAI22_X1 U9709 ( .A1(n7930), .A2(n10256), .B1(n8171), .B2(n10254), .ZN(n7931) );
  AOI21_X1 U9710 ( .B1(n7933), .B2(n7932), .A(n7931), .ZN(n10323) );
  MUX2_X1 U9711 ( .A(n7934), .B(n10323), .S(n10282), .Z(n7939) );
  INV_X1 U9712 ( .A(n7935), .ZN(n7936) );
  AOI22_X1 U9713 ( .A1(n10292), .A2(n7937), .B1(n10293), .B2(n7936), .ZN(n7938) );
  OAI211_X1 U9714 ( .C1(n10322), .C2(n8941), .A(n7939), .B(n7938), .ZN(
        P2_U3227) );
  NAND2_X1 U9715 ( .A1(n10259), .A2(n10258), .ZN(n10261) );
  NAND2_X1 U9716 ( .A1(n10261), .A2(n7940), .ZN(n7941) );
  XOR2_X1 U9717 ( .A(n7944), .B(n7941), .Z(n8187) );
  INV_X1 U9718 ( .A(n8187), .ZN(n8103) );
  NAND2_X1 U9719 ( .A1(n7943), .A2(n7942), .ZN(n7945) );
  NAND2_X1 U9720 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U9721 ( .A1(n8136), .A2(n7946), .ZN(n7947) );
  NAND2_X1 U9722 ( .A1(n7947), .A2(n10289), .ZN(n7949) );
  AOI22_X1 U9723 ( .A1(n8607), .A2(n10286), .B1(n10284), .B2(n8605), .ZN(n7948) );
  NAND2_X1 U9724 ( .A1(n7949), .A2(n7948), .ZN(n8184) );
  INV_X1 U9725 ( .A(n8163), .ZN(n8183) );
  OAI22_X1 U9726 ( .A1(n9101), .A2(n8183), .B1(n7950), .B2(n10336), .ZN(n7951)
         );
  AOI21_X1 U9727 ( .B1(n8184), .B2(n10336), .A(n7951), .ZN(n7952) );
  OAI21_X1 U9728 ( .B1(n8103), .B2(n9096), .A(n7952), .ZN(P2_U3414) );
  XOR2_X1 U9729 ( .A(n7954), .B(n7953), .Z(n7975) );
  INV_X1 U9730 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U9731 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8170) );
  OAI21_X1 U9732 ( .B1(n8721), .B2(n7955), .A(n8170), .ZN(n7963) );
  INV_X1 U9733 ( .A(n7956), .ZN(n7958) );
  NAND3_X1 U9734 ( .A1(n7959), .A2(n7958), .A3(n7957), .ZN(n7960) );
  AOI21_X1 U9735 ( .B1(n7961), .B2(n7960), .A(n8655), .ZN(n7962) );
  AOI211_X1 U9736 ( .C1(n8632), .C2(n7964), .A(n7963), .B(n7962), .ZN(n7974)
         );
  INV_X1 U9737 ( .A(n7965), .ZN(n7969) );
  INV_X1 U9738 ( .A(n7966), .ZN(n7968) );
  NOR3_X1 U9739 ( .A1(n7969), .A2(n7968), .A3(n7967), .ZN(n7972) );
  INV_X1 U9740 ( .A(n7970), .ZN(n7971) );
  OAI21_X1 U9741 ( .B1(n7972), .B2(n7971), .A(n8639), .ZN(n7973) );
  OAI211_X1 U9742 ( .C1(n7975), .C2(n8722), .A(n7974), .B(n7973), .ZN(P2_U3190) );
  INV_X1 U9743 ( .A(n7976), .ZN(n7977) );
  AOI21_X1 U9744 ( .B1(n7987), .B2(n7978), .A(n7977), .ZN(n8109) );
  OAI22_X1 U9745 ( .A1(n9893), .A2(n7979), .B1(n9155), .B2(n9891), .ZN(n7980)
         );
  AOI21_X1 U9746 ( .B1(n9898), .B2(n9178), .A(n7980), .ZN(n7981) );
  OAI21_X1 U9747 ( .B1(n9203), .B2(n9894), .A(n7981), .ZN(n7984) );
  NOR2_X1 U9748 ( .A1(n8001), .A2(n4411), .ZN(n7982) );
  OR3_X1 U9749 ( .A1(n8033), .A2(n7982), .A3(n9920), .ZN(n8107) );
  NOR2_X1 U9750 ( .A1(n8107), .A2(n9863), .ZN(n7983) );
  AOI211_X1 U9751 ( .C1(n9930), .C2(n9157), .A(n7984), .B(n7983), .ZN(n7990)
         );
  NAND2_X1 U9752 ( .A1(n7985), .A2(n7986), .ZN(n7988) );
  NAND2_X1 U9753 ( .A1(n7988), .A2(n7987), .ZN(n8030) );
  OAI21_X1 U9754 ( .B1(n7988), .B2(n7987), .A(n8030), .ZN(n8111) );
  NAND2_X1 U9755 ( .A1(n8111), .A2(n9928), .ZN(n7989) );
  OAI211_X1 U9756 ( .C1(n8109), .C2(n9871), .A(n7990), .B(n7989), .ZN(P1_U3283) );
  INV_X1 U9757 ( .A(n7991), .ZN(n7994) );
  OAI222_X1 U9758 ( .A1(P2_U3151), .A2(n7385), .B1(n9123), .B2(n7994), .C1(
        n7992), .C2(n9121), .ZN(P2_U3274) );
  INV_X1 U9759 ( .A(n7995), .ZN(n7996) );
  AOI21_X1 U9760 ( .B1(n7997), .B2(n9353), .A(n7996), .ZN(n7998) );
  XOR2_X1 U9761 ( .A(n7999), .B(n7998), .Z(n8068) );
  INV_X1 U9762 ( .A(n8068), .ZN(n8011) );
  OAI21_X1 U9763 ( .B1(n8000), .B2(n7999), .A(n7985), .ZN(n8064) );
  AOI21_X1 U9764 ( .B1(n10212), .B2(n9590), .A(n8003), .ZN(n8066) );
  OAI22_X1 U9765 ( .A1(n9893), .A2(n8004), .B1(n9258), .B2(n9891), .ZN(n8006)
         );
  INV_X1 U9766 ( .A(n8070), .ZN(n9263) );
  NOR2_X1 U9767 ( .A1(n9263), .A2(n9926), .ZN(n8005) );
  AOI211_X1 U9768 ( .C1(n9898), .C2(n8007), .A(n8006), .B(n8005), .ZN(n8008)
         );
  OAI21_X1 U9769 ( .B1(n8066), .B2(n9863), .A(n8008), .ZN(n8009) );
  AOI21_X1 U9770 ( .B1(n9928), .B2(n8064), .A(n8009), .ZN(n8010) );
  OAI21_X1 U9771 ( .B1(n8011), .B2(n9871), .A(n8010), .ZN(P1_U3284) );
  INV_X1 U9772 ( .A(n8012), .ZN(n8014) );
  XNOR2_X1 U9773 ( .A(n10331), .B(n8364), .ZN(n8015) );
  NOR2_X1 U9774 ( .A1(n8015), .A2(n8607), .ZN(n8164) );
  AOI21_X1 U9775 ( .B1(n8607), .B2(n8015), .A(n8164), .ZN(n8016) );
  OAI21_X1 U9776 ( .B1(n8017), .B2(n8016), .A(n8166), .ZN(n8018) );
  NAND2_X1 U9777 ( .A1(n8018), .A2(n8587), .ZN(n8023) );
  AOI21_X1 U9778 ( .B1(n8580), .B2(n8606), .A(n8019), .ZN(n8020) );
  OAI21_X1 U9779 ( .B1(n10257), .B2(n8577), .A(n8020), .ZN(n8021) );
  AOI21_X1 U9780 ( .B1(n10268), .B2(n8568), .A(n8021), .ZN(n8022) );
  OAI211_X1 U9781 ( .C1(n10266), .C2(n8566), .A(n8023), .B(n8022), .ZN(
        P2_U3153) );
  NAND2_X1 U9782 ( .A1(n7976), .A2(n8024), .ZN(n8027) );
  INV_X1 U9783 ( .A(n8025), .ZN(n8026) );
  AOI211_X1 U9784 ( .C1(n9461), .C2(n8027), .A(n10210), .B(n8026), .ZN(n8157)
         );
  INV_X1 U9785 ( .A(n8157), .ZN(n8041) );
  INV_X1 U9786 ( .A(n9461), .ZN(n8029) );
  NAND3_X1 U9787 ( .A1(n8030), .A2(n8029), .A3(n8028), .ZN(n8032) );
  NAND2_X1 U9788 ( .A1(n8032), .A2(n8031), .ZN(n8159) );
  OAI211_X1 U9789 ( .C1(n8033), .C2(n9308), .A(n10002), .B(n8120), .ZN(n8156)
         );
  OAI22_X1 U9790 ( .A1(n9893), .A2(n8034), .B1(n9302), .B2(n9891), .ZN(n8035)
         );
  AOI21_X1 U9791 ( .B1(n9898), .B2(n9590), .A(n8035), .ZN(n8036) );
  OAI21_X1 U9792 ( .B1(n9911), .B2(n9894), .A(n8036), .ZN(n8037) );
  AOI21_X1 U9793 ( .B1(n9930), .B2(n7027), .A(n8037), .ZN(n8038) );
  OAI21_X1 U9794 ( .B1(n8156), .B2(n9863), .A(n8038), .ZN(n8039) );
  AOI21_X1 U9795 ( .B1(n9928), .B2(n8159), .A(n8039), .ZN(n8040) );
  OAI21_X1 U9796 ( .B1(n8041), .B2(n9933), .A(n8040), .ZN(P1_U3282) );
  INV_X1 U9797 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10356) );
  INV_X1 U9798 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U9799 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8042) );
  AOI21_X1 U9800 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n8042), .ZN(n10359) );
  NOR2_X1 U9801 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8043) );
  AOI21_X1 U9802 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8043), .ZN(n10362) );
  NOR2_X1 U9803 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8044) );
  AOI21_X1 U9804 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8044), .ZN(n10365) );
  NOR2_X1 U9805 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8045) );
  AOI21_X1 U9806 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8045), .ZN(n10368) );
  NOR2_X1 U9807 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8046) );
  AOI21_X1 U9808 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8046), .ZN(n10371) );
  NOR2_X1 U9809 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8047) );
  AOI21_X1 U9810 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8047), .ZN(n10374) );
  NOR2_X1 U9811 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8048) );
  AOI21_X1 U9812 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8048), .ZN(n10377) );
  NOR2_X1 U9813 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8049) );
  AOI21_X1 U9814 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8049), .ZN(n10380) );
  NOR2_X1 U9815 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8050) );
  AOI21_X1 U9816 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n8050), .ZN(n10683) );
  NOR2_X1 U9817 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8051) );
  AOI21_X1 U9818 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n8051), .ZN(n10689) );
  NOR2_X1 U9819 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8052) );
  AOI21_X1 U9820 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n8052), .ZN(n10686) );
  NOR2_X1 U9821 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8053) );
  AOI21_X1 U9822 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n8053), .ZN(n10677) );
  NOR2_X1 U9823 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8054) );
  AOI21_X1 U9824 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n8054), .ZN(n10680) );
  AND2_X1 U9825 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n8055) );
  NOR2_X1 U9826 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n8055), .ZN(n10348) );
  INV_X1 U9827 ( .A(n10348), .ZN(n10349) );
  INV_X1 U9828 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10351) );
  NAND3_X1 U9829 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U9830 ( .A1(n10351), .A2(n10350), .ZN(n10347) );
  NAND2_X1 U9831 ( .A1(n10349), .A2(n10347), .ZN(n10692) );
  NAND2_X1 U9832 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8056) );
  OAI21_X1 U9833 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n8056), .ZN(n10691) );
  NOR2_X1 U9834 ( .A1(n10692), .A2(n10691), .ZN(n10690) );
  AOI21_X1 U9835 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10690), .ZN(n10695) );
  NAND2_X1 U9836 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8057) );
  OAI21_X1 U9837 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n8057), .ZN(n10694) );
  NOR2_X1 U9838 ( .A1(n10695), .A2(n10694), .ZN(n10693) );
  AOI21_X1 U9839 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10693), .ZN(n10698) );
  NOR2_X1 U9840 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8058) );
  AOI21_X1 U9841 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n8058), .ZN(n10697) );
  NAND2_X1 U9842 ( .A1(n10698), .A2(n10697), .ZN(n10696) );
  OAI21_X1 U9843 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10696), .ZN(n10679) );
  NAND2_X1 U9844 ( .A1(n10680), .A2(n10679), .ZN(n10678) );
  OAI21_X1 U9845 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10678), .ZN(n10676) );
  NAND2_X1 U9846 ( .A1(n10677), .A2(n10676), .ZN(n10675) );
  OAI21_X1 U9847 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10675), .ZN(n10685) );
  NAND2_X1 U9848 ( .A1(n10686), .A2(n10685), .ZN(n10684) );
  OAI21_X1 U9849 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10684), .ZN(n10688) );
  NAND2_X1 U9850 ( .A1(n10689), .A2(n10688), .ZN(n10687) );
  OAI21_X1 U9851 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10687), .ZN(n10682) );
  NAND2_X1 U9852 ( .A1(n10683), .A2(n10682), .ZN(n10681) );
  OAI21_X1 U9853 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10681), .ZN(n10379) );
  NAND2_X1 U9854 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  OAI21_X1 U9855 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10378), .ZN(n10376) );
  NAND2_X1 U9856 ( .A1(n10377), .A2(n10376), .ZN(n10375) );
  OAI21_X1 U9857 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10375), .ZN(n10373) );
  NAND2_X1 U9858 ( .A1(n10374), .A2(n10373), .ZN(n10372) );
  OAI21_X1 U9859 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10372), .ZN(n10370) );
  NAND2_X1 U9860 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  OAI21_X1 U9861 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10369), .ZN(n10367) );
  NAND2_X1 U9862 ( .A1(n10368), .A2(n10367), .ZN(n10366) );
  OAI21_X1 U9863 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10366), .ZN(n10364) );
  NAND2_X1 U9864 ( .A1(n10365), .A2(n10364), .ZN(n10363) );
  OAI21_X1 U9865 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10363), .ZN(n10361) );
  NAND2_X1 U9866 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  OAI21_X1 U9867 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10360), .ZN(n10358) );
  NAND2_X1 U9868 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  OAI21_X1 U9869 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10357), .ZN(n8059) );
  OR2_X1 U9870 ( .A1(n10206), .A2(n8059), .ZN(n10355) );
  NAND2_X1 U9871 ( .A1(n10356), .A2(n10355), .ZN(n10352) );
  NAND2_X1 U9872 ( .A1(n10206), .A2(n8059), .ZN(n10354) );
  NAND2_X1 U9873 ( .A1(n10352), .A2(n10354), .ZN(n8063) );
  NOR2_X1 U9874 ( .A1(n8060), .A2(n8061), .ZN(n8062) );
  XNOR2_X1 U9875 ( .A(n8063), .B(n8062), .ZN(ADD_1068_U4) );
  NAND2_X1 U9876 ( .A1(n8064), .A2(n10241), .ZN(n8065) );
  OAI211_X1 U9877 ( .C1(n9257), .C2(n10038), .A(n8066), .B(n8065), .ZN(n8067)
         );
  AOI21_X1 U9878 ( .B1(n8068), .B2(n9988), .A(n8067), .ZN(n8072) );
  AOI22_X1 U9879 ( .A1(n7093), .A2(n8070), .B1(P1_REG0_REG_9__SCAN_IN), .B2(
        n7144), .ZN(n8069) );
  OAI21_X1 U9880 ( .B1(n8072), .B2(n7144), .A(n8069), .ZN(P1_U3480) );
  AOI22_X1 U9881 ( .A1(n10063), .A2(n8070), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n4409), .ZN(n8071) );
  OAI21_X1 U9882 ( .B1(n8072), .B2(n4409), .A(n8071), .ZN(P1_U3531) );
  AOI21_X1 U9883 ( .B1(n10577), .B2(n8073), .A(n4432), .ZN(n8086) );
  XNOR2_X1 U9884 ( .A(n8075), .B(n8074), .ZN(n8076) );
  NAND2_X1 U9885 ( .A1(n8076), .A2(n8704), .ZN(n8085) );
  INV_X1 U9886 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8078) );
  AND2_X1 U9887 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8217) );
  INV_X1 U9888 ( .A(n8217), .ZN(n8077) );
  OAI21_X1 U9889 ( .B1(n8721), .B2(n8078), .A(n8077), .ZN(n8082) );
  NAND2_X1 U9890 ( .A1(n8079), .A2(n8231), .ZN(n8080) );
  AOI21_X1 U9891 ( .B1(n8195), .B2(n8080), .A(n8734), .ZN(n8081) );
  AOI211_X1 U9892 ( .C1(n8632), .C2(n8083), .A(n8082), .B(n8081), .ZN(n8084)
         );
  OAI211_X1 U9893 ( .C1(n8086), .C2(n8655), .A(n8085), .B(n8084), .ZN(P2_U3191) );
  XOR2_X1 U9894 ( .A(n9620), .B(P1_REG2_REG_12__SCAN_IN), .Z(n8090) );
  OAI21_X1 U9895 ( .B1(n8090), .B2(n8089), .A(n9610), .ZN(n8094) );
  NAND2_X1 U9896 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9201) );
  NAND2_X1 U9897 ( .A1(n10169), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n8091) );
  OAI211_X1 U9898 ( .C1(n10202), .C2(n8092), .A(n9201), .B(n8091), .ZN(n8093)
         );
  AOI21_X1 U9899 ( .B1(n8094), .B2(n10193), .A(n8093), .ZN(n8102) );
  XNOR2_X1 U9900 ( .A(n9620), .B(n8095), .ZN(n8099) );
  OAI21_X1 U9901 ( .B1(n8099), .B2(n8098), .A(n9619), .ZN(n8100) );
  NAND2_X1 U9902 ( .A1(n8100), .A2(n10198), .ZN(n8101) );
  NAND2_X1 U9903 ( .A1(n8102), .A2(n8101), .ZN(P1_U3255) );
  NAND2_X1 U9904 ( .A1(n10672), .A2(n10327), .ZN(n9010) );
  OAI22_X1 U9905 ( .A1(n8103), .A2(n9010), .B1(n8183), .B2(n9018), .ZN(n8105)
         );
  MUX2_X1 U9906 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n8184), .S(n10672), .Z(n8104)
         );
  OR2_X1 U9907 ( .A1(n8105), .A2(n8104), .ZN(P2_U3467) );
  OAI22_X1 U9908 ( .A1(n9152), .A2(n10038), .B1(n9203), .B2(n10057), .ZN(n8106) );
  INV_X1 U9909 ( .A(n8106), .ZN(n8108) );
  OAI211_X1 U9910 ( .C1(n8109), .C2(n10210), .A(n8108), .B(n8107), .ZN(n8110)
         );
  AOI21_X1 U9911 ( .B1(n10241), .B2(n8111), .A(n8110), .ZN(n8114) );
  AOI22_X1 U9912 ( .A1(n10063), .A2(n9157), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n4409), .ZN(n8112) );
  OAI21_X1 U9913 ( .B1(n8114), .B2(n4409), .A(n8112), .ZN(P1_U3532) );
  AOI22_X1 U9914 ( .A1(n7093), .A2(n9157), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n7144), .ZN(n8113) );
  OAI21_X1 U9915 ( .B1(n8114), .B2(n7144), .A(n8113), .ZN(P1_U3483) );
  NAND2_X1 U9916 ( .A1(n8025), .A2(n9366), .ZN(n8117) );
  INV_X1 U9917 ( .A(n8115), .ZN(n8116) );
  AOI21_X1 U9918 ( .B1(n9460), .B2(n8117), .A(n8116), .ZN(n10059) );
  OAI21_X1 U9919 ( .B1(n8119), .B2(n9460), .A(n8118), .ZN(n10062) );
  AOI21_X1 U9920 ( .B1(n8120), .B2(n10095), .A(n9920), .ZN(n8121) );
  NAND2_X1 U9921 ( .A1(n8121), .A2(n4524), .ZN(n10056) );
  OAI22_X1 U9922 ( .A1(n9893), .A2(n8122), .B1(n9200), .B2(n9891), .ZN(n8123)
         );
  AOI21_X1 U9923 ( .B1(n9898), .B2(n10054), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9924 ( .B1(n10058), .B2(n9894), .A(n8124), .ZN(n8125) );
  AOI21_X1 U9925 ( .B1(n9930), .B2(n10095), .A(n8125), .ZN(n8126) );
  OAI21_X1 U9926 ( .B1(n10056), .B2(n9863), .A(n8126), .ZN(n8127) );
  AOI21_X1 U9927 ( .B1(n9928), .B2(n10062), .A(n8127), .ZN(n8128) );
  OAI21_X1 U9928 ( .B1(n10059), .B2(n9871), .A(n8128), .ZN(P1_U3281) );
  NAND2_X1 U9929 ( .A1(n10261), .A2(n8129), .ZN(n8131) );
  NAND2_X1 U9930 ( .A1(n8131), .A2(n8130), .ZN(n8133) );
  INV_X1 U9931 ( .A(n8132), .ZN(n8137) );
  NAND2_X1 U9932 ( .A1(n8133), .A2(n8137), .ZN(n8134) );
  NAND2_X1 U9933 ( .A1(n8234), .A2(n8134), .ZN(n8229) );
  AOI22_X1 U9934 ( .A1(n8606), .A2(n10286), .B1(n10284), .B2(n8604), .ZN(n8141) );
  NAND2_X1 U9935 ( .A1(n8136), .A2(n8135), .ZN(n8138) );
  XNOR2_X1 U9936 ( .A(n8138), .B(n8137), .ZN(n8139) );
  NAND2_X1 U9937 ( .A1(n8139), .A2(n10289), .ZN(n8140) );
  OAI211_X1 U9938 ( .C1(n8229), .C2(n10262), .A(n8141), .B(n8140), .ZN(n8223)
         );
  INV_X1 U9939 ( .A(n10317), .ZN(n10332) );
  INV_X1 U9940 ( .A(n8226), .ZN(n8222) );
  OAI22_X1 U9941 ( .A1(n8229), .A2(n10332), .B1(n8222), .B2(n10330), .ZN(n8142) );
  NOR2_X1 U9942 ( .A1(n8223), .A2(n8142), .ZN(n8230) );
  NAND2_X1 U9943 ( .A1(n10337), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8143) );
  OAI21_X1 U9944 ( .B1(n8230), .B2(n10337), .A(n8143), .ZN(P2_U3417) );
  NAND2_X1 U9945 ( .A1(n9591), .A2(n10053), .ZN(n8144) );
  OAI211_X1 U9946 ( .C1(n9152), .C2(n10057), .A(n8145), .B(n8144), .ZN(n8147)
         );
  AOI211_X1 U9947 ( .C1(n10241), .C2(n8148), .A(n8147), .B(n8146), .ZN(n8154)
         );
  AOI22_X1 U9948 ( .A1(n10063), .A2(n9183), .B1(P1_REG1_REG_8__SCAN_IN), .B2(
        n4409), .ZN(n8149) );
  OAI21_X1 U9949 ( .B1(n8154), .B2(n4409), .A(n8149), .ZN(P1_U3530) );
  INV_X1 U9950 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8150) );
  OAI22_X1 U9951 ( .A1(n10090), .A2(n8151), .B1(n10243), .B2(n8150), .ZN(n8152) );
  INV_X1 U9952 ( .A(n8152), .ZN(n8153) );
  OAI21_X1 U9953 ( .B1(n8154), .B2(n7144), .A(n8153), .ZN(P1_U3477) );
  NAND2_X1 U9954 ( .A1(n9590), .A2(n10053), .ZN(n8155) );
  OAI211_X1 U9955 ( .C1(n9911), .C2(n10057), .A(n8156), .B(n8155), .ZN(n8158)
         );
  AOI211_X1 U9956 ( .C1(n10241), .C2(n8159), .A(n8158), .B(n8157), .ZN(n8162)
         );
  AOI22_X1 U9957 ( .A1(n7027), .A2(n7093), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n7144), .ZN(n8160) );
  OAI21_X1 U9958 ( .B1(n8162), .B2(n7144), .A(n8160), .ZN(P1_U3486) );
  AOI22_X1 U9959 ( .A1(n7027), .A2(n10063), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n4409), .ZN(n8161) );
  OAI21_X1 U9960 ( .B1(n8162), .B2(n4409), .A(n8161), .ZN(P1_U3533) );
  XNOR2_X1 U9961 ( .A(n8163), .B(n8364), .ZN(n8210) );
  XNOR2_X1 U9962 ( .A(n8210), .B(n8606), .ZN(n8168) );
  INV_X1 U9963 ( .A(n8164), .ZN(n8165) );
  OAI21_X1 U9964 ( .B1(n8168), .B2(n8167), .A(n8213), .ZN(n8169) );
  NAND2_X1 U9965 ( .A1(n8169), .A2(n8587), .ZN(n8175) );
  OAI21_X1 U9966 ( .B1(n8577), .B2(n8171), .A(n8170), .ZN(n8173) );
  NOR2_X1 U9967 ( .A1(n8566), .A2(n8182), .ZN(n8172) );
  AOI211_X1 U9968 ( .C1(n8580), .C2(n8605), .A(n8173), .B(n8172), .ZN(n8174)
         );
  OAI211_X1 U9969 ( .C1(n8183), .C2(n8597), .A(n8175), .B(n8174), .ZN(P2_U3161) );
  INV_X1 U9970 ( .A(n8176), .ZN(n8180) );
  OAI222_X1 U9971 ( .A1(n9121), .A2(n8181), .B1(n9123), .B2(n8180), .C1(
        P2_U3151), .C2(n8179), .ZN(P2_U3273) );
  OAI22_X1 U9972 ( .A1(n8744), .A2(n8183), .B1(n8182), .B2(n8912), .ZN(n8186)
         );
  MUX2_X1 U9973 ( .A(n8184), .B(P2_REG2_REG_8__SCAN_IN), .S(n10296), .Z(n8185)
         );
  AOI211_X1 U9974 ( .C1(n7723), .C2(n8187), .A(n8186), .B(n8185), .ZN(n8188)
         );
  INV_X1 U9975 ( .A(n8188), .ZN(P2_U3225) );
  XOR2_X1 U9976 ( .A(n8189), .B(n8190), .Z(n8209) );
  INV_X1 U9977 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U9978 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8439) );
  OAI21_X1 U9979 ( .B1(n8721), .B2(n8191), .A(n8439), .ZN(n8199) );
  INV_X1 U9980 ( .A(n8192), .ZN(n8194) );
  NAND3_X1 U9981 ( .A1(n8195), .A2(n8194), .A3(n8193), .ZN(n8196) );
  AOI21_X1 U9982 ( .B1(n8197), .B2(n8196), .A(n8734), .ZN(n8198) );
  AOI211_X1 U9983 ( .C1(n8632), .C2(n8200), .A(n8199), .B(n8198), .ZN(n8208)
         );
  INV_X1 U9984 ( .A(n8201), .ZN(n8203) );
  NOR3_X1 U9985 ( .A1(n4432), .A2(n8203), .A3(n8202), .ZN(n8206) );
  INV_X1 U9986 ( .A(n8204), .ZN(n8205) );
  OAI21_X1 U9987 ( .B1(n8206), .B2(n8205), .A(n8730), .ZN(n8207) );
  OAI211_X1 U9988 ( .C1(n8209), .C2(n8722), .A(n8208), .B(n8207), .ZN(P2_U3192) );
  NAND2_X1 U9989 ( .A1(n8210), .A2(n10255), .ZN(n8211) );
  AND2_X1 U9990 ( .A1(n8213), .A2(n8211), .ZN(n8215) );
  XNOR2_X1 U9991 ( .A(n8226), .B(n8394), .ZN(n8340) );
  XNOR2_X1 U9992 ( .A(n8340), .B(n8605), .ZN(n8214) );
  OAI211_X1 U9993 ( .C1(n8215), .C2(n8214), .A(n8587), .B(n8342), .ZN(n8221)
         );
  INV_X1 U9994 ( .A(n8216), .ZN(n8225) );
  AOI21_X1 U9995 ( .B1(n8590), .B2(n8606), .A(n8217), .ZN(n8218) );
  OAI21_X1 U9996 ( .B1(n8554), .B2(n8592), .A(n8218), .ZN(n8219) );
  AOI21_X1 U9997 ( .B1(n8225), .B2(n8594), .A(n8219), .ZN(n8220) );
  OAI211_X1 U9998 ( .C1(n8222), .C2(n8597), .A(n8221), .B(n8220), .ZN(P2_U3171) );
  MUX2_X1 U9999 ( .A(n8223), .B(P2_REG2_REG_9__SCAN_IN), .S(n10296), .Z(n8224)
         );
  INV_X1 U10000 ( .A(n8224), .ZN(n8228) );
  AOI22_X1 U10001 ( .A1(n10292), .A2(n8226), .B1(n10293), .B2(n8225), .ZN(
        n8227) );
  OAI211_X1 U10002 ( .C1(n8229), .C2(n10267), .A(n8228), .B(n8227), .ZN(
        P2_U3224) );
  MUX2_X1 U10003 ( .A(n8231), .B(n8230), .S(n10672), .Z(n8232) );
  INV_X1 U10004 ( .A(n8232), .ZN(P2_U3468) );
  NAND2_X1 U10005 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  XNOR2_X1 U10006 ( .A(n8235), .B(n8236), .ZN(n8269) );
  XOR2_X1 U10007 ( .A(n8237), .B(n8236), .Z(n8238) );
  AOI222_X1 U10008 ( .A1(n10289), .A2(n8238), .B1(n8603), .B2(n10284), .C1(
        n8605), .C2(n10286), .ZN(n8264) );
  INV_X1 U10009 ( .A(n8264), .ZN(n8239) );
  NAND2_X1 U10010 ( .A1(n8239), .A2(n10336), .ZN(n8241) );
  AOI22_X1 U10011 ( .A1(n9093), .A2(n8444), .B1(n10337), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n8240) );
  OAI211_X1 U10012 ( .C1(n8269), .C2(n9096), .A(n8241), .B(n8240), .ZN(
        P2_U3420) );
  NAND2_X1 U10013 ( .A1(n8245), .A2(n10108), .ZN(n8242) );
  OAI211_X1 U10014 ( .C1(n8243), .C2(n10116), .A(n8242), .B(n9575), .ZN(
        P1_U3332) );
  NAND2_X1 U10015 ( .A1(n8245), .A2(n8244), .ZN(n8247) );
  OAI211_X1 U10016 ( .C1(n10501), .C2(n9121), .A(n8247), .B(n8246), .ZN(
        P2_U3272) );
  XOR2_X1 U10017 ( .A(n8248), .B(n8249), .Z(n8260) );
  OAI21_X1 U10018 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n8250), .A(n8289), .ZN(
        n8255) );
  NOR2_X1 U10019 ( .A1(n8717), .A2(n8251), .ZN(n8254) );
  INV_X1 U10020 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U10021 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8552) );
  OAI21_X1 U10022 ( .B1(n8721), .B2(n8252), .A(n8552), .ZN(n8253) );
  AOI211_X1 U10023 ( .C1(n8255), .C2(n8639), .A(n8254), .B(n8253), .ZN(n8259)
         );
  OAI21_X1 U10024 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8256), .A(n8295), .ZN(
        n8257) );
  NAND2_X1 U10025 ( .A1(n8257), .A2(n8730), .ZN(n8258) );
  OAI211_X1 U10026 ( .C1(n8260), .C2(n8722), .A(n8259), .B(n8258), .ZN(
        P2_U3193) );
  INV_X1 U10027 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8261) );
  MUX2_X1 U10028 ( .A(n8261), .B(n8264), .S(n10672), .Z(n8263) );
  NAND2_X1 U10029 ( .A1(n9007), .A2(n8444), .ZN(n8262) );
  OAI211_X1 U10030 ( .C1(n8269), .C2(n9010), .A(n8263), .B(n8262), .ZN(
        P2_U3469) );
  INV_X1 U10031 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8265) );
  MUX2_X1 U10032 ( .A(n8265), .B(n8264), .S(n10282), .Z(n8268) );
  INV_X1 U10033 ( .A(n8442), .ZN(n8266) );
  AOI22_X1 U10034 ( .A1(n10292), .A2(n8444), .B1(n10293), .B2(n8266), .ZN(
        n8267) );
  OAI211_X1 U10035 ( .C1(n8269), .C2(n8941), .A(n8268), .B(n8267), .ZN(
        P2_U3223) );
  XNOR2_X1 U10036 ( .A(n8270), .B(n8347), .ZN(n8284) );
  XNOR2_X1 U10037 ( .A(n8271), .B(n8347), .ZN(n8272) );
  NAND2_X1 U10038 ( .A1(n8272), .A2(n10289), .ZN(n8274) );
  AOI22_X1 U10039 ( .A1(n10284), .A2(n8931), .B1(n8604), .B2(n10286), .ZN(
        n8273) );
  AND2_X1 U10040 ( .A1(n8274), .A2(n8273), .ZN(n8280) );
  MUX2_X1 U10041 ( .A(n8280), .B(n8275), .S(n10337), .Z(n8277) );
  NAND2_X1 U10042 ( .A1(n9093), .A2(n8548), .ZN(n8276) );
  OAI211_X1 U10043 ( .C1(n8284), .C2(n9096), .A(n8277), .B(n8276), .ZN(
        P2_U3423) );
  MUX2_X1 U10044 ( .A(n8280), .B(n4858), .S(n8960), .Z(n8279) );
  NAND2_X1 U10045 ( .A1(n8548), .A2(n9007), .ZN(n8278) );
  OAI211_X1 U10046 ( .C1(n8284), .C2(n9010), .A(n8279), .B(n8278), .ZN(
        P2_U3470) );
  MUX2_X1 U10047 ( .A(n8280), .B(n10488), .S(n10296), .Z(n8283) );
  INV_X1 U10048 ( .A(n8281), .ZN(n8556) );
  AOI22_X1 U10049 ( .A1(n8548), .A2(n10292), .B1(n10293), .B2(n8556), .ZN(
        n8282) );
  OAI211_X1 U10050 ( .C1(n8284), .C2(n8941), .A(n8283), .B(n8282), .ZN(
        P2_U3222) );
  XOR2_X1 U10051 ( .A(n8286), .B(n8285), .Z(n8304) );
  INV_X1 U10052 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10053 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8476) );
  OAI21_X1 U10054 ( .B1(n8721), .B2(n8287), .A(n8476), .ZN(n8293) );
  NAND3_X1 U10055 ( .A1(n8289), .A2(n4531), .A3(n8288), .ZN(n8290) );
  AOI21_X1 U10056 ( .B1(n8291), .B2(n8290), .A(n8734), .ZN(n8292) );
  AOI211_X1 U10057 ( .C1(n8632), .C2(n8294), .A(n8293), .B(n8292), .ZN(n8303)
         );
  INV_X1 U10058 ( .A(n8295), .ZN(n8298) );
  NOR3_X1 U10059 ( .A1(n8298), .A2(n4898), .A3(n8297), .ZN(n8301) );
  INV_X1 U10060 ( .A(n8299), .ZN(n8300) );
  OAI21_X1 U10061 ( .B1(n8301), .B2(n8300), .A(n8730), .ZN(n8302) );
  OAI211_X1 U10062 ( .C1(n8304), .C2(n8722), .A(n8303), .B(n8302), .ZN(
        P2_U3194) );
  INV_X1 U10063 ( .A(n8305), .ZN(n8309) );
  OAI222_X1 U10064 ( .A1(P2_U3151), .A2(n8307), .B1(n9123), .B2(n8309), .C1(
        n8306), .C2(n9121), .ZN(P2_U3271) );
  OAI222_X1 U10065 ( .A1(n8310), .A2(P1_U3086), .B1(n8337), .B2(n8309), .C1(
        n8308), .C2(n10116), .ZN(P1_U3331) );
  INV_X1 U10066 ( .A(n7098), .ZN(n9109) );
  NAND2_X1 U10067 ( .A1(n9675), .A2(n6933), .ZN(n8315) );
  NAND2_X1 U10068 ( .A1(n9657), .A2(n8313), .ZN(n8314) );
  NAND2_X1 U10069 ( .A1(n8315), .A2(n8314), .ZN(n8317) );
  XNOR2_X1 U10070 ( .A(n8317), .B(n8316), .ZN(n8321) );
  NOR2_X1 U10071 ( .A1(n9947), .A2(n8318), .ZN(n8319) );
  AOI21_X1 U10072 ( .B1(n9675), .B2(n8313), .A(n8319), .ZN(n8320) );
  XNOR2_X1 U10073 ( .A(n8321), .B(n8320), .ZN(n8322) );
  INV_X1 U10074 ( .A(n8322), .ZN(n8328) );
  NAND3_X1 U10075 ( .A1(n8328), .A2(n9320), .A3(n8327), .ZN(n8333) );
  INV_X1 U10076 ( .A(n9667), .ZN(n8324) );
  AOI22_X1 U10077 ( .A1(n8324), .A2(n9338), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8326) );
  NAND2_X1 U10078 ( .A1(n9669), .A2(n9332), .ZN(n8325) );
  OAI211_X1 U10079 ( .C1(n9671), .C2(n9334), .A(n8326), .B(n8325), .ZN(n8330)
         );
  NOR3_X1 U10080 ( .A1(n8328), .A2(n8327), .A3(n9340), .ZN(n8329) );
  AOI211_X1 U10081 ( .C1(n9675), .C2(n9272), .A(n8330), .B(n8329), .ZN(n8331)
         );
  OAI211_X1 U10082 ( .C1(n8334), .C2(n8333), .A(n8332), .B(n8331), .ZN(
        P1_U3220) );
  INV_X1 U10083 ( .A(n8335), .ZN(n8407) );
  XNOR2_X1 U10084 ( .A(n8444), .B(n8394), .ZN(n8436) );
  XNOR2_X1 U10085 ( .A(n8345), .B(n8381), .ZN(n8550) );
  OAI21_X1 U10086 ( .B1(n8554), .B2(n8436), .A(n8550), .ZN(n8351) );
  NAND3_X1 U10087 ( .A1(n8343), .A2(n8554), .A3(n8381), .ZN(n8344) );
  OAI211_X1 U10088 ( .C1(n8603), .C2(n8381), .A(n8345), .B(n8344), .ZN(n8349)
         );
  NAND3_X1 U10089 ( .A1(n8444), .A2(n8554), .A3(n8364), .ZN(n8346) );
  OAI211_X1 U10090 ( .C1(n8364), .C2(n8603), .A(n8347), .B(n8346), .ZN(n8348)
         );
  XNOR2_X1 U10091 ( .A(n8482), .B(n8394), .ZN(n8353) );
  XNOR2_X1 U10092 ( .A(n8353), .B(n8352), .ZN(n8475) );
  AOI21_X1 U10093 ( .B1(n8349), .B2(n8348), .A(n8475), .ZN(n8350) );
  INV_X1 U10094 ( .A(n8533), .ZN(n8356) );
  XNOR2_X1 U10095 ( .A(n9092), .B(n8394), .ZN(n8354) );
  NAND2_X1 U10096 ( .A1(n8354), .A2(n8477), .ZN(n8357) );
  OAI21_X1 U10097 ( .B1(n8354), .B2(n8477), .A(n8357), .ZN(n8532) );
  NAND2_X1 U10098 ( .A1(n8356), .A2(n8355), .ZN(n8530) );
  NAND2_X1 U10099 ( .A1(n8530), .A2(n8357), .ZN(n8419) );
  XNOR2_X1 U10100 ( .A(n4626), .B(n8394), .ZN(n8358) );
  XNOR2_X1 U10101 ( .A(n8358), .B(n8932), .ZN(n8420) );
  XNOR2_X1 U10102 ( .A(n8998), .B(n8364), .ZN(n8360) );
  XNOR2_X1 U10103 ( .A(n8360), .B(n8921), .ZN(n8588) );
  NAND2_X1 U10104 ( .A1(n8358), .A2(n8907), .ZN(n8584) );
  XNOR2_X1 U10105 ( .A(n8902), .B(n8394), .ZN(n8497) );
  NAND2_X1 U10106 ( .A1(n8497), .A2(n8908), .ZN(n8362) );
  NAND2_X1 U10107 ( .A1(n8363), .A2(n8362), .ZN(n8506) );
  XNOR2_X1 U10108 ( .A(n9071), .B(n8364), .ZN(n8365) );
  XNOR2_X1 U10109 ( .A(n8365), .B(n8865), .ZN(n8505) );
  NAND2_X1 U10110 ( .A1(n8506), .A2(n8505), .ZN(n8367) );
  XNOR2_X1 U10111 ( .A(n8871), .B(n8394), .ZN(n8368) );
  XNOR2_X1 U10112 ( .A(n8368), .B(n8601), .ZN(n8560) );
  NAND2_X1 U10113 ( .A1(n8368), .A2(n8883), .ZN(n8369) );
  XNOR2_X1 U10114 ( .A(n8987), .B(n8381), .ZN(n8448) );
  NOR2_X1 U10115 ( .A1(n8448), .A2(n8866), .ZN(n8372) );
  NAND2_X1 U10116 ( .A1(n8448), .A2(n8866), .ZN(n8371) );
  XNOR2_X1 U10117 ( .A(n9060), .B(n8394), .ZN(n8373) );
  NAND2_X1 U10118 ( .A1(n8373), .A2(n8855), .ZN(n8456) );
  OAI21_X1 U10119 ( .B1(n8373), .B2(n8855), .A(n8456), .ZN(n8524) );
  XNOR2_X1 U10120 ( .A(n9054), .B(n8394), .ZN(n8374) );
  NAND2_X1 U10121 ( .A1(n8374), .A2(n8816), .ZN(n8378) );
  INV_X1 U10122 ( .A(n8374), .ZN(n8375) );
  NAND2_X1 U10123 ( .A1(n8375), .A2(n8845), .ZN(n8376) );
  XNOR2_X1 U10124 ( .A(n8825), .B(n8394), .ZN(n8379) );
  XNOR2_X1 U10125 ( .A(n8379), .B(n8834), .ZN(n8541) );
  NAND2_X1 U10126 ( .A1(n8379), .A2(n8465), .ZN(n8380) );
  XNOR2_X1 U10127 ( .A(n9045), .B(n8381), .ZN(n8428) );
  NOR2_X1 U10128 ( .A1(n8428), .A2(n8788), .ZN(n8384) );
  XNOR2_X1 U10129 ( .A(n8792), .B(n8381), .ZN(n8382) );
  NAND2_X1 U10130 ( .A1(n8382), .A2(n8493), .ZN(n8486) );
  OAI21_X1 U10131 ( .B1(n8382), .B2(n8493), .A(n8486), .ZN(n8512) );
  AOI21_X1 U10132 ( .B1(n8788), .B2(n8428), .A(n8512), .ZN(n8383) );
  OAI21_X2 U10133 ( .B1(n8427), .B2(n8384), .A(n8383), .ZN(n8485) );
  XNOR2_X1 U10134 ( .A(n9034), .B(n8394), .ZN(n8385) );
  NAND2_X1 U10135 ( .A1(n8385), .A2(n8578), .ZN(n8389) );
  INV_X1 U10136 ( .A(n8385), .ZN(n8386) );
  NAND2_X1 U10137 ( .A1(n8386), .A2(n8789), .ZN(n8387) );
  XNOR2_X1 U10138 ( .A(n9028), .B(n8394), .ZN(n8390) );
  XNOR2_X1 U10139 ( .A(n8390), .B(n8779), .ZN(n8574) );
  XNOR2_X1 U10140 ( .A(n8392), .B(n8401), .ZN(n8411) );
  INV_X1 U10141 ( .A(n8390), .ZN(n8391) );
  NOR2_X1 U10142 ( .A1(n8391), .A2(n8779), .ZN(n8412) );
  NAND2_X1 U10143 ( .A1(n8413), .A2(n8393), .ZN(n8397) );
  XNOR2_X1 U10144 ( .A(n8395), .B(n8394), .ZN(n8396) );
  XNOR2_X1 U10145 ( .A(n8397), .B(n8396), .ZN(n8405) );
  NOR2_X1 U10146 ( .A1(n8398), .A2(n8592), .ZN(n8403) );
  AOI22_X1 U10147 ( .A1(n8399), .A2(n8594), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8400) );
  OAI21_X1 U10148 ( .B1(n8401), .B2(n8577), .A(n8400), .ZN(n8402) );
  AOI211_X1 U10149 ( .C1(n8951), .C2(n8568), .A(n8403), .B(n8402), .ZN(n8404)
         );
  OAI21_X1 U10150 ( .B1(n8405), .B2(n8570), .A(n8404), .ZN(P2_U3160) );
  OAI222_X1 U10151 ( .A1(P2_U3151), .A2(n8408), .B1(n9123), .B2(n8407), .C1(
        n8406), .C2(n9121), .ZN(P2_U3265) );
  INV_X1 U10152 ( .A(n8409), .ZN(n9112) );
  INV_X1 U10153 ( .A(n8762), .ZN(n9026) );
  NAND3_X1 U10154 ( .A1(n8414), .A2(n8587), .A3(n8413), .ZN(n8418) );
  AOI22_X1 U10155 ( .A1(n8758), .A2(n8594), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8415) );
  OAI21_X1 U10156 ( .B1(n8755), .B2(n8577), .A(n8415), .ZN(n8416) );
  AOI21_X1 U10157 ( .B1(n8580), .B2(n8757), .A(n8416), .ZN(n8417) );
  OAI211_X1 U10158 ( .C1(n9026), .C2(n8597), .A(n8418), .B(n8417), .ZN(
        P2_U3154) );
  INV_X1 U10159 ( .A(n4626), .ZN(n8426) );
  OAI21_X1 U10160 ( .B1(n8420), .B2(n8419), .A(n8585), .ZN(n8421) );
  NAND2_X1 U10161 ( .A1(n8421), .A2(n8587), .ZN(n8425) );
  AND2_X1 U10162 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8647) );
  AOI21_X1 U10163 ( .B1(n8580), .B2(n8921), .A(n8647), .ZN(n8422) );
  OAI21_X1 U10164 ( .B1(n8477), .B2(n8577), .A(n8422), .ZN(n8423) );
  AOI21_X1 U10165 ( .B1(n8923), .B2(n8594), .A(n8423), .ZN(n8424) );
  OAI211_X1 U10166 ( .C1(n8426), .C2(n8597), .A(n8425), .B(n8424), .ZN(
        P2_U3155) );
  INV_X1 U10167 ( .A(n8428), .ZN(n8429) );
  NAND2_X1 U10168 ( .A1(n8427), .A2(n8429), .ZN(n8513) );
  OAI21_X1 U10169 ( .B1(n8427), .B2(n8429), .A(n8513), .ZN(n8430) );
  NOR2_X1 U10170 ( .A1(n8430), .A2(n8788), .ZN(n8516) );
  AOI21_X1 U10171 ( .B1(n8788), .B2(n8430), .A(n8516), .ZN(n8435) );
  AND2_X1 U10172 ( .A1(P2_U3151), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U10173 ( .A1(n8465), .A2(n8577), .ZN(n8431) );
  AOI211_X1 U10174 ( .C1(n8810), .C2(n8594), .A(n10417), .B(n8431), .ZN(n8432)
         );
  OAI21_X1 U10175 ( .B1(n8493), .B2(n8592), .A(n8432), .ZN(n8433) );
  AOI21_X1 U10176 ( .B1(n9045), .B2(n8568), .A(n8433), .ZN(n8434) );
  OAI21_X1 U10177 ( .B1(n8435), .B2(n8570), .A(n8434), .ZN(P2_U3156) );
  INV_X1 U10178 ( .A(n8436), .ZN(n8438) );
  XNOR2_X1 U10179 ( .A(n8470), .B(n8604), .ZN(n8437) );
  NOR2_X1 U10180 ( .A1(n8437), .A2(n8438), .ZN(n8471) );
  AOI21_X1 U10181 ( .B1(n8438), .B2(n8437), .A(n8471), .ZN(n8446) );
  OAI21_X1 U10182 ( .B1(n8592), .B2(n8473), .A(n8439), .ZN(n8440) );
  AOI21_X1 U10183 ( .B1(n8590), .B2(n8605), .A(n8440), .ZN(n8441) );
  OAI21_X1 U10184 ( .B1(n8566), .B2(n8442), .A(n8441), .ZN(n8443) );
  AOI21_X1 U10185 ( .B1(n8444), .B2(n8568), .A(n8443), .ZN(n8445) );
  OAI21_X1 U10186 ( .B1(n8446), .B2(n8570), .A(n8445), .ZN(P2_U3157) );
  XNOR2_X1 U10187 ( .A(n8448), .B(n8866), .ZN(n8449) );
  XNOR2_X1 U10188 ( .A(n8447), .B(n8449), .ZN(n8455) );
  AOI21_X1 U10189 ( .B1(n8833), .B2(n8580), .A(n8450), .ZN(n8452) );
  NAND2_X1 U10190 ( .A1(n8594), .A2(n8859), .ZN(n8451) );
  OAI211_X1 U10191 ( .C1(n8883), .C2(n8577), .A(n8452), .B(n8451), .ZN(n8453)
         );
  AOI21_X1 U10192 ( .B1(n8987), .B2(n8568), .A(n8453), .ZN(n8454) );
  OAI21_X1 U10193 ( .B1(n8455), .B2(n8570), .A(n8454), .ZN(P2_U3159) );
  INV_X1 U10194 ( .A(n4558), .ZN(n8469) );
  INV_X1 U10195 ( .A(n8456), .ZN(n8458) );
  NOR3_X1 U10196 ( .A1(n5191), .A2(n8458), .A3(n8457), .ZN(n8463) );
  OR2_X1 U10197 ( .A1(n8523), .A2(n8459), .ZN(n8461) );
  NAND2_X1 U10198 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  OAI21_X1 U10199 ( .B1(n8463), .B2(n8462), .A(n8587), .ZN(n8468) );
  AOI22_X1 U10200 ( .A1(n8833), .A2(n8590), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8464) );
  OAI21_X1 U10201 ( .B1(n8465), .B2(n8592), .A(n8464), .ZN(n8466) );
  AOI21_X1 U10202 ( .B1(n8837), .B2(n8594), .A(n8466), .ZN(n8467) );
  OAI211_X1 U10203 ( .C1(n8469), .C2(n8597), .A(n8468), .B(n8467), .ZN(
        P2_U3163) );
  INV_X1 U10204 ( .A(n8470), .ZN(n8472) );
  AOI21_X1 U10205 ( .B1(n8472), .B2(n8554), .A(n8471), .ZN(n8551) );
  NAND2_X1 U10206 ( .A1(n8551), .A2(n8550), .ZN(n8549) );
  OAI21_X1 U10207 ( .B1(n8473), .B2(n8550), .A(n8549), .ZN(n8474) );
  XOR2_X1 U10208 ( .A(n8475), .B(n8474), .Z(n8484) );
  OAI21_X1 U10209 ( .B1(n8592), .B2(n8477), .A(n8476), .ZN(n8478) );
  AOI21_X1 U10210 ( .B1(n8590), .B2(n8603), .A(n8478), .ZN(n8479) );
  OAI21_X1 U10211 ( .B1(n8566), .B2(n8480), .A(n8479), .ZN(n8481) );
  AOI21_X1 U10212 ( .B1(n8482), .B2(n8568), .A(n8481), .ZN(n8483) );
  OAI21_X1 U10213 ( .B1(n8484), .B2(n8570), .A(n8483), .ZN(P2_U3164) );
  INV_X1 U10214 ( .A(n8485), .ZN(n8517) );
  INV_X1 U10215 ( .A(n8486), .ZN(n8488) );
  NOR3_X1 U10216 ( .A1(n8517), .A2(n8488), .A3(n8487), .ZN(n8491) );
  INV_X1 U10217 ( .A(n8489), .ZN(n8490) );
  OAI21_X1 U10218 ( .B1(n8491), .B2(n8490), .A(n8587), .ZN(n8496) );
  AOI22_X1 U10219 ( .A1(n8782), .A2(n8594), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8492) );
  OAI21_X1 U10220 ( .B1(n8493), .B2(n8577), .A(n8492), .ZN(n8494) );
  AOI21_X1 U10221 ( .B1(n8580), .B2(n8779), .A(n8494), .ZN(n8495) );
  OAI211_X1 U10222 ( .C1(n5732), .C2(n8597), .A(n8496), .B(n8495), .ZN(
        P2_U3165) );
  XNOR2_X1 U10223 ( .A(n8497), .B(n8602), .ZN(n8498) );
  XNOR2_X1 U10224 ( .A(n8499), .B(n8498), .ZN(n8504) );
  NAND2_X1 U10225 ( .A1(n8590), .A2(n8921), .ZN(n8500) );
  NAND2_X1 U10226 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8683) );
  OAI211_X1 U10227 ( .C1(n8894), .C2(n8592), .A(n8500), .B(n8683), .ZN(n8502)
         );
  INV_X1 U10228 ( .A(n8902), .ZN(n9076) );
  NOR2_X1 U10229 ( .A1(n9076), .A2(n8597), .ZN(n8501) );
  AOI211_X1 U10230 ( .C1(n8901), .C2(n8594), .A(n8502), .B(n8501), .ZN(n8503)
         );
  OAI21_X1 U10231 ( .B1(n8504), .B2(n8570), .A(n8503), .ZN(P2_U3166) );
  XOR2_X1 U10232 ( .A(n8506), .B(n8505), .Z(n8511) );
  NAND2_X1 U10233 ( .A1(n8601), .A2(n8580), .ZN(n8507) );
  NAND2_X1 U10234 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8700) );
  OAI211_X1 U10235 ( .C1(n8908), .C2(n8577), .A(n8507), .B(n8700), .ZN(n8508)
         );
  AOI21_X1 U10236 ( .B1(n8887), .B2(n8594), .A(n8508), .ZN(n8510) );
  NAND2_X1 U10237 ( .A1(n9071), .A2(n8568), .ZN(n8509) );
  OAI211_X1 U10238 ( .C1(n8511), .C2(n8570), .A(n8510), .B(n8509), .ZN(
        P2_U3168) );
  INV_X1 U10239 ( .A(n8512), .ZN(n8515) );
  INV_X1 U10240 ( .A(n8513), .ZN(n8514) );
  NOR3_X1 U10241 ( .A1(n8516), .A2(n8515), .A3(n8514), .ZN(n8518) );
  OAI21_X1 U10242 ( .B1(n8518), .B2(n8517), .A(n8587), .ZN(n8522) );
  AOI22_X1 U10243 ( .A1(n8794), .A2(n8594), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8519) );
  OAI21_X1 U10244 ( .B1(n8817), .B2(n8577), .A(n8519), .ZN(n8520) );
  AOI21_X1 U10245 ( .B1(n8789), .B2(n8580), .A(n8520), .ZN(n8521) );
  OAI211_X1 U10246 ( .C1(n8792), .C2(n8597), .A(n8522), .B(n8521), .ZN(
        P2_U3169) );
  AOI21_X1 U10247 ( .B1(n8524), .B2(n8523), .A(n5191), .ZN(n8529) );
  AOI22_X1 U10248 ( .A1(n8866), .A2(n8590), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8526) );
  NAND2_X1 U10249 ( .A1(n8594), .A2(n8848), .ZN(n8525) );
  OAI211_X1 U10250 ( .C1(n8816), .C2(n8592), .A(n8526), .B(n8525), .ZN(n8527)
         );
  AOI21_X1 U10251 ( .B1(n9060), .B2(n8568), .A(n8527), .ZN(n8528) );
  OAI21_X1 U10252 ( .B1(n8529), .B2(n8570), .A(n8528), .ZN(P2_U3173) );
  INV_X1 U10253 ( .A(n8530), .ZN(n8531) );
  AOI21_X1 U10254 ( .B1(n8533), .B2(n8532), .A(n8531), .ZN(n8538) );
  NAND2_X1 U10255 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8629) );
  OAI21_X1 U10256 ( .B1(n8592), .B2(n8907), .A(n8629), .ZN(n8534) );
  AOI21_X1 U10257 ( .B1(n8590), .B2(n8931), .A(n8534), .ZN(n8535) );
  OAI21_X1 U10258 ( .B1(n8566), .B2(n8934), .A(n8535), .ZN(n8536) );
  AOI21_X1 U10259 ( .B1(n9092), .B2(n8568), .A(n8536), .ZN(n8537) );
  OAI21_X1 U10260 ( .B1(n8538), .B2(n8570), .A(n8537), .ZN(P2_U3174) );
  INV_X1 U10261 ( .A(n8825), .ZN(n9051) );
  OAI21_X1 U10262 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8542) );
  NAND2_X1 U10263 ( .A1(n8542), .A2(n8587), .ZN(n8547) );
  INV_X1 U10264 ( .A(n8543), .ZN(n8819) );
  AOI22_X1 U10265 ( .A1(n8845), .A2(n8590), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8544) );
  OAI21_X1 U10266 ( .B1(n8819), .B2(n8566), .A(n8544), .ZN(n8545) );
  AOI21_X1 U10267 ( .B1(n8580), .B2(n8788), .A(n8545), .ZN(n8546) );
  OAI211_X1 U10268 ( .C1(n9051), .C2(n8597), .A(n8547), .B(n8546), .ZN(
        P2_U3175) );
  INV_X1 U10269 ( .A(n8548), .ZN(n8559) );
  OAI211_X1 U10270 ( .C1(n8551), .C2(n8550), .A(n8549), .B(n8587), .ZN(n8558)
         );
  NAND2_X1 U10271 ( .A1(n8580), .A2(n8931), .ZN(n8553) );
  OAI211_X1 U10272 ( .C1(n8554), .C2(n8577), .A(n8553), .B(n8552), .ZN(n8555)
         );
  AOI21_X1 U10273 ( .B1(n8556), .B2(n8594), .A(n8555), .ZN(n8557) );
  OAI211_X1 U10274 ( .C1(n8559), .C2(n8597), .A(n8558), .B(n8557), .ZN(
        P2_U3176) );
  XOR2_X1 U10275 ( .A(n8561), .B(n8560), .Z(n8571) );
  INV_X1 U10276 ( .A(n8562), .ZN(n8868) );
  NAND2_X1 U10277 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8720) );
  OAI21_X1 U10278 ( .B1(n8563), .B2(n8592), .A(n8720), .ZN(n8564) );
  AOI21_X1 U10279 ( .B1(n8590), .B2(n8865), .A(n8564), .ZN(n8565) );
  OAI21_X1 U10280 ( .B1(n8868), .B2(n8566), .A(n8565), .ZN(n8567) );
  AOI21_X1 U10281 ( .B1(n8871), .B2(n8568), .A(n8567), .ZN(n8569) );
  OAI21_X1 U10282 ( .B1(n8571), .B2(n8570), .A(n8569), .ZN(P2_U3178) );
  OAI21_X1 U10283 ( .B1(n8574), .B2(n8573), .A(n8572), .ZN(n8575) );
  NAND2_X1 U10284 ( .A1(n8575), .A2(n8587), .ZN(n8582) );
  AOI22_X1 U10285 ( .A1(n8771), .A2(n8594), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8576) );
  OAI21_X1 U10286 ( .B1(n8578), .B2(n8577), .A(n8576), .ZN(n8579) );
  AOI21_X1 U10287 ( .B1(n8768), .B2(n8580), .A(n8579), .ZN(n8581) );
  OAI211_X1 U10288 ( .C1(n8583), .C2(n8597), .A(n8582), .B(n8581), .ZN(
        P2_U3180) );
  INV_X1 U10289 ( .A(n8998), .ZN(n8598) );
  AND2_X1 U10290 ( .A1(n8585), .A2(n8584), .ZN(n8589) );
  OAI211_X1 U10291 ( .C1(n8589), .C2(n8588), .A(n8587), .B(n8586), .ZN(n8596)
         );
  NAND2_X1 U10292 ( .A1(n8590), .A2(n8932), .ZN(n8591) );
  NAND2_X1 U10293 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8667) );
  OAI211_X1 U10294 ( .C1(n8908), .C2(n8592), .A(n8591), .B(n8667), .ZN(n8593)
         );
  AOI21_X1 U10295 ( .B1(n8911), .B2(n8594), .A(n8593), .ZN(n8595) );
  OAI211_X1 U10296 ( .C1(n8598), .C2(n8597), .A(n8596), .B(n8595), .ZN(
        P2_U3181) );
  MUX2_X1 U10297 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8737), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10298 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8599), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10299 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8600), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10300 ( .A(n8757), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8718), .Z(
        P2_U3519) );
  MUX2_X1 U10301 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8768), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10302 ( .A(n8779), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8718), .Z(
        P2_U3517) );
  MUX2_X1 U10303 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8789), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10304 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8807), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10305 ( .A(n8788), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8718), .Z(
        P2_U3514) );
  MUX2_X1 U10306 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8834), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10307 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8845), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10308 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8833), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10309 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8866), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10310 ( .A(n8601), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8718), .Z(
        P2_U3509) );
  MUX2_X1 U10311 ( .A(n8602), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8718), .Z(
        P2_U3507) );
  MUX2_X1 U10312 ( .A(n8921), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8718), .Z(
        P2_U3506) );
  MUX2_X1 U10313 ( .A(n8932), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8718), .Z(
        P2_U3505) );
  MUX2_X1 U10314 ( .A(n8920), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8718), .Z(
        P2_U3504) );
  MUX2_X1 U10315 ( .A(n8931), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8718), .Z(
        P2_U3503) );
  MUX2_X1 U10316 ( .A(n8603), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8718), .Z(
        P2_U3502) );
  MUX2_X1 U10317 ( .A(n8604), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8718), .Z(
        P2_U3501) );
  MUX2_X1 U10318 ( .A(n8605), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8718), .Z(
        P2_U3500) );
  MUX2_X1 U10319 ( .A(n8606), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8718), .Z(
        P2_U3499) );
  MUX2_X1 U10320 ( .A(n8607), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8718), .Z(
        P2_U3498) );
  MUX2_X1 U10321 ( .A(n8608), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8718), .Z(
        P2_U3497) );
  MUX2_X1 U10322 ( .A(n10275), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8718), .Z(
        P2_U3496) );
  MUX2_X1 U10323 ( .A(n10285), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8718), .Z(
        P2_U3495) );
  MUX2_X1 U10324 ( .A(n10276), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8718), .Z(
        P2_U3494) );
  MUX2_X1 U10325 ( .A(n10287), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8718), .Z(
        P2_U3493) );
  MUX2_X1 U10326 ( .A(n8609), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8718), .Z(
        P2_U3492) );
  MUX2_X1 U10327 ( .A(n6109), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8718), .Z(
        P2_U3491) );
  OAI21_X1 U10328 ( .B1(n8612), .B2(n8611), .A(n8610), .ZN(n8613) );
  AOI22_X1 U10329 ( .A1(n8699), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8639), .B2(
        n8613), .ZN(n8626) );
  OAI21_X1 U10330 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8618) );
  NOR2_X1 U10331 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7621), .ZN(n8617) );
  AOI21_X1 U10332 ( .B1(n8730), .B2(n8618), .A(n8617), .ZN(n8625) );
  NAND2_X1 U10333 ( .A1(n8632), .A2(n8619), .ZN(n8624) );
  OAI211_X1 U10334 ( .C1(n8622), .C2(n8621), .A(n8704), .B(n8620), .ZN(n8623)
         );
  NAND4_X1 U10335 ( .A1(n8626), .A2(n8625), .A3(n8624), .A4(n8623), .ZN(
        P2_U3184) );
  XOR2_X1 U10336 ( .A(n8628), .B(n8627), .Z(n8642) );
  INV_X1 U10337 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8630) );
  OAI21_X1 U10338 ( .B1(n8721), .B2(n8630), .A(n8629), .ZN(n8631) );
  AOI21_X1 U10339 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(n8641) );
  OAI21_X1 U10340 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n4530), .A(n8634), .ZN(
        n8638) );
  OAI21_X1 U10341 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8636), .A(n8635), .ZN(
        n8637) );
  AOI22_X1 U10342 ( .A1(n8639), .A2(n8638), .B1(n8637), .B2(n8730), .ZN(n8640)
         );
  OAI211_X1 U10343 ( .C1(n8642), .C2(n8722), .A(n8641), .B(n8640), .ZN(
        P2_U3195) );
  XOR2_X1 U10344 ( .A(n8644), .B(n8643), .Z(n8662) );
  NOR2_X1 U10345 ( .A1(n8717), .A2(n8645), .ZN(n8646) );
  AOI211_X1 U10346 ( .C1(n8699), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8647), .B(
        n8646), .ZN(n8661) );
  INV_X1 U10347 ( .A(n8648), .ZN(n8650) );
  NAND3_X1 U10348 ( .A1(n8634), .A2(n8650), .A3(n8649), .ZN(n8651) );
  AOI21_X1 U10349 ( .B1(n8652), .B2(n8651), .A(n8734), .ZN(n8659) );
  NAND3_X1 U10350 ( .A1(n8635), .A2(n4903), .A3(n8654), .ZN(n8656) );
  AOI21_X1 U10351 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8658) );
  NOR2_X1 U10352 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  OAI211_X1 U10353 ( .C1(n8662), .C2(n8722), .A(n8661), .B(n8660), .ZN(
        P2_U3196) );
  OAI21_X1 U10354 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n4430), .A(n8663), .ZN(
        n8664) );
  INV_X1 U10355 ( .A(n8664), .ZN(n8675) );
  XNOR2_X1 U10356 ( .A(n8666), .B(n8665), .ZN(n8670) );
  NAND2_X1 U10357 ( .A1(n8699), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U10358 ( .C1(n8717), .C2(n4899), .A(n8668), .B(n8667), .ZN(n8669)
         );
  AOI21_X1 U10359 ( .B1(n8670), .B2(n8704), .A(n8669), .ZN(n8674) );
  OAI21_X1 U10360 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8671), .A(n8689), .ZN(
        n8672) );
  NAND2_X1 U10361 ( .A1(n8672), .A2(n8730), .ZN(n8673) );
  OAI211_X1 U10362 ( .C1(n8675), .C2(n8734), .A(n8674), .B(n8673), .ZN(
        P2_U3197) );
  AND3_X1 U10363 ( .A1(n8663), .A2(n8677), .A3(n8676), .ZN(n8678) );
  NOR2_X1 U10364 ( .A1(n8679), .A2(n8678), .ZN(n8693) );
  XNOR2_X1 U10365 ( .A(n8681), .B(n8680), .ZN(n8686) );
  NAND2_X1 U10366 ( .A1(n8699), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8682) );
  OAI211_X1 U10367 ( .C1(n8717), .C2(n8684), .A(n8683), .B(n8682), .ZN(n8685)
         );
  AOI21_X1 U10368 ( .B1(n8686), .B2(n8704), .A(n8685), .ZN(n8692) );
  AND3_X1 U10369 ( .A1(n8689), .A2(n8688), .A3(n8687), .ZN(n8690) );
  OAI21_X1 U10370 ( .B1(n4884), .B2(n8690), .A(n8730), .ZN(n8691) );
  OAI211_X1 U10371 ( .C1(n8693), .C2(n8734), .A(n8692), .B(n8691), .ZN(
        P2_U3198) );
  OAI21_X1 U10372 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8695), .A(n8694), .ZN(
        n8696) );
  INV_X1 U10373 ( .A(n8696), .ZN(n8709) );
  XNOR2_X1 U10374 ( .A(n8698), .B(n8697), .ZN(n8705) );
  NAND2_X1 U10375 ( .A1(n8699), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8701) );
  OAI211_X1 U10376 ( .C1(n8717), .C2(n8702), .A(n8701), .B(n8700), .ZN(n8703)
         );
  AOI21_X1 U10377 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8708) );
  OAI21_X1 U10378 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n4506), .A(n8729), .ZN(
        n8706) );
  NAND2_X1 U10379 ( .A1(n8706), .A2(n8730), .ZN(n8707) );
  OAI211_X1 U10380 ( .C1(n8709), .C2(n8734), .A(n8708), .B(n8707), .ZN(
        P2_U3199) );
  AND3_X1 U10381 ( .A1(n8694), .A2(n8711), .A3(n8710), .ZN(n8712) );
  NOR2_X1 U10382 ( .A1(n8713), .A2(n8712), .ZN(n8735) );
  INV_X1 U10383 ( .A(n8714), .ZN(n8715) );
  INV_X1 U10384 ( .A(n8723), .ZN(n8719) );
  OAI21_X1 U10385 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8726) );
  OAI21_X1 U10386 ( .B1(n8721), .B2(n10356), .A(n8720), .ZN(n8725) );
  NOR3_X1 U10387 ( .A1(n8723), .A2(n8727), .A3(n8722), .ZN(n8724) );
  AND3_X1 U10388 ( .A1(n8729), .A2(n4461), .A3(n8728), .ZN(n8731) );
  OAI21_X1 U10389 ( .B1(n8732), .B2(n8731), .A(n8730), .ZN(n8733) );
  NOR2_X1 U10390 ( .A1(n8738), .A2(n8912), .ZN(n8747) );
  AOI21_X1 U10391 ( .B1(n9019), .B2(n10282), .A(n8747), .ZN(n8741) );
  NAND2_X1 U10392 ( .A1(n10296), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8739) );
  OAI211_X1 U10393 ( .C1(n9021), .C2(n8744), .A(n8741), .B(n8739), .ZN(
        P2_U3202) );
  INV_X1 U10394 ( .A(n6085), .ZN(n8947) );
  NAND2_X1 U10395 ( .A1(n10296), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8740) );
  OAI211_X1 U10396 ( .C1(n8947), .C2(n8744), .A(n8741), .B(n8740), .ZN(
        P2_U3203) );
  INV_X1 U10397 ( .A(n8742), .ZN(n8750) );
  NAND2_X1 U10398 ( .A1(n8743), .A2(n10282), .ZN(n8749) );
  NOR2_X1 U10399 ( .A1(n8745), .A2(n8744), .ZN(n8746) );
  AOI211_X1 U10400 ( .C1(n10296), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8747), .B(
        n8746), .ZN(n8748) );
  OAI211_X1 U10401 ( .C1(n8750), .C2(n10267), .A(n8749), .B(n8748), .ZN(
        P2_U3204) );
  OAI21_X1 U10402 ( .B1(n8752), .B2(n8753), .A(n8751), .ZN(n8955) );
  XNOR2_X1 U10403 ( .A(n8754), .B(n5122), .ZN(n8756) );
  OAI21_X1 U10404 ( .B1(n8958), .B2(n8956), .A(n10282), .ZN(n8764) );
  INV_X1 U10405 ( .A(n8758), .ZN(n8760) );
  INV_X1 U10406 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8759) );
  OAI22_X1 U10407 ( .A1(n8760), .A2(n8912), .B1(n10282), .B2(n8759), .ZN(n8761) );
  AOI21_X1 U10408 ( .B1(n8762), .B2(n10292), .A(n8761), .ZN(n8763) );
  OAI211_X1 U10409 ( .C1(n8955), .C2(n8941), .A(n8764), .B(n8763), .ZN(
        P2_U3206) );
  INV_X1 U10410 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8770) );
  XOR2_X1 U10411 ( .A(n8767), .B(n8766), .Z(n8769) );
  AOI222_X1 U10412 ( .A1(n10289), .A2(n8769), .B1(n8768), .B2(n10284), .C1(
        n8789), .C2(n10286), .ZN(n9027) );
  MUX2_X1 U10413 ( .A(n8770), .B(n9027), .S(n10282), .Z(n8773) );
  AOI22_X1 U10414 ( .A1(n9028), .A2(n10292), .B1(n10293), .B2(n8771), .ZN(
        n8772) );
  OAI211_X1 U10415 ( .C1(n9031), .C2(n8941), .A(n8773), .B(n8772), .ZN(
        P2_U3207) );
  OAI21_X1 U10416 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8780) );
  AOI222_X1 U10417 ( .A1(n10289), .A2(n8780), .B1(n8779), .B2(n10284), .C1(
        n8807), .C2(n10286), .ZN(n9032) );
  OAI21_X1 U10418 ( .B1(n5732), .B2(n8791), .A(n9032), .ZN(n8781) );
  NAND2_X1 U10419 ( .A1(n8781), .A2(n10282), .ZN(n8784) );
  AOI22_X1 U10420 ( .A1(n8782), .A2(n10293), .B1(n10296), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8783) );
  OAI211_X1 U10421 ( .C1(n9037), .C2(n8941), .A(n8784), .B(n8783), .ZN(
        P2_U3208) );
  XOR2_X1 U10422 ( .A(n8785), .B(n8786), .Z(n9043) );
  XNOR2_X1 U10423 ( .A(n8787), .B(n8786), .ZN(n8790) );
  AOI222_X1 U10424 ( .A1(n10289), .A2(n8790), .B1(n8789), .B2(n10284), .C1(
        n8788), .C2(n10286), .ZN(n9038) );
  OAI21_X1 U10425 ( .B1(n8792), .B2(n8791), .A(n9038), .ZN(n8793) );
  NAND2_X1 U10426 ( .A1(n8793), .A2(n10282), .ZN(n8796) );
  AOI22_X1 U10427 ( .A1(n8794), .A2(n10293), .B1(n10296), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8795) );
  OAI211_X1 U10428 ( .C1(n9043), .C2(n8941), .A(n8796), .B(n8795), .ZN(
        P2_U3209) );
  NAND2_X1 U10429 ( .A1(n8798), .A2(n8797), .ZN(n8821) );
  NAND2_X1 U10430 ( .A1(n8821), .A2(n8820), .ZN(n8976) );
  NAND2_X1 U10431 ( .A1(n8976), .A2(n8799), .ZN(n8800) );
  XOR2_X1 U10432 ( .A(n8805), .B(n8800), .Z(n9048) );
  INV_X1 U10433 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8809) );
  AOI21_X1 U10434 ( .B1(n8802), .B2(n8801), .A(n8820), .ZN(n8814) );
  INV_X1 U10435 ( .A(n8814), .ZN(n8804) );
  NAND2_X1 U10436 ( .A1(n8804), .A2(n8803), .ZN(n8806) );
  XNOR2_X1 U10437 ( .A(n8806), .B(n8805), .ZN(n8808) );
  AOI222_X1 U10438 ( .A1(n10289), .A2(n8808), .B1(n8807), .B2(n10284), .C1(
        n8834), .C2(n10286), .ZN(n9044) );
  MUX2_X1 U10439 ( .A(n8809), .B(n9044), .S(n10282), .Z(n8812) );
  AOI22_X1 U10440 ( .A1(n9045), .A2(n10292), .B1(n10293), .B2(n8810), .ZN(
        n8811) );
  OAI211_X1 U10441 ( .C1(n9048), .C2(n8941), .A(n8812), .B(n8811), .ZN(
        P2_U3210) );
  OAI21_X1 U10442 ( .B1(n8841), .B2(n8830), .A(n8829), .ZN(n8832) );
  OAI222_X1 U10443 ( .A1(n10254), .A2(n8817), .B1(n10256), .B2(n8816), .C1(
        n8853), .C2(n8815), .ZN(n8975) );
  INV_X1 U10444 ( .A(n8975), .ZN(n8827) );
  OAI22_X1 U10445 ( .A1(n8819), .A2(n8912), .B1(n10282), .B2(n8818), .ZN(n8824) );
  NOR2_X1 U10446 ( .A1(n8821), .A2(n8820), .ZN(n8974) );
  INV_X1 U10447 ( .A(n8976), .ZN(n8822) );
  NOR3_X1 U10448 ( .A1(n8974), .A2(n8822), .A3(n8941), .ZN(n8823) );
  AOI211_X1 U10449 ( .C1(n10292), .C2(n8825), .A(n8824), .B(n8823), .ZN(n8826)
         );
  OAI21_X1 U10450 ( .B1(n8827), .B2(n10296), .A(n8826), .ZN(P2_U3211) );
  XNOR2_X1 U10451 ( .A(n8828), .B(n8829), .ZN(n9057) );
  INV_X1 U10452 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8836) );
  OR3_X1 U10453 ( .A1(n8841), .A2(n8830), .A3(n8829), .ZN(n8831) );
  NAND2_X1 U10454 ( .A1(n8832), .A2(n8831), .ZN(n8835) );
  AOI222_X1 U10455 ( .A1(n10289), .A2(n8835), .B1(n8834), .B2(n10284), .C1(
        n8833), .C2(n10286), .ZN(n9052) );
  MUX2_X1 U10456 ( .A(n8836), .B(n9052), .S(n10282), .Z(n8839) );
  AOI22_X1 U10457 ( .A1(n4558), .A2(n10292), .B1(n10293), .B2(n8837), .ZN(
        n8838) );
  OAI211_X1 U10458 ( .C1(n9057), .C2(n8941), .A(n8839), .B(n8838), .ZN(
        P2_U3212) );
  XOR2_X1 U10459 ( .A(n8843), .B(n8840), .Z(n9063) );
  INV_X1 U10460 ( .A(n8841), .ZN(n8842) );
  OAI21_X1 U10461 ( .B1(n8844), .B2(n8843), .A(n8842), .ZN(n8846) );
  AOI222_X1 U10462 ( .A1(n10289), .A2(n8846), .B1(n8845), .B2(n10284), .C1(
        n8866), .C2(n10286), .ZN(n9058) );
  MUX2_X1 U10463 ( .A(n8847), .B(n9058), .S(n10282), .Z(n8850) );
  AOI22_X1 U10464 ( .A1(n9060), .A2(n10292), .B1(n10293), .B2(n8848), .ZN(
        n8849) );
  OAI211_X1 U10465 ( .C1(n9063), .C2(n8941), .A(n8850), .B(n8849), .ZN(
        P2_U3213) );
  XNOR2_X1 U10466 ( .A(n8852), .B(n8851), .ZN(n8854) );
  OAI222_X1 U10467 ( .A1(n10254), .A2(n8855), .B1(n10256), .B2(n8883), .C1(
        n8854), .C2(n8853), .ZN(n8986) );
  OR2_X1 U10468 ( .A1(n8856), .A2(n4810), .ZN(n8857) );
  NAND2_X1 U10469 ( .A1(n4589), .A2(n8857), .ZN(n9067) );
  AOI22_X1 U10470 ( .A1(n10296), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8859), 
        .B2(n10293), .ZN(n8861) );
  NAND2_X1 U10471 ( .A1(n8987), .A2(n10292), .ZN(n8860) );
  OAI211_X1 U10472 ( .C1(n9067), .C2(n8941), .A(n8861), .B(n8860), .ZN(n8862)
         );
  AOI21_X1 U10473 ( .B1(n8986), .B2(n10282), .A(n8862), .ZN(n8863) );
  INV_X1 U10474 ( .A(n8863), .ZN(P2_U3214) );
  XOR2_X1 U10475 ( .A(n8864), .B(n8875), .Z(n8867) );
  AOI222_X1 U10476 ( .A1(n10289), .A2(n8867), .B1(n8866), .B2(n10284), .C1(
        n8865), .C2(n10286), .ZN(n8991) );
  OAI22_X1 U10477 ( .A1(n10282), .A2(n8869), .B1(n8868), .B2(n8912), .ZN(n8870) );
  AOI21_X1 U10478 ( .B1(n8871), .B2(n10292), .A(n8870), .ZN(n8877) );
  NAND2_X1 U10479 ( .A1(n8874), .A2(n8875), .ZN(n8989) );
  NAND3_X1 U10480 ( .A1(n8873), .A2(n8989), .A3(n7723), .ZN(n8876) );
  OAI211_X1 U10481 ( .C1(n8991), .C2(n10296), .A(n8877), .B(n8876), .ZN(
        P2_U3215) );
  XNOR2_X1 U10482 ( .A(n8879), .B(n8878), .ZN(n9074) );
  INV_X1 U10483 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U10484 ( .A1(n8890), .A2(n8898), .ZN(n8892) );
  NAND2_X1 U10485 ( .A1(n8892), .A2(n8880), .ZN(n8882) );
  XNOR2_X1 U10486 ( .A(n8882), .B(n8881), .ZN(n8885) );
  OAI22_X1 U10487 ( .A1(n8883), .A2(n10254), .B1(n8908), .B2(n10256), .ZN(
        n8884) );
  AOI21_X1 U10488 ( .B1(n8885), .B2(n10289), .A(n8884), .ZN(n9069) );
  MUX2_X1 U10489 ( .A(n8886), .B(n9069), .S(n10282), .Z(n8889) );
  AOI22_X1 U10490 ( .A1(n9071), .A2(n10292), .B1(n10293), .B2(n8887), .ZN(
        n8888) );
  OAI211_X1 U10491 ( .C1(n9074), .C2(n8941), .A(n8889), .B(n8888), .ZN(
        P2_U3216) );
  OR2_X1 U10492 ( .A1(n8890), .A2(n8898), .ZN(n8891) );
  NAND3_X1 U10493 ( .A1(n8892), .A2(n10289), .A3(n8891), .ZN(n8897) );
  OAI22_X1 U10494 ( .A1(n8894), .A2(n10254), .B1(n8893), .B2(n10256), .ZN(
        n8895) );
  INV_X1 U10495 ( .A(n8895), .ZN(n8896) );
  NAND2_X1 U10496 ( .A1(n8897), .A2(n8896), .ZN(n9075) );
  MUX2_X1 U10497 ( .A(n9075), .B(P2_REG2_REG_16__SCAN_IN), .S(n10296), .Z(
        n8905) );
  INV_X1 U10498 ( .A(n8898), .ZN(n8899) );
  XNOR2_X1 U10499 ( .A(n8900), .B(n8899), .ZN(n9077) );
  AOI22_X1 U10500 ( .A1(n8902), .A2(n10292), .B1(n10293), .B2(n8901), .ZN(
        n8903) );
  OAI21_X1 U10501 ( .B1(n9077), .B2(n8941), .A(n8903), .ZN(n8904) );
  XNOR2_X1 U10502 ( .A(n8906), .B(n8915), .ZN(n8910) );
  OAI22_X1 U10503 ( .A1(n8908), .A2(n10254), .B1(n8907), .B2(n10256), .ZN(
        n8909) );
  AOI21_X1 U10504 ( .B1(n8910), .B2(n10289), .A(n8909), .ZN(n9000) );
  INV_X1 U10505 ( .A(n8911), .ZN(n8913) );
  OAI22_X1 U10506 ( .A1(n10282), .A2(n10652), .B1(n8913), .B2(n8912), .ZN(
        n8914) );
  AOI21_X1 U10507 ( .B1(n8998), .B2(n10292), .A(n8914), .ZN(n8918) );
  XNOR2_X1 U10508 ( .A(n8916), .B(n8915), .ZN(n9083) );
  OR2_X1 U10509 ( .A1(n9083), .A2(n8941), .ZN(n8917) );
  OAI211_X1 U10510 ( .C1(n9000), .C2(n10296), .A(n8918), .B(n8917), .ZN(
        P2_U3218) );
  XOR2_X1 U10511 ( .A(n8919), .B(n8926), .Z(n8922) );
  AOI222_X1 U10512 ( .A1(n10289), .A2(n8922), .B1(n8921), .B2(n10284), .C1(
        n8920), .C2(n10286), .ZN(n9084) );
  AOI22_X1 U10513 ( .A1(n4626), .A2(n8936), .B1(n10293), .B2(n8923), .ZN(n8924) );
  AOI21_X1 U10514 ( .B1(n9084), .B2(n8924), .A(n10296), .ZN(n8929) );
  XOR2_X1 U10515 ( .A(n8926), .B(n8925), .Z(n9089) );
  OAI22_X1 U10516 ( .A1(n9089), .A2(n8941), .B1(n8927), .B2(n10282), .ZN(n8928) );
  OR2_X1 U10517 ( .A1(n8929), .A2(n8928), .ZN(P2_U3219) );
  XOR2_X1 U10518 ( .A(n8930), .B(n8939), .Z(n8933) );
  AOI222_X1 U10519 ( .A1(n10289), .A2(n8933), .B1(n8932), .B2(n10284), .C1(
        n8931), .C2(n10286), .ZN(n9090) );
  INV_X1 U10520 ( .A(n8934), .ZN(n8935) );
  AOI22_X1 U10521 ( .A1(n9092), .A2(n8936), .B1(n10293), .B2(n8935), .ZN(n8937) );
  AOI21_X1 U10522 ( .B1(n9090), .B2(n8937), .A(n10296), .ZN(n8943) );
  NAND2_X1 U10523 ( .A1(n9014), .A2(n8938), .ZN(n8940) );
  XNOR2_X1 U10524 ( .A(n8940), .B(n8939), .ZN(n9097) );
  OAI22_X1 U10525 ( .A1(n9097), .A2(n8941), .B1(n10520), .B2(n10282), .ZN(
        n8942) );
  OR2_X1 U10526 ( .A1(n8943), .A2(n8942), .ZN(P2_U3220) );
  NAND2_X1 U10527 ( .A1(n8960), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U10528 ( .A1(n9019), .A2(n10672), .ZN(n8946) );
  OAI211_X1 U10529 ( .C1(n9021), .C2(n9018), .A(n8944), .B(n8946), .ZN(
        P2_U3490) );
  NAND2_X1 U10530 ( .A1(n8960), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8945) );
  OAI211_X1 U10531 ( .C1(n8947), .C2(n9018), .A(n8946), .B(n8945), .ZN(
        P2_U3489) );
  NAND2_X1 U10532 ( .A1(n8960), .A2(n10506), .ZN(n8949) );
  NAND2_X1 U10533 ( .A1(n8951), .A2(n9007), .ZN(n8952) );
  OAI211_X1 U10534 ( .C1(n8954), .C2(n9010), .A(n8953), .B(n8952), .ZN(
        P2_U3487) );
  INV_X1 U10535 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U10536 ( .A1(n8960), .A2(n8959), .ZN(n8961) );
  OAI21_X1 U10537 ( .B1(n9026), .B2(n9018), .A(n8963), .ZN(P2_U3486) );
  MUX2_X1 U10538 ( .A(n10505), .B(n9027), .S(n10672), .Z(n8965) );
  NAND2_X1 U10539 ( .A1(n9028), .A2(n9007), .ZN(n8964) );
  MUX2_X1 U10540 ( .A(n10609), .B(n9032), .S(n10672), .Z(n8967) );
  NAND2_X1 U10541 ( .A1(n9034), .A2(n9007), .ZN(n8966) );
  OAI211_X1 U10542 ( .C1(n9037), .C2(n9010), .A(n8967), .B(n8966), .ZN(
        P2_U3484) );
  INV_X1 U10543 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8968) );
  MUX2_X1 U10544 ( .A(n8968), .B(n9038), .S(n10672), .Z(n8970) );
  NAND2_X1 U10545 ( .A1(n9040), .A2(n9007), .ZN(n8969) );
  OAI211_X1 U10546 ( .C1(n9010), .C2(n9043), .A(n8970), .B(n8969), .ZN(
        P2_U3483) );
  INV_X1 U10547 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8971) );
  MUX2_X1 U10548 ( .A(n8971), .B(n9044), .S(n10672), .Z(n8973) );
  NAND2_X1 U10549 ( .A1(n9045), .A2(n9007), .ZN(n8972) );
  OAI211_X1 U10550 ( .C1(n9048), .C2(n9010), .A(n8973), .B(n8972), .ZN(
        P2_U3482) );
  INV_X1 U10551 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8978) );
  INV_X1 U10552 ( .A(n10327), .ZN(n9011) );
  NOR2_X1 U10553 ( .A1(n8974), .A2(n9011), .ZN(n8977) );
  AOI21_X1 U10554 ( .B1(n8977), .B2(n8976), .A(n8975), .ZN(n9049) );
  MUX2_X1 U10555 ( .A(n8978), .B(n9049), .S(n10672), .Z(n8979) );
  OAI21_X1 U10556 ( .B1(n9051), .B2(n9018), .A(n8979), .ZN(P2_U3481) );
  INV_X1 U10557 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8980) );
  MUX2_X1 U10558 ( .A(n8980), .B(n9052), .S(n10672), .Z(n8982) );
  NAND2_X1 U10559 ( .A1(n4558), .A2(n9007), .ZN(n8981) );
  OAI211_X1 U10560 ( .C1(n9010), .C2(n9057), .A(n8982), .B(n8981), .ZN(
        P2_U3480) );
  INV_X1 U10561 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8983) );
  MUX2_X1 U10562 ( .A(n8983), .B(n9058), .S(n10672), .Z(n8985) );
  NAND2_X1 U10563 ( .A1(n9060), .A2(n9007), .ZN(n8984) );
  OAI211_X1 U10564 ( .C1(n9063), .C2(n9010), .A(n8985), .B(n8984), .ZN(
        P2_U3479) );
  AOI21_X1 U10565 ( .B1(n10316), .B2(n8987), .A(n8986), .ZN(n9064) );
  MUX2_X1 U10566 ( .A(n10545), .B(n9064), .S(n10672), .Z(n8988) );
  OAI21_X1 U10567 ( .B1(n9010), .B2(n9067), .A(n8988), .ZN(P2_U3478) );
  NAND3_X1 U10568 ( .A1(n8873), .A2(n10327), .A3(n8989), .ZN(n8990) );
  OAI211_X1 U10569 ( .C1(n8992), .C2(n10330), .A(n8991), .B(n8990), .ZN(n9068)
         );
  MUX2_X1 U10570 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9068), .S(n10672), .Z(
        P2_U3477) );
  INV_X1 U10571 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8993) );
  MUX2_X1 U10572 ( .A(n8993), .B(n9069), .S(n10672), .Z(n8995) );
  NAND2_X1 U10573 ( .A1(n9071), .A2(n9007), .ZN(n8994) );
  OAI211_X1 U10574 ( .C1(n9010), .C2(n9074), .A(n8995), .B(n8994), .ZN(
        P2_U3476) );
  MUX2_X1 U10575 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9075), .S(n10672), .Z(
        n8997) );
  OAI22_X1 U10576 ( .A1(n9077), .A2(n9010), .B1(n9076), .B2(n9018), .ZN(n8996)
         );
  NAND2_X1 U10577 ( .A1(n8998), .A2(n10316), .ZN(n8999) );
  NAND2_X1 U10578 ( .A1(n9000), .A2(n8999), .ZN(n9080) );
  MUX2_X1 U10579 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9080), .S(n10672), .Z(
        n9001) );
  INV_X1 U10580 ( .A(n9001), .ZN(n9002) );
  OAI21_X1 U10581 ( .B1(n9010), .B2(n9083), .A(n9002), .ZN(P2_U3474) );
  INV_X1 U10582 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U10583 ( .A(n9003), .B(n9084), .S(n10672), .Z(n9005) );
  NAND2_X1 U10584 ( .A1(n4626), .A2(n9007), .ZN(n9004) );
  OAI211_X1 U10585 ( .C1(n9089), .C2(n9010), .A(n9005), .B(n9004), .ZN(
        P2_U3473) );
  INV_X1 U10586 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9006) );
  MUX2_X1 U10587 ( .A(n9006), .B(n9090), .S(n10672), .Z(n9009) );
  NAND2_X1 U10588 ( .A1(n9092), .A2(n9007), .ZN(n9008) );
  OAI211_X1 U10589 ( .C1(n9010), .C2(n9097), .A(n9009), .B(n9008), .ZN(
        P2_U3472) );
  NOR2_X1 U10590 ( .A1(n9012), .A2(n9011), .ZN(n9015) );
  AOI21_X1 U10591 ( .B1(n9015), .B2(n9014), .A(n9013), .ZN(n9098) );
  MUX2_X1 U10592 ( .A(n9016), .B(n9098), .S(n10672), .Z(n9017) );
  OAI21_X1 U10593 ( .B1(n9102), .B2(n9018), .A(n9017), .ZN(P2_U3471) );
  NAND2_X1 U10594 ( .A1(n10337), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U10595 ( .A1(n9019), .A2(n10336), .ZN(n9022) );
  OAI211_X1 U10596 ( .C1(n9021), .C2(n9101), .A(n9020), .B(n9022), .ZN(
        P2_U3458) );
  NAND2_X1 U10597 ( .A1(n6085), .A2(n9093), .ZN(n9023) );
  OAI211_X1 U10598 ( .C1(n10336), .C2(n10446), .A(n9023), .B(n9022), .ZN(
        P2_U3457) );
  MUX2_X1 U10599 ( .A(n10449), .B(n9024), .S(n10336), .Z(n9025) );
  OAI21_X1 U10600 ( .B1(n9026), .B2(n9101), .A(n9025), .ZN(P2_U3454) );
  MUX2_X1 U10601 ( .A(n10590), .B(n9027), .S(n10336), .Z(n9030) );
  NAND2_X1 U10602 ( .A1(n9028), .A2(n9093), .ZN(n9029) );
  INV_X1 U10603 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9033) );
  MUX2_X1 U10604 ( .A(n9033), .B(n9032), .S(n10336), .Z(n9036) );
  NAND2_X1 U10605 ( .A1(n9034), .A2(n9093), .ZN(n9035) );
  OAI211_X1 U10606 ( .C1(n9037), .C2(n9096), .A(n9036), .B(n9035), .ZN(
        P2_U3452) );
  MUX2_X1 U10607 ( .A(n9039), .B(n9038), .S(n10336), .Z(n9042) );
  NAND2_X1 U10608 ( .A1(n9040), .A2(n9093), .ZN(n9041) );
  OAI211_X1 U10609 ( .C1(n9043), .C2(n9096), .A(n9042), .B(n9041), .ZN(
        P2_U3451) );
  MUX2_X1 U10610 ( .A(n10574), .B(n9044), .S(n10336), .Z(n9047) );
  NAND2_X1 U10611 ( .A1(n9045), .A2(n9093), .ZN(n9046) );
  OAI211_X1 U10612 ( .C1(n9048), .C2(n9096), .A(n9047), .B(n9046), .ZN(
        P2_U3450) );
  MUX2_X1 U10613 ( .A(n10655), .B(n9049), .S(n10336), .Z(n9050) );
  MUX2_X1 U10614 ( .A(n9053), .B(n9052), .S(n10336), .Z(n9056) );
  NAND2_X1 U10615 ( .A1(n4558), .A2(n9093), .ZN(n9055) );
  OAI211_X1 U10616 ( .C1(n9057), .C2(n9096), .A(n9056), .B(n9055), .ZN(
        P2_U3448) );
  INV_X1 U10617 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9059) );
  MUX2_X1 U10618 ( .A(n9059), .B(n9058), .S(n10336), .Z(n9062) );
  NAND2_X1 U10619 ( .A1(n9060), .A2(n9093), .ZN(n9061) );
  OAI211_X1 U10620 ( .C1(n9063), .C2(n9096), .A(n9062), .B(n9061), .ZN(
        P2_U3447) );
  INV_X1 U10621 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9065) );
  MUX2_X1 U10622 ( .A(n9065), .B(n9064), .S(n10336), .Z(n9066) );
  OAI21_X1 U10623 ( .B1(n9067), .B2(n9096), .A(n9066), .ZN(P2_U3446) );
  MUX2_X1 U10624 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9068), .S(n10336), .Z(
        P2_U3444) );
  INV_X1 U10625 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9070) );
  MUX2_X1 U10626 ( .A(n9070), .B(n9069), .S(n10336), .Z(n9073) );
  NAND2_X1 U10627 ( .A1(n9071), .A2(n9093), .ZN(n9072) );
  OAI211_X1 U10628 ( .C1(n9074), .C2(n9096), .A(n9073), .B(n9072), .ZN(
        P2_U3441) );
  MUX2_X1 U10629 ( .A(n9075), .B(P2_REG0_REG_16__SCAN_IN), .S(n10337), .Z(
        n9079) );
  OAI22_X1 U10630 ( .A1(n9077), .A2(n9096), .B1(n9076), .B2(n9101), .ZN(n9078)
         );
  MUX2_X1 U10631 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9080), .S(n10336), .Z(
        n9081) );
  INV_X1 U10632 ( .A(n9081), .ZN(n9082) );
  OAI21_X1 U10633 ( .B1(n9083), .B2(n9096), .A(n9082), .ZN(P2_U3435) );
  MUX2_X1 U10634 ( .A(n9085), .B(n9084), .S(n10336), .Z(n9088) );
  NAND2_X1 U10635 ( .A1(n4626), .A2(n9093), .ZN(n9087) );
  OAI211_X1 U10636 ( .C1(n9089), .C2(n9096), .A(n9088), .B(n9087), .ZN(
        P2_U3432) );
  INV_X1 U10637 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9091) );
  MUX2_X1 U10638 ( .A(n9091), .B(n9090), .S(n10336), .Z(n9095) );
  NAND2_X1 U10639 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  OAI211_X1 U10640 ( .C1(n9097), .C2(n9096), .A(n9095), .B(n9094), .ZN(
        P2_U3429) );
  INV_X1 U10641 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9099) );
  MUX2_X1 U10642 ( .A(n9099), .B(n9098), .S(n10336), .Z(n9100) );
  OAI21_X1 U10643 ( .B1(n9102), .B2(n9101), .A(n9100), .ZN(P2_U3426) );
  INV_X1 U10644 ( .A(n10109), .ZN(n9107) );
  NOR4_X1 U10645 ( .A1(n5102), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9104), .A4(
        P2_U3151), .ZN(n9105) );
  AOI21_X1 U10646 ( .B1(n9115), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9105), .ZN(
        n9106) );
  OAI21_X1 U10647 ( .B1(n9107), .B2(n9123), .A(n9106), .ZN(P2_U3264) );
  OAI222_X1 U10648 ( .A1(n9121), .A2(n10636), .B1(n9123), .B2(n9109), .C1(
        n9108), .C2(P2_U3151), .ZN(P2_U3266) );
  AOI21_X1 U10649 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9115), .A(n9110), .ZN(
        n9111) );
  OAI21_X1 U10650 ( .B1(n9112), .B2(n9123), .A(n9111), .ZN(P2_U3267) );
  INV_X1 U10651 ( .A(n9113), .ZN(n10111) );
  AOI21_X1 U10652 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9115), .A(n9114), .ZN(
        n9116) );
  OAI21_X1 U10653 ( .B1(n10111), .B2(n9123), .A(n9116), .ZN(P2_U3268) );
  INV_X1 U10654 ( .A(n9117), .ZN(n10114) );
  OAI222_X1 U10655 ( .A1(P2_U3151), .A2(n9119), .B1(n9123), .B2(n10114), .C1(
        n9118), .C2(n9121), .ZN(P2_U3269) );
  INV_X1 U10656 ( .A(n9120), .ZN(n10117) );
  OAI222_X1 U10657 ( .A1(P2_U3151), .A2(n9124), .B1(n9123), .B2(n10117), .C1(
        n9122), .C2(n9121), .ZN(P2_U3270) );
  MUX2_X1 U10658 ( .A(n9125), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10659 ( .A(n10042), .ZN(n9900) );
  INV_X1 U10660 ( .A(n9126), .ZN(n9130) );
  NAND2_X1 U10661 ( .A1(n9129), .A2(n9130), .ZN(n9221) );
  OAI21_X1 U10662 ( .B1(n9130), .B2(n9129), .A(n9221), .ZN(n9131) );
  NAND2_X1 U10663 ( .A1(n9131), .A2(n9320), .ZN(n9135) );
  NAND2_X1 U10664 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10149)
         );
  OAI21_X1 U10665 ( .B1(n9324), .B2(n10058), .A(n10149), .ZN(n9133) );
  NOR2_X1 U10666 ( .A1(n9303), .A2(n9892), .ZN(n9132) );
  AOI211_X1 U10667 ( .C1(n9326), .C2(n10023), .A(n9133), .B(n9132), .ZN(n9134)
         );
  OAI211_X1 U10668 ( .C1(n9900), .C2(n9335), .A(n9135), .B(n9134), .ZN(
        P1_U3215) );
  INV_X1 U10669 ( .A(n9136), .ZN(n9138) );
  NAND2_X1 U10670 ( .A1(n9138), .A2(n9137), .ZN(n9288) );
  NAND2_X1 U10671 ( .A1(n9288), .A2(n9286), .ZN(n9285) );
  NAND2_X1 U10672 ( .A1(n9136), .A2(n9139), .ZN(n9287) );
  AOI21_X1 U10673 ( .B1(n9285), .B2(n9287), .A(n9141), .ZN(n9242) );
  AND3_X1 U10674 ( .A1(n9285), .A2(n9287), .A3(n9141), .ZN(n9142) );
  OAI21_X1 U10675 ( .B1(n9242), .B2(n9142), .A(n9320), .ZN(n9147) );
  INV_X1 U10676 ( .A(n9747), .ZN(n9144) );
  AOI22_X1 U10677 ( .A1(n9973), .A2(n9332), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9143) );
  OAI21_X1 U10678 ( .B1(n9303), .B2(n9144), .A(n9143), .ZN(n9145) );
  AOI21_X1 U10679 ( .B1(n9974), .B2(n9326), .A(n9145), .ZN(n9146) );
  OAI211_X1 U10680 ( .C1(n9977), .C2(n9335), .A(n9147), .B(n9146), .ZN(
        P1_U3216) );
  INV_X1 U10681 ( .A(n9148), .ZN(n9298) );
  AOI21_X1 U10682 ( .B1(n9150), .B2(n9149), .A(n9298), .ZN(n9159) );
  OAI21_X1 U10683 ( .B1(n9324), .B2(n9152), .A(n9151), .ZN(n9153) );
  AOI21_X1 U10684 ( .B1(n9326), .B2(n10054), .A(n9153), .ZN(n9154) );
  OAI21_X1 U10685 ( .B1(n9303), .B2(n9155), .A(n9154), .ZN(n9156) );
  AOI21_X1 U10686 ( .B1(n9157), .B2(n9272), .A(n9156), .ZN(n9158) );
  OAI21_X1 U10687 ( .B1(n9159), .B2(n9340), .A(n9158), .ZN(P1_U3217) );
  XNOR2_X1 U10688 ( .A(n4598), .B(n9161), .ZN(n9310) );
  NOR2_X1 U10689 ( .A1(n9310), .A2(n9311), .ZN(n9309) );
  AOI21_X1 U10690 ( .B1(n4598), .B2(n9161), .A(n9309), .ZN(n9165) );
  XNOR2_X1 U10691 ( .A(n9163), .B(n9162), .ZN(n9164) );
  XNOR2_X1 U10692 ( .A(n9165), .B(n9164), .ZN(n9170) );
  NAND2_X1 U10693 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9609) );
  OAI21_X1 U10694 ( .B1(n9233), .B2(n9324), .A(n9609), .ZN(n9166) );
  AOI21_X1 U10695 ( .B1(n9779), .B2(n9326), .A(n9166), .ZN(n9167) );
  OAI21_X1 U10696 ( .B1(n9303), .B2(n9813), .A(n9167), .ZN(n9168) );
  AOI21_X1 U10697 ( .B1(n10009), .B2(n9272), .A(n9168), .ZN(n9169) );
  OAI21_X1 U10698 ( .B1(n9170), .B2(n9340), .A(n9169), .ZN(P1_U3219) );
  NAND2_X1 U10699 ( .A1(n4523), .A2(n9171), .ZN(n9249) );
  OAI21_X1 U10700 ( .B1(n4523), .B2(n9171), .A(n9249), .ZN(n9172) );
  NOR2_X1 U10701 ( .A1(n9172), .A2(n9173), .ZN(n9252) );
  AOI21_X1 U10702 ( .B1(n9173), .B2(n9172), .A(n9252), .ZN(n9185) );
  INV_X1 U10703 ( .A(n9174), .ZN(n9175) );
  AOI21_X1 U10704 ( .B1(n9332), .B2(n9591), .A(n9175), .ZN(n9181) );
  INV_X1 U10705 ( .A(n9176), .ZN(n9177) );
  NAND2_X1 U10706 ( .A1(n9338), .A2(n9177), .ZN(n9180) );
  NAND2_X1 U10707 ( .A1(n9178), .A2(n9326), .ZN(n9179) );
  NAND3_X1 U10708 ( .A1(n9181), .A2(n9180), .A3(n9179), .ZN(n9182) );
  AOI21_X1 U10709 ( .B1(n9183), .B2(n9272), .A(n9182), .ZN(n9184) );
  OAI21_X1 U10710 ( .B1(n9185), .B2(n9340), .A(n9184), .ZN(P1_U3221) );
  XOR2_X1 U10711 ( .A(n9187), .B(n9186), .Z(n9192) );
  OAI22_X1 U10712 ( .A1(n9992), .A2(n9324), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10647), .ZN(n9188) );
  AOI21_X1 U10713 ( .B1(n9973), .B2(n9326), .A(n9188), .ZN(n9189) );
  OAI21_X1 U10714 ( .B1(n9303), .B2(n9777), .A(n9189), .ZN(n9190) );
  AOI21_X1 U10715 ( .B1(n9996), .B2(n9272), .A(n9190), .ZN(n9191) );
  OAI21_X1 U10716 ( .B1(n9192), .B2(n9340), .A(n9191), .ZN(P1_U3223) );
  INV_X1 U10717 ( .A(n4415), .ZN(n9299) );
  INV_X1 U10718 ( .A(n9194), .ZN(n9196) );
  NOR3_X1 U10719 ( .A1(n9299), .A2(n9196), .A3(n9195), .ZN(n9199) );
  INV_X1 U10720 ( .A(n9197), .ZN(n9198) );
  OAI21_X1 U10721 ( .B1(n9199), .B2(n9198), .A(n9320), .ZN(n9207) );
  INV_X1 U10722 ( .A(n9200), .ZN(n9205) );
  NAND2_X1 U10723 ( .A1(n9897), .A2(n9326), .ZN(n9202) );
  OAI211_X1 U10724 ( .C1(n9203), .C2(n9324), .A(n9202), .B(n9201), .ZN(n9204)
         );
  AOI21_X1 U10725 ( .B1(n9205), .B2(n9338), .A(n9204), .ZN(n9206) );
  OAI211_X1 U10726 ( .C1(n5061), .C2(n9335), .A(n9207), .B(n9206), .ZN(
        P1_U3224) );
  AOI21_X1 U10727 ( .B1(n9210), .B2(n9209), .A(n9208), .ZN(n9216) );
  INV_X1 U10728 ( .A(n9714), .ZN(n9211) );
  AOI22_X1 U10729 ( .A1(n9211), .A2(n9338), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9213) );
  NAND2_X1 U10730 ( .A1(n9974), .A2(n9332), .ZN(n9212) );
  OAI211_X1 U10731 ( .C1(n9946), .C2(n9334), .A(n9213), .B(n9212), .ZN(n9214)
         );
  AOI21_X1 U10732 ( .B1(n9961), .B2(n9272), .A(n9214), .ZN(n9215) );
  OAI21_X1 U10733 ( .B1(n9216), .B2(n9340), .A(n9215), .ZN(P1_U3225) );
  NAND2_X1 U10734 ( .A1(n9218), .A2(n9217), .ZN(n9225) );
  INV_X1 U10735 ( .A(n9219), .ZN(n9220) );
  NAND2_X1 U10736 ( .A1(n9223), .A2(n9222), .ZN(n9224) );
  OAI21_X1 U10737 ( .B1(n9223), .B2(n9222), .A(n9224), .ZN(n9330) );
  NOR2_X1 U10738 ( .A1(n9330), .A2(n9331), .ZN(n9329) );
  AND2_X1 U10739 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10168) );
  AOI21_X1 U10740 ( .B1(n10024), .B2(n9326), .A(n10168), .ZN(n9227) );
  NAND2_X1 U10741 ( .A1(n9338), .A2(n9858), .ZN(n9226) );
  OAI211_X1 U10742 ( .C1(n10039), .C2(n9324), .A(n9227), .B(n9226), .ZN(n9228)
         );
  AOI21_X1 U10743 ( .B1(n9866), .B2(n9272), .A(n9228), .ZN(n9229) );
  OAI21_X1 U10744 ( .B1(n9230), .B2(n9340), .A(n9229), .ZN(P1_U3226) );
  XOR2_X1 U10745 ( .A(n9232), .B(n9231), .Z(n9238) );
  NAND2_X1 U10746 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10186)
         );
  OAI21_X1 U10747 ( .B1(n9233), .B2(n9334), .A(n10186), .ZN(n9234) );
  AOI21_X1 U10748 ( .B1(n9332), .B2(n9587), .A(n9234), .ZN(n9235) );
  OAI21_X1 U10749 ( .B1(n9303), .B2(n9848), .A(n9235), .ZN(n9236) );
  AOI21_X1 U10750 ( .B1(n10020), .B2(n9272), .A(n9236), .ZN(n9237) );
  OAI21_X1 U10751 ( .B1(n9238), .B2(n9340), .A(n9237), .ZN(P1_U3228) );
  INV_X1 U10752 ( .A(n4426), .ZN(n9969) );
  INV_X1 U10753 ( .A(n9239), .ZN(n9240) );
  NOR3_X1 U10754 ( .A1(n9242), .A2(n9241), .A3(n9240), .ZN(n9244) );
  OAI21_X1 U10755 ( .B1(n9244), .B2(n9243), .A(n9320), .ZN(n9248) );
  AOI22_X1 U10756 ( .A1(n9728), .A2(n9338), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9245) );
  OAI21_X1 U10757 ( .B1(n9953), .B2(n9334), .A(n9245), .ZN(n9246) );
  AOI21_X1 U10758 ( .B1(n9332), .B2(n9983), .A(n9246), .ZN(n9247) );
  OAI211_X1 U10759 ( .C1(n9969), .C2(n9335), .A(n9248), .B(n9247), .ZN(
        P1_U3229) );
  INV_X1 U10760 ( .A(n9249), .ZN(n9251) );
  NOR3_X1 U10761 ( .A1(n9252), .A2(n9251), .A3(n9250), .ZN(n9255) );
  INV_X1 U10762 ( .A(n9253), .ZN(n9254) );
  OAI21_X1 U10763 ( .B1(n9255), .B2(n9254), .A(n9320), .ZN(n9262) );
  OAI21_X1 U10764 ( .B1(n9324), .B2(n9257), .A(n9256), .ZN(n9260) );
  NOR2_X1 U10765 ( .A1(n9303), .A2(n9258), .ZN(n9259) );
  AOI211_X1 U10766 ( .C1(n9326), .C2(n9590), .A(n9260), .B(n9259), .ZN(n9261)
         );
  OAI211_X1 U10767 ( .C1(n9263), .C2(n9335), .A(n9262), .B(n9261), .ZN(
        P1_U3231) );
  INV_X1 U10768 ( .A(n9264), .ZN(n9266) );
  NOR2_X1 U10769 ( .A1(n9266), .A2(n9265), .ZN(n9267) );
  XNOR2_X1 U10770 ( .A(n9268), .B(n9267), .ZN(n9275) );
  OAI22_X1 U10771 ( .A1(n9822), .A2(n9324), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9269), .ZN(n9271) );
  NOR2_X1 U10772 ( .A1(n9792), .A2(n9334), .ZN(n9270) );
  AOI211_X1 U10773 ( .C1(n9797), .C2(n9338), .A(n9271), .B(n9270), .ZN(n9274)
         );
  NAND2_X1 U10774 ( .A1(n10001), .A2(n9272), .ZN(n9273) );
  OAI211_X1 U10775 ( .C1(n9275), .C2(n9340), .A(n9274), .B(n9273), .ZN(
        P1_U3233) );
  OAI21_X1 U10776 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(n9279) );
  NAND2_X1 U10777 ( .A1(n9279), .A2(n9320), .ZN(n9283) );
  NAND2_X1 U10778 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10137)
         );
  OAI21_X1 U10779 ( .B1(n9324), .B2(n9911), .A(n10137), .ZN(n9281) );
  NOR2_X1 U10780 ( .A1(n9303), .A2(n9922), .ZN(n9280) );
  AOI211_X1 U10781 ( .C1(n9326), .C2(n9588), .A(n9281), .B(n9280), .ZN(n9282)
         );
  OAI211_X1 U10782 ( .C1(n7076), .C2(n9335), .A(n9283), .B(n9282), .ZN(
        P1_U3234) );
  INV_X1 U10783 ( .A(n9287), .ZN(n9284) );
  NOR2_X1 U10784 ( .A1(n9285), .A2(n9284), .ZN(n9290) );
  AOI21_X1 U10785 ( .B1(n9288), .B2(n9287), .A(n9286), .ZN(n9289) );
  OAI21_X1 U10786 ( .B1(n9290), .B2(n9289), .A(n9320), .ZN(n9294) );
  AOI22_X1 U10787 ( .A1(n9982), .A2(n9332), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9291) );
  OAI21_X1 U10788 ( .B1(n9303), .B2(n9765), .A(n9291), .ZN(n9292) );
  AOI21_X1 U10789 ( .B1(n9326), .B2(n9983), .A(n9292), .ZN(n9293) );
  OAI211_X1 U10790 ( .C1(n9985), .C2(n9335), .A(n9294), .B(n9293), .ZN(
        P1_U3235) );
  INV_X1 U10791 ( .A(n9295), .ZN(n9297) );
  NOR3_X1 U10792 ( .A1(n9298), .A2(n9297), .A3(n9296), .ZN(n9300) );
  OAI21_X1 U10793 ( .B1(n9300), .B2(n9299), .A(n9320), .ZN(n9307) );
  OAI21_X1 U10794 ( .B1(n9334), .B2(n9911), .A(n9301), .ZN(n9305) );
  NOR2_X1 U10795 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  AOI211_X1 U10796 ( .C1(n9332), .C2(n9590), .A(n9305), .B(n9304), .ZN(n9306)
         );
  OAI211_X1 U10797 ( .C1(n9308), .C2(n9335), .A(n9307), .B(n9306), .ZN(
        P1_U3236) );
  AOI21_X1 U10798 ( .B1(n9311), .B2(n9310), .A(n9309), .ZN(n9316) );
  NAND2_X1 U10799 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10204)
         );
  NAND2_X1 U10800 ( .A1(n10024), .A2(n9332), .ZN(n9312) );
  OAI211_X1 U10801 ( .C1(n9822), .C2(n9334), .A(n10204), .B(n9312), .ZN(n9314)
         );
  NOR2_X1 U10802 ( .A1(n9831), .A2(n9335), .ZN(n9313) );
  AOI211_X1 U10803 ( .C1(n9828), .C2(n9338), .A(n9314), .B(n9313), .ZN(n9315)
         );
  OAI21_X1 U10804 ( .B1(n9316), .B2(n9340), .A(n9315), .ZN(P1_U3238) );
  INV_X1 U10805 ( .A(n9959), .ZN(n10074) );
  OAI21_X1 U10806 ( .B1(n9208), .B2(n9318), .A(n9317), .ZN(n9319) );
  NAND3_X1 U10807 ( .A1(n9321), .A2(n9320), .A3(n9319), .ZN(n9328) );
  INV_X1 U10808 ( .A(n9699), .ZN(n9322) );
  AOI22_X1 U10809 ( .A1(n9322), .A2(n9338), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9323) );
  OAI21_X1 U10810 ( .B1(n9953), .B2(n9324), .A(n9323), .ZN(n9325) );
  AOI21_X1 U10811 ( .B1(n9669), .B2(n9326), .A(n9325), .ZN(n9327) );
  OAI211_X1 U10812 ( .C1(n10074), .C2(n9335), .A(n9328), .B(n9327), .ZN(
        P1_U3240) );
  AOI21_X1 U10813 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9341) );
  NAND2_X1 U10814 ( .A1(n9332), .A2(n9588), .ZN(n9333) );
  NAND2_X1 U10815 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10161)
         );
  OAI211_X1 U10816 ( .C1(n9881), .C2(n9334), .A(n9333), .B(n10161), .ZN(n9337)
         );
  NOR2_X1 U10817 ( .A1(n9877), .A2(n9335), .ZN(n9336) );
  AOI211_X1 U10818 ( .C1(n9875), .C2(n9338), .A(n9337), .B(n9336), .ZN(n9339)
         );
  OAI21_X1 U10819 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(P1_U3241) );
  NOR2_X1 U10820 ( .A1(n9509), .A2(n9629), .ZN(n9446) );
  NAND2_X1 U10821 ( .A1(n9345), .A2(n9344), .ZN(n9358) );
  NAND3_X1 U10822 ( .A1(n9358), .A2(n9346), .A3(n9533), .ZN(n9348) );
  AND2_X1 U10823 ( .A1(n9347), .A2(n9537), .ZN(n9356) );
  NAND2_X1 U10824 ( .A1(n9348), .A2(n9356), .ZN(n9349) );
  INV_X1 U10825 ( .A(n9350), .ZN(n9355) );
  INV_X1 U10826 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U10827 ( .A1(n9353), .A2(n9352), .ZN(n9354) );
  INV_X1 U10828 ( .A(n9533), .ZN(n9357) );
  NAND3_X1 U10829 ( .A1(n9361), .A2(n9360), .A3(n9359), .ZN(n9363) );
  NAND2_X1 U10830 ( .A1(n9366), .A2(n9373), .ZN(n9367) );
  OAI211_X1 U10831 ( .C1(n9368), .C2(n9367), .A(n9380), .B(n9376), .ZN(n9369)
         );
  NAND3_X1 U10832 ( .A1(n9369), .A2(n9449), .A3(n9370), .ZN(n9386) );
  INV_X1 U10833 ( .A(n9370), .ZN(n9372) );
  NOR2_X1 U10834 ( .A1(n9372), .A2(n9371), .ZN(n9379) );
  NAND2_X1 U10835 ( .A1(n9379), .A2(n9373), .ZN(n9539) );
  AOI21_X1 U10836 ( .B1(n9375), .B2(n9374), .A(n9539), .ZN(n9383) );
  INV_X1 U10837 ( .A(n9376), .ZN(n9378) );
  NOR2_X1 U10838 ( .A1(n9378), .A2(n9377), .ZN(n9382) );
  INV_X1 U10839 ( .A(n9379), .ZN(n9381) );
  OAI21_X1 U10840 ( .B1(n9382), .B2(n9381), .A(n9380), .ZN(n9542) );
  NOR2_X1 U10841 ( .A1(n9383), .A2(n9542), .ZN(n9384) );
  NAND2_X1 U10842 ( .A1(n9384), .A2(n9342), .ZN(n9385) );
  INV_X1 U10843 ( .A(n9387), .ZN(n9902) );
  OAI211_X1 U10844 ( .C1(n9390), .C2(n9902), .A(n9462), .B(n9543), .ZN(n9388)
         );
  AND2_X1 U10845 ( .A1(n9397), .A2(n9393), .ZN(n9525) );
  OAI21_X1 U10846 ( .B1(n9390), .B2(n9389), .A(n9550), .ZN(n9396) );
  NAND2_X1 U10847 ( .A1(n9838), .A2(n9391), .ZN(n9398) );
  INV_X1 U10848 ( .A(n9462), .ZN(n9392) );
  NOR2_X1 U10849 ( .A1(n9398), .A2(n9392), .ZN(n9547) );
  INV_X1 U10850 ( .A(n9838), .ZN(n9394) );
  OAI21_X1 U10851 ( .B1(n9394), .B2(n9393), .A(n9397), .ZN(n9395) );
  INV_X1 U10852 ( .A(n9840), .ZN(n9836) );
  NAND2_X1 U10853 ( .A1(n9410), .A2(n9399), .ZN(n9552) );
  NOR2_X1 U10854 ( .A1(n9413), .A2(n9552), .ZN(n9417) );
  NAND2_X1 U10855 ( .A1(n9402), .A2(n9401), .ZN(n9400) );
  INV_X1 U10856 ( .A(n9400), .ZN(n9492) );
  NAND4_X1 U10857 ( .A1(n9492), .A2(n9449), .A3(n9561), .A4(n9409), .ZN(n9416)
         );
  OR2_X1 U10858 ( .A1(n9996), .A2(n9792), .ZN(n9487) );
  NAND2_X1 U10859 ( .A1(n9487), .A2(n9403), .ZN(n9501) );
  NAND3_X1 U10860 ( .A1(n9501), .A2(n9342), .A3(n9402), .ZN(n9407) );
  NAND3_X1 U10861 ( .A1(n9400), .A2(n9449), .A3(n9487), .ZN(n9406) );
  NAND4_X1 U10862 ( .A1(n9402), .A2(n9342), .A3(n9401), .A4(n9561), .ZN(n9405)
         );
  NAND4_X1 U10863 ( .A1(n9487), .A2(n9449), .A3(n9403), .A4(n9411), .ZN(n9404)
         );
  NAND4_X1 U10864 ( .A1(n9407), .A2(n9406), .A3(n9405), .A4(n9404), .ZN(n9415)
         );
  NAND2_X1 U10865 ( .A1(n10020), .A2(n9861), .ZN(n9408) );
  NAND2_X1 U10866 ( .A1(n9409), .A2(n9408), .ZN(n9556) );
  NAND2_X1 U10867 ( .A1(n9411), .A2(n9410), .ZN(n9554) );
  NOR3_X1 U10868 ( .A1(n9501), .A2(n9449), .A3(n9554), .ZN(n9412) );
  NAND2_X1 U10869 ( .A1(n9480), .A2(n9419), .ZN(n9488) );
  OR2_X1 U10870 ( .A1(n9763), .A2(n9993), .ZN(n9420) );
  NAND2_X1 U10871 ( .A1(n9421), .A2(n9420), .ZN(n9481) );
  MUX2_X1 U10872 ( .A(n9488), .B(n9481), .S(n9449), .Z(n9423) );
  MUX2_X1 U10873 ( .A(n9421), .B(n9480), .S(n9449), .Z(n9422) );
  INV_X1 U10874 ( .A(n9486), .ZN(n9425) );
  AND2_X1 U10875 ( .A1(n9434), .A2(n9431), .ZN(n9493) );
  NAND2_X1 U10876 ( .A1(n9427), .A2(n9426), .ZN(n9433) );
  OAI211_X1 U10877 ( .C1(n9432), .C2(n4734), .A(n9497), .B(n9486), .ZN(n9435)
         );
  INV_X1 U10878 ( .A(n9433), .ZN(n9499) );
  MUX2_X1 U10879 ( .A(n9505), .B(n9507), .S(n9449), .Z(n9436) );
  AOI21_X1 U10880 ( .B1(n9509), .B2(n9585), .A(n9567), .ZN(n9440) );
  INV_X1 U10881 ( .A(n9585), .ZN(n9476) );
  OR2_X1 U10882 ( .A1(n9945), .A2(n9476), .ZN(n9510) );
  OAI211_X1 U10883 ( .C1(n9449), .C2(n9510), .A(n9442), .B(n9509), .ZN(n9443)
         );
  NOR3_X1 U10884 ( .A1(n9575), .A2(n9521), .A3(n9447), .ZN(n9448) );
  OAI21_X1 U10885 ( .B1(n9516), .B2(n9629), .A(n9448), .ZN(n9583) );
  NAND2_X1 U10886 ( .A1(n9522), .A2(n9635), .ZN(n9573) );
  AOI211_X1 U10887 ( .C1(n9451), .C2(n9449), .A(n9573), .B(n9575), .ZN(n9478)
         );
  NOR2_X1 U10888 ( .A1(n10067), .A2(n9509), .ZN(n9514) );
  INV_X1 U10889 ( .A(n9510), .ZN(n9450) );
  NOR2_X1 U10890 ( .A1(n9514), .A2(n9450), .ZN(n9569) );
  INV_X1 U10891 ( .A(n9552), .ZN(n9471) );
  NOR4_X1 U10892 ( .A1(n9461), .A2(n9460), .A3(n9459), .A4(n9458), .ZN(n9467)
         );
  INV_X1 U10893 ( .A(n9916), .ZN(n9466) );
  INV_X1 U10894 ( .A(n9464), .ZN(n9465) );
  NAND4_X1 U10895 ( .A1(n9467), .A2(n9466), .A3(n9903), .A4(n9465), .ZN(n9468)
         );
  NAND4_X1 U10896 ( .A1(n9789), .A2(n9471), .A3(n9806), .A4(n9470), .ZN(n9472)
         );
  NAND4_X1 U10897 ( .A1(n9693), .A2(n9736), .A3(n7070), .A4(n9473), .ZN(n9474)
         );
  NAND2_X1 U10898 ( .A1(n9945), .A2(n9476), .ZN(n9508) );
  NAND4_X1 U10899 ( .A1(n9477), .A2(n9569), .A3(n9516), .A4(n9508), .ZN(n9523)
         );
  NAND2_X1 U10900 ( .A1(n9481), .A2(n9480), .ZN(n9482) );
  NAND2_X1 U10901 ( .A1(n9483), .A2(n9482), .ZN(n9484) );
  NAND2_X1 U10902 ( .A1(n9484), .A2(n9490), .ZN(n9485) );
  NAND2_X1 U10903 ( .A1(n9486), .A2(n9485), .ZN(n9502) );
  INV_X1 U10904 ( .A(n9502), .ZN(n9496) );
  INV_X1 U10905 ( .A(n9487), .ZN(n9491) );
  INV_X1 U10906 ( .A(n9488), .ZN(n9489) );
  OAI211_X1 U10907 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9495)
         );
  INV_X1 U10908 ( .A(n9493), .ZN(n9494) );
  AOI21_X1 U10909 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9500) );
  NAND2_X1 U10910 ( .A1(n9498), .A2(n9497), .ZN(n9558) );
  OAI21_X1 U10911 ( .B1(n9500), .B2(n9558), .A(n9499), .ZN(n9562) );
  OR2_X1 U10912 ( .A1(n9502), .A2(n9501), .ZN(n9559) );
  NOR3_X1 U10913 ( .A1(n9558), .A2(n9788), .A3(n9559), .ZN(n9503) );
  NOR2_X1 U10914 ( .A1(n9562), .A2(n9503), .ZN(n9506) );
  NAND2_X1 U10915 ( .A1(n9505), .A2(n9504), .ZN(n9565) );
  OAI22_X1 U10916 ( .A1(n9506), .A2(n9565), .B1(n5034), .B2(n9509), .ZN(n9513)
         );
  AND2_X1 U10917 ( .A1(n9508), .A2(n9507), .ZN(n9564) );
  INV_X1 U10918 ( .A(n9564), .ZN(n9512) );
  INV_X1 U10919 ( .A(n9509), .ZN(n9511) );
  OAI22_X1 U10920 ( .A1(n9513), .A2(n9512), .B1(n9511), .B2(n9510), .ZN(n9517)
         );
  AOI211_X1 U10921 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9580)
         );
  NAND2_X1 U10922 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  OAI211_X1 U10923 ( .C1(n9521), .C2(n9575), .A(n9520), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9574) );
  NAND3_X1 U10924 ( .A1(n9523), .A2(n9522), .A3(n9574), .ZN(n9579) );
  NAND2_X1 U10925 ( .A1(n9574), .A2(n9635), .ZN(n9572) );
  NAND2_X1 U10926 ( .A1(n9574), .A2(n9524), .ZN(n9571) );
  INV_X1 U10927 ( .A(n9525), .ZN(n9553) );
  INV_X1 U10928 ( .A(n7658), .ZN(n9534) );
  AOI21_X1 U10929 ( .B1(n7073), .B2(n6400), .A(n9526), .ZN(n9531) );
  NAND4_X1 U10930 ( .A1(n9531), .A2(n9530), .A3(n9529), .A4(n9528), .ZN(n9532)
         );
  NAND3_X1 U10931 ( .A1(n9534), .A2(n9533), .A3(n9532), .ZN(n9538) );
  INV_X1 U10932 ( .A(n9535), .ZN(n9536) );
  AOI21_X1 U10933 ( .B1(n9538), .B2(n9537), .A(n9536), .ZN(n9546) );
  INV_X1 U10934 ( .A(n9539), .ZN(n9541) );
  NAND2_X1 U10935 ( .A1(n9541), .A2(n9540), .ZN(n9545) );
  INV_X1 U10936 ( .A(n9542), .ZN(n9544) );
  OAI211_X1 U10937 ( .C1(n9546), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9549)
         );
  INV_X1 U10938 ( .A(n9547), .ZN(n9548) );
  AOI21_X1 U10939 ( .B1(n9550), .B2(n9549), .A(n9548), .ZN(n9551) );
  AOI211_X1 U10940 ( .C1(n9838), .C2(n9553), .A(n9552), .B(n9551), .ZN(n9557)
         );
  INV_X1 U10941 ( .A(n9554), .ZN(n9555) );
  OAI21_X1 U10942 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n9560) );
  AOI211_X1 U10943 ( .C1(n9561), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9563)
         );
  NOR2_X1 U10944 ( .A1(n9563), .A2(n9562), .ZN(n9566) );
  OAI21_X1 U10945 ( .B1(n9566), .B2(n9565), .A(n9564), .ZN(n9568) );
  AOI21_X1 U10946 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9570) );
  MUX2_X1 U10947 ( .A(n9572), .B(n9571), .S(n9570), .Z(n9578) );
  INV_X1 U10948 ( .A(n9573), .ZN(n9576) );
  OAI21_X1 U10949 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9577) );
  OAI211_X1 U10950 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9577), .ZN(n9581)
         );
  OAI211_X1 U10951 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9581), .ZN(
        P1_U3242) );
  MUX2_X1 U10952 ( .A(n9585), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9596), .Z(
        P1_U3584) );
  MUX2_X1 U10953 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9657), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10954 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9669), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10955 ( .A(n9712), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9596), .Z(
        P1_U3580) );
  MUX2_X1 U10956 ( .A(n9701), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9596), .Z(
        P1_U3579) );
  MUX2_X1 U10957 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9974), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10958 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9983), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10959 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9973), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10960 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9982), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10961 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9779), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10962 ( .A(n9586), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9596), .Z(
        P1_U3573) );
  MUX2_X1 U10963 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9842), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10964 ( .A(n10024), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9596), .Z(
        P1_U3571) );
  MUX2_X1 U10965 ( .A(n9587), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9596), .Z(
        P1_U3570) );
  MUX2_X1 U10966 ( .A(n10023), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9596), .Z(
        P1_U3569) );
  MUX2_X1 U10967 ( .A(n9588), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9596), .Z(
        P1_U3568) );
  MUX2_X1 U10968 ( .A(n9897), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9596), .Z(
        P1_U3567) );
  MUX2_X1 U10969 ( .A(n9589), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9596), .Z(
        P1_U3566) );
  MUX2_X1 U10970 ( .A(n10054), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9596), .Z(
        P1_U3565) );
  MUX2_X1 U10971 ( .A(n9590), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9596), .Z(
        P1_U3564) );
  MUX2_X1 U10972 ( .A(n9591), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9596), .Z(
        P1_U3561) );
  MUX2_X1 U10973 ( .A(n9592), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9596), .Z(
        P1_U3560) );
  MUX2_X1 U10974 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9593), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10975 ( .A(n9594), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9596), .Z(
        P1_U3558) );
  MUX2_X1 U10976 ( .A(n9595), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9596), .Z(
        P1_U3557) );
  MUX2_X1 U10977 ( .A(n7009), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9596), .Z(
        P1_U3556) );
  OAI211_X1 U10978 ( .C1(n9599), .C2(n9598), .A(n10193), .B(n9597), .ZN(n9608)
         );
  OAI211_X1 U10979 ( .C1(n9602), .C2(n9601), .A(n10198), .B(n9600), .ZN(n9607)
         );
  AOI22_X1 U10980 ( .A1(n10169), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9606) );
  NAND2_X1 U10981 ( .A1(n10183), .A2(n9604), .ZN(n9605) );
  NAND4_X1 U10982 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(
        P1_U3244) );
  INV_X1 U10983 ( .A(n9609), .ZN(n9638) );
  NOR2_X1 U10984 ( .A1(n10184), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9614) );
  AOI21_X1 U10985 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10184), .A(n9614), .ZN(
        n10177) );
  XNOR2_X1 U10986 ( .A(n10136), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U10987 ( .A1(n10148), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9611) );
  OAI21_X1 U10988 ( .B1(n10148), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9611), .ZN(
        n10141) );
  XNOR2_X1 U10989 ( .A(n9621), .B(n9612), .ZN(n10157) );
  NAND2_X1 U10990 ( .A1(n10172), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9613) );
  OAI21_X1 U10991 ( .B1(n10172), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9613), .ZN(
        n10166) );
  NAND2_X1 U10992 ( .A1(n10177), .A2(n10178), .ZN(n10176) );
  NAND2_X1 U10993 ( .A1(n9625), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9616) );
  OAI21_X1 U10994 ( .B1(n9625), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9616), .ZN(
        n10190) );
  XNOR2_X1 U10995 ( .A(n9617), .B(n9812), .ZN(n9632) );
  INV_X1 U10996 ( .A(n9632), .ZN(n9628) );
  OR2_X1 U10997 ( .A1(n10184), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9624) );
  AOI22_X1 U10998 ( .A1(n10172), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n10030), 
        .B2(n9618), .ZN(n10171) );
  OAI21_X1 U10999 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9620), .A(n9619), .ZN(
        n10129) );
  XNOR2_X1 U11000 ( .A(n10136), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10130) );
  XNOR2_X1 U11001 ( .A(n10148), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10144) );
  XOR2_X1 U11002 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10184), .Z(n10180) );
  NAND2_X1 U11003 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U11004 ( .A1(n9624), .A2(n10179), .ZN(n10194) );
  NAND2_X1 U11005 ( .A1(n9625), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9626) );
  OAI21_X1 U11006 ( .B1(n9625), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9626), .ZN(
        n10195) );
  NAND2_X1 U11007 ( .A1(n10197), .A2(n9626), .ZN(n9627) );
  XNOR2_X1 U11008 ( .A(n9627), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9631) );
  OAI22_X1 U11009 ( .A1(n9628), .A2(n10164), .B1(n10152), .B2(n9631), .ZN(
        n9630) );
  AOI21_X1 U11010 ( .B1(n10198), .B2(n9631), .A(n10183), .ZN(n9634) );
  NAND2_X1 U11011 ( .A1(n9634), .A2(n9633), .ZN(n9636) );
  NOR2_X1 U11012 ( .A1(n9863), .A2(n9920), .ZN(n9931) );
  NAND2_X1 U11013 ( .A1(n9639), .A2(n9931), .ZN(n9642) );
  INV_X1 U11014 ( .A(n9640), .ZN(n9941) );
  NOR2_X1 U11015 ( .A1(n9933), .A2(n9941), .ZN(n9645) );
  AOI21_X1 U11016 ( .B1(n9933), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9645), .ZN(
        n9641) );
  OAI211_X1 U11017 ( .C1(n10067), .C2(n9926), .A(n9642), .B(n9641), .ZN(
        P1_U3263) );
  NOR2_X1 U11018 ( .A1(n9854), .A2(n9644), .ZN(n9646) );
  AOI211_X1 U11019 ( .C1(n9945), .C2(n9930), .A(n9646), .B(n9645), .ZN(n9647)
         );
  OAI21_X1 U11020 ( .B1(n9942), .B2(n9863), .A(n9647), .ZN(P1_U3264) );
  NOR2_X1 U11021 ( .A1(n9652), .A2(n9863), .ZN(n9661) );
  NOR2_X1 U11022 ( .A1(n9653), .A2(n9891), .ZN(n9656) );
  MUX2_X1 U11023 ( .A(P1_REG2_REG_29__SCAN_IN), .B(n9654), .S(n9854), .Z(n9655) );
  AOI211_X1 U11024 ( .C1(n9657), .C2(n9898), .A(n9656), .B(n9655), .ZN(n9658)
         );
  OAI21_X1 U11025 ( .B1(n9659), .B2(n9926), .A(n9658), .ZN(n9660) );
  OAI21_X1 U11026 ( .B1(n9648), .B2(n9871), .A(n9664), .ZN(P1_U3356) );
  NAND2_X1 U11027 ( .A1(n9665), .A2(n9759), .ZN(n9677) );
  OAI22_X1 U11028 ( .A1(n9667), .A2(n9891), .B1(n9666), .B2(n9893), .ZN(n9668)
         );
  AOI21_X1 U11029 ( .B1(n9898), .B2(n9669), .A(n9668), .ZN(n9670) );
  OAI21_X1 U11030 ( .B1(n9671), .B2(n9894), .A(n9670), .ZN(n9674) );
  NOR2_X1 U11031 ( .A1(n9672), .A2(n9863), .ZN(n9673) );
  AOI211_X1 U11032 ( .C1(n9930), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  OAI211_X1 U11033 ( .C1(n9909), .C2(n9678), .A(n9677), .B(n9676), .ZN(
        P1_U3265) );
  XOR2_X1 U11034 ( .A(n9686), .B(n9679), .Z(n9951) );
  AOI211_X1 U11035 ( .C1(n9680), .C2(n4454), .A(n9920), .B(n7077), .ZN(n9949)
         );
  NOR2_X1 U11036 ( .A1(n10072), .A2(n9926), .ZN(n9685) );
  AOI22_X1 U11037 ( .A1(n9681), .A2(n9932), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9933), .ZN(n9683) );
  NAND2_X1 U11038 ( .A1(n9712), .A2(n9898), .ZN(n9682) );
  OAI211_X1 U11039 ( .C1(n9947), .C2(n9894), .A(n9683), .B(n9682), .ZN(n9684)
         );
  AOI211_X1 U11040 ( .C1(n9949), .C2(n9921), .A(n9685), .B(n9684), .ZN(n9689)
         );
  XNOR2_X1 U11041 ( .A(n9687), .B(n9686), .ZN(n9950) );
  NAND2_X1 U11042 ( .A1(n9950), .A2(n9928), .ZN(n9688) );
  OAI211_X1 U11043 ( .C1(n9951), .C2(n9871), .A(n9689), .B(n9688), .ZN(
        P1_U3266) );
  NAND2_X1 U11044 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  XNOR2_X1 U11045 ( .A(n9693), .B(n9692), .ZN(n9956) );
  INV_X1 U11046 ( .A(n9956), .ZN(n9707) );
  OR2_X1 U11047 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  NAND2_X1 U11048 ( .A1(n9696), .A2(n9695), .ZN(n9952) );
  AOI21_X1 U11049 ( .B1(n4469), .B2(n9959), .A(n9920), .ZN(n9697) );
  NAND2_X1 U11050 ( .A1(n4454), .A2(n9697), .ZN(n9957) );
  OAI22_X1 U11051 ( .A1(n9699), .A2(n9891), .B1(n9698), .B2(n9893), .ZN(n9700)
         );
  AOI21_X1 U11052 ( .B1(n9701), .B2(n9898), .A(n9700), .ZN(n9702) );
  OAI21_X1 U11053 ( .B1(n9954), .B2(n9894), .A(n9702), .ZN(n9703) );
  AOI21_X1 U11054 ( .B1(n9959), .B2(n9930), .A(n9703), .ZN(n9704) );
  OAI21_X1 U11055 ( .B1(n9957), .B2(n9863), .A(n9704), .ZN(n9705) );
  AOI21_X1 U11056 ( .B1(n9952), .B2(n9759), .A(n9705), .ZN(n9706) );
  OAI21_X1 U11057 ( .B1(n9909), .B2(n9707), .A(n9706), .ZN(P1_U3267) );
  XNOR2_X1 U11058 ( .A(n9708), .B(n9709), .ZN(n9965) );
  OAI22_X1 U11059 ( .A1(n9714), .A2(n9891), .B1(n9713), .B2(n9893), .ZN(n9715)
         );
  AOI21_X1 U11060 ( .B1(n9961), .B2(n9930), .A(n9715), .ZN(n9718) );
  NAND2_X1 U11061 ( .A1(n9731), .A2(n9961), .ZN(n9716) );
  NAND2_X1 U11062 ( .A1(n9962), .A2(n9931), .ZN(n9717) );
  OAI211_X1 U11063 ( .C1(n9964), .C2(n9933), .A(n9718), .B(n9717), .ZN(n9719)
         );
  INV_X1 U11064 ( .A(n9719), .ZN(n9720) );
  OAI21_X1 U11065 ( .B1(n9909), .B2(n9965), .A(n9720), .ZN(P1_U3268) );
  NAND2_X1 U11066 ( .A1(n9722), .A2(n9721), .ZN(n9723) );
  NAND3_X1 U11067 ( .A1(n9724), .A2(n9988), .A3(n9723), .ZN(n9727) );
  OAI22_X1 U11068 ( .A1(n9953), .A2(n10057), .B1(n9769), .B2(n10038), .ZN(
        n9725) );
  INV_X1 U11069 ( .A(n9725), .ZN(n9726) );
  NAND2_X1 U11070 ( .A1(n9727), .A2(n9726), .ZN(n9972) );
  INV_X1 U11071 ( .A(n9972), .ZN(n9740) );
  INV_X1 U11072 ( .A(n9728), .ZN(n9730) );
  OAI22_X1 U11073 ( .A1(n9730), .A2(n9891), .B1(n9729), .B2(n9854), .ZN(n9734)
         );
  AOI21_X1 U11074 ( .B1(n9744), .B2(n4426), .A(n9920), .ZN(n9732) );
  NAND2_X1 U11075 ( .A1(n9732), .A2(n9731), .ZN(n9968) );
  NOR2_X1 U11076 ( .A1(n9968), .A2(n9863), .ZN(n9733) );
  AOI211_X1 U11077 ( .C1(n9930), .C2(n4426), .A(n9734), .B(n9733), .ZN(n9739)
         );
  NAND2_X1 U11078 ( .A1(n9737), .A2(n9736), .ZN(n9966) );
  NAND3_X1 U11079 ( .A1(n9967), .A2(n9966), .A3(n9928), .ZN(n9738) );
  OAI211_X1 U11080 ( .C1(n9740), .C2(n9933), .A(n9739), .B(n9738), .ZN(
        P1_U3269) );
  XNOR2_X1 U11081 ( .A(n9741), .B(n4692), .ZN(n9981) );
  XNOR2_X1 U11082 ( .A(n9742), .B(n9743), .ZN(n9979) );
  OAI211_X1 U11083 ( .C1(n9761), .C2(n9977), .A(n10002), .B(n9744), .ZN(n9976)
         );
  NOR2_X1 U11084 ( .A1(n9854), .A2(n9745), .ZN(n9746) );
  AOI21_X1 U11085 ( .B1(n9973), .B2(n9898), .A(n9746), .ZN(n9749) );
  NAND2_X1 U11086 ( .A1(n9747), .A2(n9932), .ZN(n9748) );
  OAI211_X1 U11087 ( .C1(n9750), .C2(n9894), .A(n9749), .B(n9748), .ZN(n9751)
         );
  AOI21_X1 U11088 ( .B1(n4611), .B2(n9930), .A(n9751), .ZN(n9753) );
  OAI21_X1 U11089 ( .B1(n9976), .B2(n9863), .A(n9753), .ZN(n9754) );
  AOI21_X1 U11090 ( .B1(n9979), .B2(n9759), .A(n9754), .ZN(n9755) );
  OAI21_X1 U11091 ( .B1(n9909), .B2(n9981), .A(n9755), .ZN(P1_U3270) );
  XNOR2_X1 U11092 ( .A(n9756), .B(n4663), .ZN(n9991) );
  XNOR2_X1 U11093 ( .A(n9757), .B(n9758), .ZN(n9989) );
  NAND2_X1 U11094 ( .A1(n9989), .A2(n9759), .ZN(n9772) );
  OAI21_X1 U11095 ( .B1(n9760), .B2(n9985), .A(n10002), .ZN(n9762) );
  NOR2_X1 U11096 ( .A1(n9762), .A2(n9761), .ZN(n9987) );
  NAND2_X1 U11097 ( .A1(n9763), .A2(n9930), .ZN(n9768) );
  OAI22_X1 U11098 ( .A1(n9765), .A2(n9891), .B1(n9764), .B2(n9893), .ZN(n9766)
         );
  AOI21_X1 U11099 ( .B1(n9982), .B2(n9898), .A(n9766), .ZN(n9767) );
  OAI211_X1 U11100 ( .C1(n9769), .C2(n9894), .A(n9768), .B(n9767), .ZN(n9770)
         );
  AOI21_X1 U11101 ( .B1(n9987), .B2(n9921), .A(n9770), .ZN(n9771) );
  OAI211_X1 U11102 ( .C1(n9991), .C2(n9909), .A(n9772), .B(n9771), .ZN(
        P1_U3271) );
  INV_X1 U11103 ( .A(n9773), .ZN(n9774) );
  AOI21_X1 U11104 ( .B1(n9783), .B2(n9775), .A(n9774), .ZN(n10000) );
  AOI211_X1 U11105 ( .C1(n9996), .C2(n5175), .A(n9920), .B(n9760), .ZN(n9994)
         );
  NAND2_X1 U11106 ( .A1(n9996), .A2(n9930), .ZN(n9781) );
  OAI22_X1 U11107 ( .A1(n9777), .A2(n9891), .B1(n9776), .B2(n9893), .ZN(n9778)
         );
  AOI21_X1 U11108 ( .B1(n9898), .B2(n9779), .A(n9778), .ZN(n9780) );
  OAI211_X1 U11109 ( .C1(n9993), .C2(n9894), .A(n9781), .B(n9780), .ZN(n9782)
         );
  AOI21_X1 U11110 ( .B1(n9994), .B2(n9921), .A(n9782), .ZN(n9786) );
  XNOR2_X1 U11111 ( .A(n9784), .B(n9783), .ZN(n9997) );
  NAND2_X1 U11112 ( .A1(n9997), .A2(n9928), .ZN(n9785) );
  OAI211_X1 U11113 ( .C1(n10000), .C2(n9871), .A(n9786), .B(n9785), .ZN(
        P1_U3272) );
  XOR2_X1 U11114 ( .A(n4584), .B(n9789), .Z(n10006) );
  INV_X1 U11115 ( .A(n9788), .ZN(n9791) );
  INV_X1 U11116 ( .A(n9789), .ZN(n9790) );
  AOI21_X1 U11117 ( .B1(n9791), .B2(n9790), .A(n10210), .ZN(n9795) );
  OAI22_X1 U11118 ( .A1(n9792), .A2(n10057), .B1(n9822), .B2(n10038), .ZN(
        n9793) );
  AOI21_X1 U11119 ( .B1(n9795), .B2(n4580), .A(n9793), .ZN(n10005) );
  INV_X1 U11120 ( .A(n10005), .ZN(n9801) );
  NAND2_X1 U11121 ( .A1(n9810), .A2(n10001), .ZN(n9796) );
  AND2_X1 U11122 ( .A1(n5175), .A2(n9796), .ZN(n10003) );
  NAND2_X1 U11123 ( .A1(n10003), .A2(n9931), .ZN(n9799) );
  AOI22_X1 U11124 ( .A1(n9797), .A2(n9932), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9933), .ZN(n9798) );
  OAI211_X1 U11125 ( .C1(n5054), .C2(n9926), .A(n9799), .B(n9798), .ZN(n9800)
         );
  AOI21_X1 U11126 ( .B1(n9801), .B2(n9854), .A(n9800), .ZN(n9802) );
  OAI21_X1 U11127 ( .B1(n9909), .B2(n10006), .A(n9802), .ZN(P1_U3273) );
  XNOR2_X1 U11128 ( .A(n9803), .B(n9806), .ZN(n10011) );
  OAI211_X1 U11129 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n9988), .ZN(n9808)
         );
  NAND2_X1 U11130 ( .A1(n9842), .A2(n10053), .ZN(n9807) );
  OAI211_X1 U11131 ( .C1(n9992), .C2(n10057), .A(n9808), .B(n9807), .ZN(n10007) );
  NAND2_X1 U11132 ( .A1(n10007), .A2(n9854), .ZN(n9817) );
  OR2_X1 U11133 ( .A1(n9826), .A2(n9811), .ZN(n9809) );
  AND3_X1 U11134 ( .A1(n9810), .A2(n9809), .A3(n10002), .ZN(n10008) );
  NOR2_X1 U11135 ( .A1(n9811), .A2(n9926), .ZN(n9815) );
  OAI22_X1 U11136 ( .A1(n9813), .A2(n9891), .B1(n9812), .B2(n9893), .ZN(n9814)
         );
  AOI211_X1 U11137 ( .C1(n10008), .C2(n9921), .A(n9815), .B(n9814), .ZN(n9816)
         );
  OAI211_X1 U11138 ( .C1(n10011), .C2(n9909), .A(n9817), .B(n9816), .ZN(
        P1_U3274) );
  XNOR2_X1 U11139 ( .A(n9818), .B(n9820), .ZN(n10012) );
  INV_X1 U11140 ( .A(n10012), .ZN(n9834) );
  OAI211_X1 U11141 ( .C1(n9821), .C2(n9820), .A(n4413), .B(n9988), .ZN(n9825)
         );
  OAI22_X1 U11142 ( .A1(n9822), .A2(n10057), .B1(n9861), .B2(n10038), .ZN(
        n9823) );
  INV_X1 U11143 ( .A(n9823), .ZN(n9824) );
  NAND2_X1 U11144 ( .A1(n9825), .A2(n9824), .ZN(n10015) );
  OAI21_X1 U11145 ( .B1(n9847), .B2(n9831), .A(n10002), .ZN(n9827) );
  NOR2_X1 U11146 ( .A1(n9827), .A2(n9826), .ZN(n10013) );
  NAND2_X1 U11147 ( .A1(n10013), .A2(n9921), .ZN(n9830) );
  AOI22_X1 U11148 ( .A1(n9933), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9828), .B2(
        n9932), .ZN(n9829) );
  OAI211_X1 U11149 ( .C1(n9831), .C2(n9926), .A(n9830), .B(n9829), .ZN(n9832)
         );
  AOI21_X1 U11150 ( .B1(n10015), .B2(n9854), .A(n9832), .ZN(n9833) );
  OAI21_X1 U11151 ( .B1(n9909), .B2(n9834), .A(n9833), .ZN(P1_U3275) );
  XNOR2_X1 U11152 ( .A(n9835), .B(n9836), .ZN(n10022) );
  AND2_X1 U11153 ( .A1(n9837), .A2(n9838), .ZN(n9841) );
  OAI211_X1 U11154 ( .C1(n9841), .C2(n9840), .A(n9839), .B(n9988), .ZN(n9844)
         );
  NAND2_X1 U11155 ( .A1(n9842), .A2(n10212), .ZN(n9843) );
  OAI211_X1 U11156 ( .C1(n9881), .C2(n10038), .A(n9844), .B(n9843), .ZN(n10018) );
  NAND2_X1 U11157 ( .A1(n4449), .A2(n10020), .ZN(n9845) );
  NAND2_X1 U11158 ( .A1(n9845), .A2(n10002), .ZN(n9846) );
  NOR2_X1 U11159 ( .A1(n9847), .A2(n9846), .ZN(n10019) );
  NAND2_X1 U11160 ( .A1(n10019), .A2(n9921), .ZN(n9852) );
  INV_X1 U11161 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9849) );
  OAI22_X1 U11162 ( .A1(n9893), .A2(n9849), .B1(n9848), .B2(n9891), .ZN(n9850)
         );
  AOI21_X1 U11163 ( .B1(n10020), .B2(n9930), .A(n9850), .ZN(n9851) );
  NAND2_X1 U11164 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  AOI21_X1 U11165 ( .B1(n10018), .B2(n9854), .A(n9853), .ZN(n9855) );
  OAI21_X1 U11166 ( .B1(n10022), .B2(n9909), .A(n9855), .ZN(P1_U3276) );
  OAI21_X1 U11167 ( .B1(n9856), .B2(n9868), .A(n9837), .ZN(n9857) );
  INV_X1 U11168 ( .A(n9857), .ZN(n10027) );
  AOI22_X1 U11169 ( .A1(n9933), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9858), .B2(
        n9932), .ZN(n9860) );
  NAND2_X1 U11170 ( .A1(n9898), .A2(n10023), .ZN(n9859) );
  OAI211_X1 U11171 ( .C1(n9861), .C2(n9894), .A(n9860), .B(n9859), .ZN(n9865)
         );
  INV_X1 U11172 ( .A(n9866), .ZN(n10091) );
  INV_X1 U11173 ( .A(n9862), .ZN(n9873) );
  OAI211_X1 U11174 ( .C1(n10091), .C2(n9873), .A(n4449), .B(n10002), .ZN(
        n10025) );
  NOR2_X1 U11175 ( .A1(n10025), .A2(n9863), .ZN(n9864) );
  AOI211_X1 U11176 ( .C1(n9930), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9870)
         );
  XNOR2_X1 U11177 ( .A(n9867), .B(n9868), .ZN(n10029) );
  NAND2_X1 U11178 ( .A1(n10029), .A2(n9928), .ZN(n9869) );
  OAI211_X1 U11179 ( .C1(n10027), .C2(n9871), .A(n9870), .B(n9869), .ZN(
        P1_U3277) );
  XOR2_X1 U11180 ( .A(n9872), .B(n9878), .Z(n10037) );
  INV_X1 U11181 ( .A(n9890), .ZN(n9874) );
  AOI211_X1 U11182 ( .C1(n10034), .C2(n9874), .A(n9920), .B(n9873), .ZN(n10033) );
  AOI22_X1 U11183 ( .A1(n9933), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9875), .B2(
        n9932), .ZN(n9876) );
  OAI21_X1 U11184 ( .B1(n9877), .B2(n9926), .A(n9876), .ZN(n9885) );
  AOI21_X1 U11185 ( .B1(n9879), .B2(n9878), .A(n10210), .ZN(n9883) );
  OAI22_X1 U11186 ( .A1(n9881), .A2(n10057), .B1(n9912), .B2(n10038), .ZN(
        n9882) );
  AOI21_X1 U11187 ( .B1(n9883), .B2(n9880), .A(n9882), .ZN(n10035) );
  NOR2_X1 U11188 ( .A1(n10035), .A2(n9933), .ZN(n9884) );
  AOI211_X1 U11189 ( .C1(n10033), .C2(n9921), .A(n9885), .B(n9884), .ZN(n9886)
         );
  OAI21_X1 U11190 ( .B1(n10037), .B2(n9909), .A(n9886), .ZN(P1_U3278) );
  XNOR2_X1 U11191 ( .A(n9887), .B(n9903), .ZN(n10045) );
  NAND2_X1 U11192 ( .A1(n9918), .A2(n10042), .ZN(n9888) );
  NAND2_X1 U11193 ( .A1(n9888), .A2(n10002), .ZN(n9889) );
  NOR2_X1 U11194 ( .A1(n9890), .A2(n9889), .ZN(n10040) );
  OAI22_X1 U11195 ( .A1(n9893), .A2(n10461), .B1(n9892), .B2(n9891), .ZN(n9896) );
  NOR2_X1 U11196 ( .A1(n9894), .A2(n10039), .ZN(n9895) );
  AOI211_X1 U11197 ( .C1(n9898), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9899)
         );
  OAI21_X1 U11198 ( .B1(n9900), .B2(n9926), .A(n9899), .ZN(n9907) );
  NOR2_X1 U11199 ( .A1(n9901), .A2(n9916), .ZN(n9910) );
  NOR2_X1 U11200 ( .A1(n9910), .A2(n9902), .ZN(n9904) );
  XNOR2_X1 U11201 ( .A(n9904), .B(n9903), .ZN(n9905) );
  NAND2_X1 U11202 ( .A1(n9905), .A2(n9988), .ZN(n10044) );
  NOR2_X1 U11203 ( .A1(n10044), .A2(n9933), .ZN(n9906) );
  AOI211_X1 U11204 ( .C1(n10040), .C2(n9921), .A(n9907), .B(n9906), .ZN(n9908)
         );
  OAI21_X1 U11205 ( .B1(n10045), .B2(n9909), .A(n9908), .ZN(P1_U3279) );
  AOI211_X1 U11206 ( .C1(n9916), .C2(n9901), .A(n10210), .B(n9910), .ZN(n9914)
         );
  OAI22_X1 U11207 ( .A1(n9912), .A2(n10057), .B1(n9911), .B2(n10038), .ZN(
        n9913) );
  NOR2_X1 U11208 ( .A1(n9914), .A2(n9913), .ZN(n10051) );
  OAI21_X1 U11209 ( .B1(n9917), .B2(n9916), .A(n9915), .ZN(n10046) );
  INV_X1 U11210 ( .A(n9918), .ZN(n9919) );
  AOI211_X1 U11211 ( .C1(n10048), .C2(n4524), .A(n9920), .B(n9919), .ZN(n10047) );
  NAND2_X1 U11212 ( .A1(n10047), .A2(n9921), .ZN(n9925) );
  INV_X1 U11213 ( .A(n9922), .ZN(n9923) );
  AOI22_X1 U11214 ( .A1(n9933), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9923), .B2(
        n9932), .ZN(n9924) );
  OAI211_X1 U11215 ( .C1(n7076), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9927)
         );
  AOI21_X1 U11216 ( .B1(n9928), .B2(n10046), .A(n9927), .ZN(n9929) );
  OAI21_X1 U11217 ( .B1(n10051), .B2(n9933), .A(n9929), .ZN(P1_U3280) );
  OAI21_X1 U11218 ( .B1(n9931), .B2(n9930), .A(n5016), .ZN(n9940) );
  AOI22_X1 U11219 ( .A1(n9933), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9932), .ZN(n9939) );
  NAND4_X1 U11220 ( .A1(n10213), .A2(n9935), .A3(n9934), .A4(n9854), .ZN(n9938) );
  NAND2_X1 U11221 ( .A1(n9936), .A2(n6400), .ZN(n9937) );
  NAND4_X1 U11222 ( .A1(n9940), .A2(n9939), .A3(n9938), .A4(n9937), .ZN(
        P1_U3293) );
  OAI22_X1 U11223 ( .A1(n9947), .A2(n10057), .B1(n9946), .B2(n10038), .ZN(
        n9948) );
  OAI22_X1 U11224 ( .A1(n9954), .A2(n10057), .B1(n9953), .B2(n10038), .ZN(
        n9955) );
  INV_X1 U11225 ( .A(n9955), .ZN(n9958) );
  INV_X1 U11226 ( .A(n9960), .ZN(P1_U3548) );
  AOI22_X1 U11227 ( .A1(n9962), .A2(n10002), .B1(n10049), .B2(n9961), .ZN(
        n9963) );
  OAI211_X1 U11228 ( .C1(n10211), .C2(n9965), .A(n9964), .B(n9963), .ZN(n10075) );
  MUX2_X1 U11229 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10075), .S(n10252), .Z(
        P1_U3547) );
  AND3_X1 U11230 ( .A1(n9967), .A2(n10241), .A3(n9966), .ZN(n9971) );
  OAI21_X1 U11231 ( .B1(n9969), .B2(n10237), .A(n9968), .ZN(n9970) );
  MUX2_X1 U11232 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10076), .S(n10252), .Z(
        P1_U3546) );
  AOI22_X1 U11233 ( .A1(n9974), .A2(n10212), .B1(n10053), .B2(n9973), .ZN(
        n9975) );
  OAI211_X1 U11234 ( .C1(n9977), .C2(n10237), .A(n9976), .B(n9975), .ZN(n9978)
         );
  AOI21_X1 U11235 ( .B1(n9979), .B2(n9988), .A(n9978), .ZN(n9980) );
  OAI21_X1 U11236 ( .B1(n10211), .B2(n9981), .A(n9980), .ZN(n10077) );
  MUX2_X1 U11237 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10077), .S(n10252), .Z(
        P1_U3545) );
  AOI22_X1 U11238 ( .A1(n9983), .A2(n10212), .B1(n10053), .B2(n9982), .ZN(
        n9984) );
  OAI21_X1 U11239 ( .B1(n9985), .B2(n10237), .A(n9984), .ZN(n9986) );
  AOI211_X1 U11240 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9990)
         );
  OAI21_X1 U11241 ( .B1(n10211), .B2(n9991), .A(n9990), .ZN(n10078) );
  MUX2_X1 U11242 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10078), .S(n10252), .Z(
        P1_U3544) );
  OAI22_X1 U11243 ( .A1(n9993), .A2(n10057), .B1(n9992), .B2(n10038), .ZN(
        n9995) );
  AOI211_X1 U11244 ( .C1(n10049), .C2(n9996), .A(n9995), .B(n9994), .ZN(n9999)
         );
  NAND2_X1 U11245 ( .A1(n9997), .A2(n10241), .ZN(n9998) );
  OAI211_X1 U11246 ( .C1(n10000), .C2(n10210), .A(n9999), .B(n9998), .ZN(
        n10079) );
  MUX2_X1 U11247 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10079), .S(n10252), .Z(
        P1_U3543) );
  AOI22_X1 U11248 ( .A1(n10003), .A2(n10002), .B1(n10049), .B2(n10001), .ZN(
        n10004) );
  OAI211_X1 U11249 ( .C1(n10211), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        n10080) );
  MUX2_X1 U11250 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10080), .S(n10252), .Z(
        P1_U3542) );
  AOI211_X1 U11251 ( .C1(n10049), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10010) );
  OAI21_X1 U11252 ( .B1(n10211), .B2(n10011), .A(n10010), .ZN(n10081) );
  MUX2_X1 U11253 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10081), .S(n10252), .Z(
        P1_U3541) );
  AND2_X1 U11254 ( .A1(n10012), .A2(n10241), .ZN(n10014) );
  MUX2_X1 U11255 ( .A(n10082), .B(P1_REG1_REG_18__SCAN_IN), .S(n4409), .Z(
        n10016) );
  AOI21_X1 U11256 ( .B1(n10063), .B2(n10084), .A(n10016), .ZN(n10017) );
  INV_X1 U11257 ( .A(n10017), .ZN(P1_U3540) );
  AOI211_X1 U11258 ( .C1(n10049), .C2(n10020), .A(n10019), .B(n10018), .ZN(
        n10021) );
  OAI21_X1 U11259 ( .B1(n10211), .B2(n10022), .A(n10021), .ZN(n10086) );
  MUX2_X1 U11260 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10086), .S(n10252), .Z(
        P1_U3539) );
  AOI22_X1 U11261 ( .A1(n10024), .A2(n10212), .B1(n10023), .B2(n10053), .ZN(
        n10026) );
  OAI211_X1 U11262 ( .C1(n10027), .C2(n10210), .A(n10026), .B(n10025), .ZN(
        n10028) );
  AOI21_X1 U11263 ( .B1(n10029), .B2(n10241), .A(n10028), .ZN(n10087) );
  MUX2_X1 U11264 ( .A(n10030), .B(n10087), .S(n10252), .Z(n10031) );
  OAI21_X1 U11265 ( .B1(n10091), .B2(n10032), .A(n10031), .ZN(P1_U3538) );
  AOI21_X1 U11266 ( .B1(n10049), .B2(n10034), .A(n10033), .ZN(n10036) );
  OAI211_X1 U11267 ( .C1(n10211), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10092) );
  MUX2_X1 U11268 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10092), .S(n10252), .Z(
        P1_U3537) );
  OAI22_X1 U11269 ( .A1(n10039), .A2(n10057), .B1(n10058), .B2(n10038), .ZN(
        n10041) );
  AOI211_X1 U11270 ( .C1(n10049), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10043) );
  OAI211_X1 U11271 ( .C1(n10211), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10093) );
  MUX2_X1 U11272 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10093), .S(n10252), .Z(
        P1_U3536) );
  INV_X1 U11273 ( .A(n10046), .ZN(n10052) );
  AOI21_X1 U11274 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(n10050) );
  OAI211_X1 U11275 ( .C1(n10211), .C2(n10052), .A(n10051), .B(n10050), .ZN(
        n10094) );
  MUX2_X1 U11276 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10094), .S(n10252), .Z(
        P1_U3535) );
  NAND2_X1 U11277 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  OAI211_X1 U11278 ( .C1(n10058), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        n10061) );
  NOR2_X1 U11279 ( .A1(n10059), .A2(n10210), .ZN(n10060) );
  AOI211_X1 U11280 ( .C1(n10241), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        n10097) );
  AOI22_X1 U11281 ( .A1(n10095), .A2(n10063), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n4409), .ZN(n10064) );
  OAI21_X1 U11282 ( .B1(n10097), .B2(n4409), .A(n10064), .ZN(P1_U3534) );
  OAI21_X1 U11283 ( .B1(n10067), .B2(n10090), .A(n10066), .ZN(P1_U3521) );
  INV_X1 U11284 ( .A(n10069), .ZN(n10070) );
  OAI21_X1 U11285 ( .B1(n5034), .B2(n10090), .A(n10070), .ZN(P1_U3520) );
  MUX2_X1 U11286 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10075), .S(n10243), .Z(
        P1_U3515) );
  MUX2_X1 U11287 ( .A(n10076), .B(P1_REG0_REG_24__SCAN_IN), .S(n7144), .Z(
        P1_U3514) );
  MUX2_X1 U11288 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10077), .S(n10243), .Z(
        P1_U3513) );
  MUX2_X1 U11289 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10078), .S(n10243), .Z(
        P1_U3512) );
  MUX2_X1 U11290 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10079), .S(n10243), .Z(
        P1_U3511) );
  MUX2_X1 U11291 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10080), .S(n10243), .Z(
        P1_U3510) );
  MUX2_X1 U11292 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10081), .S(n10243), .Z(
        P1_U3509) );
  MUX2_X1 U11293 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10082), .S(n10243), .Z(
        n10083) );
  AOI21_X1 U11294 ( .B1(n7093), .B2(n10084), .A(n10083), .ZN(n10085) );
  INV_X1 U11295 ( .A(n10085), .ZN(P1_U3507) );
  MUX2_X1 U11296 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10086), .S(n10243), .Z(
        P1_U3504) );
  INV_X1 U11297 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10088) );
  MUX2_X1 U11298 ( .A(n10088), .B(n10087), .S(n10243), .Z(n10089) );
  OAI21_X1 U11299 ( .B1(n10091), .B2(n10090), .A(n10089), .ZN(P1_U3501) );
  MUX2_X1 U11300 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10092), .S(n10243), .Z(
        P1_U3498) );
  MUX2_X1 U11301 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10093), .S(n10243), .Z(
        P1_U3495) );
  MUX2_X1 U11302 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10094), .S(n10243), .Z(
        P1_U3492) );
  AOI22_X1 U11303 ( .A1(n10095), .A2(n7093), .B1(P1_REG0_REG_12__SCAN_IN), 
        .B2(n7144), .ZN(n10096) );
  OAI21_X1 U11304 ( .B1(n10097), .B2(n7144), .A(n10096), .ZN(P1_U3489) );
  MUX2_X1 U11305 ( .A(P1_D_REG_1__SCAN_IN), .B(n10100), .S(n10208), .Z(
        P1_U3440) );
  MUX2_X1 U11306 ( .A(P1_D_REG_0__SCAN_IN), .B(n10101), .S(n10208), .Z(
        P1_U3439) );
  NOR2_X1 U11307 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n10104) );
  NAND4_X1 U11308 ( .A1(n10104), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n10103), .ZN(n10106) );
  OAI22_X1 U11309 ( .A1(n10102), .A2(n10106), .B1(n10105), .B2(n10116), .ZN(
        n10107) );
  AOI21_X1 U11310 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(n10110) );
  INV_X1 U11311 ( .A(n10110), .ZN(P1_U3324) );
  OAI222_X1 U11312 ( .A1(n10115), .A2(P1_U3086), .B1(n8337), .B2(n10114), .C1(
        n10113), .C2(n10116), .ZN(P1_U3329) );
  OAI222_X1 U11313 ( .A1(n10118), .A2(P1_U3086), .B1(n8337), .B2(n10117), .C1(
        n10563), .C2(n10116), .ZN(P1_U3330) );
  XNOR2_X1 U11314 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U11315 ( .A(n10119), .ZN(n10124) );
  INV_X1 U11316 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10383) );
  NAND2_X1 U11317 ( .A1(n10120), .A2(n10122), .ZN(n10121) );
  MUX2_X1 U11318 ( .A(n10122), .B(n10121), .S(P1_IR_REG_0__SCAN_IN), .Z(n10123) );
  NAND2_X1 U11319 ( .A1(n10124), .A2(n10123), .ZN(n10126) );
  AOI22_X1 U11320 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10169), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10125) );
  OAI21_X1 U11321 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(P1_U3243) );
  INV_X1 U11322 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10139) );
  AOI211_X1 U11323 ( .C1(n10130), .C2(n10129), .A(n10152), .B(n10128), .ZN(
        n10135) );
  AOI211_X1 U11324 ( .C1(n10133), .C2(n10132), .A(n10164), .B(n10131), .ZN(
        n10134) );
  AOI211_X1 U11325 ( .C1(n10183), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10138) );
  OAI211_X1 U11326 ( .C1(n10207), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        P1_U3256) );
  INV_X1 U11327 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10151) );
  AOI211_X1 U11328 ( .C1(n10142), .C2(n10141), .A(n10140), .B(n10164), .ZN(
        n10147) );
  AOI211_X1 U11329 ( .C1(n10145), .C2(n10144), .A(n10152), .B(n10143), .ZN(
        n10146) );
  AOI211_X1 U11330 ( .C1(n10183), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10150) );
  OAI211_X1 U11331 ( .C1(n10207), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        P1_U3257) );
  INV_X1 U11332 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10163) );
  AOI211_X1 U11333 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10159) );
  AOI211_X1 U11334 ( .C1(n10157), .C2(n6701), .A(n10156), .B(n10164), .ZN(
        n10158) );
  AOI211_X1 U11335 ( .C1(n10183), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        n10162) );
  OAI211_X1 U11336 ( .C1(n10207), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        P1_U3258) );
  AOI211_X1 U11337 ( .C1(n4515), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        n10167) );
  AOI211_X1 U11338 ( .C1(n10169), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10168), 
        .B(n10167), .ZN(n10175) );
  OAI21_X1 U11339 ( .B1(n10171), .B2(n4518), .A(n10170), .ZN(n10173) );
  AOI22_X1 U11340 ( .A1(n10173), .A2(n10198), .B1(n10172), .B2(n10183), .ZN(
        n10174) );
  NAND2_X1 U11341 ( .A1(n10175), .A2(n10174), .ZN(P1_U3259) );
  INV_X1 U11342 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10188) );
  OAI21_X1 U11343 ( .B1(n10178), .B2(n10177), .A(n10176), .ZN(n10185) );
  OAI21_X1 U11344 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(n10182) );
  AOI222_X1 U11345 ( .A1(n10185), .A2(n10193), .B1(n10184), .B2(n10183), .C1(
        n10182), .C2(n10198), .ZN(n10187) );
  OAI211_X1 U11346 ( .C1(n10207), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        P1_U3260) );
  NAND2_X1 U11347 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  NAND3_X1 U11348 ( .A1(n10193), .A2(n10192), .A3(n10191), .ZN(n10200) );
  NAND2_X1 U11349 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  NAND3_X1 U11350 ( .A1(n10198), .A2(n10197), .A3(n10196), .ZN(n10199) );
  OAI211_X1 U11351 ( .C1(n10202), .C2(n10201), .A(n10200), .B(n10199), .ZN(
        n10203) );
  INV_X1 U11352 ( .A(n10203), .ZN(n10205) );
  OAI211_X1 U11353 ( .C1(n10207), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        P1_U3261) );
  AND2_X1 U11354 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10209), .ZN(P1_U3294) );
  AND2_X1 U11355 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10209), .ZN(P1_U3295) );
  NOR2_X1 U11356 ( .A1(n10208), .A2(n10650), .ZN(P1_U3296) );
  NOR2_X1 U11357 ( .A1(n10208), .A2(n10445), .ZN(P1_U3297) );
  AND2_X1 U11358 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10209), .ZN(P1_U3298) );
  AND2_X1 U11359 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10209), .ZN(P1_U3299) );
  AND2_X1 U11360 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10209), .ZN(P1_U3300) );
  INV_X1 U11361 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10448) );
  NOR2_X1 U11362 ( .A1(n10208), .A2(n10448), .ZN(P1_U3301) );
  AND2_X1 U11363 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10209), .ZN(P1_U3302) );
  AND2_X1 U11364 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10209), .ZN(P1_U3303) );
  NOR2_X1 U11365 ( .A1(n10208), .A2(n10576), .ZN(P1_U3304) );
  AND2_X1 U11366 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10209), .ZN(P1_U3305) );
  AND2_X1 U11367 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10209), .ZN(P1_U3306) );
  INV_X1 U11368 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U11369 ( .A1(n10208), .A2(n10566), .ZN(P1_U3307) );
  AND2_X1 U11370 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10209), .ZN(P1_U3308) );
  AND2_X1 U11371 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10209), .ZN(P1_U3309) );
  INV_X1 U11372 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10525) );
  NOR2_X1 U11373 ( .A1(n10208), .A2(n10525), .ZN(P1_U3310) );
  INV_X1 U11374 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10625) );
  NOR2_X1 U11375 ( .A1(n10208), .A2(n10625), .ZN(P1_U3311) );
  INV_X1 U11376 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10610) );
  NOR2_X1 U11377 ( .A1(n10208), .A2(n10610), .ZN(P1_U3312) );
  INV_X1 U11378 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U11379 ( .A1(n10208), .A2(n10649), .ZN(P1_U3313) );
  AND2_X1 U11380 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10209), .ZN(P1_U3314) );
  AND2_X1 U11381 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10209), .ZN(P1_U3315) );
  AND2_X1 U11382 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10209), .ZN(P1_U3316) );
  AND2_X1 U11383 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10209), .ZN(P1_U3317) );
  AND2_X1 U11384 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10209), .ZN(P1_U3318) );
  NOR2_X1 U11385 ( .A1(n10208), .A2(n10552), .ZN(P1_U3319) );
  AND2_X1 U11386 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10209), .ZN(P1_U3320) );
  AND2_X1 U11387 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10209), .ZN(P1_U3321) );
  AND2_X1 U11388 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10209), .ZN(P1_U3322) );
  AND2_X1 U11389 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10209), .ZN(P1_U3323) );
  NAND2_X1 U11390 ( .A1(n10211), .A2(n10210), .ZN(n10214) );
  AOI222_X1 U11391 ( .A1(n10214), .A2(n10213), .B1(n5016), .B2(n5181), .C1(
        n6400), .C2(n10212), .ZN(n10244) );
  AOI22_X1 U11392 ( .A1(n10243), .A2(n10244), .B1(n6328), .B2(n7144), .ZN(
        P1_U3453) );
  INV_X1 U11393 ( .A(n10215), .ZN(n10216) );
  NAND2_X1 U11394 ( .A1(n10217), .A2(n10216), .ZN(n10219) );
  OAI211_X1 U11395 ( .C1(n7073), .C2(n10237), .A(n10219), .B(n10218), .ZN(
        n10220) );
  NOR2_X1 U11396 ( .A1(n10221), .A2(n10220), .ZN(n10246) );
  INV_X1 U11397 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U11398 ( .A1(n10243), .A2(n10246), .B1(n10222), .B2(n7144), .ZN(
        P1_U3456) );
  INV_X1 U11399 ( .A(n10223), .ZN(n10224) );
  OAI21_X1 U11400 ( .B1(n10225), .B2(n10237), .A(n10224), .ZN(n10226) );
  AOI211_X1 U11401 ( .C1(n10241), .C2(n10228), .A(n10227), .B(n10226), .ZN(
        n10248) );
  INV_X1 U11402 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U11403 ( .A1(n10243), .A2(n10248), .B1(n10229), .B2(n7144), .ZN(
        P1_U3459) );
  OAI21_X1 U11404 ( .B1(n10231), .B2(n10237), .A(n10230), .ZN(n10233) );
  AOI211_X1 U11405 ( .C1(n10241), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        n10250) );
  INV_X1 U11406 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U11407 ( .A1(n10243), .A2(n10250), .B1(n10235), .B2(n7144), .ZN(
        P1_U3462) );
  OAI21_X1 U11408 ( .B1(n5051), .B2(n10237), .A(n10236), .ZN(n10239) );
  AOI211_X1 U11409 ( .C1(n10241), .C2(n10240), .A(n10239), .B(n10238), .ZN(
        n10251) );
  INV_X1 U11410 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U11411 ( .A1(n10243), .A2(n10251), .B1(n10242), .B2(n7144), .ZN(
        P1_U3468) );
  AOI22_X1 U11412 ( .A1(n10252), .A2(n10244), .B1(n10383), .B2(n4409), .ZN(
        P1_U3522) );
  INV_X1 U11413 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U11414 ( .A1(n10252), .A2(n10246), .B1(n10245), .B2(n4409), .ZN(
        P1_U3523) );
  AOI22_X1 U11415 ( .A1(n10252), .A2(n10248), .B1(n10247), .B2(n4409), .ZN(
        P1_U3524) );
  INV_X1 U11416 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U11417 ( .A1(n10252), .A2(n10250), .B1(n10249), .B2(n4409), .ZN(
        P1_U3525) );
  AOI22_X1 U11418 ( .A1(n10252), .A2(n10251), .B1(n6470), .B2(n4409), .ZN(
        P1_U3527) );
  XNOR2_X1 U11419 ( .A(n10253), .B(n10258), .ZN(n10265) );
  OAI22_X1 U11420 ( .A1(n10257), .A2(n10256), .B1(n10255), .B2(n10254), .ZN(
        n10264) );
  OR2_X1 U11421 ( .A1(n10259), .A2(n10258), .ZN(n10260) );
  NAND2_X1 U11422 ( .A1(n10261), .A2(n10260), .ZN(n10333) );
  NOR2_X1 U11423 ( .A1(n10333), .A2(n10262), .ZN(n10263) );
  AOI211_X1 U11424 ( .C1(n10265), .C2(n10289), .A(n10264), .B(n10263), .ZN(
        n10329) );
  INV_X1 U11425 ( .A(n10266), .ZN(n10271) );
  INV_X1 U11426 ( .A(n10333), .ZN(n10270) );
  INV_X1 U11427 ( .A(n10267), .ZN(n10269) );
  AOI222_X1 U11428 ( .A1(n10271), .A2(n10293), .B1(n10270), .B2(n10269), .C1(
        n10268), .C2(n10292), .ZN(n10272) );
  OAI221_X1 U11429 ( .B1(n10296), .B2(n10329), .C1(n10282), .C2(n10273), .A(
        n10272), .ZN(P2_U3226) );
  XNOR2_X1 U11430 ( .A(n10274), .B(n10279), .ZN(n10277) );
  AOI222_X1 U11431 ( .A1(n10289), .A2(n10277), .B1(n10276), .B2(n10286), .C1(
        n10275), .C2(n10284), .ZN(n10314) );
  XNOR2_X1 U11432 ( .A(n10278), .B(n10279), .ZN(n10312) );
  AOI222_X1 U11433 ( .A1(n10312), .A2(n7723), .B1(n10280), .B2(n10293), .C1(
        n10311), .C2(n10292), .ZN(n10281) );
  OAI221_X1 U11434 ( .B1(n10296), .B2(n10314), .C1(n10282), .C2(n5983), .A(
        n10281), .ZN(P2_U3229) );
  XOR2_X1 U11435 ( .A(n10291), .B(n10283), .Z(n10288) );
  AOI222_X1 U11436 ( .A1(n10289), .A2(n10288), .B1(n10287), .B2(n10286), .C1(
        n10285), .C2(n10284), .ZN(n10309) );
  XNOR2_X1 U11437 ( .A(n10290), .B(n10291), .ZN(n10307) );
  AOI222_X1 U11438 ( .A1(n10307), .A2(n7723), .B1(n10294), .B2(n10293), .C1(
        n6121), .C2(n10292), .ZN(n10295) );
  OAI221_X1 U11439 ( .B1(n10296), .B2(n10309), .C1(n10282), .C2(n4889), .A(
        n10295), .ZN(P2_U3230) );
  INV_X1 U11440 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10301) );
  NOR2_X1 U11441 ( .A1(n10297), .A2(n10330), .ZN(n10299) );
  AOI211_X1 U11442 ( .C1(n10327), .C2(n10300), .A(n10299), .B(n10298), .ZN(
        n10671) );
  AOI22_X1 U11443 ( .A1(n10337), .A2(n10301), .B1(n10671), .B2(n10336), .ZN(
        P2_U3393) );
  INV_X1 U11444 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10306) );
  OAI22_X1 U11445 ( .A1(n10303), .A2(n10332), .B1(n10302), .B2(n10330), .ZN(
        n10304) );
  NOR2_X1 U11446 ( .A1(n10305), .A2(n10304), .ZN(n10339) );
  AOI22_X1 U11447 ( .A1(n10337), .A2(n10306), .B1(n10339), .B2(n10336), .ZN(
        P2_U3396) );
  INV_X1 U11448 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U11449 ( .A1(n10307), .A2(n10327), .B1(n10316), .B2(n6121), .ZN(
        n10308) );
  AND2_X1 U11450 ( .A1(n10309), .A2(n10308), .ZN(n10341) );
  AOI22_X1 U11451 ( .A1(n10337), .A2(n10310), .B1(n10341), .B2(n10336), .ZN(
        P2_U3399) );
  AOI22_X1 U11452 ( .A1(n10312), .A2(n10327), .B1(n10316), .B2(n10311), .ZN(
        n10313) );
  AND2_X1 U11453 ( .A1(n10314), .A2(n10313), .ZN(n10342) );
  AOI22_X1 U11454 ( .A1(n10337), .A2(n5295), .B1(n10342), .B2(n10336), .ZN(
        P2_U3402) );
  INV_X1 U11455 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U11456 ( .A1(n10318), .A2(n10317), .B1(n10316), .B2(n10315), .ZN(
        n10319) );
  AND2_X1 U11457 ( .A1(n10320), .A2(n10319), .ZN(n10343) );
  AOI22_X1 U11458 ( .A1(n10337), .A2(n10321), .B1(n10343), .B2(n10336), .ZN(
        P2_U3405) );
  INV_X1 U11459 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10328) );
  INV_X1 U11460 ( .A(n10322), .ZN(n10326) );
  OAI21_X1 U11461 ( .B1(n10324), .B2(n10330), .A(n10323), .ZN(n10325) );
  AOI21_X1 U11462 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10344) );
  AOI22_X1 U11463 ( .A1(n10337), .A2(n10328), .B1(n10344), .B2(n10336), .ZN(
        P2_U3408) );
  INV_X1 U11464 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10529) );
  INV_X1 U11465 ( .A(n10329), .ZN(n10335) );
  OAI22_X1 U11466 ( .A1(n10333), .A2(n10332), .B1(n10331), .B2(n10330), .ZN(
        n10334) );
  NOR2_X1 U11467 ( .A1(n10335), .A2(n10334), .ZN(n10346) );
  AOI22_X1 U11468 ( .A1(n10337), .A2(n10529), .B1(n10346), .B2(n10336), .ZN(
        P2_U3411) );
  INV_X1 U11469 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U11470 ( .A1(n10672), .A2(n10339), .B1(n10338), .B2(n8960), .ZN(
        P2_U3461) );
  AOI22_X1 U11471 ( .A1(n10672), .A2(n10341), .B1(n10340), .B2(n8960), .ZN(
        P2_U3462) );
  AOI22_X1 U11472 ( .A1(n10672), .A2(n10342), .B1(n5953), .B2(n8960), .ZN(
        P2_U3463) );
  AOI22_X1 U11473 ( .A1(n10672), .A2(n10343), .B1(n4863), .B2(n8960), .ZN(
        P2_U3464) );
  AOI22_X1 U11474 ( .A1(n10672), .A2(n10344), .B1(n10546), .B2(n8960), .ZN(
        P2_U3465) );
  AOI22_X1 U11475 ( .A1(n10672), .A2(n10346), .B1(n10345), .B2(n8960), .ZN(
        P2_U3466) );
  OAI222_X1 U11476 ( .A1(n10351), .A2(n10350), .B1(n10351), .B2(n10349), .C1(
        n10348), .C2(n10347), .ZN(ADD_1068_U5) );
  XOR2_X1 U11477 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11478 ( .A(n10354), .ZN(n10353) );
  OAI222_X1 U11479 ( .A1(n10356), .A2(n10355), .B1(n10356), .B2(n10354), .C1(
        n10353), .C2(n10352), .ZN(ADD_1068_U55) );
  OAI21_X1 U11480 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(ADD_1068_U56) );
  OAI21_X1 U11481 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(ADD_1068_U57) );
  OAI21_X1 U11482 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(ADD_1068_U58) );
  OAI21_X1 U11483 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(ADD_1068_U59) );
  OAI21_X1 U11484 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(ADD_1068_U60) );
  OAI21_X1 U11485 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(ADD_1068_U61) );
  OAI21_X1 U11486 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(ADD_1068_U62) );
  OAI21_X1 U11487 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(ADD_1068_U63) );
  NAND4_X1 U11488 ( .A1(n4846), .A2(SI_12_), .A3(SI_7_), .A4(
        P2_REG0_REG_30__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U11489 ( .A1(n10449), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10381) );
  NOR4_X1 U11490 ( .A1(n10382), .A2(n10381), .A3(P1_IR_REG_8__SCAN_IN), .A4(
        P1_IR_REG_4__SCAN_IN), .ZN(n10389) );
  NOR4_X1 U11491 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(P2_REG0_REG_23__SCAN_IN), 
        .A3(P2_REG2_REG_1__SCAN_IN), .A4(n10573), .ZN(n10385) );
  NOR4_X1 U11492 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(P1_REG1_REG_7__SCAN_IN), 
        .A3(P1_REG1_REG_6__SCAN_IN), .A4(P2_IR_REG_11__SCAN_IN), .ZN(n10384)
         );
  NAND3_X1 U11493 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n10385), .A3(n10384), 
        .ZN(n10386) );
  NOR4_X1 U11494 ( .A1(n10387), .A2(P2_IR_REG_15__SCAN_IN), .A3(
        P2_IR_REG_16__SCAN_IN), .A4(n10386), .ZN(n10388) );
  NAND4_X1 U11495 ( .A1(n10389), .A2(P1_D_REG_24__SCAN_IN), .A3(n10388), .A4(
        n10461), .ZN(n10397) );
  NAND4_X1 U11496 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), 
        .A3(P2_REG2_REG_11__SCAN_IN), .A4(n9745), .ZN(n10396) );
  INV_X1 U11497 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10390) );
  NAND4_X1 U11498 ( .A1(n10391), .A2(n10390), .A3(n10460), .A4(
        P1_IR_REG_18__SCAN_IN), .ZN(n10395) );
  NAND4_X1 U11499 ( .A1(n10393), .A2(n10392), .A3(P1_REG2_REG_1__SCAN_IN), 
        .A4(P2_DATAO_REG_19__SCAN_IN), .ZN(n10394) );
  NOR4_X1 U11500 ( .A1(n10397), .A2(n10396), .A3(n10395), .A4(n10394), .ZN(
        n10400) );
  NAND4_X1 U11501 ( .A1(P1_B_REG_SCAN_IN), .A2(P2_DATAO_REG_15__SCAN_IN), .A3(
        P1_REG2_REG_19__SCAN_IN), .A4(P2_REG2_REG_22__SCAN_IN), .ZN(n10398) );
  NOR3_X1 U11502 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .A3(n10398), .ZN(n10399) );
  NAND2_X1 U11503 ( .A1(n10400), .A2(n10399), .ZN(n10409) );
  NOR4_X1 U11504 ( .A1(SI_28_), .A2(n10501), .A3(n10500), .A4(n10506), .ZN(
        n10407) );
  NOR4_X1 U11505 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(P1_DATAO_REG_5__SCAN_IN), 
        .A3(P1_REG0_REG_30__SCAN_IN), .A4(n5597), .ZN(n10406) );
  NAND4_X1 U11506 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_REG1_REG_28__SCAN_IN), 
        .A3(P2_REG2_REG_13__SCAN_IN), .A4(n10519), .ZN(n10404) );
  NAND4_X1 U11507 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), 
        .A3(n10505), .A4(n10517), .ZN(n10403) );
  INV_X1 U11508 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10532) );
  NAND4_X1 U11509 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(n10532), .A3(n10535), .A4(
        n8770), .ZN(n10402) );
  NAND4_X1 U11510 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(n6012), .ZN(n10401) );
  NOR4_X1 U11511 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10405) );
  NAND3_X1 U11512 ( .A1(n10407), .A2(n10406), .A3(n10405), .ZN(n10408) );
  NOR2_X1 U11513 ( .A1(n10409), .A2(n10408), .ZN(n10433) );
  INV_X1 U11514 ( .A(n10410), .ZN(n10430) );
  INV_X1 U11515 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10596) );
  NOR4_X1 U11516 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .A3(n10470), .A4(n10596), .ZN(n10416) );
  NAND4_X1 U11517 ( .A1(SI_13_), .A2(SI_3_), .A3(P1_REG0_REG_15__SCAN_IN), 
        .A4(n10623), .ZN(n10414) );
  NAND4_X1 U11518 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), 
        .A3(SI_15_), .A4(P2_IR_REG_7__SCAN_IN), .ZN(n10413) );
  NAND4_X1 U11519 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), 
        .A3(P2_REG0_REG_22__SCAN_IN), .A4(n10656), .ZN(n10412) );
  NAND4_X1 U11520 ( .A1(P2_REG0_REG_28__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_25__SCAN_IN), .A4(n10613), .ZN(n10411) );
  NOR4_X1 U11521 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10415) );
  NAND4_X1 U11522 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10534), .ZN(
        n10429) );
  NAND4_X1 U11523 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), 
        .A3(n10563), .A4(n5983), .ZN(n10418) );
  NOR3_X1 U11524 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n5367), .A3(n10418), .ZN(
        n10427) );
  NAND4_X1 U11525 ( .A1(SI_27_), .A2(P1_REG2_REG_4__SCAN_IN), .A3(
        P2_REG1_REG_19__SCAN_IN), .A4(P2_REG1_REG_6__SCAN_IN), .ZN(n10425) );
  NAND4_X1 U11526 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), 
        .A3(P1_REG1_REG_14__SCAN_IN), .A4(n10565), .ZN(n10424) );
  NOR4_X1 U11527 ( .A1(P1_RD_REG_SCAN_IN), .A2(P1_REG0_REG_10__SCAN_IN), .A3(
        P1_REG0_REG_0__SCAN_IN), .A4(P2_REG3_REG_3__SCAN_IN), .ZN(n10422) );
  NOR4_X1 U11528 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(P2_D_REG_1__SCAN_IN), 
        .A3(P2_REG2_REG_15__SCAN_IN), .A4(n10636), .ZN(n10421) );
  NOR4_X1 U11529 ( .A1(SI_25_), .A2(P1_REG0_REG_22__SCAN_IN), .A3(
        P2_IR_REG_25__SCAN_IN), .A4(P2_REG3_REG_21__SCAN_IN), .ZN(n10420) );
  INV_X1 U11530 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10551) );
  NOR4_X1 U11531 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(SI_30_), .A3(n10551), 
        .A4(n10590), .ZN(n10419) );
  NAND4_X1 U11532 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10423) );
  NOR3_X1 U11533 ( .A1(n10425), .A2(n10424), .A3(n10423), .ZN(n10426) );
  NAND4_X1 U11534 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_REG2_REG_10__SCAN_IN), 
        .A3(n10427), .A4(n10426), .ZN(n10428) );
  NOR4_X1 U11535 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10432) );
  AOI21_X1 U11536 ( .B1(n10433), .B2(n10432), .A(P1_IR_REG_24__SCAN_IN), .ZN(
        n10670) );
  INV_X1 U11537 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U11538 ( .A1(P2_U3151), .A2(keyinput116), .B1(n10435), .B2(
        keyinput112), .ZN(n10434) );
  OAI221_X1 U11539 ( .B1(P2_U3151), .B2(keyinput116), .C1(n10435), .C2(
        keyinput112), .A(n10434), .ZN(n10443) );
  XOR2_X1 U11540 ( .A(P1_REG1_REG_7__SCAN_IN), .B(keyinput118), .Z(n10442) );
  XNOR2_X1 U11541 ( .A(keyinput8), .B(n7260), .ZN(n10441) );
  XNOR2_X1 U11542 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput121), .ZN(n10439)
         );
  XNOR2_X1 U11543 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput58), .ZN(n10438)
         );
  XNOR2_X1 U11544 ( .A(SI_7_), .B(keyinput87), .ZN(n10437) );
  XNOR2_X1 U11545 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput100), .ZN(n10436) );
  NAND4_X1 U11546 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        n10440) );
  NOR4_X1 U11547 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10483) );
  AOI22_X1 U11548 ( .A1(n10446), .A2(keyinput49), .B1(n10445), .B2(keyinput2), 
        .ZN(n10444) );
  OAI221_X1 U11549 ( .B1(n10446), .B2(keyinput49), .C1(n10445), .C2(keyinput2), 
        .A(n10444), .ZN(n10456) );
  AOI22_X1 U11550 ( .A1(n10449), .A2(keyinput96), .B1(n10448), .B2(keyinput34), 
        .ZN(n10447) );
  OAI221_X1 U11551 ( .B1(n10449), .B2(keyinput96), .C1(n10448), .C2(keyinput34), .A(n10447), .ZN(n10455) );
  XNOR2_X1 U11552 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput53), .ZN(n10453) );
  XNOR2_X1 U11553 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput93), .ZN(n10452)
         );
  XNOR2_X1 U11554 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput45), .ZN(n10451) );
  XNOR2_X1 U11555 ( .A(keyinput24), .B(P1_REG1_REG_0__SCAN_IN), .ZN(n10450) );
  NAND4_X1 U11556 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  NOR3_X1 U11557 ( .A1(n10456), .A2(n10455), .A3(n10454), .ZN(n10482) );
  INV_X1 U11558 ( .A(P1_B_REG_SCAN_IN), .ZN(n10458) );
  AOI22_X1 U11559 ( .A1(n8818), .A2(keyinput20), .B1(n10458), .B2(keyinput75), 
        .ZN(n10457) );
  OAI221_X1 U11560 ( .B1(n8818), .B2(keyinput20), .C1(n10458), .C2(keyinput75), 
        .A(n10457), .ZN(n10468) );
  AOI22_X1 U11561 ( .A1(n10461), .A2(keyinput83), .B1(n10460), .B2(keyinput104), .ZN(n10459) );
  OAI221_X1 U11562 ( .B1(n10461), .B2(keyinput83), .C1(n10460), .C2(
        keyinput104), .A(n10459), .ZN(n10467) );
  XNOR2_X1 U11563 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput85), .ZN(n10465)
         );
  XNOR2_X1 U11564 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput3), .ZN(n10464) );
  XNOR2_X1 U11565 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput122), .ZN(n10463)
         );
  XNOR2_X1 U11566 ( .A(P1_REG3_REG_19__SCAN_IN), .B(keyinput84), .ZN(n10462)
         );
  NAND4_X1 U11567 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10466) );
  NOR3_X1 U11568 ( .A1(n10468), .A2(n10467), .A3(n10466), .ZN(n10481) );
  AOI22_X1 U11569 ( .A1(n9812), .A2(keyinput54), .B1(keyinput72), .B2(n10470), 
        .ZN(n10469) );
  OAI221_X1 U11570 ( .B1(n9812), .B2(keyinput54), .C1(n10470), .C2(keyinput72), 
        .A(n10469), .ZN(n10479) );
  AOI22_X1 U11571 ( .A1(n9269), .A2(keyinput52), .B1(keyinput21), .B2(n9745), 
        .ZN(n10471) );
  OAI221_X1 U11572 ( .B1(n9269), .B2(keyinput52), .C1(n9745), .C2(keyinput21), 
        .A(n10471), .ZN(n10478) );
  XNOR2_X1 U11573 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput126), .ZN(n10474) );
  XNOR2_X1 U11574 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput37), .ZN(n10473) );
  XNOR2_X1 U11575 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput31), .ZN(n10472)
         );
  NAND3_X1 U11576 ( .A1(n10474), .A2(n10473), .A3(n10472), .ZN(n10477) );
  XNOR2_X1 U11577 ( .A(n10475), .B(keyinput125), .ZN(n10476) );
  NOR4_X1 U11578 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10480) );
  NAND4_X1 U11579 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10668) );
  AOI22_X1 U11580 ( .A1(n10486), .A2(keyinput113), .B1(keyinput94), .B2(n10485), .ZN(n10484) );
  OAI221_X1 U11581 ( .B1(n10486), .B2(keyinput113), .C1(n10485), .C2(
        keyinput94), .A(n10484), .ZN(n10498) );
  AOI22_X1 U11582 ( .A1(n10489), .A2(keyinput111), .B1(keyinput70), .B2(n10488), .ZN(n10487) );
  OAI221_X1 U11583 ( .B1(n10489), .B2(keyinput111), .C1(n10488), .C2(
        keyinput70), .A(n10487), .ZN(n10497) );
  AOI22_X1 U11584 ( .A1(n10492), .A2(keyinput50), .B1(keyinput18), .B2(n10491), 
        .ZN(n10490) );
  OAI221_X1 U11585 ( .B1(n10492), .B2(keyinput50), .C1(n10491), .C2(keyinput18), .A(n10490), .ZN(n10496) );
  XNOR2_X1 U11586 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput89), .ZN(n10494)
         );
  XNOR2_X1 U11587 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput47), .ZN(n10493)
         );
  NAND2_X1 U11588 ( .A1(n10494), .A2(n10493), .ZN(n10495) );
  NOR4_X1 U11589 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10543) );
  AOI22_X1 U11590 ( .A1(n10501), .A2(keyinput98), .B1(keyinput29), .B2(n10500), 
        .ZN(n10499) );
  OAI221_X1 U11591 ( .B1(n10501), .B2(keyinput98), .C1(n10500), .C2(keyinput29), .A(n10499), .ZN(n10512) );
  INV_X1 U11592 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U11593 ( .A1(n10503), .A2(keyinput17), .B1(n5597), .B2(keyinput86), 
        .ZN(n10502) );
  OAI221_X1 U11594 ( .B1(n10503), .B2(keyinput17), .C1(n5597), .C2(keyinput86), 
        .A(n10502), .ZN(n10511) );
  AOI22_X1 U11595 ( .A1(n10506), .A2(keyinput77), .B1(keyinput103), .B2(n10505), .ZN(n10504) );
  OAI221_X1 U11596 ( .B1(n10506), .B2(keyinput77), .C1(n10505), .C2(
        keyinput103), .A(n10504), .ZN(n10510) );
  XNOR2_X1 U11597 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput68), .ZN(n10508)
         );
  XNOR2_X1 U11598 ( .A(SI_28_), .B(keyinput41), .ZN(n10507) );
  NAND2_X1 U11599 ( .A1(n10508), .A2(n10507), .ZN(n10509) );
  NOR4_X1 U11600 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10542) );
  AOI22_X1 U11601 ( .A1(n10515), .A2(keyinput14), .B1(n10514), .B2(keyinput67), 
        .ZN(n10513) );
  OAI221_X1 U11602 ( .B1(n10515), .B2(keyinput14), .C1(n10514), .C2(keyinput67), .A(n10513), .ZN(n10524) );
  AOI22_X1 U11603 ( .A1(n5936), .A2(keyinput88), .B1(keyinput9), .B2(n10517), 
        .ZN(n10516) );
  OAI221_X1 U11604 ( .B1(n5936), .B2(keyinput88), .C1(n10517), .C2(keyinput9), 
        .A(n10516), .ZN(n10523) );
  AOI22_X1 U11605 ( .A1(n10520), .A2(keyinput66), .B1(n10519), .B2(keyinput10), 
        .ZN(n10518) );
  OAI221_X1 U11606 ( .B1(n10520), .B2(keyinput66), .C1(n10519), .C2(keyinput10), .A(n10518), .ZN(n10522) );
  XOR2_X1 U11607 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput43), .Z(n10521) );
  NOR4_X1 U11608 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10527) );
  XOR2_X1 U11609 ( .A(keyinput123), .B(n10525), .Z(n10526) );
  AND2_X1 U11610 ( .A1(n10527), .A2(n10526), .ZN(n10541) );
  AOI22_X1 U11611 ( .A1(n10529), .A2(keyinput82), .B1(n6012), .B2(keyinput59), 
        .ZN(n10528) );
  OAI221_X1 U11612 ( .B1(n10529), .B2(keyinput82), .C1(n6012), .C2(keyinput59), 
        .A(n10528), .ZN(n10539) );
  AOI22_X1 U11613 ( .A1(n8847), .A2(keyinput127), .B1(n5138), .B2(keyinput6), 
        .ZN(n10530) );
  OAI221_X1 U11614 ( .B1(n8847), .B2(keyinput127), .C1(n5138), .C2(keyinput6), 
        .A(n10530), .ZN(n10538) );
  AOI22_X1 U11615 ( .A1(n10532), .A2(keyinput46), .B1(keyinput63), .B2(n8770), 
        .ZN(n10531) );
  OAI221_X1 U11616 ( .B1(n10532), .B2(keyinput46), .C1(n8770), .C2(keyinput63), 
        .A(n10531), .ZN(n10537) );
  AOI22_X1 U11617 ( .A1(n10535), .A2(keyinput27), .B1(keyinput39), .B2(n10534), 
        .ZN(n10533) );
  OAI221_X1 U11618 ( .B1(n10535), .B2(keyinput27), .C1(n10534), .C2(keyinput39), .A(n10533), .ZN(n10536) );
  NOR4_X1 U11619 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10540) );
  NAND4_X1 U11620 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10667) );
  AOI22_X1 U11621 ( .A1(n10546), .A2(keyinput71), .B1(n10545), .B2(keyinput62), 
        .ZN(n10544) );
  OAI221_X1 U11622 ( .B1(n10546), .B2(keyinput71), .C1(n10545), .C2(keyinput62), .A(n10544), .ZN(n10558) );
  AOI22_X1 U11623 ( .A1(n10549), .A2(keyinput4), .B1(keyinput124), .B2(n10548), 
        .ZN(n10547) );
  OAI221_X1 U11624 ( .B1(n10549), .B2(keyinput4), .C1(n10548), .C2(keyinput124), .A(n10547), .ZN(n10557) );
  AOI22_X1 U11625 ( .A1(n10552), .A2(keyinput16), .B1(keyinput90), .B2(n10551), 
        .ZN(n10550) );
  OAI221_X1 U11626 ( .B1(n10552), .B2(keyinput16), .C1(n10551), .C2(keyinput90), .A(n10550), .ZN(n10556) );
  AOI22_X1 U11627 ( .A1(n7244), .A2(keyinput32), .B1(n10554), .B2(keyinput42), 
        .ZN(n10553) );
  OAI221_X1 U11628 ( .B1(n7244), .B2(keyinput32), .C1(n10554), .C2(keyinput42), 
        .A(n10553), .ZN(n10555) );
  NOR4_X1 U11629 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10604) );
  AOI22_X1 U11630 ( .A1(n10560), .A2(keyinput105), .B1(keyinput76), .B2(n5983), 
        .ZN(n10559) );
  OAI221_X1 U11631 ( .B1(n10560), .B2(keyinput105), .C1(n5983), .C2(keyinput76), .A(n10559), .ZN(n10571) );
  AOI22_X1 U11632 ( .A1(n10563), .A2(keyinput78), .B1(keyinput57), .B2(n10562), 
        .ZN(n10561) );
  OAI221_X1 U11633 ( .B1(n10563), .B2(keyinput78), .C1(n10562), .C2(keyinput57), .A(n10561), .ZN(n10570) );
  AOI22_X1 U11634 ( .A1(n10566), .A2(keyinput48), .B1(keyinput30), .B2(n10565), 
        .ZN(n10564) );
  OAI221_X1 U11635 ( .B1(n10566), .B2(keyinput48), .C1(n10565), .C2(keyinput30), .A(n10564), .ZN(n10569) );
  AOI22_X1 U11636 ( .A1(n6344), .A2(keyinput36), .B1(keyinput25), .B2(n7979), 
        .ZN(n10567) );
  OAI221_X1 U11637 ( .B1(n6344), .B2(keyinput36), .C1(n7979), .C2(keyinput25), 
        .A(n10567), .ZN(n10568) );
  NOR4_X1 U11638 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10603) );
  AOI22_X1 U11639 ( .A1(n10574), .A2(keyinput101), .B1(n10573), .B2(keyinput99), .ZN(n10572) );
  OAI221_X1 U11640 ( .B1(n10574), .B2(keyinput101), .C1(n10573), .C2(
        keyinput99), .A(n10572), .ZN(n10584) );
  AOI22_X1 U11641 ( .A1(n10577), .A2(keyinput7), .B1(n10576), .B2(keyinput92), 
        .ZN(n10575) );
  OAI221_X1 U11642 ( .B1(n10577), .B2(keyinput7), .C1(n10576), .C2(keyinput92), 
        .A(n10575), .ZN(n10583) );
  XOR2_X1 U11643 ( .A(n10391), .B(keyinput65), .Z(n10581) );
  XNOR2_X1 U11644 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput19), .ZN(n10580) );
  XNOR2_X1 U11645 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput56), .ZN(n10579)
         );
  XNOR2_X1 U11646 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput44), .ZN(n10578) );
  NAND4_X1 U11647 ( .A1(n10581), .A2(n10580), .A3(n10579), .A4(n10578), .ZN(
        n10582) );
  NOR3_X1 U11648 ( .A1(n10584), .A2(n10583), .A3(n10582), .ZN(n10602) );
  INV_X1 U11649 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U11650 ( .A1(n10587), .A2(keyinput80), .B1(n10586), .B2(keyinput69), 
        .ZN(n10585) );
  OAI221_X1 U11651 ( .B1(n10587), .B2(keyinput80), .C1(n10586), .C2(keyinput69), .A(n10585), .ZN(n10600) );
  AOI22_X1 U11652 ( .A1(n10590), .A2(keyinput74), .B1(n10589), .B2(keyinput55), 
        .ZN(n10588) );
  OAI221_X1 U11653 ( .B1(n10590), .B2(keyinput74), .C1(n10589), .C2(keyinput55), .A(n10588), .ZN(n10599) );
  AOI22_X1 U11654 ( .A1(n10593), .A2(keyinput51), .B1(keyinput35), .B2(n10592), 
        .ZN(n10591) );
  OAI221_X1 U11655 ( .B1(n10593), .B2(keyinput51), .C1(n10592), .C2(keyinput35), .A(n10591), .ZN(n10598) );
  AOI22_X1 U11656 ( .A1(n10596), .A2(keyinput110), .B1(n10595), .B2(keyinput0), 
        .ZN(n10594) );
  OAI221_X1 U11657 ( .B1(n10596), .B2(keyinput110), .C1(n10595), .C2(keyinput0), .A(n10594), .ZN(n10597) );
  NOR4_X1 U11658 ( .A1(n10600), .A2(n10599), .A3(n10598), .A4(n10597), .ZN(
        n10601) );
  NAND4_X1 U11659 ( .A1(n10604), .A2(n10603), .A3(n10602), .A4(n10601), .ZN(
        n10666) );
  AOI22_X1 U11660 ( .A1(n10607), .A2(keyinput33), .B1(n10606), .B2(keyinput61), 
        .ZN(n10605) );
  OAI221_X1 U11661 ( .B1(n10607), .B2(keyinput33), .C1(n10606), .C2(keyinput61), .A(n10605), .ZN(n10619) );
  AOI22_X1 U11662 ( .A1(n10610), .A2(keyinput115), .B1(keyinput60), .B2(n10609), .ZN(n10608) );
  OAI221_X1 U11663 ( .B1(n10610), .B2(keyinput115), .C1(n10609), .C2(
        keyinput60), .A(n10608), .ZN(n10618) );
  AOI22_X1 U11664 ( .A1(n10613), .A2(keyinput102), .B1(n10612), .B2(keyinput64), .ZN(n10611) );
  OAI221_X1 U11665 ( .B1(n10613), .B2(keyinput102), .C1(n10612), .C2(
        keyinput64), .A(n10611), .ZN(n10617) );
  XNOR2_X1 U11666 ( .A(SI_3_), .B(keyinput28), .ZN(n10615) );
  XNOR2_X1 U11667 ( .A(SI_13_), .B(keyinput11), .ZN(n10614) );
  NAND2_X1 U11668 ( .A1(n10615), .A2(n10614), .ZN(n10616) );
  NOR4_X1 U11669 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10664) );
  AOI22_X1 U11670 ( .A1(keyinput119), .A2(n10621), .B1(keyinput114), .B2(n6341), .ZN(n10620) );
  OAI21_X1 U11671 ( .B1(n10621), .B2(keyinput119), .A(n10620), .ZN(n10632) );
  AOI22_X1 U11672 ( .A1(n10624), .A2(keyinput73), .B1(n10623), .B2(keyinput15), 
        .ZN(n10622) );
  OAI221_X1 U11673 ( .B1(n10624), .B2(keyinput73), .C1(n10623), .C2(keyinput15), .A(n10622), .ZN(n10631) );
  XNOR2_X1 U11674 ( .A(n10625), .B(keyinput26), .ZN(n10630) );
  XNOR2_X1 U11675 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput95), .ZN(n10628) );
  XNOR2_X1 U11676 ( .A(P1_REG0_REG_26__SCAN_IN), .B(keyinput109), .ZN(n10627)
         );
  XNOR2_X1 U11677 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput79), .ZN(n10626) );
  NAND3_X1 U11678 ( .A1(n10628), .A2(n10627), .A3(n10626), .ZN(n10629) );
  NOR4_X1 U11679 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10663) );
  AOI22_X1 U11680 ( .A1(n10634), .A2(keyinput108), .B1(keyinput97), .B2(n6328), 
        .ZN(n10633) );
  OAI221_X1 U11681 ( .B1(n10634), .B2(keyinput108), .C1(n6328), .C2(keyinput97), .A(n10633), .ZN(n10644) );
  AOI22_X1 U11682 ( .A1(n10637), .A2(keyinput5), .B1(keyinput38), .B2(n10636), 
        .ZN(n10635) );
  OAI221_X1 U11683 ( .B1(n10637), .B2(keyinput5), .C1(n10636), .C2(keyinput38), 
        .A(n10635), .ZN(n10643) );
  XOR2_X1 U11684 ( .A(n10294), .B(keyinput107), .Z(n10641) );
  XOR2_X1 U11685 ( .A(n5367), .B(keyinput12), .Z(n10640) );
  XNOR2_X1 U11686 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput1), .ZN(n10639) );
  XNOR2_X1 U11687 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput22), .ZN(n10638)
         );
  NAND4_X1 U11688 ( .A1(n10641), .A2(n10640), .A3(n10639), .A4(n10638), .ZN(
        n10642) );
  NOR3_X1 U11689 ( .A1(n10644), .A2(n10643), .A3(n10642), .ZN(n10662) );
  AOI22_X1 U11690 ( .A1(n10647), .A2(keyinput91), .B1(keyinput40), .B2(n10646), 
        .ZN(n10645) );
  OAI221_X1 U11691 ( .B1(n10647), .B2(keyinput91), .C1(n10646), .C2(keyinput40), .A(n10645), .ZN(n10660) );
  AOI22_X1 U11692 ( .A1(n10650), .A2(keyinput117), .B1(keyinput120), .B2(
        n10649), .ZN(n10648) );
  OAI221_X1 U11693 ( .B1(n10650), .B2(keyinput117), .C1(n10649), .C2(
        keyinput120), .A(n10648), .ZN(n10659) );
  AOI22_X1 U11694 ( .A1(n10653), .A2(keyinput106), .B1(keyinput81), .B2(n10652), .ZN(n10651) );
  OAI221_X1 U11695 ( .B1(n10653), .B2(keyinput106), .C1(n10652), .C2(
        keyinput81), .A(n10651), .ZN(n10658) );
  AOI22_X1 U11696 ( .A1(n10656), .A2(keyinput23), .B1(keyinput13), .B2(n10655), 
        .ZN(n10654) );
  OAI221_X1 U11697 ( .B1(n10656), .B2(keyinput23), .C1(n10655), .C2(keyinput13), .A(n10654), .ZN(n10657) );
  NOR4_X1 U11698 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10661) );
  NAND4_X1 U11699 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10665) );
  NOR4_X1 U11700 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10669) );
  OAI21_X1 U11701 ( .B1(keyinput114), .B2(n10670), .A(n10669), .ZN(n10674) );
  AOI22_X1 U11702 ( .A1(n10672), .A2(n10671), .B1(n4588), .B2(n8960), .ZN(
        n10673) );
  XNOR2_X1 U11703 ( .A(n10674), .B(n10673), .ZN(P2_U3460) );
  OAI21_X1 U11704 ( .B1(n10677), .B2(n10676), .A(n10675), .ZN(ADD_1068_U50) );
  OAI21_X1 U11705 ( .B1(n10680), .B2(n10679), .A(n10678), .ZN(ADD_1068_U51) );
  OAI21_X1 U11706 ( .B1(n10683), .B2(n10682), .A(n10681), .ZN(ADD_1068_U47) );
  OAI21_X1 U11707 ( .B1(n10686), .B2(n10685), .A(n10684), .ZN(ADD_1068_U49) );
  OAI21_X1 U11708 ( .B1(n10689), .B2(n10688), .A(n10687), .ZN(ADD_1068_U48) );
  AOI21_X1 U11709 ( .B1(n10692), .B2(n10691), .A(n10690), .ZN(ADD_1068_U54) );
  AOI21_X1 U11710 ( .B1(n10695), .B2(n10694), .A(n10693), .ZN(ADD_1068_U53) );
  OAI21_X1 U11711 ( .B1(n10698), .B2(n10697), .A(n10696), .ZN(ADD_1068_U52) );
  OR2_X1 U5007 ( .A1(n9735), .A2(n9750), .ZN(n9483) );
  OR2_X2 U5086 ( .A1(n9744), .A2(n4426), .ZN(n9731) );
  CLKBUF_X1 U5147 ( .A(n8370), .Z(n4579) );
  CLKBUF_X1 U5468 ( .A(n9160), .Z(n4598) );
  CLKBUF_X2 U5581 ( .A(n6512), .Z(n7122) );
  CLKBUF_X1 U6434 ( .A(n9787), .Z(n4584) );
endmodule

