

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291;

  NAND2_X1 U4906 ( .A1(n5328), .A2(n8694), .ZN(n7540) );
  CLKBUF_X1 U4907 ( .A(n5460), .Z(n5657) );
  INV_X1 U4908 ( .A(n7589), .ZN(n5639) );
  CLKBUF_X2 U4909 ( .A(n5210), .Z(n5631) );
  INV_X1 U4910 ( .A(n5889), .ZN(n6244) );
  INV_X1 U4912 ( .A(n7885), .ZN(n4660) );
  CLKBUF_X2 U4913 ( .A(n6734), .Z(n7118) );
  OR2_X1 U4915 ( .A1(n6136), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6146) );
  INV_X1 U4916 ( .A(n8078), .ZN(n8083) );
  NAND2_X1 U4917 ( .A1(n5594), .A2(n8614), .ZN(n8617) );
  OAI21_X1 U4918 ( .B1(n8730), .B2(n8732), .A(n5450), .ZN(n8646) );
  OR2_X1 U4919 ( .A1(n9479), .A2(n4798), .ZN(n4797) );
  AND4_X1 U4920 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), .ZN(n7086)
         );
  AND2_X1 U4921 ( .A1(n7473), .A2(n7472), .ZN(n4400) );
  NAND2_X1 U4923 ( .A1(n5135), .A2(n6433), .ZN(n4401) );
  NAND2_X1 U4924 ( .A1(n5135), .A2(n6433), .ZN(n7589) );
  OR2_X2 U4925 ( .A1(n9173), .A2(n4846), .ZN(n4844) );
  NAND2_X1 U4926 ( .A1(n5719), .A2(n4401), .ZN(n5165) );
  NAND2_X2 U4927 ( .A1(n5327), .A2(n5326), .ZN(n8694) );
  AOI21_X2 U4928 ( .B1(n8563), .B2(n8665), .A(n5675), .ZN(n5676) );
  NAND2_X2 U4929 ( .A1(n4960), .A2(n4481), .ZN(n8563) );
  OAI21_X2 U4930 ( .B1(n4447), .B2(n9147), .A(n9141), .ZN(n9331) );
  XOR2_X2 U4931 ( .A(n6370), .B(n6890), .Z(n4502) );
  NAND4_X2 U4932 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n9569)
         );
  AND2_X1 U4933 ( .A1(n6433), .A2(n5083), .ZN(n4402) );
  NAND4_X2 U4934 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n8990)
         );
  OAI22_X2 U4935 ( .A1(n8319), .A2(n6048), .B1(n7926), .B2(n8514), .ZN(n8306)
         );
  BUF_X1 U4936 ( .A(n6694), .Z(n4403) );
  AND2_X4 U4937 ( .A1(n4564), .A2(n4565), .ZN(n7885) );
  OAI21_X2 U4938 ( .B1(n9108), .B2(n5038), .A(n9107), .ZN(n9228) );
  NAND2_X2 U4939 ( .A1(n4787), .A2(n4786), .ZN(n9108) );
  NOR2_X2 U4940 ( .A1(n5966), .A2(n4408), .ZN(n5996) );
  NOR2_X2 U4941 ( .A1(n7091), .A2(n4691), .ZN(n4694) );
  AND2_X4 U4942 ( .A1(n5815), .A2(n7685), .ZN(n5889) );
  NAND2_X1 U4943 ( .A1(n7855), .A2(n7856), .ZN(n7854) );
  NAND2_X1 U4944 ( .A1(n7867), .A2(n5002), .ZN(n7777) );
  OAI22_X1 U4945 ( .A1(n7814), .A2(n7813), .B1(n7647), .B2(n8371), .ZN(n7708)
         );
  NAND2_X1 U4946 ( .A1(n6135), .A2(n6134), .ZN(n8474) );
  NAND2_X1 U4947 ( .A1(n5019), .A2(n7752), .ZN(n7814) );
  OR2_X1 U4948 ( .A1(n8713), .A2(n5190), .ZN(n4954) );
  INV_X1 U4949 ( .A(n5165), .ZN(n5666) );
  INV_X1 U4950 ( .A(n9594), .ZN(n7148) );
  INV_X1 U4951 ( .A(n9585), .ZN(n7085) );
  AND4_X1 U4952 ( .A1(n5233), .A2(n5232), .A3(n5231), .A4(n5230), .ZN(n9605)
         );
  INV_X1 U4953 ( .A(n6880), .ZN(n7141) );
  INV_X1 U4954 ( .A(n6433), .ZN(n5754) );
  NAND4_X1 U4955 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n8111)
         );
  CLKBUF_X2 U4956 ( .A(n5159), .Z(n8992) );
  CLKBUF_X2 U4957 ( .A(n5862), .Z(n5896) );
  INV_X1 U4958 ( .A(n7913), .ZN(n4512) );
  BUF_X1 U4959 ( .A(n5060), .Z(n7620) );
  XNOR2_X1 U4960 ( .A(n5088), .B(n5087), .ZN(n5159) );
  XNOR2_X1 U4961 ( .A(n5059), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5060) );
  OR2_X1 U4962 ( .A1(n6365), .A2(n9724), .ZN(n4713) );
  NAND2_X1 U4963 ( .A1(n8812), .A2(n8811), .ZN(n8827) );
  NAND2_X1 U4964 ( .A1(n7854), .A2(n4446), .ZN(n7700) );
  AND2_X1 U4965 ( .A1(n4532), .A2(n4533), .ZN(n4531) );
  NAND2_X1 U4966 ( .A1(n4736), .A2(n4735), .ZN(n8172) );
  NOR3_X1 U4967 ( .A1(n8070), .A2(n8069), .A3(n8068), .ZN(n8071) );
  AOI21_X1 U4968 ( .B1(n7742), .B2(n5006), .A(n5004), .ZN(n5003) );
  OAI21_X1 U4969 ( .B1(n8194), .B2(n6232), .A(n6233), .ZN(n8181) );
  NAND2_X1 U4970 ( .A1(n5005), .A2(n7770), .ZN(n5004) );
  NAND2_X1 U4971 ( .A1(n6231), .A2(n6230), .ZN(n8194) );
  NAND2_X1 U4972 ( .A1(n5006), .A2(n5008), .ZN(n5005) );
  OAI21_X1 U4973 ( .B1(n8273), .B2(n4762), .A(n4760), .ZN(n6124) );
  OR2_X1 U4974 ( .A1(n8130), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U4975 ( .A1(n7869), .A2(n7868), .ZN(n7867) );
  INV_X1 U4976 ( .A(n4761), .ZN(n4760) );
  XNOR2_X1 U4977 ( .A(n5649), .B(n5648), .ZN(n7509) );
  NAND2_X1 U4978 ( .A1(n7397), .A2(n4528), .ZN(n5327) );
  NAND2_X1 U4979 ( .A1(n4766), .A2(n4764), .ZN(n8343) );
  NAND2_X1 U4980 ( .A1(n7362), .A2(n7363), .ZN(n7473) );
  NAND2_X1 U4981 ( .A1(n5512), .A2(n5511), .ZN(n5579) );
  NAND2_X1 U4982 ( .A1(n7376), .A2(n7638), .ZN(n8361) );
  OR2_X1 U4983 ( .A1(n7485), .A2(n6376), .ZN(n6379) );
  NAND2_X1 U4984 ( .A1(n7278), .A2(n7976), .ZN(n9911) );
  AOI21_X1 U4985 ( .B1(n6221), .B2(n6220), .A(n6219), .ZN(n7278) );
  NAND2_X1 U4986 ( .A1(n4954), .A2(n4950), .ZN(n4952) );
  NAND2_X1 U4987 ( .A1(n5430), .A2(n5429), .ZN(n5432) );
  AND2_X1 U4988 ( .A1(n4721), .A2(n4722), .ZN(n6373) );
  AND2_X1 U4989 ( .A1(n7238), .A2(n7235), .ZN(n5018) );
  NAND2_X1 U4990 ( .A1(n5755), .A2(n8970), .ZN(n8742) );
  INV_X2 U4991 ( .A(n5666), .ZN(n8593) );
  INV_X2 U4992 ( .A(n9672), .ZN(n4404) );
  OR2_X1 U4993 ( .A1(n6029), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6042) );
  INV_X2 U4994 ( .A(n6508), .ZN(n6674) );
  INV_X1 U4995 ( .A(n5666), .ZN(n4405) );
  INV_X1 U4996 ( .A(n9565), .ZN(n8919) );
  AND2_X1 U4997 ( .A1(n5133), .A2(n5132), .ZN(n5719) );
  AND3_X1 U4998 ( .A1(n5199), .A2(n5198), .A3(n5197), .ZN(n9579) );
  NAND4_X2 U4999 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n9586)
         );
  NAND3_X1 U5000 ( .A1(n6727), .A2(n6728), .A3(n4511), .ZN(n6734) );
  INV_X1 U5001 ( .A(n6947), .ZN(n9560) );
  OR2_X1 U5002 ( .A1(n5754), .A2(n8969), .ZN(n5133) );
  AND2_X1 U5003 ( .A1(n5175), .A2(n4657), .ZN(n7026) );
  NAND2_X1 U5004 ( .A1(n5461), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5152) );
  NAND2_X2 U5005 ( .A1(n6437), .A2(n7885), .ZN(n8823) );
  CLKBUF_X3 U5006 ( .A(n5461), .Z(n5661) );
  AND3_X1 U5007 ( .A1(n5883), .A2(n5882), .A3(n5881), .ZN(n7263) );
  OR2_X2 U5008 ( .A1(n8092), .A2(n7913), .ZN(n8078) );
  NAND2_X1 U5009 ( .A1(n6204), .A2(n6269), .ZN(n8092) );
  NAND2_X1 U5010 ( .A1(n6090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U5011 ( .A1(n5076), .A2(n5725), .ZN(n6433) );
  NAND2_X2 U5012 ( .A1(n5159), .A2(n5160), .ZN(n6437) );
  AND2_X1 U5013 ( .A1(n5070), .A2(n5086), .ZN(n5725) );
  NAND4_X1 U5014 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n8112)
         );
  NAND4_X2 U5015 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n9884)
         );
  NAND2_X1 U5016 ( .A1(n5546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U5017 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5082) );
  NOR2_X1 U5018 ( .A1(n5356), .A2(n4936), .ZN(n4935) );
  NAND2_X1 U5019 ( .A1(n5128), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U5020 ( .A1(n5073), .A2(n5069), .ZN(n7574) );
  NAND2_X1 U5021 ( .A1(n5075), .A2(n4437), .ZN(n7568) );
  NAND2_X1 U5022 ( .A1(n6239), .A2(n6240), .ZN(n5862) );
  XNOR2_X1 U5023 ( .A(n6206), .B(n6205), .ZN(n7913) );
  CLKBUF_X3 U5024 ( .A(n6240), .Z(n8548) );
  OR2_X1 U5025 ( .A1(n9404), .A2(n9406), .ZN(n5056) );
  OR2_X1 U5026 ( .A1(n4436), .A2(n5813), .ZN(n6206) );
  XNOR2_X1 U5027 ( .A(n6257), .B(n6256), .ZN(n7571) );
  MUX2_X1 U5028 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5832), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5833) );
  NAND2_X1 U5029 ( .A1(n5057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5085) );
  INV_X1 U5030 ( .A(n5816), .ZN(n7685) );
  AND2_X1 U5031 ( .A1(n4536), .A2(n4535), .ZN(n5838) );
  NOR2_X1 U5032 ( .A1(n6199), .A2(n6198), .ZN(n6207) );
  OR2_X1 U5033 ( .A1(n5831), .A2(n5813), .ZN(n5814) );
  AND2_X1 U5034 ( .A1(n5996), .A2(n5995), .ZN(n6013) );
  AND2_X1 U5035 ( .A1(n5359), .A2(n10227), .ZN(n5361) );
  INV_X1 U5036 ( .A(n7885), .ZN(n5104) );
  CLKBUF_X1 U5037 ( .A(n5089), .Z(n5255) );
  NAND2_X1 U5038 ( .A1(n5917), .A2(n4783), .ZN(n5966) );
  AND2_X1 U5039 ( .A1(n4434), .A2(n5052), .ZN(n5071) );
  NAND2_X1 U5040 ( .A1(n4870), .A2(n5860), .ZN(n9703) );
  NAND3_X1 U5041 ( .A1(n4949), .A2(n5174), .A3(n5040), .ZN(n5089) );
  AND2_X2 U5042 ( .A1(n5897), .A2(n5913), .ZN(n5917) );
  AND3_X1 U5043 ( .A1(n5802), .A2(n5804), .A3(n5803), .ZN(n4537) );
  AND3_X1 U5044 ( .A1(n5801), .A2(n6050), .A3(n5800), .ZN(n5805) );
  AND2_X1 U5045 ( .A1(n4784), .A2(n5798), .ZN(n4783) );
  AND3_X1 U5046 ( .A1(n4772), .A2(n4771), .A3(n5855), .ZN(n5897) );
  NAND2_X1 U5047 ( .A1(n5809), .A2(n5024), .ZN(n5023) );
  NOR2_X1 U5048 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9415) );
  INV_X1 U5049 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5275) );
  INV_X4 U5050 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X2 U5051 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5174) );
  INV_X1 U5052 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4947) );
  NOR2_X1 U5053 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5041) );
  NOR2_X1 U5054 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5042) );
  NOR2_X1 U5055 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5043) );
  INV_X1 U5056 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5798) );
  INV_X1 U5057 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5129) );
  INV_X1 U5058 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6205) );
  NOR2_X1 U5059 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4784) );
  NOR2_X1 U5060 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4772) );
  INV_X1 U5061 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6200) );
  NOR2_X1 U5062 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4771) );
  INV_X1 U5063 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5055) );
  OAI21_X2 U5064 ( .B1(n9228), .B2(n4823), .A(n4821), .ZN(n9187) );
  AND2_X1 U5065 ( .A1(n7117), .A2(n7116), .ZN(n4406) );
  BUF_X1 U5066 ( .A(n7742), .Z(n4407) );
  OR2_X1 U5067 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4408) );
  CLKBUF_X1 U5068 ( .A(n6089), .Z(n4409) );
  OAI21_X1 U5069 ( .B1(n7787), .B2(n7786), .A(n7785), .ZN(n4410) );
  OAI22_X1 U5070 ( .A1(n7814), .A2(n7813), .B1(n7647), .B2(n8371), .ZN(n4411)
         );
  AOI21_X2 U5071 ( .B1(n6991), .B2(n6990), .A(n6989), .ZN(n7117) );
  NAND2_X1 U5072 ( .A1(n7741), .A2(n7743), .ZN(n7742) );
  OAI21_X1 U5073 ( .B1(n7787), .B2(n7786), .A(n7785), .ZN(n7784) );
  NAND2_X1 U5074 ( .A1(n6906), .A2(n6905), .ZN(n6984) );
  NAND2_X1 U5075 ( .A1(n6852), .A2(n6851), .ZN(n6906) );
  AND3_X1 U5076 ( .A1(n4782), .A2(n5808), .A3(n5917), .ZN(n6259) );
  XNOR2_X2 U5077 ( .A(n5812), .B(n5811), .ZN(n5815) );
  NAND2_X1 U5078 ( .A1(n6736), .A2(n6737), .ZN(n6798) );
  AND2_X1 U5079 ( .A1(n6733), .A2(n6797), .ZN(n6736) );
  XNOR2_X1 U5080 ( .A(n5856), .B(n5855), .ZN(n9724) );
  NOR2_X1 U5081 ( .A1(n5966), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5982) );
  NOR2_X2 U5082 ( .A1(n6053), .A2(n6052), .ZN(n6067) );
  XNOR2_X2 U5083 ( .A(n7668), .B(n7669), .ZN(n7855) );
  NAND2_X2 U5084 ( .A1(n7773), .A2(n7666), .ZN(n7668) );
  XNOR2_X1 U5085 ( .A(n6734), .B(n6880), .ZN(n6732) );
  OAI21_X2 U5086 ( .B1(n6077), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6089) );
  NAND2_X2 U5087 ( .A1(n6237), .A2(n8088), .ZN(n6728) );
  XNOR2_X2 U5088 ( .A(n6091), .B(n5800), .ZN(n6237) );
  AOI21_X1 U5089 ( .B1(n8034), .B2(n8078), .A(n8039), .ZN(n4525) );
  INV_X1 U5090 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U5091 ( .A1(n5681), .A2(n5680), .ZN(n5703) );
  OR2_X1 U5092 ( .A1(n6757), .A2(n4855), .ZN(n4851) );
  NAND2_X1 U5093 ( .A1(n5862), .A2(n7885), .ZN(n5865) );
  NAND2_X1 U5094 ( .A1(n8827), .A2(n4438), .ZN(n4539) );
  INV_X1 U5095 ( .A(n8769), .ZN(n4684) );
  NAND2_X1 U5096 ( .A1(n4523), .A2(n8038), .ZN(n8043) );
  NAND2_X1 U5097 ( .A1(n4525), .A2(n4524), .ZN(n4523) );
  AND2_X1 U5098 ( .A1(n8071), .A2(n8072), .ZN(n8082) );
  NOR2_X1 U5099 ( .A1(n8101), .A2(n4908), .ZN(n4907) );
  INV_X1 U5100 ( .A(n6190), .ZN(n4908) );
  INV_X1 U5101 ( .A(n4986), .ZN(n4985) );
  INV_X1 U5102 ( .A(n4995), .ZN(n4993) );
  NAND2_X1 U5103 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  OR2_X1 U5104 ( .A1(n5988), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6004) );
  OR2_X1 U5105 ( .A1(n5972), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U5106 ( .A1(n4752), .A2(n4749), .ZN(n4748) );
  INV_X1 U5107 ( .A(n4741), .ZN(n4740) );
  OR2_X1 U5108 ( .A1(n8468), .A2(n7764), .ZN(n8047) );
  OR2_X1 U5109 ( .A1(n8279), .A2(n8284), .ZN(n8028) );
  INV_X1 U5110 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U5111 ( .A1(n6013), .A2(n6012), .ZN(n6053) );
  OR2_X1 U5112 ( .A1(n9335), .A2(n9325), .ZN(n8952) );
  AND2_X1 U5113 ( .A1(n4845), .A2(n4843), .ZN(n4842) );
  OR2_X1 U5114 ( .A1(n9322), .A2(n8809), .ZN(n8899) );
  NAND2_X1 U5115 ( .A1(n4612), .A2(n5830), .ZN(n4611) );
  INV_X1 U5116 ( .A(n6187), .ZN(n4612) );
  NAND2_X1 U5117 ( .A1(n5825), .A2(n5824), .ZN(n6172) );
  NAND2_X1 U5118 ( .A1(n5823), .A2(n5822), .ZN(n5825) );
  AND3_X1 U5119 ( .A1(n4989), .A2(n5045), .A3(n4988), .ZN(n4415) );
  INV_X1 U5120 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4988) );
  INV_X1 U5121 ( .A(n5048), .ZN(n4989) );
  NAND2_X1 U5122 ( .A1(n4590), .A2(n4588), .ZN(n5679) );
  AOI21_X1 U5123 ( .B1(n4591), .B2(n4596), .A(n4589), .ZN(n4588) );
  INV_X1 U5124 ( .A(n5650), .ZN(n4589) );
  OAI21_X1 U5125 ( .B1(n5501), .B2(n5500), .A(n5502), .ZN(n5542) );
  AOI21_X1 U5126 ( .B1(n4466), .B2(n5451), .A(n4928), .ZN(n4927) );
  NOR2_X1 U5127 ( .A1(n5431), .A2(SI_15_), .ZN(n4928) );
  AOI21_X1 U5128 ( .B1(n4586), .B2(n4931), .A(n5403), .ZN(n4585) );
  AOI21_X1 U5129 ( .B1(n5332), .B2(n4935), .A(n4934), .ZN(n4933) );
  INV_X1 U5130 ( .A(n5358), .ZN(n4934) );
  NAND2_X1 U5131 ( .A1(n5310), .A2(n5309), .ZN(n5333) );
  AND2_X1 U5132 ( .A1(n7734), .A2(n4443), .ZN(n4998) );
  AND2_X1 U5133 ( .A1(n7722), .A2(n8106), .ZN(n5022) );
  NAND2_X1 U5134 ( .A1(n4754), .A2(n5816), .ZN(n5868) );
  XNOR2_X1 U5135 ( .A(n6367), .B(n4855), .ZN(n9738) );
  NAND2_X1 U5136 ( .A1(n6397), .A2(n6754), .ZN(n6757) );
  AND2_X1 U5137 ( .A1(n6367), .A2(n6462), .ZN(n4734) );
  NAND2_X1 U5138 ( .A1(n4892), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4889) );
  INV_X1 U5139 ( .A(n7489), .ZN(n4892) );
  INV_X1 U5140 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U5141 ( .A1(n4621), .A2(n4624), .ZN(n8239) );
  AOI21_X1 U5142 ( .B1(n8036), .B2(n4626), .A(n4625), .ZN(n4624) );
  NAND2_X1 U5143 ( .A1(n6225), .A2(n4622), .ZN(n4621) );
  INV_X1 U5144 ( .A(n8035), .ZN(n4626) );
  NAND2_X1 U5145 ( .A1(n8368), .A2(n6010), .ZN(n4766) );
  NAND2_X1 U5146 ( .A1(n9911), .A2(n7972), .ZN(n4619) );
  NAND2_X1 U5147 ( .A1(n7271), .A2(n7907), .ZN(n4768) );
  NAND2_X1 U5148 ( .A1(n8450), .A2(n8185), .ZN(n6183) );
  XNOR2_X1 U5149 ( .A(n8444), .B(n8174), .ZN(n8165) );
  AND2_X1 U5150 ( .A1(n5037), .A2(n6133), .ZN(n4769) );
  AND4_X1 U5151 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n8310)
         );
  INV_X1 U5152 ( .A(n5865), .ZN(n7890) );
  AND2_X1 U5153 ( .A1(n4783), .A2(n4785), .ZN(n4782) );
  NOR2_X1 U5154 ( .A1(n5023), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4785) );
  NAND3_X1 U5155 ( .A1(n4967), .A2(n4965), .A3(n4964), .ZN(n8552) );
  NOR2_X1 U5156 ( .A1(n4966), .A2(n8555), .ZN(n4965) );
  INV_X1 U5157 ( .A(n4969), .ZN(n4966) );
  NAND2_X1 U5158 ( .A1(n5302), .A2(n4529), .ZN(n4528) );
  INV_X1 U5159 ( .A(n5305), .ZN(n4529) );
  NAND2_X1 U5160 ( .A1(n5647), .A2(n8686), .ZN(n4959) );
  INV_X1 U5161 ( .A(n8823), .ZN(n5548) );
  INV_X1 U5162 ( .A(n6437), .ZN(n5547) );
  OAI21_X1 U5163 ( .B1(n8827), .B2(n9098), .A(n4599), .ZN(n4598) );
  AND2_X1 U5164 ( .A1(n8973), .A2(n4600), .ZN(n4599) );
  AOI21_X1 U5165 ( .B1(n9098), .B2(n8831), .A(n4504), .ZN(n4600) );
  AND2_X1 U5166 ( .A1(n5737), .A2(n8918), .ZN(n8904) );
  NAND2_X1 U5167 ( .A1(n7697), .A2(n5061), .ZN(n8820) );
  NAND2_X1 U5168 ( .A1(n8816), .A2(n8815), .ZN(n8829) );
  OR2_X1 U5169 ( .A1(n9187), .A2(n9111), .ZN(n9113) );
  NAND2_X1 U5170 ( .A1(n9260), .A2(n9276), .ZN(n4786) );
  OR2_X1 U5171 ( .A1(n9255), .A2(n4788), .ZN(n4787) );
  AND2_X1 U5172 ( .A1(n9377), .A2(n9370), .ZN(n4788) );
  NAND2_X1 U5173 ( .A1(n9503), .A2(n9275), .ZN(n4796) );
  AND2_X1 U5174 ( .A1(n9488), .A2(n9299), .ZN(n4798) );
  NAND2_X1 U5175 ( .A1(n4467), .A2(n4818), .ZN(n4816) );
  NAND2_X1 U5176 ( .A1(n9619), .A2(n9627), .ZN(n7249) );
  AOI21_X1 U5177 ( .B1(n4694), .B2(n4690), .A(n4689), .ZN(n4692) );
  AND2_X1 U5178 ( .A1(n6449), .A2(n8904), .ZN(n9626) );
  NOR2_X1 U5179 ( .A1(n4946), .A2(n5618), .ZN(n4945) );
  INV_X1 U5180 ( .A(n5602), .ZN(n4946) );
  NAND2_X1 U5181 ( .A1(n4594), .A2(n5577), .ZN(n5581) );
  OR2_X1 U5182 ( .A1(n5579), .A2(n5578), .ZN(n4594) );
  NAND2_X1 U5183 ( .A1(n9414), .A2(n5093), .ZN(n4564) );
  INV_X1 U5184 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5093) );
  NAND2_X1 U5185 ( .A1(n6250), .A2(n6249), .ZN(n8156) );
  INV_X1 U5186 ( .A(n9356), .ZN(n9242) );
  NAND2_X1 U5187 ( .A1(n8755), .A2(n8826), .ZN(n4688) );
  AND2_X1 U5188 ( .A1(n8027), .A2(n8020), .ZN(n4521) );
  NAND2_X1 U5189 ( .A1(n4681), .A2(n4679), .ZN(n8771) );
  NAND2_X1 U5190 ( .A1(n4470), .A2(n4682), .ZN(n4681) );
  NOR2_X1 U5191 ( .A1(n4699), .A2(n8831), .ZN(n4698) );
  INV_X1 U5192 ( .A(n8943), .ZN(n4699) );
  NOR2_X1 U5193 ( .A1(n4490), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U5194 ( .A1(n8033), .A2(n8083), .ZN(n4524) );
  NAND2_X1 U5195 ( .A1(n8788), .A2(n4439), .ZN(n4678) );
  INV_X1 U5196 ( .A(n4916), .ZN(n4915) );
  OAI21_X1 U5197 ( .B1(n6171), .B2(n4917), .A(n6187), .ZN(n4916) );
  NOR2_X1 U5198 ( .A1(n4638), .A2(n8066), .ZN(n4636) );
  NAND2_X1 U5199 ( .A1(n4641), .A2(n4639), .ZN(n4638) );
  NAND2_X1 U5200 ( .A1(n7891), .A2(n4640), .ZN(n4639) );
  INV_X1 U5201 ( .A(n8081), .ZN(n4641) );
  INV_X1 U5202 ( .A(n6236), .ZN(n4640) );
  NAND2_X1 U5203 ( .A1(n7107), .A2(n7105), .ZN(n4986) );
  OR2_X1 U5204 ( .A1(n7107), .A2(n7105), .ZN(n4987) );
  NAND2_X1 U5205 ( .A1(n4582), .A2(n4581), .ZN(n4580) );
  NOR2_X1 U5206 ( .A1(n8803), .A2(n4706), .ZN(n4581) );
  NAND2_X1 U5207 ( .A1(n4541), .A2(n4455), .ZN(n4582) );
  NAND2_X1 U5208 ( .A1(n4708), .A2(n4707), .ZN(n4706) );
  AOI21_X1 U5209 ( .B1(n8804), .B2(n8889), .A(n8810), .ZN(n4705) );
  AND2_X1 U5210 ( .A1(n8805), .A2(n8831), .ZN(n8810) );
  NAND2_X1 U5211 ( .A1(n7183), .A2(n8850), .ZN(n8925) );
  AOI21_X1 U5212 ( .B1(n4595), .B2(n4593), .A(n4592), .ZN(n4591) );
  NOR2_X1 U5213 ( .A1(n5577), .A2(n5578), .ZN(n4593) );
  INV_X1 U5214 ( .A(n4940), .ZN(n4592) );
  INV_X1 U5215 ( .A(SI_11_), .ZN(n5334) );
  INV_X1 U5216 ( .A(SI_10_), .ZN(n10054) );
  NAND2_X1 U5217 ( .A1(n5012), .A2(n7824), .ZN(n5011) );
  INV_X1 U5218 ( .A(n5015), .ZN(n5012) );
  NAND2_X1 U5219 ( .A1(n8088), .A2(n4512), .ZN(n4511) );
  AOI21_X1 U5220 ( .B1(n5007), .B2(n5014), .A(n4462), .ZN(n5006) );
  OR2_X1 U5221 ( .A1(n8106), .A2(n9929), .ZN(n7989) );
  INV_X1 U5222 ( .A(n4739), .ZN(n4738) );
  OAI21_X1 U5223 ( .B1(n4740), .B2(n4742), .A(n6170), .ZN(n4739) );
  NAND2_X1 U5224 ( .A1(n7865), .A2(n7856), .ZN(n6170) );
  NAND2_X1 U5225 ( .A1(n4468), .A2(n4743), .ZN(n4741) );
  AND2_X1 U5226 ( .A1(n6227), .A2(n8208), .ZN(n6228) );
  OR2_X1 U5227 ( .A1(n8403), .A2(n8237), .ZN(n8040) );
  AND2_X1 U5228 ( .A1(n8261), .A2(n6104), .ZN(n4763) );
  OR2_X1 U5229 ( .A1(n8287), .A2(n7736), .ZN(n8027) );
  OR2_X1 U5230 ( .A1(n8508), .A2(n8321), .ZN(n8018) );
  INV_X1 U5231 ( .A(n4632), .ZN(n4631) );
  OAI21_X1 U5232 ( .B1(n6222), .B2(n4633), .A(n8002), .ZN(n4632) );
  INV_X1 U5233 ( .A(n7999), .ZN(n4633) );
  INV_X1 U5234 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U5235 ( .A1(n6259), .A2(n5031), .ZN(n5837) );
  INV_X1 U5236 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5809) );
  INV_X1 U5237 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5024) );
  INV_X1 U5238 ( .A(n5402), .ZN(n4971) );
  NOR2_X1 U5239 ( .A1(n4978), .A2(n4974), .ZN(n4973) );
  INV_X1 U5240 ( .A(n8657), .ZN(n4974) );
  INV_X1 U5241 ( .A(n5565), .ZN(n4978) );
  AND2_X1 U5242 ( .A1(n5574), .A2(n8616), .ZN(n5575) );
  OR2_X1 U5243 ( .A1(n5039), .A2(n5569), .ZN(n5574) );
  NAND2_X1 U5244 ( .A1(n5565), .A2(n4977), .ZN(n4976) );
  INV_X1 U5245 ( .A(n5499), .ZN(n4977) );
  AND2_X1 U5246 ( .A1(n5669), .A2(n5668), .ZN(n5671) );
  NAND2_X1 U5247 ( .A1(n8617), .A2(n5598), .ZN(n4962) );
  NAND2_X1 U5249 ( .A1(n8552), .A2(n5426), .ZN(n5448) );
  NAND2_X1 U5250 ( .A1(n4968), .A2(n5425), .ZN(n5426) );
  NAND2_X1 U5251 ( .A1(n7624), .A2(n5402), .ZN(n4968) );
  NOR2_X1 U5252 ( .A1(n9240), .A2(n4874), .ZN(n4873) );
  INV_X1 U5253 ( .A(n4876), .ZN(n4874) );
  NOR2_X1 U5254 ( .A1(n9489), .A2(n9488), .ZN(n9278) );
  AOI21_X1 U5255 ( .B1(n4814), .B2(n4816), .A(n4464), .ZN(n4813) );
  INV_X1 U5256 ( .A(n4431), .ZN(n4814) );
  INV_X1 U5257 ( .A(n4816), .ZN(n4815) );
  AND2_X1 U5258 ( .A1(n4562), .A2(n8859), .ZN(n4560) );
  AND2_X1 U5259 ( .A1(n4669), .A2(n4668), .ZN(n4667) );
  NOR2_X1 U5260 ( .A1(n7558), .A2(n7517), .ZN(n4669) );
  NAND2_X1 U5261 ( .A1(n7517), .A2(n8982), .ZN(n4818) );
  NAND2_X1 U5262 ( .A1(n7169), .A2(n4572), .ZN(n4575) );
  NOR2_X1 U5263 ( .A1(n8850), .A2(n4573), .ZN(n4572) );
  INV_X1 U5264 ( .A(n7168), .ZN(n4573) );
  NAND2_X1 U5265 ( .A1(n8925), .A2(n4571), .ZN(n8928) );
  NAND2_X1 U5266 ( .A1(n8847), .A2(n7186), .ZN(n4571) );
  INV_X1 U5267 ( .A(n6483), .ZN(n4906) );
  NOR2_X1 U5268 ( .A1(n6471), .A2(n7885), .ZN(n4658) );
  NAND2_X1 U5269 ( .A1(n7692), .A2(n7691), .ZN(n7884) );
  OR2_X1 U5270 ( .A1(n7690), .A2(n7689), .ZN(n7691) );
  AND2_X1 U5271 ( .A1(n6187), .A2(n6171), .ZN(n4610) );
  AOI21_X1 U5272 ( .B1(n4609), .B2(n4608), .A(n4497), .ZN(n4607) );
  INV_X1 U5273 ( .A(n6171), .ZN(n4608) );
  INV_X1 U5274 ( .A(n4611), .ZN(n4609) );
  AND2_X1 U5275 ( .A1(n5680), .A2(n5654), .ZN(n5678) );
  NAND2_X1 U5276 ( .A1(n4613), .A2(n4926), .ZN(n5501) );
  AOI21_X1 U5277 ( .B1(n4927), .B2(n4417), .A(n4494), .ZN(n4926) );
  NAND2_X1 U5278 ( .A1(n5432), .A2(n4925), .ZN(n4613) );
  AOI21_X1 U5279 ( .B1(n4930), .B2(n4587), .A(n4459), .ZN(n4586) );
  INV_X1 U5280 ( .A(n4935), .ZN(n4587) );
  INV_X1 U5281 ( .A(n5113), .ZN(n4553) );
  NAND2_X1 U5282 ( .A1(n5788), .A2(n5787), .ZN(n6117) );
  OR2_X1 U5283 ( .A1(n6907), .A2(n9885), .ZN(n6987) );
  AOI21_X1 U5284 ( .B1(n4998), .B2(n4996), .A(n4454), .ZN(n4995) );
  INV_X1 U5285 ( .A(n7844), .ZN(n4996) );
  XNOR2_X1 U5286 ( .A(n6271), .B(n6270), .ZN(n7505) );
  NAND2_X1 U5287 ( .A1(n6269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6271) );
  INV_X1 U5288 ( .A(n4921), .ZN(n4920) );
  INV_X1 U5289 ( .A(n8085), .ZN(n4922) );
  AOI21_X1 U5290 ( .B1(n7938), .B2(n7937), .A(n7936), .ZN(n8089) );
  AND3_X1 U5291 ( .A1(n6150), .A2(n6149), .A3(n6148), .ZN(n7764) );
  OR2_X1 U5292 ( .A1(n9701), .A2(n6393), .ZN(n6395) );
  NAND2_X1 U5293 ( .A1(n6606), .A2(n6605), .ZN(n6604) );
  NAND2_X1 U5294 ( .A1(n6604), .A2(n4836), .ZN(n4835) );
  NOR2_X1 U5295 ( .A1(n4837), .A2(n9724), .ZN(n4836) );
  INV_X1 U5296 ( .A(n6396), .ZN(n4837) );
  AND2_X1 U5297 ( .A1(n4849), .A2(n4850), .ZN(n4848) );
  NOR2_X1 U5298 ( .A1(n4854), .A2(n5908), .ZN(n4850) );
  NAND2_X1 U5299 ( .A1(n4732), .A2(n4731), .ZN(n9760) );
  NAND2_X1 U5300 ( .A1(n4734), .A2(n4733), .ZN(n4731) );
  NAND2_X1 U5301 ( .A1(n4538), .A2(n6315), .ZN(n6888) );
  INV_X1 U5302 ( .A(n9757), .ZN(n4538) );
  AND2_X1 U5303 ( .A1(n6399), .A2(n4864), .ZN(n4861) );
  NAND2_X1 U5304 ( .A1(n4725), .A2(n4724), .ZN(n4723) );
  INV_X1 U5305 ( .A(n9778), .ZN(n4724) );
  INV_X1 U5306 ( .A(n6371), .ZN(n4725) );
  NAND2_X1 U5307 ( .A1(n4502), .A2(n4419), .ZN(n4722) );
  NAND2_X1 U5308 ( .A1(n4502), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6885) );
  OR2_X1 U5309 ( .A1(n7488), .A2(n6407), .ZN(n6409) );
  AOI21_X1 U5310 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6507), .A(n7525), .ZN(
        n6411) );
  OAI21_X1 U5311 ( .B1(n9820), .B2(n4894), .A(n4893), .ZN(n8123) );
  NAND2_X1 U5312 ( .A1(n4897), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U5313 ( .A1(n6412), .A2(n4897), .ZN(n4893) );
  INV_X1 U5314 ( .A(n8124), .ZN(n4897) );
  OR2_X1 U5315 ( .A1(n8141), .A2(n8140), .ZN(n4869) );
  INV_X1 U5316 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6066) );
  AND2_X1 U5317 ( .A1(n8165), .A2(n4644), .ZN(n4643) );
  AND4_X1 U5318 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n8252)
         );
  NOR2_X1 U5319 ( .A1(n8285), .A2(n4653), .ZN(n4652) );
  INV_X1 U5320 ( .A(n8025), .ZN(n4653) );
  INV_X1 U5321 ( .A(n6004), .ZN(n5781) );
  NOR2_X1 U5322 ( .A1(n8353), .A2(n4765), .ZN(n4764) );
  INV_X1 U5323 ( .A(n6011), .ZN(n4765) );
  NAND2_X1 U5324 ( .A1(n4617), .A2(n7989), .ZN(n7376) );
  OAI21_X1 U5325 ( .B1(n9911), .B2(n4615), .A(n4614), .ZN(n4617) );
  AND2_X1 U5326 ( .A1(n4616), .A2(n7986), .ZN(n4614) );
  NAND2_X1 U5327 ( .A1(n7920), .A2(n4422), .ZN(n4616) );
  INV_X1 U5328 ( .A(n4615), .ZN(n4618) );
  AND2_X1 U5329 ( .A1(n7985), .A2(n7980), .ZN(n7920) );
  AND2_X1 U5330 ( .A1(n5958), .A2(n5945), .ZN(n4767) );
  AND3_X1 U5331 ( .A1(n5944), .A2(n5943), .A3(n5942), .ZN(n7275) );
  NOR2_X1 U5332 ( .A1(n7963), .A2(n4647), .ZN(n4646) );
  INV_X1 U5333 ( .A(n7964), .ZN(n4647) );
  INV_X1 U5334 ( .A(n4747), .ZN(n4746) );
  INV_X1 U5335 ( .A(n4748), .ZN(n4744) );
  INV_X1 U5336 ( .A(n6929), .ZN(n4751) );
  AND2_X1 U5337 ( .A1(n6267), .A2(n8078), .ZN(n6922) );
  NAND2_X1 U5338 ( .A1(n7619), .A2(n7890), .ZN(n4909) );
  INV_X1 U5339 ( .A(n8067), .ZN(n4644) );
  INV_X1 U5340 ( .A(n8181), .ZN(n6234) );
  NAND2_X1 U5341 ( .A1(n6126), .A2(n6125), .ZN(n7822) );
  OR2_X1 U5342 ( .A1(n8487), .A2(n8252), .ZN(n8035) );
  NAND2_X1 U5343 ( .A1(n6225), .A2(n8031), .ZN(n8259) );
  INV_X1 U5344 ( .A(n8270), .ZN(n6102) );
  AOI21_X1 U5345 ( .B1(n8295), .B2(n4652), .A(n4649), .ZN(n8269) );
  INV_X1 U5346 ( .A(n4650), .ZN(n4649) );
  AOI21_X1 U5347 ( .B1(n4652), .B2(n7905), .A(n4651), .ZN(n4650) );
  INV_X1 U5348 ( .A(n8027), .ZN(n4651) );
  OAI21_X1 U5349 ( .B1(n8327), .B2(n8006), .A(n7927), .ZN(n8317) );
  NAND2_X1 U5350 ( .A1(n6719), .A2(n8083), .ZN(n8351) );
  OR2_X1 U5351 ( .A1(n8533), .A2(n8350), .ZN(n7999) );
  INV_X1 U5352 ( .A(n5864), .ZN(n7889) );
  INV_X1 U5353 ( .A(n5896), .ZN(n6092) );
  NAND2_X1 U5354 ( .A1(n8361), .A2(n6222), .ZN(n8365) );
  OR2_X1 U5355 ( .A1(n6728), .A2(n8078), .ZN(n6720) );
  AND2_X1 U5356 ( .A1(n6711), .A2(n6709), .ZN(n6743) );
  AOI21_X1 U5357 ( .B1(n4436), .B2(n6205), .A(n6200), .ZN(n6201) );
  INV_X1 U5358 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5800) );
  AND2_X1 U5359 ( .A1(n6038), .A2(n6026), .ZN(n8119) );
  INV_X1 U5360 ( .A(n5639), .ZN(n8588) );
  AND2_X1 U5361 ( .A1(n8665), .A2(n5645), .ZN(n8564) );
  OR2_X1 U5362 ( .A1(n7604), .A2(n7602), .ZN(n8599) );
  INV_X1 U5363 ( .A(n6788), .ZN(n4950) );
  XNOR2_X1 U5364 ( .A(n5227), .B(n5226), .ZN(n6826) );
  NAND2_X1 U5365 ( .A1(n4981), .A2(n4979), .ZN(n7397) );
  AND2_X1 U5366 ( .A1(n4980), .A2(n5036), .ZN(n4979) );
  NAND2_X1 U5367 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  INV_X1 U5368 ( .A(n5677), .ZN(n4957) );
  AND2_X1 U5369 ( .A1(n4878), .A2(n4428), .ZN(n9121) );
  AND4_X1 U5370 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n8809)
         );
  AND4_X1 U5371 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n7162)
         );
  NOR3_X1 U5372 ( .A1(n9192), .A2(n4664), .A3(n9322), .ZN(n9132) );
  NAND2_X1 U5373 ( .A1(n4469), .A2(n9127), .ZN(n4845) );
  NAND2_X1 U5374 ( .A1(n9166), .A2(n9126), .ZN(n4847) );
  NAND2_X1 U5375 ( .A1(n9127), .A2(n9126), .ZN(n4846) );
  NAND2_X1 U5376 ( .A1(n9173), .A2(n9174), .ZN(n9172) );
  OR2_X1 U5377 ( .A1(n9353), .A2(n9191), .ZN(n9182) );
  AND2_X1 U5378 ( .A1(n8836), .A2(n9125), .ZN(n9188) );
  AND2_X1 U5379 ( .A1(n9182), .A2(n8885), .ZN(n9199) );
  AOI21_X1 U5380 ( .B1(n4825), .B2(n9110), .A(n4449), .ZN(n4824) );
  OR2_X1 U5381 ( .A1(n9364), .A2(n9242), .ZN(n9109) );
  AND2_X1 U5382 ( .A1(n8837), .A2(n8875), .ZN(n9217) );
  AND2_X1 U5383 ( .A1(n8790), .A2(n9123), .ZN(n9225) );
  OR2_X1 U5384 ( .A1(n9120), .A2(n8896), .ZN(n4877) );
  OR2_X1 U5385 ( .A1(n4428), .A2(n9120), .ZN(n4876) );
  NAND2_X1 U5386 ( .A1(n9106), .A2(n5030), .ZN(n9255) );
  OR2_X1 U5387 ( .A1(n9283), .A2(n9105), .ZN(n5030) );
  OR2_X1 U5388 ( .A1(n9384), .A2(n9484), .ZN(n9104) );
  AND2_X1 U5389 ( .A1(n4549), .A2(n4548), .ZN(n9272) );
  AND2_X1 U5390 ( .A1(n9101), .A2(n9298), .ZN(n4799) );
  NAND2_X1 U5391 ( .A1(n7463), .A2(n4667), .ZN(n9288) );
  INV_X1 U5392 ( .A(n4563), .ZN(n4562) );
  OAI21_X1 U5393 ( .B1(n8857), .B2(n8937), .A(n8761), .ZN(n4563) );
  NAND2_X1 U5394 ( .A1(n7463), .A2(n4669), .ZN(n7552) );
  AOI21_X1 U5395 ( .B1(n4882), .B2(n4885), .A(n7455), .ZN(n4881) );
  INV_X1 U5396 ( .A(n4882), .ZN(n4879) );
  NAND2_X1 U5397 ( .A1(n5385), .A2(n5384), .ZN(n7621) );
  NOR2_X1 U5398 ( .A1(n7352), .A2(n7621), .ZN(n7463) );
  NAND2_X1 U5399 ( .A1(n4887), .A2(n4884), .ZN(n7347) );
  OR2_X1 U5400 ( .A1(n7338), .A2(n8852), .ZN(n4887) );
  AOI21_X1 U5401 ( .B1(n4793), .B2(n7251), .A(n4452), .ZN(n4792) );
  OAI21_X1 U5402 ( .B1(n9534), .B2(n9532), .A(n7181), .ZN(n7248) );
  NAND2_X1 U5403 ( .A1(n7079), .A2(n7060), .ZN(n7061) );
  NAND2_X1 U5404 ( .A1(n7059), .A2(n7058), .ZN(n4695) );
  AND2_X1 U5405 ( .A1(n5160), .A2(n8904), .ZN(n9535) );
  OR2_X1 U5406 ( .A1(n7002), .A2(n6957), .ZN(n9487) );
  INV_X1 U5407 ( .A(n9098), .ZN(n9316) );
  AND2_X1 U5408 ( .A1(n9322), .A2(n9625), .ZN(n4567) );
  AND2_X1 U5409 ( .A1(n5294), .A2(n4475), .ZN(n4576) );
  OR2_X1 U5410 ( .A1(n6480), .A2(n5311), .ZN(n4577) );
  INV_X1 U5411 ( .A(n9626), .ZN(n9656) );
  NAND2_X1 U5412 ( .A1(n5382), .A2(n4518), .ZN(n5057) );
  AND2_X1 U5413 ( .A1(n5054), .A2(n4478), .ZN(n4518) );
  XNOR2_X1 U5414 ( .A(n7884), .B(n7883), .ZN(n8821) );
  NAND2_X1 U5415 ( .A1(n5086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5088) );
  AND2_X1 U5416 ( .A1(n5650), .A2(n5623), .ZN(n5648) );
  INV_X1 U5417 ( .A(n5617), .ZN(n4944) );
  OR2_X1 U5418 ( .A1(n5527), .A2(n5526), .ZN(n5512) );
  OAI21_X1 U5419 ( .B1(n5432), .B2(n4929), .A(n4927), .ZN(n5476) );
  NAND2_X1 U5420 ( .A1(n5432), .A2(n5431), .ZN(n5453) );
  NAND2_X1 U5421 ( .A1(n4932), .A2(n4933), .ZN(n5380) );
  NAND2_X1 U5422 ( .A1(n5333), .A2(n4935), .ZN(n4932) );
  AND2_X1 U5423 ( .A1(n5121), .A2(n5120), .ZN(n5292) );
  NAND2_X1 U5424 ( .A1(n5237), .A2(n5236), .ZN(n5111) );
  INV_X1 U5425 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4948) );
  AND4_X1 U5426 ( .A1(n6132), .A2(n6131), .A3(n6130), .A4(n6129), .ZN(n8251)
         );
  OR2_X1 U5427 ( .A1(n7649), .A2(n7926), .ZN(n5002) );
  AND4_X1 U5428 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(n7273)
         );
  OR2_X1 U5429 ( .A1(n7832), .A2(n5022), .ZN(n5021) );
  INV_X1 U5430 ( .A(n7645), .ZN(n5020) );
  INV_X1 U5431 ( .A(n8215), .ZN(n8236) );
  INV_X1 U5432 ( .A(n8105), .ZN(n8350) );
  OAI21_X2 U5433 ( .B1(n7653), .B2(n8102), .A(n7784), .ZN(n7843) );
  NAND2_X1 U5434 ( .A1(n8355), .A2(n6716), .ZN(n7850) );
  INV_X1 U5435 ( .A(n8104), .ZN(n8348) );
  AOI21_X1 U5436 ( .B1(n7708), .B2(n7709), .A(n4510), .ZN(n7869) );
  AND2_X1 U5437 ( .A1(n7648), .A2(n8348), .ZN(n4510) );
  NAND2_X1 U5438 ( .A1(n4755), .A2(n4759), .ZN(n6731) );
  NAND2_X1 U5439 ( .A1(n5815), .A2(n4758), .ZN(n4759) );
  AOI22_X1 U5440 ( .A1(n4756), .A2(n4754), .B1(n5815), .B2(n4416), .ZN(n4755)
         );
  AND2_X1 U5441 ( .A1(n7685), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4758) );
  NAND2_X1 U5442 ( .A1(n4866), .A2(n6401), .ZN(n6884) );
  AND2_X1 U5443 ( .A1(n6401), .A2(n4867), .ZN(n9772) );
  OR2_X1 U5444 ( .A1(n9788), .A2(n6302), .ZN(n4891) );
  XNOR2_X1 U5445 ( .A(n6404), .B(n6403), .ZN(n9788) );
  OR2_X1 U5446 ( .A1(n9820), .A2(n9821), .ZN(n4896) );
  INV_X1 U5447 ( .A(P2_U3893), .ZN(n8113) );
  AND3_X1 U5448 ( .A1(n4901), .A2(n4900), .A3(n4898), .ZN(n4532) );
  AND2_X1 U5449 ( .A1(n5027), .A2(n5026), .ZN(n4900) );
  OAI21_X1 U5450 ( .B1(n9457), .B2(n4420), .A(n4902), .ZN(n4901) );
  NAND2_X1 U5451 ( .A1(n4899), .A2(n9863), .ZN(n4898) );
  NAND2_X1 U5452 ( .A1(n6357), .A2(n9460), .ZN(n4533) );
  OR2_X1 U5453 ( .A1(n8373), .A2(n8168), .ZN(n4779) );
  OR2_X1 U5454 ( .A1(n6919), .A2(n9933), .ZN(n8336) );
  OAI21_X2 U5455 ( .B1(n6927), .B2(n7262), .A(n8373), .ZN(n8378) );
  OR2_X1 U5456 ( .A1(n6715), .A2(n6714), .ZN(n8355) );
  AND2_X1 U5457 ( .A1(n8155), .A2(n6821), .ZN(n6251) );
  AOI21_X1 U5458 ( .B1(n4776), .B2(n6212), .A(n4775), .ZN(n8442) );
  INV_X1 U5459 ( .A(n4780), .ZN(n4775) );
  AOI21_X1 U5460 ( .B1(n8167), .B2(n8370), .A(n4781), .ZN(n4780) );
  NAND2_X1 U5461 ( .A1(n6152), .A2(n6151), .ZN(n8462) );
  AND3_X1 U5462 ( .A1(n5917), .A2(n4424), .A3(n4656), .ZN(n4655) );
  INV_X1 U5463 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4656) );
  OR2_X1 U5464 ( .A1(n5921), .A2(n5920), .ZN(n9756) );
  NOR2_X1 U5465 ( .A1(n7574), .A2(n7568), .ZN(n5076) );
  INV_X1 U5466 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U5467 ( .A1(n7582), .A2(n7581), .ZN(n9335) );
  AND4_X1 U5468 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n7546)
         );
  AND4_X1 U5469 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n8633)
         );
  AND2_X1 U5470 ( .A1(n5610), .A2(n5609), .ZN(n9235) );
  AND2_X1 U5471 ( .A1(n7604), .A2(n5712), .ZN(n9169) );
  AND4_X1 U5472 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n8738)
         );
  AOI21_X1 U5473 ( .B1(n8834), .B2(n9306), .A(n8833), .ZN(n8968) );
  NAND2_X1 U5474 ( .A1(n4598), .A2(n4539), .ZN(n8832) );
  CLKBUF_X1 U5475 ( .A(n5736), .Z(n5737) );
  INV_X1 U5476 ( .A(n4803), .ZN(n4802) );
  NAND2_X1 U5477 ( .A1(n4568), .A2(n9131), .ZN(n9320) );
  NAND2_X1 U5478 ( .A1(n4569), .A2(n9486), .ZN(n4568) );
  XNOR2_X1 U5479 ( .A(n4570), .B(n9118), .ZN(n4569) );
  AND4_X1 U5480 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n9356)
         );
  AND4_X1 U5481 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n9232)
         );
  AND4_X1 U5482 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n7254)
         );
  MUX2_X1 U5483 ( .A(n7970), .B(n7969), .S(n8078), .Z(n7977) );
  OAI21_X1 U5484 ( .B1(n8769), .B2(n8764), .A(n4423), .ZN(n4683) );
  INV_X1 U5485 ( .A(n4688), .ZN(n4687) );
  INV_X1 U5486 ( .A(n4680), .ZN(n4679) );
  OAI21_X1 U5487 ( .B1(n4686), .B2(n4683), .A(n8770), .ZN(n4680) );
  AOI21_X1 U5488 ( .B1(n4688), .B2(n8826), .A(n7185), .ZN(n4686) );
  NAND2_X1 U5489 ( .A1(n4520), .A2(n8078), .ZN(n4519) );
  NAND2_X1 U5490 ( .A1(n8023), .A2(n8083), .ZN(n4522) );
  NAND2_X1 U5491 ( .A1(n4701), .A2(n8895), .ZN(n8783) );
  NOR2_X1 U5492 ( .A1(n4445), .A2(n4421), .ZN(n4700) );
  NAND2_X1 U5493 ( .A1(n4872), .A2(n8831), .ZN(n4674) );
  NAND2_X1 U5494 ( .A1(n4677), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U5495 ( .A1(n8914), .A2(n8831), .ZN(n4676) );
  INV_X1 U5496 ( .A(n8802), .ZN(n4707) );
  NOR2_X1 U5497 ( .A1(n8889), .A2(n8805), .ZN(n4708) );
  AOI21_X1 U5498 ( .B1(n4943), .B2(n4942), .A(n4941), .ZN(n4940) );
  INV_X1 U5499 ( .A(n5648), .ZN(n4941) );
  INV_X1 U5500 ( .A(n4945), .ZN(n4942) );
  INV_X1 U5501 ( .A(n7904), .ZN(n4743) );
  INV_X1 U5502 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5801) );
  NOR2_X1 U5503 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5803) );
  NOR2_X1 U5504 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5804) );
  INV_X1 U5505 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6051) );
  OR2_X1 U5506 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  OR2_X1 U5507 ( .A1(n8753), .A2(n7182), .ZN(n8850) );
  NOR2_X1 U5508 ( .A1(n7185), .A2(n8752), .ZN(n8847) );
  NOR2_X1 U5509 ( .A1(n7165), .A2(n4663), .ZN(n4661) );
  NAND2_X1 U5510 ( .A1(n4914), .A2(n4913), .ZN(n7690) );
  AOI21_X1 U5511 ( .B1(n4915), .B2(n4917), .A(n4500), .ZN(n4913) );
  NAND2_X1 U5512 ( .A1(n5577), .A2(n5578), .ZN(n4597) );
  INV_X1 U5513 ( .A(n5474), .ZN(n5475) );
  AND2_X1 U5514 ( .A1(n4927), .A2(n4435), .ZN(n4925) );
  INV_X1 U5515 ( .A(SI_17_), .ZN(n5477) );
  INV_X1 U5516 ( .A(n5011), .ZN(n5009) );
  AOI21_X1 U5517 ( .B1(n5018), .B2(n7120), .A(n4453), .ZN(n5016) );
  INV_X1 U5518 ( .A(n5018), .ZN(n5017) );
  NOR2_X1 U5519 ( .A1(n6488), .A2(n6286), .ZN(n6702) );
  OR2_X1 U5520 ( .A1(n8080), .A2(n8444), .ZN(n8074) );
  OR2_X1 U5521 ( .A1(n8081), .A2(n8083), .ZN(n4924) );
  OR2_X1 U5522 ( .A1(n4638), .A2(n4642), .ZN(n4635) );
  AND2_X1 U5523 ( .A1(n4643), .A2(n7891), .ZN(n4642) );
  INV_X1 U5524 ( .A(n9761), .ZN(n4733) );
  INV_X1 U5525 ( .A(n6114), .ZN(n4762) );
  OAI21_X1 U5526 ( .B1(n4763), .B2(n4762), .A(n8249), .ZN(n4761) );
  NOR2_X1 U5527 ( .A1(n4627), .A2(n4623), .ZN(n4622) );
  INV_X1 U5528 ( .A(n8031), .ZN(n4623) );
  INV_X1 U5529 ( .A(n8036), .ZN(n4627) );
  INV_X1 U5530 ( .A(n8040), .ZN(n4625) );
  NAND2_X1 U5531 ( .A1(n7920), .A2(n7978), .ZN(n4615) );
  NAND2_X1 U5532 ( .A1(n6731), .A2(n7141), .ZN(n7912) );
  AND2_X1 U5533 ( .A1(n4743), .A2(n8210), .ZN(n4742) );
  OR2_X1 U5534 ( .A1(n8456), .A2(n7856), .ZN(n8061) );
  OR2_X1 U5535 ( .A1(n8048), .A2(n8207), .ZN(n6229) );
  OR2_X1 U5536 ( .A1(n7822), .A2(n8251), .ZN(n8045) );
  AND2_X1 U5537 ( .A1(n8095), .A2(n6351), .ZN(n6717) );
  INV_X1 U5538 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6260) );
  INV_X1 U5539 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6050) );
  INV_X1 U5540 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5995) );
  INV_X1 U5541 ( .A(n5598), .ZN(n4958) );
  NAND2_X1 U5542 ( .A1(n4982), .A2(n4986), .ZN(n7394) );
  NAND2_X1 U5543 ( .A1(n4515), .A2(n4987), .ZN(n4982) );
  INV_X1 U5544 ( .A(n4984), .ZN(n4983) );
  OAI21_X1 U5545 ( .B1(n4987), .B2(n4985), .A(n5301), .ZN(n4984) );
  NAND2_X1 U5546 ( .A1(n4983), .A2(n4985), .ZN(n4980) );
  AND2_X1 U5547 ( .A1(n5570), .A2(n5571), .ZN(n5039) );
  NAND2_X1 U5548 ( .A1(n8655), .A2(n5499), .ZN(n8571) );
  NAND2_X1 U5549 ( .A1(n4704), .A2(n9118), .ZN(n8812) );
  NAND2_X1 U5550 ( .A1(n4580), .A2(n4705), .ZN(n4704) );
  OR2_X1 U5551 ( .A1(n9328), .A2(n4665), .ZN(n4664) );
  OR2_X1 U5552 ( .A1(n9335), .A2(n9339), .ZN(n4665) );
  NOR2_X1 U5553 ( .A1(n9364), .A2(n9371), .ZN(n4672) );
  AOI21_X1 U5554 ( .B1(n4884), .B2(n8852), .A(n4883), .ZN(n4882) );
  INV_X1 U5555 ( .A(n8936), .ZN(n4883) );
  NOR2_X1 U5556 ( .A1(n4794), .A2(n4791), .ZN(n4790) );
  INV_X1 U5557 ( .A(n7191), .ZN(n4791) );
  INV_X1 U5558 ( .A(n7251), .ZN(n4794) );
  INV_X1 U5559 ( .A(n7193), .ZN(n4793) );
  INV_X1 U5560 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5282) );
  OR2_X1 U5561 ( .A1(n5283), .A2(n5282), .ZN(n5285) );
  NAND2_X1 U5562 ( .A1(n7169), .A2(n7168), .ZN(n8931) );
  INV_X1 U5563 ( .A(n4610), .ZN(n4605) );
  OR2_X1 U5564 ( .A1(n6172), .A2(n4606), .ZN(n4602) );
  NAND2_X1 U5565 ( .A1(n4607), .A2(n4611), .ZN(n4606) );
  AND2_X1 U5566 ( .A1(n9256), .A2(n4670), .ZN(n9204) );
  AND2_X1 U5567 ( .A1(n4412), .A2(n9208), .ZN(n4670) );
  NAND2_X1 U5568 ( .A1(n9256), .A2(n9250), .ZN(n9249) );
  NAND3_X1 U5569 ( .A1(n7099), .A2(n9619), .A3(n4661), .ZN(n7255) );
  NAND2_X1 U5570 ( .A1(n7099), .A2(n4661), .ZN(n9547) );
  XNOR2_X1 U5571 ( .A(n7690), .B(n7689), .ZN(n7688) );
  AND2_X1 U5572 ( .A1(n5830), .A2(n5829), .ZN(n6171) );
  NAND2_X1 U5573 ( .A1(n4509), .A2(n4508), .ZN(n5086) );
  INV_X1 U5574 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4508) );
  INV_X1 U5575 ( .A(n5069), .ZN(n4509) );
  NAND2_X1 U5576 ( .A1(n4579), .A2(n5704), .ZN(n5823) );
  NAND2_X1 U5577 ( .A1(n5703), .A2(n5702), .ZN(n4579) );
  AND2_X1 U5578 ( .A1(n5824), .A2(n5708), .ZN(n5822) );
  INV_X1 U5579 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5052) );
  INV_X1 U5580 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5081) );
  INV_X1 U5581 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5543) );
  INV_X1 U5582 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5045) );
  NOR2_X1 U5583 ( .A1(n5451), .A2(n5452), .ZN(n4929) );
  INV_X1 U5584 ( .A(SI_14_), .ZN(n5408) );
  INV_X1 U5585 ( .A(n5331), .ZN(n4936) );
  INV_X1 U5586 ( .A(n4552), .ZN(n4551) );
  NOR2_X1 U5587 ( .A1(n4429), .A2(n4911), .ZN(n4910) );
  INV_X1 U5588 ( .A(n5100), .ZN(n4911) );
  INV_X1 U5589 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5092) );
  INV_X1 U5590 ( .A(SI_12_), .ZN(n10241) );
  NAND2_X1 U5591 ( .A1(n7843), .A2(n7844), .ZN(n4999) );
  AOI21_X1 U5592 ( .B1(n4992), .B2(n4997), .A(n4485), .ZN(n4990) );
  NOR2_X1 U5593 ( .A1(n4993), .A2(n7804), .ZN(n4992) );
  NOR2_X1 U5594 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  NAND2_X1 U5595 ( .A1(n5792), .A2(n5791), .ZN(n6153) );
  INV_X1 U5596 ( .A(n4998), .ZN(n4997) );
  NAND2_X1 U5597 ( .A1(n5790), .A2(n5789), .ZN(n6127) );
  XNOR2_X1 U5598 ( .A(n7118), .B(n7263), .ZN(n6846) );
  OR2_X1 U5599 ( .A1(n9707), .A2(n9706), .ZN(n9709) );
  OAI21_X1 U5600 ( .B1(n9703), .B2(n6392), .A(n6394), .ZN(n9701) );
  NAND2_X1 U5601 ( .A1(n4507), .A2(n4713), .ZN(n9720) );
  NAND2_X1 U5602 ( .A1(n4831), .A2(n4835), .ZN(n9730) );
  AOI21_X1 U5603 ( .B1(n4833), .B2(n9724), .A(n4832), .ZN(n4831) );
  OAI21_X1 U5604 ( .B1(n4838), .B2(n6396), .A(P2_REG1_REG_3__SCAN_IN), .ZN(
        n4832) );
  NOR2_X1 U5605 ( .A1(n4860), .A2(n6462), .ZN(n4852) );
  AND2_X1 U5606 ( .A1(n9738), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U5607 ( .A1(n4864), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4863) );
  INV_X1 U5608 ( .A(n6317), .ZN(n9775) );
  NOR2_X1 U5609 ( .A1(n9775), .A2(n9774), .ZN(n9773) );
  NOR2_X1 U5610 ( .A1(n6320), .A2(n9773), .ZN(n9794) );
  AND2_X1 U5611 ( .A1(n4723), .A2(n4426), .ZN(n4721) );
  OAI21_X1 U5612 ( .B1(n6379), .B2(n9806), .A(n6378), .ZN(n9808) );
  NOR2_X1 U5613 ( .A1(n6410), .A2(n9803), .ZN(n7527) );
  NOR2_X1 U5614 ( .A1(n7527), .A2(n7526), .ZN(n7525) );
  AOI21_X1 U5615 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6507), .A(n7521), .ZN(
        n6381) );
  AOI21_X1 U5616 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6662), .A(n8123), .ZN(
        n6414) );
  AOI21_X1 U5617 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6662), .A(n8114), .ZN(
        n6384) );
  XNOR2_X1 U5618 ( .A(n6384), .B(n6413), .ZN(n9843) );
  NOR2_X1 U5619 ( .A1(n10128), .A2(n9860), .ZN(n9859) );
  NAND2_X1 U5620 ( .A1(n4714), .A2(n4715), .ZN(n9472) );
  INV_X1 U5621 ( .A(n6390), .ZN(n4715) );
  OR2_X1 U5622 ( .A1(n6177), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8150) );
  OR2_X1 U5623 ( .A1(n6127), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U5624 ( .A1(n5786), .A2(n5785), .ZN(n6095) );
  INV_X1 U5625 ( .A(n6080), .ZN(n5786) );
  OR2_X1 U5626 ( .A1(n6095), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6107) );
  AND4_X1 U5627 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n8284)
         );
  NAND2_X1 U5628 ( .A1(n5784), .A2(n10237), .ZN(n6058) );
  INV_X1 U5629 ( .A(n6042), .ZN(n5784) );
  OR2_X1 U5630 ( .A1(n6058), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U5631 ( .A1(n5783), .A2(n5782), .ZN(n6029) );
  NAND2_X1 U5632 ( .A1(n5780), .A2(n5779), .ZN(n5972) );
  INV_X1 U5633 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5777) );
  OR2_X1 U5634 ( .A1(n7129), .A2(n7137), .ZN(n5931) );
  OR2_X1 U5635 ( .A1(n5924), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U5636 ( .A1(n4620), .A2(n7942), .ZN(n9888) );
  NAND2_X1 U5637 ( .A1(n6897), .A2(n6896), .ZN(n4620) );
  NAND2_X1 U5638 ( .A1(n6840), .A2(n5879), .ZN(n9879) );
  AND2_X1 U5639 ( .A1(n7286), .A2(n6238), .ZN(n6927) );
  OR2_X2 U5640 ( .A1(n6731), .A2(n7141), .ZN(n7945) );
  AND2_X1 U5641 ( .A1(n6726), .A2(n6494), .ZN(n6699) );
  INV_X1 U5642 ( .A(n6494), .ZN(n6920) );
  AND2_X1 U5643 ( .A1(n6919), .A2(n8092), .ZN(n6821) );
  AND2_X1 U5644 ( .A1(n8185), .A2(n9883), .ZN(n4781) );
  AOI21_X1 U5645 ( .B1(n4738), .B2(n4740), .A(n4461), .ZN(n4735) );
  OR2_X1 U5646 ( .A1(n8067), .A2(n8066), .ZN(n8173) );
  NAND2_X1 U5647 ( .A1(n4737), .A2(n4741), .ZN(n8184) );
  NAND2_X1 U5648 ( .A1(n8212), .A2(n4742), .ZN(n4737) );
  AND2_X1 U5649 ( .A1(n7902), .A2(n8061), .ZN(n8183) );
  INV_X1 U5650 ( .A(n8183), .ZN(n8180) );
  OR2_X1 U5651 ( .A1(n7904), .A2(n4440), .ZN(n8196) );
  OR2_X1 U5652 ( .A1(n8474), .A2(n8236), .ZN(n8207) );
  NAND2_X1 U5653 ( .A1(n8233), .A2(n8238), .ZN(n4770) );
  AND2_X1 U5654 ( .A1(n8207), .A2(n8208), .ZN(n8225) );
  AND2_X1 U5655 ( .A1(n8028), .A2(n8031), .ZN(n8270) );
  AND4_X1 U5656 ( .A1(n6063), .A2(n6062), .A3(n6061), .A4(n6060), .ZN(n8321)
         );
  OR2_X1 U5657 ( .A1(n8006), .A2(n8007), .ZN(n8329) );
  AOI21_X1 U5658 ( .B1(n4631), .B2(n4633), .A(n4630), .ZN(n4629) );
  INV_X1 U5659 ( .A(n8003), .ZN(n4630) );
  INV_X1 U5660 ( .A(n8351), .ZN(n9883) );
  AND2_X1 U5661 ( .A1(n6428), .A2(n6699), .ZN(n6739) );
  OR2_X1 U5662 ( .A1(n6425), .A2(n6724), .ZN(n6741) );
  NAND2_X1 U5663 ( .A1(n7389), .A2(n9925), .ZN(n9938) );
  OR2_X1 U5664 ( .A1(n6487), .A2(n6297), .ZN(n6714) );
  INV_X1 U5665 ( .A(n5836), .ZN(n4535) );
  OR2_X1 U5666 ( .A1(n6259), .A2(n4477), .ZN(n4536) );
  NAND2_X1 U5667 ( .A1(n6203), .A2(n6202), .ZN(n6269) );
  NOR2_X1 U5668 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4774) );
  INV_X1 U5669 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4773) );
  INV_X1 U5670 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5846) );
  OAI21_X1 U5671 ( .B1(n5128), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U5672 ( .A1(n4971), .A2(n5425), .ZN(n4969) );
  NAND2_X1 U5673 ( .A1(n4963), .A2(n5425), .ZN(n4967) );
  NOR2_X1 U5674 ( .A1(n5425), .A2(n4971), .ZN(n4970) );
  AND2_X1 U5675 ( .A1(n5575), .A2(n4976), .ZN(n4975) );
  AND2_X1 U5676 ( .A1(n5396), .A2(n5378), .ZN(n8626) );
  INV_X1 U5677 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U5678 ( .A1(n8656), .A2(n8657), .ZN(n8655) );
  INV_X1 U5679 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10081) );
  OR2_X1 U5680 ( .A1(n5463), .A2(n5462), .ZN(n5487) );
  AND2_X1 U5681 ( .A1(n5677), .A2(n5674), .ZN(n8666) );
  NAND2_X1 U5682 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n5586), .ZN(n5629) );
  INV_X1 U5683 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5248) );
  XNOR2_X1 U5684 ( .A(n5741), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5736) );
  AND2_X1 U5685 ( .A1(n6873), .A2(n6872), .ZN(n6970) );
  NOR2_X1 U5686 ( .A1(n4807), .A2(n9174), .ZN(n4804) );
  OAI21_X1 U5687 ( .B1(n4807), .B2(n4809), .A(n4805), .ZN(n4803) );
  AOI21_X1 U5688 ( .B1(n4806), .B2(n9159), .A(n4460), .ZN(n4805) );
  NAND2_X1 U5689 ( .A1(n4839), .A2(n4840), .ZN(n4570) );
  AOI21_X1 U5690 ( .B1(n4842), .B2(n4846), .A(n4841), .ZN(n4840) );
  INV_X1 U5691 ( .A(n9128), .ZN(n4841) );
  NOR2_X1 U5692 ( .A1(n9167), .A2(n9335), .ZN(n9155) );
  OR2_X1 U5693 ( .A1(n9192), .A2(n9339), .ZN(n9167) );
  NAND2_X1 U5694 ( .A1(n4824), .A2(n4482), .ZN(n4823) );
  AND2_X1 U5695 ( .A1(n4822), .A2(n4830), .ZN(n4821) );
  NAND2_X1 U5696 ( .A1(n9256), .A2(n4672), .ZN(n9233) );
  NAND2_X1 U5697 ( .A1(n4545), .A2(n9225), .ZN(n9223) );
  AOI21_X1 U5698 ( .B1(n4873), .B2(n4877), .A(n4872), .ZN(n4871) );
  OR2_X1 U5699 ( .A1(n9272), .A2(n8896), .ZN(n4878) );
  AND2_X1 U5700 ( .A1(n9278), .A2(n9283), .ZN(n9279) );
  AND2_X1 U5701 ( .A1(n9279), .A2(n9260), .ZN(n9256) );
  NOR2_X1 U5702 ( .A1(n5552), .A2(n5531), .ZN(n5530) );
  NOR2_X1 U5703 ( .A1(n5487), .A2(n10081), .ZN(n5551) );
  NAND2_X1 U5704 ( .A1(n5550), .A2(n5549), .ZN(n9488) );
  OAI21_X1 U5705 ( .B1(n9287), .B2(n9103), .A(n4458), .ZN(n9479) );
  AND2_X1 U5706 ( .A1(n8839), .A2(n9269), .ZN(n9482) );
  OAI21_X1 U5707 ( .B1(n4559), .B2(n8892), .A(n4555), .ZN(n9297) );
  INV_X1 U5708 ( .A(n4556), .ZN(n4555) );
  NAND2_X1 U5709 ( .A1(n7463), .A2(n4666), .ZN(n9489) );
  AND2_X1 U5710 ( .A1(n4667), .A2(n9509), .ZN(n4666) );
  NAND2_X1 U5711 ( .A1(n4811), .A2(n4810), .ZN(n7559) );
  AOI21_X1 U5712 ( .B1(n4813), .B2(n4815), .A(n4465), .ZN(n4810) );
  AOI21_X1 U5713 ( .B1(n4560), .B2(n8857), .A(n4558), .ZN(n4557) );
  INV_X1 U5714 ( .A(n4456), .ZN(n4558) );
  NAND2_X1 U5715 ( .A1(n7457), .A2(n4560), .ZN(n4559) );
  AND2_X1 U5716 ( .A1(n7463), .A2(n9666), .ZN(n7513) );
  INV_X1 U5717 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U5718 ( .A1(n5364), .A2(n5363), .ZN(n7354) );
  OR2_X1 U5719 ( .A1(n7351), .A2(n7354), .ZN(n7352) );
  NOR2_X1 U5720 ( .A1(n7256), .A2(n7548), .ZN(n7214) );
  AND2_X1 U5721 ( .A1(n5317), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U5722 ( .A1(n8928), .A2(n4575), .ZN(n7187) );
  INV_X1 U5723 ( .A(n8851), .ZN(n4574) );
  AND2_X1 U5724 ( .A1(n4904), .A2(n4903), .ZN(n7194) );
  AND2_X1 U5725 ( .A1(n5127), .A2(n4472), .ZN(n4903) );
  NAND2_X1 U5726 ( .A1(n4906), .A2(n4905), .ZN(n4904) );
  NAND2_X1 U5727 ( .A1(n4540), .A2(n7247), .ZN(n8751) );
  INV_X1 U5728 ( .A(n7248), .ZN(n4540) );
  AND4_X1 U5729 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n7443)
         );
  NAND2_X1 U5730 ( .A1(n7099), .A2(n7148), .ZN(n7153) );
  OR3_X1 U5731 ( .A1(n9570), .A2(n9560), .A3(n8919), .ZN(n7073) );
  NOR2_X1 U5732 ( .A1(n7073), .A2(n7060), .ZN(n7066) );
  OAI21_X1 U5733 ( .B1(n4658), .B2(n4659), .A(n6437), .ZN(n4657) );
  NOR2_X1 U5734 ( .A1(n4660), .A2(n6472), .ZN(n4659) );
  INV_X1 U5735 ( .A(n9487), .ZN(n9546) );
  NAND2_X1 U5736 ( .A1(n5515), .A2(n5514), .ZN(n9377) );
  NAND2_X1 U5737 ( .A1(n5529), .A2(n5528), .ZN(n9384) );
  AND2_X1 U5738 ( .A1(n5316), .A2(n5315), .ZN(n9636) );
  OR2_X1 U5739 ( .A1(n8823), .A2(n6470), .ZN(n5199) );
  AND2_X1 U5740 ( .A1(n9561), .A2(n5738), .ZN(n9625) );
  INV_X1 U5741 ( .A(n9625), .ZN(n9665) );
  NAND2_X1 U5742 ( .A1(n6172), .A2(n4610), .ZN(n4603) );
  OR2_X1 U5743 ( .A1(n6172), .A2(n4611), .ZN(n4604) );
  XNOR2_X1 U5744 ( .A(n5823), .B(n5822), .ZN(n7575) );
  AND2_X2 U5745 ( .A1(n5361), .A2(n4415), .ZN(n5456) );
  OAI21_X1 U5746 ( .B1(n5604), .B2(n5603), .A(n5602), .ZN(n5619) );
  INV_X1 U5747 ( .A(SI_20_), .ZN(n5578) );
  INV_X1 U5748 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U5749 ( .A1(n5382), .A2(n5045), .ZN(n5412) );
  NAND2_X1 U5750 ( .A1(n4584), .A2(n4586), .ZN(n5404) );
  OR2_X1 U5751 ( .A1(n5333), .A2(n4931), .ZN(n4584) );
  NAND2_X1 U5752 ( .A1(n4937), .A2(n5331), .ZN(n5357) );
  NAND2_X1 U5753 ( .A1(n4938), .A2(n5329), .ZN(n4937) );
  INV_X1 U5754 ( .A(n5333), .ZN(n4938) );
  INV_X1 U5755 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10146) );
  AND2_X1 U5756 ( .A1(n7236), .A2(n7235), .ZN(n7239) );
  INV_X1 U5757 ( .A(n7699), .ZN(n5000) );
  NAND2_X1 U5758 ( .A1(n7854), .A2(n7671), .ZN(n5001) );
  INV_X1 U5759 ( .A(n8298), .ZN(n7736) );
  AND2_X1 U5760 ( .A1(n4999), .A2(n4443), .ZN(n7735) );
  NAND2_X1 U5761 ( .A1(n4999), .A2(n4998), .ZN(n7733) );
  XNOR2_X1 U5762 ( .A(n8165), .B(n7664), .ZN(n7675) );
  AND4_X1 U5763 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8237)
         );
  NAND2_X1 U5764 ( .A1(n4994), .A2(n4995), .ZN(n7806) );
  OR2_X1 U5765 ( .A1(n7843), .A2(n4997), .ZN(n4994) );
  AOI21_X1 U5766 ( .B1(n4407), .B2(n7823), .A(n7824), .ZN(n7826) );
  NAND2_X1 U5767 ( .A1(n6079), .A2(n6078), .ZN(n8287) );
  INV_X1 U5768 ( .A(n8185), .ZN(n7861) );
  NAND2_X1 U5769 ( .A1(n6721), .A2(n6743), .ZN(n7860) );
  INV_X1 U5770 ( .A(n7852), .ZN(n7866) );
  NAND2_X1 U5771 ( .A1(n4918), .A2(n4920), .ZN(n4526) );
  INV_X1 U5772 ( .A(n7764), .ZN(n8226) );
  OAI211_X1 U5773 ( .C1(n5870), .C2(n10240), .A(n6141), .B(n6140), .ZN(n8215)
         );
  INV_X1 U5774 ( .A(n8284), .ZN(n8262) );
  INV_X1 U5775 ( .A(n8310), .ZN(n8102) );
  AND4_X1 U5776 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n7728)
         );
  NAND4_X1 U5777 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n8106)
         );
  INV_X1 U5778 ( .A(n7273), .ZN(n8110) );
  NAND2_X1 U5779 ( .A1(n6753), .A2(n4835), .ZN(n9731) );
  AND2_X1 U5780 ( .A1(n4857), .A2(n4856), .ZN(n9755) );
  NAND2_X1 U5781 ( .A1(n6757), .A2(n4859), .ZN(n4858) );
  NOR2_X1 U5782 ( .A1(n9740), .A2(n4734), .ZN(n9762) );
  NOR2_X1 U5783 ( .A1(n9772), .A2(n9771), .ZN(n9770) );
  NAND2_X1 U5784 ( .A1(n4722), .A2(n4723), .ZN(n9777) );
  AND2_X1 U5785 ( .A1(n6885), .A2(n6371), .ZN(n9779) );
  INV_X1 U5786 ( .A(n6405), .ZN(n4890) );
  NOR2_X1 U5787 ( .A1(n9826), .A2(n8357), .ZN(n9825) );
  INV_X1 U5788 ( .A(n6412), .ZN(n4895) );
  OAI21_X1 U5789 ( .B1(n9826), .B2(n4729), .A(n4728), .ZN(n8114) );
  NAND2_X1 U5790 ( .A1(n4730), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5791 ( .A1(n6382), .A2(n4730), .ZN(n4728) );
  INV_X1 U5792 ( .A(n8115), .ZN(n4730) );
  NOR2_X1 U5793 ( .A1(n9843), .A2(n8322), .ZN(n9842) );
  INV_X1 U5794 ( .A(n4869), .ZN(n8139) );
  OAI21_X1 U5795 ( .B1(n9843), .B2(n4719), .A(n4718), .ZN(n8130) );
  NAND2_X1 U5796 ( .A1(n4720), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5797 ( .A1(n6385), .A2(n4720), .ZN(n4718) );
  INV_X1 U5798 ( .A(n8131), .ZN(n4720) );
  AND2_X1 U5799 ( .A1(P2_U3893), .A2(n8544), .ZN(n9868) );
  NAND2_X1 U5800 ( .A1(n4637), .A2(n6236), .ZN(n7893) );
  NAND2_X1 U5801 ( .A1(n4645), .A2(n4643), .ZN(n4637) );
  NAND2_X1 U5802 ( .A1(n8260), .A2(n6114), .ZN(n8248) );
  NAND2_X1 U5803 ( .A1(n6116), .A2(n6115), .ZN(n8403) );
  NAND2_X1 U5804 ( .A1(n6094), .A2(n6093), .ZN(n8279) );
  NAND2_X1 U5805 ( .A1(n4654), .A2(n8025), .ZN(n8286) );
  OR2_X1 U5806 ( .A1(n8295), .A2(n7905), .ZN(n4654) );
  NAND2_X1 U5807 ( .A1(n4766), .A2(n6011), .ZN(n8345) );
  AND2_X1 U5808 ( .A1(n4619), .A2(n7978), .ZN(n7384) );
  AND3_X1 U5809 ( .A1(n5957), .A2(n5956), .A3(n5955), .ZN(n9919) );
  OR2_X1 U5810 ( .A1(n5865), .A2(n6480), .ZN(n5957) );
  NAND2_X1 U5811 ( .A1(n4750), .A2(n4752), .ZN(n7047) );
  NAND2_X1 U5812 ( .A1(n4751), .A2(n4503), .ZN(n4750) );
  NAND2_X1 U5813 ( .A1(n4648), .A2(n7964), .ZN(n7046) );
  AND3_X1 U5814 ( .A1(n5904), .A2(n5903), .A3(n5902), .ZN(n9901) );
  INV_X1 U5815 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9891) );
  INV_X1 U5816 ( .A(n8378), .ZN(n9892) );
  NAND2_X1 U5817 ( .A1(n6932), .A2(n8352), .ZN(n8288) );
  INV_X1 U5818 ( .A(n8355), .ZN(n9890) );
  NAND2_X1 U5819 ( .A1(n6041), .A2(n6040), .ZN(n8421) );
  NAND2_X1 U5820 ( .A1(n7881), .A2(n7880), .ZN(n8439) );
  NAND2_X1 U5821 ( .A1(n6174), .A2(n6173), .ZN(n8450) );
  NAND2_X1 U5822 ( .A1(n6145), .A2(n6144), .ZN(n8468) );
  NAND2_X1 U5823 ( .A1(n8259), .A2(n8035), .ZN(n8246) );
  NAND2_X1 U5824 ( .A1(n6106), .A2(n6105), .ZN(n8487) );
  NAND2_X1 U5825 ( .A1(n6070), .A2(n6069), .ZN(n8502) );
  NAND2_X1 U5826 ( .A1(n6057), .A2(n6056), .ZN(n8508) );
  NAND2_X1 U5827 ( .A1(n6028), .A2(n6027), .ZN(n8520) );
  NAND2_X1 U5828 ( .A1(n8365), .A2(n7999), .ZN(n8354) );
  NAND2_X1 U5829 ( .A1(n6003), .A2(n6002), .ZN(n8533) );
  INV_X1 U5830 ( .A(n6808), .ZN(n7291) );
  NAND2_X1 U5831 ( .A1(n8539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  CLKBUF_X1 U5832 ( .A(n6239), .Z(n8544) );
  INV_X1 U5833 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6256) );
  OR2_X1 U5834 ( .A1(n6252), .A2(n5813), .ZN(n6253) );
  INV_X1 U5835 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7507) );
  INV_X1 U5836 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7437) );
  INV_X1 U5837 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10110) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7683) );
  INV_X1 U5839 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6088) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10172) );
  INV_X1 U5841 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6866) );
  INV_X1 U5842 ( .A(n9857), .ZN(n6864) );
  INV_X1 U5843 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10114) );
  INV_X1 U5844 ( .A(n8119), .ZN(n6662) );
  INV_X1 U5845 ( .A(n7528), .ZN(n6507) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6504) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6482) );
  INV_X1 U5848 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6479) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10052) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6463) );
  CLKBUF_X1 U5851 ( .A(n7109), .Z(n4515) );
  NAND2_X1 U5852 ( .A1(n8684), .A2(n8686), .ZN(n8565) );
  XNOR2_X1 U5853 ( .A(n5207), .B(n4953), .ZN(n6788) );
  INV_X1 U5854 ( .A(n4952), .ZN(n6828) );
  AND2_X1 U5855 ( .A1(n7592), .A2(n7591), .ZN(n8607) );
  AND2_X1 U5856 ( .A1(n8599), .A2(n7605), .ZN(n9144) );
  AND4_X1 U5857 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n7447)
         );
  NAND2_X1 U5858 ( .A1(n4952), .A2(n4951), .ZN(n6830) );
  INV_X1 U5859 ( .A(n8986), .ZN(n7404) );
  INV_X1 U5860 ( .A(n9413), .ZN(n4709) );
  CLKBUF_X1 U5861 ( .A(n7538), .Z(n8698) );
  INV_X1 U5862 ( .A(n9483), .ZN(n9102) );
  NAND2_X1 U5863 ( .A1(n5247), .A2(n6938), .ZN(n7038) );
  AOI21_X1 U5864 ( .B1(n4957), .B2(n8639), .A(n4463), .ZN(n4955) );
  AND2_X1 U5865 ( .A1(n5767), .A2(n5745), .ZN(n8722) );
  NAND2_X1 U5866 ( .A1(n5762), .A2(n9626), .ZN(n8737) );
  OR4_X1 U5868 ( .A1(n8960), .A2(n8905), .A3(n8870), .A4(n8869), .ZN(n8908) );
  NAND2_X1 U5869 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  INV_X1 U5870 ( .A(n9232), .ZN(n9363) );
  OR2_X1 U5871 ( .A1(n6450), .A2(n6449), .ZN(n9070) );
  INV_X1 U5872 ( .A(n8829), .ZN(n9306) );
  NAND2_X1 U5873 ( .A1(n8825), .A2(n8824), .ZN(n9098) );
  NAND2_X1 U5874 ( .A1(n4844), .A2(n4845), .ZN(n9148) );
  AND4_X1 U5875 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n9325)
         );
  NAND2_X1 U5876 ( .A1(n4808), .A2(n4806), .ZN(n9141) );
  NAND2_X1 U5877 ( .A1(n4801), .A2(n4418), .ZN(n4808) );
  NAND2_X1 U5878 ( .A1(n9172), .A2(n9126), .ZN(n9160) );
  AND4_X1 U5879 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(n9332)
         );
  AND2_X1 U5880 ( .A1(n4801), .A2(n4809), .ZN(n9154) );
  NAND2_X1 U5881 ( .A1(n5687), .A2(n5686), .ZN(n9346) );
  NAND2_X1 U5882 ( .A1(n4820), .A2(n4824), .ZN(n9198) );
  NAND2_X1 U5883 ( .A1(n9228), .A2(n4825), .ZN(n4820) );
  NAND2_X1 U5884 ( .A1(n4827), .A2(n9109), .ZN(n9211) );
  NAND2_X1 U5885 ( .A1(n4829), .A2(n4828), .ZN(n4827) );
  INV_X1 U5886 ( .A(n9235), .ZN(n9364) );
  INV_X1 U5887 ( .A(n9370), .ZN(n9276) );
  INV_X1 U5888 ( .A(n9108), .ZN(n9245) );
  NAND2_X1 U5889 ( .A1(n4875), .A2(n4876), .ZN(n9241) );
  OR2_X1 U5890 ( .A1(n9272), .A2(n4877), .ZN(n4875) );
  INV_X1 U5891 ( .A(n9488), .ZN(n9503) );
  AND2_X1 U5892 ( .A1(n7553), .A2(n9288), .ZN(n9516) );
  OR2_X1 U5893 ( .A1(n7457), .A2(n8857), .ZN(n4561) );
  NAND2_X1 U5894 ( .A1(n4812), .A2(n4816), .ZN(n7557) );
  NAND2_X1 U5895 ( .A1(n7456), .A2(n4431), .ZN(n4812) );
  AND2_X1 U5896 ( .A1(n4817), .A2(n4819), .ZN(n7518) );
  NAND2_X1 U5897 ( .A1(n7456), .A2(n7455), .ZN(n4817) );
  AND4_X1 U5898 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n9657)
         );
  NAND2_X1 U5899 ( .A1(n4887), .A2(n8767), .ZN(n7349) );
  OR2_X1 U5900 ( .A1(n9553), .A2(n9493), .ZN(n9295) );
  INV_X1 U5901 ( .A(n9286), .ZN(n9480) );
  INV_X1 U5902 ( .A(n9636), .ZN(n7548) );
  NAND2_X1 U5903 ( .A1(n4795), .A2(n7193), .ZN(n7246) );
  NAND2_X1 U5904 ( .A1(n7192), .A2(n7191), .ZN(n4795) );
  INV_X1 U5905 ( .A(n7194), .ZN(n9624) );
  NAND2_X1 U5906 ( .A1(n4695), .A2(n4694), .ZN(n7096) );
  OR2_X1 U5907 ( .A1(n9553), .A2(n9492), .ZN(n9544) );
  NAND2_X1 U5908 ( .A1(n4695), .A2(n7061), .ZN(n7092) );
  OR2_X1 U5909 ( .A1(n9553), .A2(n9656), .ZN(n9248) );
  INV_X1 U5910 ( .A(n9295), .ZN(n9549) );
  INV_X1 U5911 ( .A(n7026), .ZN(n9570) );
  INV_X1 U5912 ( .A(n9544), .ZN(n9291) );
  INV_X1 U5913 ( .A(n9499), .ZN(n9541) );
  NOR2_X1 U5914 ( .A1(n9320), .A2(n4566), .ZN(n9323) );
  OR2_X1 U5915 ( .A1(n9321), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U5916 ( .A1(n5084), .A2(n4517), .ZN(n4516) );
  INV_X1 U5917 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4517) );
  INV_X1 U5918 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9406) );
  INV_X1 U5919 ( .A(n5725), .ZN(n7579) );
  INV_X1 U5920 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U5921 ( .A1(n4939), .A2(n4943), .ZN(n5649) );
  NAND2_X1 U5922 ( .A1(n5604), .A2(n4945), .ZN(n4939) );
  INV_X1 U5923 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7439) );
  INV_X1 U5924 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7294) );
  INV_X1 U5925 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7617) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6918) );
  INV_X1 U5927 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6863) );
  INV_X1 U5928 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6820) );
  INV_X1 U5929 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10143) );
  INV_X1 U5930 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10206) );
  INV_X1 U5931 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6484) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U5933 ( .A1(n4550), .A2(n5113), .ZN(n5278) );
  NAND2_X1 U5934 ( .A1(n5259), .A2(n5258), .ZN(n4550) );
  INV_X1 U5935 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6477) );
  INV_X1 U5936 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U5937 ( .A1(n4949), .A2(n5174), .ZN(n5216) );
  AND2_X1 U5938 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9414) );
  AND2_X2 U5939 ( .A1(n6359), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  NAND2_X1 U5940 ( .A1(n4514), .A2(n4488), .ZN(P2_U3165) );
  INV_X1 U5941 ( .A(n7775), .ZN(n4514) );
  AND2_X1 U5942 ( .A1(n8462), .A2(n7850), .ZN(n4513) );
  INV_X1 U5943 ( .A(n4891), .ZN(n9787) );
  INV_X1 U5944 ( .A(n4896), .ZN(n9819) );
  NAND2_X1 U5945 ( .A1(n6358), .A2(n6420), .ZN(n4534) );
  OAI21_X1 U5946 ( .B1(n8442), .B2(n8340), .A(n4777), .ZN(P2_U3205) );
  INV_X1 U5947 ( .A(n4778), .ZN(n4777) );
  NAND2_X1 U5948 ( .A1(n6293), .A2(n8432), .ZN(n6295) );
  NAND2_X1 U5949 ( .A1(n6293), .A2(n8534), .ZN(n6432) );
  NAND2_X1 U5950 ( .A1(n4868), .A2(n6890), .ZN(n6401) );
  AND2_X1 U5951 ( .A1(n4672), .A2(n4671), .ZN(n4412) );
  AND2_X1 U5952 ( .A1(n5150), .A2(n8969), .ZN(n4413) );
  AND2_X1 U5953 ( .A1(n8468), .A2(n8226), .ZN(n4414) );
  INV_X1 U5954 ( .A(n4931), .ZN(n4930) );
  NAND2_X1 U5955 ( .A1(n4933), .A2(n5379), .ZN(n4931) );
  NAND2_X1 U5956 ( .A1(n6437), .A2(n4660), .ZN(n5311) );
  INV_X1 U5957 ( .A(n7165), .ZN(n9612) );
  AND2_X1 U5958 ( .A1(n5816), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U5959 ( .A1(n8273), .A2(n4763), .ZN(n8260) );
  INV_X1 U5960 ( .A(n7120), .ZN(n7121) );
  AND2_X1 U5961 ( .A1(n4929), .A2(n4435), .ZN(n4417) );
  AND2_X1 U5962 ( .A1(n9114), .A2(n4809), .ZN(n4418) );
  NOR2_X1 U5963 ( .A1(n9778), .A2(n4726), .ZN(n4419) );
  INV_X1 U5964 ( .A(n9110), .ZN(n4828) );
  NOR2_X1 U5965 ( .A1(n9235), .A2(n9356), .ZN(n9110) );
  AND2_X1 U5966 ( .A1(n6422), .A2(n6421), .ZN(n4420) );
  INV_X1 U5967 ( .A(n4885), .ZN(n4884) );
  NAND2_X1 U5968 ( .A1(n4886), .A2(n8767), .ZN(n4885) );
  NOR2_X1 U5969 ( .A1(n8891), .A2(n8831), .ZN(n4421) );
  AND2_X1 U5970 ( .A1(n7978), .A2(n7973), .ZN(n4422) );
  INV_X1 U5971 ( .A(n5014), .ZN(n5013) );
  OR2_X1 U5972 ( .A1(n5015), .A2(n7658), .ZN(n5014) );
  AND2_X1 U5973 ( .A1(n8768), .A2(n8936), .ZN(n4423) );
  NAND2_X1 U5974 ( .A1(n4448), .A2(n9109), .ZN(n4826) );
  NAND2_X1 U5975 ( .A1(n4717), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U5976 ( .A1(n7194), .A2(n8987), .ZN(n8765) );
  AND2_X1 U5977 ( .A1(n5031), .A2(n10094), .ZN(n4424) );
  NOR2_X1 U5978 ( .A1(n8087), .A2(n6729), .ZN(n4425) );
  OR2_X1 U5979 ( .A1(n4727), .A2(n5946), .ZN(n4426) );
  AND2_X1 U5980 ( .A1(n5656), .A2(n5655), .ZN(n9208) );
  INV_X1 U5981 ( .A(n9208), .ZN(n9353) );
  INV_X1 U5982 ( .A(n9514), .ZN(n8981) );
  AND4_X1 U5983 ( .A1(n5443), .A2(n5442), .A3(n5441), .A4(n5440), .ZN(n9514)
         );
  OR2_X1 U5984 ( .A1(n6400), .A2(n9945), .ZN(n4427) );
  INV_X1 U5985 ( .A(n5830), .ZN(n4917) );
  NAND2_X1 U5986 ( .A1(n4909), .A2(n4907), .ZN(n7891) );
  OR2_X2 U5987 ( .A1(n5815), .A2(n5816), .ZN(n5869) );
  INV_X1 U5988 ( .A(n6462), .ZN(n4855) );
  NAND2_X1 U5989 ( .A1(n5917), .A2(n5798), .ZN(n5919) );
  OR2_X1 U5990 ( .A1(n9377), .A2(n9276), .ZN(n4428) );
  AND2_X1 U5991 ( .A1(n5103), .A2(SI_3_), .ZN(n4429) );
  OR2_X1 U5992 ( .A1(n9335), .A2(n9175), .ZN(n4430) );
  AND2_X1 U5993 ( .A1(n4818), .A2(n7455), .ZN(n4431) );
  NAND2_X1 U5994 ( .A1(n6169), .A2(n6168), .ZN(n8197) );
  INV_X1 U5995 ( .A(n8197), .ZN(n7856) );
  INV_X1 U5996 ( .A(n4807), .ZN(n4806) );
  NAND2_X1 U5997 ( .A1(n9147), .A2(n4430), .ZN(n4807) );
  OR2_X1 U5998 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4432) );
  NOR2_X1 U5999 ( .A1(n8106), .A2(n7730), .ZN(n4433) );
  AND4_X1 U6000 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5077), .ZN(n4434)
         );
  NAND2_X1 U6001 ( .A1(n8808), .A2(n8807), .ZN(n9322) );
  OR2_X1 U6002 ( .A1(n5475), .A2(SI_16_), .ZN(n4435) );
  INV_X1 U6003 ( .A(n9267), .ZN(n4548) );
  AND2_X1 U6004 ( .A1(n6207), .A2(n6209), .ZN(n4436) );
  NAND2_X1 U6005 ( .A1(n5456), .A2(n5071), .ZN(n4437) );
  INV_X1 U6006 ( .A(n9724), .ZN(n4838) );
  NAND2_X1 U6007 ( .A1(n4770), .A2(n6133), .ZN(n8224) );
  INV_X1 U6008 ( .A(n9228), .ZN(n4829) );
  AND3_X1 U6009 ( .A1(n8829), .A2(n9130), .A3(n9098), .ZN(n4438) );
  NAND4_X1 U6010 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n9885)
         );
  INV_X1 U6011 ( .A(n9885), .ZN(n4753) );
  AND2_X1 U6012 ( .A1(n8899), .A2(n8871), .ZN(n9118) );
  OR2_X1 U6013 ( .A1(n8881), .A2(n8831), .ZN(n4439) );
  AND2_X1 U6014 ( .A1(n8462), .A2(n8214), .ZN(n4440) );
  OR2_X1 U6015 ( .A1(n5919), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4441) );
  AND2_X1 U6016 ( .A1(n4873), .A2(n4548), .ZN(n4442) );
  NAND2_X1 U6017 ( .A1(n7654), .A2(n7736), .ZN(n4443) );
  OAI21_X1 U6018 ( .B1(n4406), .B2(n5017), .A(n5016), .ZN(n7469) );
  AND2_X1 U6019 ( .A1(n9666), .A2(n8738), .ZN(n4444) );
  NAND2_X1 U6020 ( .A1(n5845), .A2(n5846), .ZN(n5854) );
  NOR2_X1 U6021 ( .A1(n8779), .A2(n8778), .ZN(n4445) );
  INV_X1 U6022 ( .A(n4860), .ZN(n4859) );
  AND2_X1 U6023 ( .A1(n7671), .A2(n5000), .ZN(n4446) );
  AND2_X1 U6024 ( .A1(n4808), .A2(n4430), .ZN(n4447) );
  AND2_X1 U6025 ( .A1(n8893), .A2(n8780), .ZN(n8895) );
  AND2_X1 U6026 ( .A1(n8456), .A2(n7856), .ZN(n8062) );
  NAND2_X1 U6027 ( .A1(n6161), .A2(n6160), .ZN(n8456) );
  OR2_X1 U6028 ( .A1(n9213), .A2(n9226), .ZN(n4448) );
  INV_X1 U6029 ( .A(n9122), .ZN(n4872) );
  AND2_X1 U6030 ( .A1(n9213), .A2(n9226), .ZN(n4449) );
  AND2_X1 U6031 ( .A1(n8003), .A2(n8002), .ZN(n8353) );
  INV_X1 U6032 ( .A(n4854), .ZN(n4853) );
  NOR2_X1 U6033 ( .A1(n4859), .A2(n4855), .ZN(n4854) );
  NOR2_X1 U6034 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4450) );
  OR2_X1 U6035 ( .A1(n5870), .A2(n6391), .ZN(n4451) );
  AND2_X1 U6036 ( .A1(n7447), .A2(n7194), .ZN(n4452) );
  NOR2_X1 U6037 ( .A1(n7360), .A2(n8109), .ZN(n4453) );
  XNOR2_X1 U6038 ( .A(n7688), .B(SI_29_), .ZN(n7619) );
  NOR2_X1 U6039 ( .A1(n7655), .A2(n8284), .ZN(n4454) );
  NAND2_X1 U6040 ( .A1(n8796), .A2(n8797), .ZN(n4455) );
  INV_X1 U6041 ( .A(n5008), .ZN(n5007) );
  OR2_X1 U6042 ( .A1(n7663), .A2(n5009), .ZN(n5008) );
  INV_X1 U6043 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10094) );
  INV_X1 U6044 ( .A(n9619), .ZN(n7177) );
  AND2_X1 U6045 ( .A1(n4577), .A2(n4576), .ZN(n9619) );
  INV_X1 U6046 ( .A(n9522), .ZN(n7558) );
  AND2_X1 U6047 ( .A1(n5437), .A2(n5436), .ZN(n9522) );
  OR2_X1 U6048 ( .A1(n7558), .A2(n9514), .ZN(n4456) );
  NAND2_X1 U6049 ( .A1(n5456), .A2(n4434), .ZN(n4457) );
  XNOR2_X1 U6050 ( .A(n6172), .B(n6171), .ZN(n7580) );
  OR2_X1 U6051 ( .A1(n9509), .A2(n9102), .ZN(n4458) );
  INV_X1 U6052 ( .A(n4663), .ZN(n4662) );
  NAND2_X1 U6053 ( .A1(n7148), .A2(n9604), .ZN(n4663) );
  AND2_X1 U6054 ( .A1(n5381), .A2(SI_12_), .ZN(n4459) );
  AND2_X1 U6055 ( .A1(n9328), .A2(n9117), .ZN(n4460) );
  AND2_X1 U6056 ( .A1(n6264), .A2(n6263), .ZN(n6274) );
  INV_X1 U6057 ( .A(n6274), .ZN(n4527) );
  AND2_X1 U6058 ( .A1(n8456), .A2(n8197), .ZN(n4461) );
  NAND2_X1 U6059 ( .A1(n7662), .A2(n7771), .ZN(n4462) );
  NAND2_X1 U6060 ( .A1(n5748), .A2(n5746), .ZN(n4463) );
  NOR2_X1 U6061 ( .A1(n9522), .A2(n9514), .ZN(n4464) );
  AND2_X1 U6062 ( .A1(n9522), .A2(n9514), .ZN(n4465) );
  NAND2_X1 U6063 ( .A1(n5431), .A2(SI_15_), .ZN(n4466) );
  INV_X1 U6064 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6065 ( .A1(n4444), .A2(n7454), .ZN(n4467) );
  OR2_X1 U6066 ( .A1(n4414), .A2(n4440), .ZN(n4468) );
  NAND2_X1 U6067 ( .A1(n9159), .A2(n4847), .ZN(n4469) );
  NAND2_X1 U6068 ( .A1(n4687), .A2(n4684), .ZN(n4470) );
  NAND2_X1 U6069 ( .A1(n7891), .A2(n7892), .ZN(n8068) );
  NAND2_X1 U6070 ( .A1(n8898), .A2(n9128), .ZN(n9147) );
  INV_X1 U6071 ( .A(n9147), .ZN(n4843) );
  AND2_X1 U6072 ( .A1(n8273), .A2(n6104), .ZN(n4471) );
  NAND2_X1 U6073 ( .A1(n8587), .A2(n8586), .ZN(n9328) );
  AND2_X1 U6074 ( .A1(n7327), .A2(n7979), .ZN(n7972) );
  OR2_X1 U6075 ( .A1(n6437), .A2(n6595), .ZN(n4472) );
  AND2_X1 U6076 ( .A1(n8077), .A2(n7891), .ZN(n4473) );
  NOR2_X1 U6077 ( .A1(n4961), .A2(n4958), .ZN(n4474) );
  OR2_X1 U6078 ( .A1(n6437), .A2(n6582), .ZN(n4475) );
  AND2_X1 U6079 ( .A1(n8089), .A2(n6729), .ZN(n4476) );
  NAND2_X1 U6080 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4477) );
  OR2_X1 U6081 ( .A1(n9101), .A2(n8661), .ZN(n8891) );
  AND2_X1 U6082 ( .A1(n4415), .A2(n4450), .ZN(n4478) );
  AND2_X1 U6083 ( .A1(n4716), .A2(n6387), .ZN(n4479) );
  AND2_X1 U6084 ( .A1(n4733), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4480) );
  AND2_X1 U6085 ( .A1(n8564), .A2(n4959), .ZN(n4481) );
  AND2_X1 U6086 ( .A1(n8891), .A2(n8942), .ZN(n8861) );
  INV_X1 U6087 ( .A(n7664), .ZN(n7667) );
  INV_X1 U6088 ( .A(n9301), .ZN(n9494) );
  NAND2_X1 U6089 ( .A1(n5625), .A2(n5624), .ZN(n9213) );
  INV_X1 U6090 ( .A(n9213), .ZN(n4671) );
  INV_X1 U6091 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5047) );
  XNOR2_X1 U6092 ( .A(n6381), .B(n9822), .ZN(n9826) );
  OR2_X1 U6093 ( .A1(n9208), .A2(n9191), .ZN(n4482) );
  INV_X1 U6094 ( .A(n8854), .ZN(n4886) );
  AND2_X1 U6095 ( .A1(n4561), .A2(n4562), .ZN(n4483) );
  AND2_X1 U6096 ( .A1(n4559), .A2(n4557), .ZN(n4484) );
  NAND2_X1 U6097 ( .A1(n6159), .A2(n6158), .ZN(n8214) );
  AND2_X1 U6098 ( .A1(n8912), .A2(n9493), .ZN(n8826) );
  AND2_X1 U6099 ( .A1(n7656), .A2(n8252), .ZN(n4485) );
  NOR2_X1 U6100 ( .A1(n9825), .A2(n6382), .ZN(n4486) );
  NOR2_X1 U6101 ( .A1(n9842), .A2(n6385), .ZN(n4487) );
  NOR2_X1 U6102 ( .A1(n7776), .A2(n4513), .ZN(n4488) );
  NAND2_X1 U6103 ( .A1(n9256), .A2(n4412), .ZN(n4673) );
  AND2_X1 U6104 ( .A1(n5416), .A2(n5415), .ZN(n9666) );
  INV_X1 U6105 ( .A(n9666), .ZN(n7517) );
  AND2_X1 U6106 ( .A1(n4654), .A2(n4652), .ZN(n4489) );
  NAND2_X1 U6107 ( .A1(n8891), .A2(n4456), .ZN(n4490) );
  NAND2_X1 U6108 ( .A1(n5710), .A2(n5709), .ZN(n9339) );
  INV_X1 U6109 ( .A(n4596), .ZN(n4595) );
  NAND2_X1 U6110 ( .A1(n4943), .A2(n4597), .ZN(n4596) );
  AND2_X1 U6111 ( .A1(n4896), .A2(n4895), .ZN(n4491) );
  NAND2_X1 U6112 ( .A1(n5840), .A2(n5839), .ZN(n8444) );
  NAND2_X1 U6113 ( .A1(n5486), .A2(n5485), .ZN(n9292) );
  INV_X1 U6114 ( .A(n9292), .ZN(n9509) );
  INV_X1 U6115 ( .A(n4826), .ZN(n4825) );
  NAND2_X1 U6116 ( .A1(n5459), .A2(n5458), .ZN(n9101) );
  INV_X1 U6117 ( .A(n9101), .ZN(n4668) );
  AOI21_X1 U6118 ( .B1(n4945), .B2(n5603), .A(n4944), .ZN(n4943) );
  OR2_X1 U6119 ( .A1(n5412), .A2(n5048), .ZN(n4492) );
  INV_X1 U6120 ( .A(SI_15_), .ZN(n5452) );
  NAND2_X1 U6121 ( .A1(n8629), .A2(n8628), .ZN(n4493) );
  AND2_X1 U6122 ( .A1(n5475), .A2(SI_16_), .ZN(n4494) );
  NAND2_X1 U6123 ( .A1(n9339), .A2(n9185), .ZN(n4809) );
  INV_X1 U6124 ( .A(n6293), .ZN(n8157) );
  NAND2_X1 U6125 ( .A1(n4909), .A2(n6190), .ZN(n6293) );
  AND2_X1 U6126 ( .A1(n8170), .A2(n4779), .ZN(n4495) );
  AND2_X1 U6127 ( .A1(n6265), .A2(n6489), .ZN(n6726) );
  NOR2_X1 U6128 ( .A1(n6361), .A2(n8548), .ZN(n9863) );
  AOI21_X1 U6129 ( .B1(n6258), .B2(n7571), .A(n4527), .ZN(n6275) );
  NAND2_X1 U6130 ( .A1(n4619), .A2(n4618), .ZN(n7383) );
  AND2_X1 U6131 ( .A1(n7099), .A2(n4662), .ZN(n4496) );
  NAND2_X1 U6132 ( .A1(n4789), .A2(n4792), .ZN(n7207) );
  NAND2_X1 U6133 ( .A1(n4746), .A2(n4745), .ZN(n7129) );
  AND2_X1 U6134 ( .A1(n6187), .A2(n4917), .ZN(n4497) );
  AND2_X1 U6135 ( .A1(n4768), .A2(n5945), .ZN(n4498) );
  NAND2_X1 U6136 ( .A1(n7236), .A2(n5018), .ZN(n7361) );
  NAND2_X1 U6137 ( .A1(n4406), .A2(n7121), .ZN(n7236) );
  AND2_X1 U6138 ( .A1(n4891), .A2(n4890), .ZN(n4499) );
  AND2_X1 U6139 ( .A1(n6189), .A2(n6188), .ZN(n4500) );
  AND2_X1 U6140 ( .A1(n7978), .A2(n7979), .ZN(n7918) );
  AND2_X1 U6141 ( .A1(n4607), .A2(n4605), .ZN(n4501) );
  INV_X1 U6142 ( .A(n7454), .ZN(n4819) );
  OR2_X1 U6143 ( .A1(n9388), .A2(n9313), .ZN(n9697) );
  INV_X1 U6144 ( .A(n9697), .ZN(n9381) );
  INV_X1 U6145 ( .A(n5768), .ZN(n6957) );
  INV_X1 U6146 ( .A(n9872), .ZN(n4902) );
  NAND2_X1 U6147 ( .A1(n7945), .A2(n7912), .ZN(n6838) );
  OR2_X1 U6148 ( .A1(n4753), .A2(n9901), .ZN(n4503) );
  AND2_X1 U6149 ( .A1(n7006), .A2(n8969), .ZN(n9557) );
  INV_X1 U6150 ( .A(n9557), .ZN(n9486) );
  AND2_X1 U6151 ( .A1(n8828), .A2(n9130), .ZN(n4504) );
  OR2_X1 U6152 ( .A1(n6416), .A2(n8417), .ZN(n4505) );
  NAND2_X1 U6153 ( .A1(n7085), .A2(n9595), .ZN(n8923) );
  XNOR2_X1 U6154 ( .A(n6210), .B(n6209), .ZN(n8088) );
  AND3_X1 U6155 ( .A1(n4851), .A2(n4853), .A3(n4849), .ZN(n4506) );
  AOI21_X1 U6156 ( .B1(n6604), .B2(n6396), .A(n4838), .ZN(n4834) );
  AND2_X1 U6157 ( .A1(n6759), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4507) );
  INV_X1 U6158 ( .A(n4834), .ZN(n6753) );
  NOR2_X1 U6159 ( .A1(n5057), .A2(n4516), .ZN(n9404) );
  INV_X1 U6160 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4710) );
  INV_X1 U6161 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4726) );
  INV_X1 U6162 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5811) );
  AOI21_X1 U6163 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n9780), .A(n9770), .ZN(
        n6404) );
  INV_X1 U6164 ( .A(n5845), .ZN(n4870) );
  NAND2_X1 U6165 ( .A1(n4713), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4711) );
  INV_X1 U6166 ( .A(n9472), .ZN(n9470) );
  NAND2_X1 U6167 ( .A1(n4712), .A2(n6758), .ZN(n6762) );
  NOR2_X1 U6168 ( .A1(n9807), .A2(n6380), .ZN(n7523) );
  INV_X1 U6169 ( .A(n6423), .ZN(n4899) );
  OAI21_X1 U6170 ( .B1(n9861), .B2(n10211), .A(n6387), .ZN(n4714) );
  NAND2_X1 U6171 ( .A1(n8646), .A2(n8647), .ZN(n8645) );
  NAND2_X1 U6172 ( .A1(n4991), .A2(n4990), .ZN(n7741) );
  NAND2_X1 U6173 ( .A1(n4956), .A2(n4955), .ZN(n7600) );
  AOI21_X1 U6174 ( .B1(n4526), .B2(n4425), .A(n4476), .ZN(n8091) );
  NAND2_X1 U6175 ( .A1(n4542), .A2(n5107), .ZN(n5237) );
  NAND2_X1 U6176 ( .A1(n4919), .A2(n8086), .ZN(n4918) );
  NAND2_X1 U6177 ( .A1(n4554), .A2(n5116), .ZN(n5293) );
  OAI21_X1 U6178 ( .B1(n7983), .B2(n7984), .A(n7988), .ZN(n7993) );
  NAND2_X1 U6179 ( .A1(n4522), .A2(n4519), .ZN(n8030) );
  OAI21_X1 U6180 ( .B1(n8022), .B2(n8021), .A(n4521), .ZN(n4520) );
  NAND2_X1 U6181 ( .A1(n4869), .A2(n4505), .ZN(n6418) );
  NOR2_X1 U6182 ( .A1(n9755), .A2(n9754), .ZN(n9753) );
  NAND2_X1 U6183 ( .A1(n4534), .A2(n4531), .ZN(P2_U3200) );
  NOR2_X1 U6184 ( .A1(n9804), .A2(n6300), .ZN(n9803) );
  NAND2_X1 U6185 ( .A1(n6229), .A2(n8047), .ZN(n8054) );
  OAI21_X1 U6186 ( .B1(n5259), .B2(n4553), .A(n4551), .ZN(n4554) );
  OAI21_X1 U6187 ( .B1(n5258), .B2(n4553), .A(n5277), .ZN(n4552) );
  AOI21_X1 U6188 ( .B1(n8060), .B2(n8059), .A(n8180), .ZN(n8065) );
  NOR2_X4 U6189 ( .A1(n7777), .A2(n7778), .ZN(n7787) );
  NAND2_X1 U6190 ( .A1(n5010), .A2(n5011), .ZN(n7767) );
  AOI21_X2 U6191 ( .B1(n7038), .B2(n7035), .A(n7034), .ZN(n7109) );
  NAND2_X1 U6192 ( .A1(n8638), .A2(n8639), .ZN(n5747) );
  NAND2_X1 U6193 ( .A1(n6418), .A2(n6864), .ZN(n6417) );
  NAND2_X1 U6194 ( .A1(n4848), .A2(n4851), .ZN(n4857) );
  NAND2_X1 U6195 ( .A1(n4866), .A2(n4865), .ZN(n4867) );
  NOR2_X1 U6196 ( .A1(n9836), .A2(n6415), .ZN(n8141) );
  NAND2_X1 U6197 ( .A1(n6405), .A2(n4892), .ZN(n4888) );
  OAI21_X1 U6198 ( .B1(n9788), .B2(n4889), .A(n4888), .ZN(n7488) );
  NAND2_X1 U6199 ( .A1(n5101), .A2(n5100), .ZN(n5192) );
  AND2_X1 U6200 ( .A1(n7964), .A2(n7957), .ZN(n7950) );
  OAI21_X1 U6201 ( .B1(n8084), .B2(n4923), .A(n4922), .ZN(n4921) );
  INV_X1 U6202 ( .A(n4912), .ZN(n5219) );
  NOR2_X1 U6203 ( .A1(n9828), .A2(n9829), .ZN(n9827) );
  NOR2_X1 U6204 ( .A1(n9759), .A2(n9758), .ZN(n9757) );
  NOR2_X1 U6205 ( .A1(n9727), .A2(n9728), .ZN(n9726) );
  NOR2_X1 U6206 ( .A1(n7493), .A2(n7494), .ZN(n7492) );
  NOR2_X1 U6207 ( .A1(n8117), .A2(n8118), .ZN(n8116) );
  OAI21_X1 U6208 ( .B1(n8132), .B2(n8134), .A(n6345), .ZN(n9867) );
  NAND2_X1 U6209 ( .A1(n4537), .A2(n5805), .ZN(n6198) );
  NAND2_X1 U6210 ( .A1(n4678), .A2(n8897), .ZN(n4677) );
  NAND2_X1 U6211 ( .A1(n4685), .A2(n4688), .ZN(n8766) );
  INV_X1 U6212 ( .A(n4694), .ZN(n4693) );
  INV_X1 U6213 ( .A(n8783), .ZN(n8784) );
  AOI21_X1 U6214 ( .B1(n4675), .B2(n4674), .A(n9229), .ZN(n8793) );
  NAND3_X1 U6215 ( .A1(n8795), .A2(n8794), .A3(n9126), .ZN(n4541) );
  NAND2_X1 U6216 ( .A1(n4578), .A2(n4543), .ZN(n4542) );
  INV_X1 U6217 ( .A(n4544), .ZN(n4543) );
  OAI21_X1 U6218 ( .B1(n5191), .B2(n4429), .A(n5218), .ZN(n4544) );
  NAND2_X1 U6219 ( .A1(n4546), .A2(n4871), .ZN(n4545) );
  NAND2_X1 U6220 ( .A1(n4549), .A2(n4442), .ZN(n4546) );
  NAND2_X1 U6221 ( .A1(n9271), .A2(n9269), .ZN(n4549) );
  NAND2_X1 U6222 ( .A1(n4547), .A2(n4871), .ZN(n9224) );
  NAND2_X1 U6223 ( .A1(n4549), .A2(n4442), .ZN(n4547) );
  OAI21_X1 U6224 ( .B1(n4557), .B2(n8892), .A(n8891), .ZN(n4556) );
  AOI21_X1 U6225 ( .B1(n7457), .B2(n8937), .A(n8857), .ZN(n7511) );
  MUX2_X1 U6226 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7885), .Z(n5103) );
  NAND2_X1 U6227 ( .A1(n9415), .A2(n5092), .ZN(n4565) );
  NAND3_X1 U6228 ( .A1(n4575), .A2(n4574), .A3(n8928), .ZN(n7210) );
  NAND2_X1 U6229 ( .A1(n7151), .A2(n8924), .ZN(n7169) );
  NAND2_X1 U6230 ( .A1(n4910), .A2(n5101), .ZN(n4578) );
  NAND2_X1 U6231 ( .A1(n5333), .A2(n4586), .ZN(n4583) );
  NAND2_X1 U6232 ( .A1(n4583), .A2(n4585), .ZN(n5407) );
  MUX2_X1 U6233 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n7885), .Z(n5156) );
  NAND2_X1 U6234 ( .A1(n5579), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U6235 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  NAND3_X1 U6236 ( .A1(n4602), .A2(n4601), .A3(n4905), .ZN(n8587) );
  NAND2_X1 U6237 ( .A1(n6172), .A2(n4501), .ZN(n4601) );
  NAND3_X1 U6238 ( .A1(n4604), .A2(n4603), .A3(n4607), .ZN(n8585) );
  INV_X1 U6239 ( .A(n6896), .ZN(n9878) );
  AND2_X2 U6240 ( .A1(n7942), .A2(n7940), .ZN(n6896) );
  NAND2_X1 U6241 ( .A1(n8361), .A2(n4631), .ZN(n4628) );
  NAND2_X1 U6242 ( .A1(n4628), .A2(n4629), .ZN(n8327) );
  NAND2_X1 U6243 ( .A1(n8171), .A2(n7903), .ZN(n4645) );
  NAND2_X1 U6244 ( .A1(n4634), .A2(n4635), .ZN(n7899) );
  NAND2_X1 U6245 ( .A1(n8171), .A2(n4636), .ZN(n4634) );
  AND2_X1 U6246 ( .A1(n4645), .A2(n4644), .ZN(n8164) );
  NAND2_X1 U6247 ( .A1(n6928), .A2(n7957), .ZN(n4648) );
  NAND2_X1 U6248 ( .A1(n4648), .A2(n4646), .ZN(n6218) );
  AND4_X1 U6249 ( .A1(n5808), .A2(n4782), .A3(n5917), .A4(n4424), .ZN(n5831)
         );
  NAND3_X1 U6250 ( .A1(n4782), .A2(n5808), .A3(n4655), .ZN(n8539) );
  NOR2_X1 U6251 ( .A1(n9192), .A2(n4664), .ZN(n9142) );
  INV_X1 U6252 ( .A(n4673), .ZN(n9212) );
  AOI21_X1 U6253 ( .B1(n8756), .B2(n4684), .A(n4683), .ZN(n4682) );
  NAND2_X1 U6254 ( .A1(n8756), .A2(n8831), .ZN(n4685) );
  INV_X1 U6255 ( .A(n8923), .ZN(n4689) );
  INV_X1 U6256 ( .A(n7058), .ZN(n4690) );
  INV_X1 U6257 ( .A(n7061), .ZN(n4691) );
  OAI21_X1 U6258 ( .B1(n4693), .B2(n7059), .A(n4692), .ZN(n7093) );
  NAND2_X1 U6259 ( .A1(n8763), .A2(n4702), .ZN(n4696) );
  NAND2_X1 U6260 ( .A1(n8776), .A2(n4698), .ZN(n4697) );
  NAND3_X1 U6261 ( .A1(n4697), .A2(n4700), .A3(n4696), .ZN(n4701) );
  NAND2_X1 U6262 ( .A1(n8938), .A2(n8831), .ZN(n4703) );
  NAND2_X1 U6263 ( .A1(n8931), .A2(n7186), .ZN(n9534) );
  MUX2_X1 U6264 ( .A(n4710), .B(n4709), .S(n6437), .Z(n6947) );
  NOR2_X2 U6265 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5845) );
  NAND2_X1 U6266 ( .A1(n4711), .A2(n6759), .ZN(n4712) );
  NAND2_X1 U6267 ( .A1(n4713), .A2(n6759), .ZN(n9718) );
  INV_X1 U6268 ( .A(n9861), .ZN(n4717) );
  INV_X1 U6269 ( .A(n9780), .ZN(n4727) );
  NAND2_X1 U6270 ( .A1(n9738), .A2(n4480), .ZN(n4732) );
  NAND2_X1 U6271 ( .A1(n8212), .A2(n4738), .ZN(n4736) );
  AOI21_X1 U6272 ( .B1(n8212), .B2(n8210), .A(n4414), .ZN(n8195) );
  NAND2_X1 U6273 ( .A1(n6929), .A2(n4744), .ZN(n4745) );
  OAI21_X1 U6274 ( .B1(n4748), .B2(n4503), .A(n7043), .ZN(n4747) );
  INV_X1 U6275 ( .A(n7045), .ZN(n4749) );
  NAND2_X1 U6276 ( .A1(n4753), .A2(n9901), .ZN(n4752) );
  INV_X1 U6277 ( .A(n5815), .ZN(n4754) );
  NAND2_X2 U6278 ( .A1(n5815), .A2(n5816), .ZN(n5870) );
  OAI21_X1 U6279 ( .B1(n5816), .B2(n9706), .A(n4757), .ZN(n4756) );
  NAND2_X1 U6280 ( .A1(n5816), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4757) );
  NAND2_X1 U6281 ( .A1(n4768), .A2(n4767), .ZN(n7324) );
  NAND2_X1 U6282 ( .A1(n4770), .A2(n4769), .ZN(n6143) );
  NAND3_X1 U6283 ( .A1(n4774), .A2(n5855), .A3(n4773), .ZN(n5898) );
  XNOR2_X1 U6284 ( .A(n8166), .B(n8165), .ZN(n4776) );
  OAI21_X1 U6285 ( .B1(n8447), .B2(n8378), .A(n4495), .ZN(n4778) );
  INV_X1 U6286 ( .A(n5808), .ZN(n5025) );
  NOR2_X2 U6287 ( .A1(n6198), .A2(n5807), .ZN(n5808) );
  NAND2_X1 U6288 ( .A1(n7192), .A2(n4790), .ZN(n4789) );
  AND2_X2 U6289 ( .A1(n4797), .A2(n4796), .ZN(n9268) );
  NOR2_X2 U6290 ( .A1(n9513), .A2(n4799), .ZN(n9287) );
  NAND2_X1 U6291 ( .A1(n9165), .A2(n9166), .ZN(n4801) );
  NAND2_X1 U6292 ( .A1(n4800), .A2(n4802), .ZN(n9119) );
  NAND2_X1 U6293 ( .A1(n9165), .A2(n4804), .ZN(n4800) );
  NAND2_X1 U6294 ( .A1(n7456), .A2(n4813), .ZN(n4811) );
  NAND3_X1 U6295 ( .A1(n4824), .A2(n4826), .A3(n4482), .ZN(n4822) );
  OR2_X1 U6296 ( .A1(n9353), .A2(n9345), .ZN(n4830) );
  NAND2_X1 U6297 ( .A1(n5456), .A2(n5054), .ZN(n5069) );
  INV_X1 U6298 ( .A(n6604), .ZN(n4833) );
  NAND2_X1 U6299 ( .A1(n9730), .A2(n6753), .ZN(n6397) );
  NAND2_X1 U6300 ( .A1(n9173), .A2(n4842), .ZN(n4839) );
  NAND2_X1 U6301 ( .A1(n6757), .A2(n4852), .ZN(n4849) );
  INV_X1 U6302 ( .A(n4857), .ZN(n9748) );
  NAND2_X1 U6303 ( .A1(n4858), .A2(n6462), .ZN(n4856) );
  NOR2_X1 U6304 ( .A1(n6764), .A2(n6398), .ZN(n4860) );
  NAND2_X1 U6305 ( .A1(n4862), .A2(n6399), .ZN(n4868) );
  NAND2_X1 U6306 ( .A1(n4862), .A2(n4861), .ZN(n4866) );
  INV_X1 U6307 ( .A(n9753), .ZN(n4862) );
  OAI21_X1 U6308 ( .B1(n9753), .B2(n4427), .A(n4863), .ZN(n4865) );
  INV_X1 U6309 ( .A(n6890), .ZN(n4864) );
  INV_X1 U6310 ( .A(n4867), .ZN(n6883) );
  INV_X1 U6311 ( .A(n4878), .ZN(n9262) );
  OR2_X1 U6312 ( .A1(n7338), .A2(n4879), .ZN(n4880) );
  NAND2_X1 U6313 ( .A1(n4880), .A2(n4881), .ZN(n7457) );
  XNOR2_X1 U6314 ( .A(n6411), .B(n9822), .ZN(n9820) );
  INV_X2 U6315 ( .A(n5311), .ZN(n4905) );
  AOI21_X1 U6316 ( .B1(n5192), .B2(n5191), .A(n4429), .ZN(n4912) );
  NAND2_X1 U6317 ( .A1(n6172), .A2(n4915), .ZN(n4914) );
  NAND3_X1 U6318 ( .A1(n8074), .A2(n8075), .A3(n4473), .ZN(n4919) );
  OR2_X1 U6319 ( .A1(n8082), .A2(n4924), .ZN(n4923) );
  NAND2_X1 U6320 ( .A1(n5581), .A2(n5580), .ZN(n5604) );
  AND2_X2 U6321 ( .A1(n4948), .A2(n4947), .ZN(n4949) );
  INV_X1 U6322 ( .A(n4954), .ZN(n6789) );
  NOR2_X1 U6323 ( .A1(n6827), .A2(n6826), .ZN(n4951) );
  INV_X1 U6324 ( .A(n5208), .ZN(n4953) );
  NAND2_X1 U6325 ( .A1(n5676), .A2(n8639), .ZN(n4956) );
  OR2_X1 U6326 ( .A1(n5676), .A2(n4957), .ZN(n8638) );
  NAND2_X1 U6327 ( .A1(n8617), .A2(n4474), .ZN(n4960) );
  OR2_X1 U6328 ( .A1(n4962), .A2(n5646), .ZN(n8685) );
  NOR2_X1 U6329 ( .A1(n5647), .A2(n8686), .ZN(n4961) );
  NAND2_X1 U6330 ( .A1(n4962), .A2(n5646), .ZN(n8684) );
  NAND2_X1 U6331 ( .A1(n7624), .A2(n4970), .ZN(n4964) );
  INV_X1 U6332 ( .A(n7624), .ZN(n4963) );
  NAND3_X1 U6333 ( .A1(n4967), .A2(n4969), .A3(n4964), .ZN(n8554) );
  NAND2_X1 U6334 ( .A1(n8656), .A2(n4973), .ZN(n4972) );
  NAND2_X1 U6335 ( .A1(n4972), .A2(n4975), .ZN(n5594) );
  NAND2_X1 U6336 ( .A1(n7109), .A2(n4983), .ZN(n4981) );
  NAND2_X1 U6337 ( .A1(n7843), .A2(n4992), .ZN(n4991) );
  AOI21_X1 U6338 ( .B1(n5001), .B2(n7699), .A(n7852), .ZN(n7701) );
  INV_X1 U6339 ( .A(n5003), .ZN(n7773) );
  NAND2_X1 U6340 ( .A1(n7742), .A2(n5013), .ZN(n5010) );
  AND2_X1 U6341 ( .A1(n7659), .A2(n8251), .ZN(n5015) );
  OAI21_X2 U6342 ( .B1(n7750), .B2(n5021), .A(n5020), .ZN(n5019) );
  NAND2_X2 U6343 ( .A1(n7637), .A2(n7636), .ZN(n7750) );
  NAND2_X2 U6344 ( .A1(n4400), .A2(n7476), .ZN(n7637) );
  NOR3_X1 U6345 ( .A1(n5966), .A2(n5025), .A3(P2_IR_REG_9__SCAN_IN), .ZN(n6252) );
  OR3_X1 U6346 ( .A1(n5966), .A2(n5025), .A3(n5023), .ZN(n6254) );
  NAND2_X1 U6347 ( .A1(n7167), .A2(n7166), .ZN(n7192) );
  INV_X1 U6348 ( .A(n7086), .ZN(n9595) );
  INV_X1 U6349 ( .A(n5456), .ZN(n5481) );
  NAND2_X1 U6350 ( .A1(n5456), .A2(n5077), .ZN(n5483) );
  OR2_X1 U6351 ( .A1(n8305), .A2(n8021), .ZN(n6224) );
  OR2_X1 U6352 ( .A1(n7688), .A2(n7687), .ZN(n7692) );
  NAND2_X1 U6353 ( .A1(n6234), .A2(n7902), .ZN(n6235) );
  CLKBUF_X1 U6354 ( .A(n5361), .Z(n5382) );
  OAI21_X1 U6355 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8974) );
  NAND2_X1 U6356 ( .A1(n8972), .A2(n5768), .ZN(n5738) );
  NAND2_X1 U6357 ( .A1(n5446), .A2(n5445), .ZN(n5449) );
  CLKBUF_X1 U6358 ( .A(n7624), .Z(n7625) );
  NAND2_X1 U6359 ( .A1(n6838), .A2(n6841), .ZN(n6840) );
  CLKBUF_X1 U6360 ( .A(n5739), .Z(n8918) );
  INV_X1 U6361 ( .A(n5739), .ZN(n8835) );
  AND2_X4 U6362 ( .A1(n5063), .A2(n7620), .ZN(n5461) );
  NAND2_X1 U6363 ( .A1(n5171), .A2(n5170), .ZN(n8710) );
  INV_X1 U6364 ( .A(n6207), .ZN(n6208) );
  NAND2_X1 U6365 ( .A1(n5838), .A2(n5837), .ZN(n6240) );
  NAND2_X1 U6366 ( .A1(n7913), .A2(n6729), .ZN(n6724) );
  NAND2_X1 U6367 ( .A1(n8092), .A2(n7913), .ZN(n9933) );
  XNOR2_X1 U6368 ( .A(n7469), .B(n7470), .ZN(n7362) );
  NOR2_X1 U6369 ( .A1(n7559), .A2(n8861), .ZN(n9513) );
  NAND2_X2 U6370 ( .A1(n7337), .A2(n7336), .ZN(n7456) );
  OR2_X1 U6371 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7845), .ZN(n5026) );
  OR2_X1 U6372 ( .A1(n9839), .A2(n9452), .ZN(n5027) );
  AND2_X1 U6373 ( .A1(n6431), .A2(n6430), .ZN(n9941) );
  INV_X1 U6374 ( .A(n8513), .ZN(n8534) );
  NAND2_X2 U6375 ( .A1(n8355), .A2(n6931), .ZN(n8373) );
  INV_X1 U6376 ( .A(n9951), .ZN(n6296) );
  INV_X1 U6377 ( .A(n8414), .ZN(n8432) );
  OR2_X1 U6378 ( .A1(n9939), .A2(n10093), .ZN(n5028) );
  AND2_X1 U6379 ( .A1(n7707), .A2(n7861), .ZN(n5029) );
  AND2_X1 U6380 ( .A1(n6260), .A2(n5810), .ZN(n5031) );
  INV_X1 U6381 ( .A(n8347), .ZN(n6212) );
  AND2_X1 U6382 ( .A1(n6432), .A2(n5028), .ZN(n5032) );
  AND2_X1 U6383 ( .A1(n6295), .A2(n6294), .ZN(n5033) );
  NOR2_X1 U6384 ( .A1(n5887), .A2(n5886), .ZN(n5034) );
  NOR2_X1 U6385 ( .A1(n5397), .A2(n7623), .ZN(n5035) );
  INV_X1 U6386 ( .A(n6237), .ZN(n8090) );
  INV_X1 U6387 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5799) );
  INV_X1 U6388 ( .A(n7959), .ZN(n6219) );
  INV_X1 U6389 ( .A(n7955), .ZN(n6220) );
  INV_X1 U6390 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5779) );
  AND4_X1 U6391 ( .A1(n7609), .A2(n7608), .A3(n7607), .A4(n7606), .ZN(n9116)
         );
  INV_X1 U6392 ( .A(n8370), .ZN(n8349) );
  OR2_X1 U6393 ( .A1(n9388), .A2(n9387), .ZN(n9672) );
  INV_X1 U6394 ( .A(n5737), .ZN(n8912) );
  AND2_X1 U6395 ( .A1(n7395), .A2(n5304), .ZN(n5036) );
  OR2_X1 U6396 ( .A1(n8474), .A2(n8215), .ZN(n5037) );
  AND2_X1 U6397 ( .A1(n9250), .A2(n9232), .ZN(n5038) );
  INV_X1 U6398 ( .A(n7393), .ZN(n5300) );
  INV_X1 U6399 ( .A(n8739), .ZN(n5770) );
  NOR3_X1 U6400 ( .A1(n8065), .A2(n8064), .A3(n8173), .ZN(n8070) );
  AOI21_X1 U6401 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8080) );
  INV_X1 U6402 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U6403 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5802) );
  NOR2_X1 U6404 ( .A1(n5039), .A2(n5564), .ZN(n5565) );
  NAND2_X1 U6405 ( .A1(n7393), .A2(n5303), .ZN(n5304) );
  NAND2_X1 U6406 ( .A1(n5165), .A2(n8919), .ZN(n5166) );
  NAND2_X1 U6407 ( .A1(n5047), .A2(n5046), .ZN(n5048) );
  NAND2_X1 U6408 ( .A1(n6370), .A2(n6890), .ZN(n6371) );
  INV_X1 U6409 ( .A(n6107), .ZN(n5788) );
  INV_X1 U6410 ( .A(n8088), .ZN(n6729) );
  INV_X1 U6411 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6012) );
  OR2_X1 U6412 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NAND2_X1 U6413 ( .A1(n5616), .A2(n8991), .ZN(n5148) );
  INV_X1 U6414 ( .A(n8666), .ZN(n5675) );
  NAND2_X1 U6415 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  INV_X1 U6416 ( .A(n9116), .ZN(n9117) );
  NOR2_X1 U6417 ( .A1(n5285), .A2(n6594), .ZN(n5317) );
  INV_X1 U6418 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5053) );
  INV_X1 U6419 ( .A(SI_19_), .ZN(n5507) );
  INV_X1 U6420 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5040) );
  XNOR2_X1 U6421 ( .A(n7939), .B(n7118), .ZN(n6904) );
  INV_X1 U6422 ( .A(n6146), .ZN(n5792) );
  AND2_X1 U6423 ( .A1(n6718), .A2(n6743), .ZN(n7858) );
  NAND2_X1 U6424 ( .A1(n5794), .A2(n5793), .ZN(n6162) );
  NAND2_X1 U6425 ( .A1(n5781), .A2(n7524), .ZN(n6016) );
  INV_X1 U6426 ( .A(n8214), .ZN(n8187) );
  OR2_X1 U6427 ( .A1(n8108), .A2(n9919), .ZN(n7978) );
  INV_X1 U6428 ( .A(n6717), .ZN(n6719) );
  AND2_X1 U6429 ( .A1(n6427), .A2(n6920), .ZN(n6711) );
  INV_X1 U6430 ( .A(n5585), .ZN(n5586) );
  INV_X1 U6431 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10195) );
  OR2_X1 U6432 ( .A1(n6774), .A2(n6773), .ZN(n6873) );
  NAND2_X1 U6433 ( .A1(n9371), .A2(n9363), .ZN(n9107) );
  OR2_X1 U6434 ( .A1(n5750), .A2(n5738), .ZN(n7003) );
  AND2_X1 U6435 ( .A1(n5053), .A2(n5071), .ZN(n5054) );
  INV_X1 U6436 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10227) );
  INV_X1 U6437 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6270) );
  INV_X1 U6438 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5775) );
  INV_X1 U6439 ( .A(n7475), .ZN(n7476) );
  OR2_X1 U6440 ( .A1(n6162), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6175) );
  INV_X1 U6441 ( .A(n6109), .ZN(n6191) );
  INV_X1 U6442 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10237) );
  AND2_X1 U6443 ( .A1(n6354), .A2(n6353), .ZN(n9841) );
  OR2_X1 U6444 ( .A1(P2_U3150), .A2(n6359), .ZN(n9839) );
  INV_X1 U6445 ( .A(n7907), .ZN(n7976) );
  AND2_X1 U6446 ( .A1(n8090), .A2(n8088), .ZN(n6919) );
  INV_X1 U6447 ( .A(n8330), .ZN(n7926) );
  INV_X1 U6448 ( .A(n8054), .ZN(n6230) );
  AND2_X1 U6449 ( .A1(n6717), .A2(n8083), .ZN(n8370) );
  INV_X1 U6450 ( .A(n7730), .ZN(n9929) );
  AND2_X1 U6451 ( .A1(n6425), .A2(n6211), .ZN(n8347) );
  NOR2_X1 U6452 ( .A1(n5418), .A2(n5417), .ZN(n5438) );
  INV_X1 U6453 ( .A(n9328), .ZN(n9115) );
  OR2_X1 U6454 ( .A1(n5366), .A2(n5365), .ZN(n5386) );
  OR2_X1 U6455 ( .A1(n5689), .A2(n5688), .ZN(n5711) );
  NAND2_X1 U6456 ( .A1(n5244), .A2(n5243), .ZN(n6937) );
  AND2_X1 U6457 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5229) );
  OR2_X1 U6458 ( .A1(n5386), .A2(n10195), .ZN(n5418) );
  NAND2_X1 U6459 ( .A1(n5762), .A2(n9535), .ZN(n8704) );
  OR2_X1 U6460 ( .A1(n5711), .A2(n5763), .ZN(n7604) );
  NAND2_X1 U6461 ( .A1(n5449), .A2(n5450), .ZN(n8730) );
  INV_X1 U6462 ( .A(n5060), .ZN(n5061) );
  INV_X1 U6463 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6594) );
  INV_X1 U6464 ( .A(n9299), .ZN(n9275) );
  INV_X1 U6465 ( .A(n8895), .ZN(n9296) );
  AND2_X1 U6466 ( .A1(n5704), .A2(n5685), .ZN(n5702) );
  INV_X1 U6467 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5077) );
  AND3_X1 U6468 ( .A1(n6274), .A2(n6273), .A3(n6272), .ZN(n6297) );
  OR2_X1 U6469 ( .A1(n5947), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5960) );
  OR2_X1 U6470 ( .A1(n6713), .A2(n6712), .ZN(n7875) );
  AND2_X1 U6471 ( .A1(n7896), .A2(n6196), .ZN(n8101) );
  AND4_X1 U6472 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n8332)
         );
  INV_X1 U6473 ( .A(n9839), .ZN(n9856) );
  XNOR2_X1 U6474 ( .A(n7893), .B(n8073), .ZN(n8155) );
  INV_X1 U6475 ( .A(n8288), .ZN(n9889) );
  AND2_X1 U6476 ( .A1(n6926), .A2(n6290), .ZN(n6291) );
  INV_X1 U6477 ( .A(n7905), .ZN(n8297) );
  INV_X1 U6478 ( .A(n9933), .ZN(n9918) );
  AND2_X1 U6479 ( .A1(n6288), .A2(n6287), .ZN(n6494) );
  INV_X1 U6480 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6209) );
  INV_X1 U6481 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5913) );
  INV_X1 U6482 ( .A(n9579), .ZN(n7060) );
  AND2_X1 U6483 ( .A1(n5747), .A2(n5746), .ZN(n5749) );
  AND4_X1 U6484 ( .A1(n5665), .A2(n5664), .A3(n5663), .A4(n5662), .ZN(n9191)
         );
  AND4_X1 U6485 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n8661)
         );
  INV_X1 U6486 ( .A(n7300), .ZN(n9075) );
  INV_X1 U6487 ( .A(n6640), .ZN(n6659) );
  INV_X1 U6488 ( .A(n7221), .ZN(n7227) );
  AND2_X1 U6489 ( .A1(n6672), .A2(n8992), .ZN(n9084) );
  INV_X1 U6490 ( .A(n8972), .ZN(n9493) );
  INV_X1 U6491 ( .A(n9114), .ZN(n9159) );
  NAND3_X1 U6492 ( .A1(n6435), .A2(P1_STATE_REG_SCAN_IN), .A3(n6433), .ZN(
        n9307) );
  OAI21_X1 U6493 ( .B1(n6950), .B2(P1_D_REG_0__SCAN_IN), .A(n9403), .ZN(n9313)
         );
  INV_X1 U6494 ( .A(n9652), .ZN(n9654) );
  NAND2_X1 U6495 ( .A1(n9318), .A2(n9317), .ZN(n9652) );
  AND2_X1 U6496 ( .A1(n8826), .A2(n5768), .ZN(n9668) );
  NAND2_X1 U6497 ( .A1(n5724), .A2(n5725), .ZN(n6950) );
  AND2_X1 U6498 ( .A1(n5434), .A2(n5414), .ZN(n6780) );
  INV_X1 U6499 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10185) );
  INV_X1 U6500 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10145) );
  INV_X1 U6501 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10238) );
  AND2_X1 U6502 ( .A1(n7505), .A2(n6297), .ZN(n6359) );
  AND2_X1 U6503 ( .A1(n6745), .A2(n6744), .ZN(n7852) );
  INV_X1 U6504 ( .A(n7850), .ZN(n7878) );
  NAND2_X1 U6505 ( .A1(n5821), .A2(n5820), .ZN(n8174) );
  INV_X1 U6506 ( .A(n8237), .ZN(n8263) );
  INV_X1 U6507 ( .A(n9868), .ZN(n9847) );
  INV_X1 U6508 ( .A(n9863), .ZN(n9849) );
  NAND2_X1 U6509 ( .A1(n6527), .A2(n8548), .ZN(n9872) );
  INV_X1 U6510 ( .A(n8373), .ZN(n8340) );
  NAND2_X1 U6511 ( .A1(n9951), .A2(n9918), .ZN(n8414) );
  NAND2_X1 U6512 ( .A1(n9938), .A2(n9951), .ZN(n8435) );
  AND2_X2 U6513 ( .A1(n6292), .A2(n6291), .ZN(n9951) );
  INV_X1 U6514 ( .A(n7822), .ZN(n8481) );
  OR2_X1 U6515 ( .A1(n9941), .A2(n9933), .ZN(n8513) );
  NAND2_X1 U6516 ( .A1(n9939), .A2(n9938), .ZN(n8537) );
  INV_X2 U6517 ( .A(n9941), .ZN(n9939) );
  INV_X1 U6518 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6664) );
  XNOR2_X1 U6519 ( .A(n5744), .B(n5743), .ZN(n6435) );
  INV_X1 U6520 ( .A(n9384), .ZN(n9283) );
  INV_X1 U6521 ( .A(n9346), .ZN(n9193) );
  INV_X1 U6522 ( .A(n9377), .ZN(n9260) );
  AND2_X1 U6523 ( .A1(n5769), .A2(n9499), .ZN(n8739) );
  INV_X1 U6524 ( .A(n8722), .ZN(n8745) );
  INV_X1 U6525 ( .A(n9191), .ZN(n9345) );
  INV_X1 U6526 ( .A(n8661), .ZN(n9298) );
  INV_X1 U6527 ( .A(n7254), .ZN(n9627) );
  INV_X1 U6528 ( .A(n9084), .ZN(n7429) );
  OR2_X1 U6529 ( .A1(n6438), .A2(n6440), .ZN(n9026) );
  OR2_X1 U6530 ( .A1(n9309), .A2(n9307), .ZN(n9499) );
  AND2_X1 U6531 ( .A1(n6956), .A2(n9499), .ZN(n9301) );
  INV_X1 U6532 ( .A(n9494), .ZN(n9553) );
  OR2_X1 U6533 ( .A1(n9553), .A2(n7018), .ZN(n9286) );
  INV_X1 U6534 ( .A(n9697), .ZN(n9700) );
  INV_X1 U6535 ( .A(n9555), .ZN(n9554) );
  NAND2_X1 U6536 ( .A1(n6951), .A2(n6950), .ZN(n9555) );
  OR2_X1 U6537 ( .A1(n6435), .A2(P1_U3086), .ZN(n8970) );
  INV_X1 U6538 ( .A(n7418), .ZN(n7315) );
  INV_X1 U6539 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6530) );
  OAI21_X1 U6540 ( .B1(n6424), .B2(n6296), .A(n5033), .ZN(P2_U3488) );
  AND2_X2 U6541 ( .A1(n6434), .A2(n6435), .ZN(P1_U3973) );
  INV_X2 U6542 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND4_X1 U6543 ( .A1(n5043), .A2(n5042), .A3(n5041), .A4(n5275), .ZN(n5044)
         );
  NOR2_X2 U6544 ( .A1(n5089), .A2(n5044), .ZN(n5359) );
  NOR2_X1 U6545 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5051) );
  NOR2_X1 U6546 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5050) );
  NOR2_X1 U6547 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5049) );
  XNOR2_X2 U6548 ( .A(n5056), .B(n5055), .ZN(n7697) );
  NAND2_X1 U6549 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5058) );
  NAND2_X1 U6550 ( .A1(n5085), .A2(n5058), .ZN(n5059) );
  INV_X4 U6551 ( .A(n8820), .ZN(n6497) );
  NAND2_X1 U6552 ( .A1(n6497), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5067) );
  AND2_X2 U6553 ( .A1(n7697), .A2(n7620), .ZN(n5460) );
  NAND2_X1 U6554 ( .A1(n5460), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5066) );
  INV_X1 U6555 ( .A(n7697), .ZN(n5063) );
  AND2_X2 U6556 ( .A1(n5063), .A2(n5061), .ZN(n5210) );
  NAND2_X1 U6557 ( .A1(n5229), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5249) );
  NOR2_X1 U6558 ( .A1(n5249), .A2(n5248), .ZN(n5268) );
  NAND2_X1 U6559 ( .A1(n5268), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5283) );
  AND2_X1 U6560 ( .A1(n5285), .A2(n6594), .ZN(n5062) );
  NOR2_X1 U6561 ( .A1(n5317), .A2(n5062), .ZN(n7401) );
  NAND2_X1 U6562 ( .A1(n5631), .A2(n7401), .ZN(n5065) );
  NAND2_X1 U6563 ( .A1(n5461), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6564 ( .A1(n5069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5068) );
  MUX2_X1 U6565 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5068), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5070) );
  NAND2_X1 U6566 ( .A1(n4437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5072) );
  MUX2_X1 U6567 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5072), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5073) );
  NAND2_X1 U6568 ( .A1(n4457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5074) );
  MUX2_X1 U6569 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5074), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5075) );
  NOR2_X2 U6570 ( .A1(n5483), .A2(n4432), .ZN(n5079) );
  NAND2_X1 U6571 ( .A1(n5079), .A2(n5081), .ZN(n5128) );
  INV_X1 U6573 ( .A(n5079), .ZN(n5080) );
  XNOR2_X2 U6574 ( .A(n5082), .B(n5081), .ZN(n5768) );
  NAND2_X1 U6575 ( .A1(n5739), .A2(n5768), .ZN(n6999) );
  INV_X1 U6576 ( .A(n6999), .ZN(n5083) );
  AND2_X4 U6577 ( .A1(n6433), .A2(n5083), .ZN(n5616) );
  XNOR2_X2 U6578 ( .A(n5085), .B(n5084), .ZN(n5160) );
  INV_X1 U6579 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5087) );
  INV_X1 U6580 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5234) );
  NAND3_X1 U6581 ( .A1(n10146), .A2(n5234), .A3(n5275), .ZN(n5090) );
  OR2_X1 U6582 ( .A1(n5255), .A2(n5090), .ZN(n5290) );
  NOR2_X1 U6583 ( .A1(n5290), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5313) );
  NOR2_X1 U6584 ( .A1(n5313), .A2(n9406), .ZN(n5091) );
  INV_X1 U6585 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6586 ( .A(n5091), .B(n5312), .ZN(n6580) );
  INV_X1 U6587 ( .A(n6580), .ZN(n6595) );
  CLKBUF_X3 U6588 ( .A(n5104), .Z(n5876) );
  AND2_X1 U6589 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6590 ( .A1(n7885), .A2(n5094), .ZN(n5878) );
  AND2_X1 U6591 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6592 ( .A1(n5104), .A2(n5095), .ZN(n5141) );
  NAND2_X1 U6593 ( .A1(n5878), .A2(n5141), .ZN(n5155) );
  OAI21_X1 U6594 ( .B1(n5156), .B2(SI_1_), .A(n5155), .ZN(n5097) );
  NAND2_X1 U6595 ( .A1(n5156), .A2(SI_1_), .ZN(n5096) );
  NAND2_X1 U6596 ( .A1(n5097), .A2(n5096), .ZN(n5173) );
  INV_X1 U6597 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6472) );
  INV_X1 U6598 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6455) );
  MUX2_X1 U6599 ( .A(n6472), .B(n6455), .S(n7885), .Z(n5098) );
  XNOR2_X1 U6600 ( .A(n5098), .B(SI_2_), .ZN(n5172) );
  NAND2_X1 U6601 ( .A1(n5173), .A2(n5172), .ZN(n5101) );
  INV_X1 U6602 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6603 ( .A1(n5099), .A2(SI_2_), .ZN(n5100) );
  INV_X1 U6604 ( .A(SI_3_), .ZN(n5102) );
  XNOR2_X1 U6605 ( .A(n5103), .B(n5102), .ZN(n5191) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6461) );
  INV_X1 U6607 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6474) );
  MUX2_X1 U6608 ( .A(n6461), .B(n6474), .S(n5104), .Z(n5105) );
  XNOR2_X1 U6609 ( .A(n5105), .B(SI_4_), .ZN(n5218) );
  INV_X1 U6610 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6611 ( .A1(n5106), .A2(SI_4_), .ZN(n5107) );
  MUX2_X1 U6612 ( .A(n6463), .B(n6476), .S(n5876), .Z(n5108) );
  XNOR2_X1 U6613 ( .A(n5108), .B(SI_5_), .ZN(n5236) );
  INV_X1 U6614 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6615 ( .A1(n5109), .A2(SI_5_), .ZN(n5110) );
  NAND2_X1 U6616 ( .A1(n5111), .A2(n5110), .ZN(n5259) );
  MUX2_X1 U6617 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5876), .Z(n5112) );
  INV_X1 U6618 ( .A(SI_6_), .ZN(n10160) );
  XNOR2_X1 U6619 ( .A(n5112), .B(n10160), .ZN(n5258) );
  NAND2_X1 U6620 ( .A1(n5112), .A2(SI_6_), .ZN(n5113) );
  MUX2_X1 U6621 ( .A(n10052), .B(n6477), .S(n5876), .Z(n5114) );
  XNOR2_X1 U6622 ( .A(n5114), .B(SI_7_), .ZN(n5277) );
  INV_X1 U6623 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6624 ( .A1(n5115), .A2(SI_7_), .ZN(n5116) );
  MUX2_X1 U6625 ( .A(n6479), .B(n6481), .S(n5876), .Z(n5118) );
  INV_X1 U6626 ( .A(SI_8_), .ZN(n5117) );
  NAND2_X1 U6627 ( .A1(n5118), .A2(n5117), .ZN(n5121) );
  INV_X1 U6628 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6629 ( .A1(n5119), .A2(SI_8_), .ZN(n5120) );
  INV_X1 U6630 ( .A(n5292), .ZN(n5122) );
  OAI21_X2 U6631 ( .B1(n5293), .B2(n5122), .A(n5121), .ZN(n5308) );
  MUX2_X1 U6632 ( .A(n6482), .B(n6484), .S(n5876), .Z(n5124) );
  INV_X1 U6633 ( .A(SI_9_), .ZN(n5123) );
  NAND2_X1 U6634 ( .A1(n5124), .A2(n5123), .ZN(n5309) );
  INV_X1 U6635 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6636 ( .A1(n5125), .A2(SI_9_), .ZN(n5126) );
  NAND2_X1 U6637 ( .A1(n5309), .A2(n5126), .ZN(n5306) );
  XNOR2_X1 U6638 ( .A(n5308), .B(n5306), .ZN(n6483) );
  OR2_X1 U6639 ( .A1(n8823), .A2(n6484), .ZN(n5127) );
  NAND2_X1 U6640 ( .A1(n5739), .A2(n6957), .ZN(n8969) );
  NAND2_X1 U6641 ( .A1(n5483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U6642 ( .A1(n5544), .A2(n5543), .ZN(n5546) );
  XNOR2_X2 U6643 ( .A(n5130), .B(n5129), .ZN(n8972) );
  NAND2_X1 U6644 ( .A1(n5736), .A2(n8972), .ZN(n7000) );
  AND2_X1 U6645 ( .A1(n8835), .A2(n6433), .ZN(n5131) );
  NAND2_X1 U6646 ( .A1(n7000), .A2(n5131), .ZN(n5132) );
  NAND2_X1 U6647 ( .A1(n6999), .A2(n5738), .ZN(n5134) );
  NAND2_X1 U6648 ( .A1(n5134), .A2(n7000), .ZN(n5135) );
  NAND2_X1 U6649 ( .A1(n9624), .A2(n8593), .ZN(n5136) );
  OAI21_X1 U6650 ( .B1(n7447), .B2(n5493), .A(n5136), .ZN(n5137) );
  INV_X2 U6651 ( .A(n5719), .ZN(n8591) );
  XNOR2_X1 U6652 ( .A(n5137), .B(n8591), .ZN(n5302) );
  OR2_X1 U6653 ( .A1(n7447), .A2(n8588), .ZN(n5139) );
  NAND2_X1 U6654 ( .A1(n9624), .A2(n5616), .ZN(n5138) );
  NAND2_X1 U6655 ( .A1(n5139), .A2(n5138), .ZN(n5305) );
  INV_X1 U6656 ( .A(SI_0_), .ZN(n5875) );
  INV_X1 U6657 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5140) );
  OAI21_X1 U6658 ( .B1(n7885), .B2(n5875), .A(n5140), .ZN(n5142) );
  AND2_X1 U6659 ( .A1(n5142), .A2(n5141), .ZN(n9413) );
  NAND2_X1 U6660 ( .A1(n5461), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6661 ( .A1(n5210), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6662 ( .A1(n5460), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5144) );
  INV_X2 U6663 ( .A(n8820), .ZN(n8598) );
  NAND2_X1 U6664 ( .A1(n8598), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6665 ( .A1(n5754), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5147) );
  AOI21_X1 U6666 ( .B1(n5165), .B2(n9560), .A(n5149), .ZN(n6693) );
  AOI222_X1 U6667 ( .A1(n8991), .A2(n5639), .B1(n9560), .B2(n4402), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(n5754), .ZN(n6694) );
  NAND2_X1 U6668 ( .A1(n7000), .A2(n8835), .ZN(n5150) );
  OAI22_X1 U6669 ( .A1(n6693), .A2(n4403), .B1(n9560), .B2(n4413), .ZN(n6815)
         );
  NAND2_X1 U6670 ( .A1(n5460), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6671 ( .A1(n5210), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6672 ( .A1(n8598), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6673 ( .A1(n9569), .A2(n4402), .ZN(n5167) );
  INV_X1 U6674 ( .A(n5160), .ZN(n6449) );
  XNOR2_X1 U6675 ( .A(n5155), .B(SI_1_), .ZN(n5157) );
  XNOR2_X1 U6676 ( .A(n5157), .B(n5156), .ZN(n6457) );
  MUX2_X1 U6677 ( .A(n6457), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7885), .Z(n5161)
         );
  NAND2_X1 U6678 ( .A1(n6449), .A2(n5161), .ZN(n5164) );
  NAND2_X1 U6679 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5158) );
  XNOR2_X1 U6680 ( .A(n5158), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6549) );
  NAND3_X1 U6681 ( .A1(n5160), .A2(n6549), .A3(n8992), .ZN(n5163) );
  INV_X1 U6682 ( .A(n8992), .ZN(n9089) );
  NAND2_X1 U6683 ( .A1(n9089), .A2(n5161), .ZN(n5162) );
  AND3_X2 U6684 ( .A1(n5164), .A2(n5163), .A3(n5162), .ZN(n9565) );
  XNOR2_X1 U6685 ( .A(n5168), .B(n8591), .ZN(n5171) );
  NOR2_X1 U6686 ( .A1(n9565), .A2(n5593), .ZN(n5169) );
  AOI21_X1 U6687 ( .B1(n9569), .B2(n5639), .A(n5169), .ZN(n5170) );
  OAI21_X1 U6688 ( .B1(n5171), .B2(n5170), .A(n8710), .ZN(n6813) );
  OR2_X2 U6689 ( .A1(n6815), .A2(n6813), .ZN(n8711) );
  XNOR2_X1 U6690 ( .A(n5173), .B(n5172), .ZN(n6471) );
  OR2_X1 U6691 ( .A1(n5174), .A2(n9406), .ZN(n5194) );
  INV_X1 U6692 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5193) );
  XNOR2_X1 U6693 ( .A(n5194), .B(n5193), .ZN(n6547) );
  OR2_X1 U6694 ( .A1(n6437), .A2(n6547), .ZN(n5175) );
  NAND2_X1 U6695 ( .A1(n5460), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6696 ( .A1(n5210), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6697 ( .A1(n5461), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6698 ( .A1(n6497), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6699 ( .A1(n8990), .A2(n5616), .ZN(n5180) );
  OAI21_X1 U6700 ( .B1(n7026), .B2(n5666), .A(n5180), .ZN(n5181) );
  XNOR2_X1 U6701 ( .A(n5181), .B(n8591), .ZN(n5184) );
  OR2_X1 U6702 ( .A1(n7026), .A2(n5493), .ZN(n5183) );
  NAND2_X1 U6703 ( .A1(n8990), .A2(n5639), .ZN(n5182) );
  AND2_X1 U6704 ( .A1(n5183), .A2(n5182), .ZN(n5185) );
  NAND2_X1 U6705 ( .A1(n5184), .A2(n5185), .ZN(n5189) );
  INV_X1 U6706 ( .A(n5184), .ZN(n5187) );
  INV_X1 U6707 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6708 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6709 ( .A1(n5189), .A2(n5188), .ZN(n8709) );
  AOI21_X1 U6710 ( .B1(n8711), .B2(n8710), .A(n8709), .ZN(n8713) );
  INV_X1 U6711 ( .A(n5189), .ZN(n5190) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6470) );
  XNOR2_X1 U6713 ( .A(n5192), .B(n5191), .ZN(n6469) );
  OR2_X1 U6714 ( .A1(n5311), .A2(n6469), .ZN(n5198) );
  NAND2_X1 U6715 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  NAND2_X1 U6716 ( .A1(n5195), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5196) );
  XNOR2_X1 U6717 ( .A(n5196), .B(n4947), .ZN(n9016) );
  OR2_X1 U6718 ( .A1(n6437), .A2(n9016), .ZN(n5197) );
  OR2_X1 U6719 ( .A1(n9579), .A2(n5493), .ZN(n5205) );
  NAND2_X1 U6720 ( .A1(n5460), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5203) );
  INV_X1 U6721 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U6722 ( .A1(n5210), .A2(n6791), .ZN(n5202) );
  NAND2_X1 U6723 ( .A1(n5661), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6724 ( .A1(n6497), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6725 ( .A1(n9586), .A2(n5639), .ZN(n5204) );
  NAND2_X1 U6726 ( .A1(n5205), .A2(n5204), .ZN(n5208) );
  AOI22_X1 U6727 ( .A1(n7060), .A2(n4405), .B1(n5616), .B2(n9586), .ZN(n5206)
         );
  XNOR2_X1 U6728 ( .A(n5206), .B(n4413), .ZN(n5207) );
  INV_X1 U6729 ( .A(n5207), .ZN(n5209) );
  NOR2_X1 U6730 ( .A1(n5209), .A2(n5208), .ZN(n6827) );
  NAND2_X1 U6731 ( .A1(n5460), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6732 ( .A1(n6497), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5214) );
  NOR2_X1 U6733 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5211) );
  NOR2_X1 U6734 ( .A1(n5229), .A2(n5211), .ZN(n7063) );
  NAND2_X1 U6735 ( .A1(n5631), .A2(n7063), .ZN(n5213) );
  NAND2_X1 U6736 ( .A1(n5661), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6737 ( .A1(n5216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U6738 ( .A(n5217), .B(n5040), .ZN(n9032) );
  OR2_X1 U6739 ( .A1(n8823), .A2(n6474), .ZN(n5221) );
  XNOR2_X1 U6740 ( .A(n5219), .B(n5218), .ZN(n6473) );
  OR2_X1 U6741 ( .A1(n5311), .A2(n6473), .ZN(n5220) );
  OAI211_X1 U6742 ( .C1(n6437), .C2(n9032), .A(n5221), .B(n5220), .ZN(n9585)
         );
  NAND2_X1 U6743 ( .A1(n9585), .A2(n4405), .ZN(n5222) );
  OAI21_X1 U6744 ( .B1(n7086), .B2(n5493), .A(n5222), .ZN(n5223) );
  XNOR2_X1 U6745 ( .A(n5223), .B(n4530), .ZN(n5227) );
  OR2_X1 U6746 ( .A1(n7086), .A2(n7589), .ZN(n5225) );
  NAND2_X1 U6747 ( .A1(n9585), .A2(n5616), .ZN(n5224) );
  NAND2_X1 U6748 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6749 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  NAND2_X1 U6750 ( .A1(n6830), .A2(n5228), .ZN(n5244) );
  INV_X1 U6751 ( .A(n5244), .ZN(n5241) );
  NAND2_X1 U6752 ( .A1(n6497), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6753 ( .A1(n5460), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5232) );
  OAI21_X1 U6754 ( .B1(n5229), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5249), .ZN(
        n7098) );
  INV_X1 U6755 ( .A(n7098), .ZN(n6943) );
  NAND2_X1 U6756 ( .A1(n5631), .A2(n6943), .ZN(n5231) );
  NAND2_X1 U6757 ( .A1(n5661), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5230) );
  INV_X1 U6758 ( .A(n9605), .ZN(n8989) );
  NAND2_X1 U6759 ( .A1(n5255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5235) );
  XNOR2_X1 U6760 ( .A(n5235), .B(n5234), .ZN(n9041) );
  OR2_X1 U6761 ( .A1(n8823), .A2(n6476), .ZN(n5239) );
  XNOR2_X1 U6762 ( .A(n5237), .B(n5236), .ZN(n6475) );
  OR2_X1 U6763 ( .A1(n5311), .A2(n6475), .ZN(n5238) );
  OAI211_X1 U6764 ( .C1(n6437), .C2(n9041), .A(n5239), .B(n5238), .ZN(n9594)
         );
  AOI22_X1 U6765 ( .A1(n8989), .A2(n5616), .B1(n9594), .B2(n8593), .ZN(n5240)
         );
  XNOR2_X1 U6766 ( .A(n5240), .B(n4530), .ZN(n5242) );
  NAND2_X1 U6767 ( .A1(n5241), .A2(n5242), .ZN(n6938) );
  INV_X1 U6768 ( .A(n5242), .ZN(n5243) );
  OR2_X1 U6769 ( .A1(n9605), .A2(n8588), .ZN(n5246) );
  NAND2_X1 U6770 ( .A1(n9594), .A2(n5616), .ZN(n5245) );
  AND2_X1 U6771 ( .A1(n5246), .A2(n5245), .ZN(n6939) );
  NAND2_X1 U6772 ( .A1(n6937), .A2(n6939), .ZN(n5247) );
  NAND2_X1 U6773 ( .A1(n6497), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6774 ( .A1(n5460), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5253) );
  AND2_X1 U6775 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  NOR2_X1 U6776 ( .A1(n5268), .A2(n5250), .ZN(n7154) );
  NAND2_X1 U6777 ( .A1(n5631), .A2(n7154), .ZN(n5252) );
  NAND2_X1 U6778 ( .A1(n5461), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5251) );
  OAI21_X1 U6779 ( .B1(n5255), .B2(P1_IR_REG_5__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6780 ( .A1(n5256), .A2(n10146), .ZN(n5274) );
  OR2_X1 U6781 ( .A1(n5256), .A2(n10146), .ZN(n5257) );
  NAND2_X1 U6782 ( .A1(n5274), .A2(n5257), .ZN(n9061) );
  XNOR2_X1 U6783 ( .A(n5259), .B(n5258), .ZN(n6467) );
  OR2_X1 U6784 ( .A1(n5311), .A2(n6467), .ZN(n5261) );
  INV_X1 U6785 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6466) );
  OR2_X1 U6786 ( .A1(n8823), .A2(n6466), .ZN(n5260) );
  OAI211_X1 U6787 ( .C1(n6437), .C2(n9061), .A(n5261), .B(n5260), .ZN(n7155)
         );
  NAND2_X1 U6788 ( .A1(n7155), .A2(n8593), .ZN(n5262) );
  OAI21_X1 U6789 ( .B1(n7162), .B2(n5493), .A(n5262), .ZN(n5263) );
  XNOR2_X1 U6790 ( .A(n5263), .B(n4413), .ZN(n5267) );
  OR2_X1 U6791 ( .A1(n7162), .A2(n8588), .ZN(n5265) );
  NAND2_X1 U6792 ( .A1(n7155), .A2(n5616), .ZN(n5264) );
  NAND2_X1 U6793 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6794 ( .A1(n5267), .A2(n5266), .ZN(n7035) );
  NOR2_X1 U6795 ( .A1(n5267), .A2(n5266), .ZN(n7034) );
  NAND2_X1 U6796 ( .A1(n5657), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6797 ( .A1(n6497), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5272) );
  OR2_X1 U6798 ( .A1(n5268), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5269) );
  AND2_X1 U6799 ( .A1(n5283), .A2(n5269), .ZN(n9542) );
  NAND2_X1 U6800 ( .A1(n5631), .A2(n9542), .ZN(n5271) );
  NAND2_X1 U6801 ( .A1(n5461), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6802 ( .A1(n5274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5276) );
  XNOR2_X1 U6803 ( .A(n5276), .B(n5275), .ZN(n9069) );
  XNOR2_X1 U6804 ( .A(n5278), .B(n5277), .ZN(n6478) );
  OR2_X1 U6805 ( .A1(n5311), .A2(n6478), .ZN(n5280) );
  OR2_X1 U6806 ( .A1(n8823), .A2(n6477), .ZN(n5279) );
  OAI211_X1 U6807 ( .C1(n6437), .C2(n9069), .A(n5280), .B(n5279), .ZN(n7165)
         );
  OAI22_X1 U6808 ( .A1(n7443), .A2(n8588), .B1(n9612), .B2(n5493), .ZN(n7105)
         );
  INV_X1 U6809 ( .A(n7443), .ZN(n8988) );
  AOI22_X1 U6810 ( .A1(n8988), .A2(n5616), .B1(n7165), .B2(n8593), .ZN(n5281)
         );
  XOR2_X1 U6811 ( .A(n4413), .B(n5281), .Z(n7107) );
  NAND2_X1 U6812 ( .A1(n6497), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6813 ( .A1(n5460), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6814 ( .A1(n5283), .A2(n5282), .ZN(n5284) );
  AND2_X1 U6815 ( .A1(n5285), .A2(n5284), .ZN(n7173) );
  NAND2_X1 U6816 ( .A1(n5631), .A2(n7173), .ZN(n5287) );
  NAND2_X1 U6817 ( .A1(n5461), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6818 ( .A1(n5290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U6819 ( .A(n5291), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6572) );
  INV_X1 U6820 ( .A(n6572), .ZN(n6582) );
  XNOR2_X1 U6821 ( .A(n5293), .B(n5292), .ZN(n6480) );
  OR2_X1 U6822 ( .A1(n8823), .A2(n6481), .ZN(n5294) );
  NAND2_X1 U6823 ( .A1(n7177), .A2(n8593), .ZN(n5295) );
  OAI21_X1 U6824 ( .B1(n7254), .B2(n5493), .A(n5295), .ZN(n5296) );
  XNOR2_X1 U6825 ( .A(n5296), .B(n4413), .ZN(n7393) );
  OR2_X1 U6826 ( .A1(n7254), .A2(n8588), .ZN(n5298) );
  NAND2_X1 U6827 ( .A1(n7177), .A2(n5616), .ZN(n5297) );
  NAND2_X1 U6828 ( .A1(n5298), .A2(n5297), .ZN(n5303) );
  INV_X1 U6829 ( .A(n5303), .ZN(n5299) );
  NAND2_X1 U6830 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  XNOR2_X1 U6831 ( .A(n5302), .B(n5305), .ZN(n7395) );
  INV_X1 U6832 ( .A(n5327), .ZN(n5325) );
  INV_X1 U6833 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6834 ( .A1(n5308), .A2(n5307), .ZN(n5310) );
  MUX2_X1 U6835 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5876), .Z(n5330) );
  XNOR2_X1 U6836 ( .A(n5330), .B(n10054), .ZN(n5329) );
  XNOR2_X1 U6837 ( .A(n5333), .B(n5329), .ZN(n6485) );
  NAND2_X1 U6838 ( .A1(n6485), .A2(n4905), .ZN(n5316) );
  NAND2_X1 U6839 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  NAND2_X1 U6840 ( .A1(n5314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U6841 ( .A(n5339), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6579) );
  AOI22_X1 U6842 ( .A1(n5548), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5547), .B2(
        n6579), .ZN(n5315) );
  NAND2_X1 U6843 ( .A1(n6497), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6844 ( .A1(n5657), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5321) );
  NOR2_X1 U6845 ( .A1(n5317), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5318) );
  OR2_X1 U6846 ( .A1(n5344), .A2(n5318), .ZN(n7195) );
  INV_X1 U6847 ( .A(n7195), .ZN(n7543) );
  NAND2_X1 U6848 ( .A1(n5631), .A2(n7543), .ZN(n5320) );
  NAND2_X1 U6849 ( .A1(n5661), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5319) );
  NAND4_X1 U6850 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n8986)
         );
  AOI22_X1 U6851 ( .A1(n7548), .A2(n8593), .B1(n5616), .B2(n8986), .ZN(n5323)
         );
  XNOR2_X1 U6852 ( .A(n5323), .B(n4530), .ZN(n5326) );
  INV_X1 U6853 ( .A(n5326), .ZN(n5324) );
  NAND2_X1 U6854 ( .A1(n5325), .A2(n5324), .ZN(n5328) );
  INV_X1 U6855 ( .A(n5616), .ZN(n5493) );
  OAI22_X1 U6856 ( .A1(n9636), .A2(n5493), .B1(n7404), .B2(n8588), .ZN(n7541)
         );
  OR2_X2 U6857 ( .A1(n7540), .A2(n7541), .ZN(n7538) );
  NAND2_X2 U6858 ( .A1(n7538), .A2(n8694), .ZN(n8624) );
  INV_X1 U6859 ( .A(n5329), .ZN(n5332) );
  NAND2_X1 U6860 ( .A1(n5330), .A2(SI_10_), .ZN(n5331) );
  MUX2_X1 U6861 ( .A(n6504), .B(n6530), .S(n5876), .Z(n5335) );
  NAND2_X1 U6862 ( .A1(n5335), .A2(n5334), .ZN(n5358) );
  INV_X1 U6863 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6864 ( .A1(n5336), .A2(SI_11_), .ZN(n5337) );
  NAND2_X1 U6865 ( .A1(n5358), .A2(n5337), .ZN(n5356) );
  XNOR2_X1 U6866 ( .A(n5357), .B(n5356), .ZN(n6502) );
  NAND2_X1 U6867 ( .A1(n6502), .A2(n4905), .ZN(n5343) );
  INV_X1 U6868 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6869 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  NAND2_X1 U6870 ( .A1(n5340), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U6871 ( .A(n5341), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U6872 ( .A1(n5548), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5547), .B2(
        n6578), .ZN(n5342) );
  NAND2_X1 U6873 ( .A1(n5343), .A2(n5342), .ZN(n8706) );
  NAND2_X1 U6874 ( .A1(n8706), .A2(n8593), .ZN(n5351) );
  NAND2_X1 U6875 ( .A1(n5657), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6876 ( .A1(n6497), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6877 ( .A1(n5344), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5366) );
  OR2_X1 U6878 ( .A1(n5344), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5345) );
  AND2_X1 U6879 ( .A1(n5366), .A2(n5345), .ZN(n8701) );
  NAND2_X1 U6880 ( .A1(n5631), .A2(n8701), .ZN(n5347) );
  NAND2_X1 U6881 ( .A1(n5661), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5346) );
  OR2_X1 U6882 ( .A1(n7546), .A2(n5493), .ZN(n5350) );
  NAND2_X1 U6883 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  XNOR2_X1 U6884 ( .A(n5352), .B(n8591), .ZN(n5354) );
  INV_X1 U6885 ( .A(n7546), .ZN(n8985) );
  AOI22_X1 U6886 ( .A1(n8706), .A2(n5616), .B1(n8985), .B2(n5639), .ZN(n5353)
         );
  NAND2_X1 U6887 ( .A1(n5354), .A2(n5353), .ZN(n8625) );
  OR2_X1 U6888 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  AND2_X1 U6889 ( .A1(n8625), .A2(n5355), .ZN(n8695) );
  MUX2_X1 U6890 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5876), .Z(n5381) );
  XNOR2_X1 U6891 ( .A(n5381), .B(n10241), .ZN(n5379) );
  XNOR2_X1 U6892 ( .A(n5380), .B(n5379), .ZN(n6505) );
  NAND2_X1 U6893 ( .A1(n6505), .A2(n4905), .ZN(n5364) );
  NOR2_X1 U6894 ( .A1(n5359), .A2(n9406), .ZN(n5360) );
  MUX2_X1 U6895 ( .A(n9406), .B(n5360), .S(P1_IR_REG_12__SCAN_IN), .Z(n5362)
         );
  OR2_X1 U6896 ( .A1(n5362), .A2(n5382), .ZN(n6640) );
  AOI22_X1 U6897 ( .A1(n5548), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5547), .B2(
        n6659), .ZN(n5363) );
  NAND2_X1 U6898 ( .A1(n7354), .A2(n8593), .ZN(n5373) );
  NAND2_X1 U6899 ( .A1(n5657), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6900 ( .A1(n5661), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6901 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  AND2_X1 U6902 ( .A1(n5386), .A2(n5367), .ZN(n8635) );
  NAND2_X1 U6903 ( .A1(n5631), .A2(n8635), .ZN(n5369) );
  NAND2_X1 U6904 ( .A1(n6497), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5368) );
  OR2_X1 U6905 ( .A1(n9657), .A2(n5493), .ZN(n5372) );
  NAND2_X1 U6906 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  XNOR2_X1 U6907 ( .A(n5374), .B(n8591), .ZN(n5377) );
  NOR2_X1 U6908 ( .A1(n9657), .A2(n8588), .ZN(n5375) );
  AOI21_X1 U6909 ( .B1(n7354), .B2(n5616), .A(n5375), .ZN(n5376) );
  NAND2_X1 U6910 ( .A1(n5377), .A2(n5376), .ZN(n5396) );
  OR2_X1 U6911 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  AND2_X1 U6912 ( .A1(n8695), .A2(n8626), .ZN(n7622) );
  MUX2_X1 U6913 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5876), .Z(n5405) );
  XNOR2_X1 U6914 ( .A(n5405), .B(SI_13_), .ZN(n5403) );
  XNOR2_X1 U6915 ( .A(n5404), .B(n5403), .ZN(n6522) );
  NAND2_X1 U6916 ( .A1(n6522), .A2(n4905), .ZN(n5385) );
  OR2_X1 U6917 ( .A1(n5382), .A2(n9406), .ZN(n5383) );
  XNOR2_X1 U6918 ( .A(n5383), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U6919 ( .A1(n5548), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5547), .B2(
        n6777), .ZN(n5384) );
  NAND2_X1 U6920 ( .A1(n7621), .A2(n8593), .ZN(n5393) );
  NAND2_X1 U6921 ( .A1(n6497), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6922 ( .A1(n5657), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6923 ( .A1(n5386), .A2(n10195), .ZN(n5387) );
  AND2_X1 U6924 ( .A1(n5418), .A2(n5387), .ZN(n7632) );
  NAND2_X1 U6925 ( .A1(n5631), .A2(n7632), .ZN(n5389) );
  NAND2_X1 U6926 ( .A1(n5661), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5388) );
  OR2_X1 U6927 ( .A1(n8633), .A2(n5493), .ZN(n5392) );
  NAND2_X1 U6928 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  XNOR2_X1 U6929 ( .A(n5394), .B(n4530), .ZN(n5401) );
  INV_X1 U6930 ( .A(n8633), .ZN(n8983) );
  AOI22_X1 U6931 ( .A1(n7621), .A2(n5616), .B1(n5639), .B2(n8983), .ZN(n5399)
         );
  XNOR2_X1 U6932 ( .A(n5401), .B(n5399), .ZN(n7627) );
  AND2_X1 U6933 ( .A1(n7622), .A2(n7627), .ZN(n5398) );
  INV_X1 U6934 ( .A(n7627), .ZN(n5397) );
  INV_X1 U6935 ( .A(n8626), .ZN(n5395) );
  OR2_X1 U6936 ( .A1(n5395), .A2(n8625), .ZN(n8628) );
  AND2_X1 U6937 ( .A1(n8628), .A2(n5396), .ZN(n7623) );
  AOI21_X2 U6938 ( .B1(n8624), .B2(n5398), .A(n5035), .ZN(n7624) );
  INV_X1 U6939 ( .A(n5399), .ZN(n5400) );
  NAND2_X1 U6940 ( .A1(n5405), .A2(SI_13_), .ZN(n5406) );
  NAND2_X1 U6941 ( .A1(n5407), .A2(n5406), .ZN(n5427) );
  MUX2_X1 U6942 ( .A(n6664), .B(n10206), .S(n4660), .Z(n5409) );
  NAND2_X1 U6943 ( .A1(n5409), .A2(n5408), .ZN(n5431) );
  INV_X1 U6944 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U6945 ( .A1(n5410), .A2(SI_14_), .ZN(n5411) );
  NAND2_X1 U6946 ( .A1(n5431), .A2(n5411), .ZN(n5428) );
  XNOR2_X1 U6947 ( .A(n5427), .B(n5428), .ZN(n6661) );
  NAND2_X1 U6948 ( .A1(n6661), .A2(n4905), .ZN(n5416) );
  NAND2_X1 U6949 ( .A1(n5412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6950 ( .A1(n5413), .A2(n5047), .ZN(n5434) );
  OR2_X1 U6951 ( .A1(n5413), .A2(n5047), .ZN(n5414) );
  AOI22_X1 U6952 ( .A1(n5548), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5547), .B2(
        n6780), .ZN(n5415) );
  NAND2_X1 U6953 ( .A1(n6497), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6954 ( .A1(n5657), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5422) );
  AND2_X1 U6955 ( .A1(n5418), .A2(n5417), .ZN(n5419) );
  NOR2_X1 U6956 ( .A1(n5438), .A2(n5419), .ZN(n8560) );
  NAND2_X1 U6957 ( .A1(n5631), .A2(n8560), .ZN(n5421) );
  NAND2_X1 U6958 ( .A1(n5661), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5420) );
  INV_X1 U6959 ( .A(n8738), .ZN(n8982) );
  AOI22_X1 U6960 ( .A1(n7517), .A2(n8593), .B1(n5616), .B2(n8982), .ZN(n5424)
         );
  XNOR2_X1 U6961 ( .A(n5424), .B(n4413), .ZN(n5425) );
  OAI22_X1 U6962 ( .A1(n9666), .A2(n5493), .B1(n8738), .B2(n8588), .ZN(n8555)
         );
  INV_X1 U6963 ( .A(n5448), .ZN(n5446) );
  INV_X1 U6964 ( .A(n5427), .ZN(n5430) );
  INV_X1 U6965 ( .A(n5428), .ZN(n5429) );
  INV_X1 U6966 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6691) );
  MUX2_X1 U6967 ( .A(n6691), .B(n10143), .S(n5876), .Z(n5451) );
  XNOR2_X1 U6968 ( .A(n5451), .B(SI_15_), .ZN(n5433) );
  XNOR2_X1 U6969 ( .A(n5453), .B(n5433), .ZN(n6690) );
  NAND2_X1 U6970 ( .A1(n6690), .A2(n4905), .ZN(n5437) );
  NAND2_X1 U6971 ( .A1(n5434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U6972 ( .A(n5435), .B(P1_IR_REG_15__SCAN_IN), .ZN(n6962) );
  AOI22_X1 U6973 ( .A1(n5548), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5547), .B2(
        n6962), .ZN(n5436) );
  NAND2_X1 U6974 ( .A1(n6497), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6975 ( .A1(n5460), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5442) );
  OR2_X1 U6976 ( .A1(n5438), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6977 ( .A1(n5438), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5463) );
  AND2_X1 U6978 ( .A1(n5439), .A2(n5463), .ZN(n8743) );
  NAND2_X1 U6979 ( .A1(n5631), .A2(n8743), .ZN(n5441) );
  NAND2_X1 U6980 ( .A1(n5461), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5440) );
  AOI22_X1 U6981 ( .A1(n7558), .A2(n8593), .B1(n5616), .B2(n8981), .ZN(n5444)
         );
  XNOR2_X1 U6982 ( .A(n5444), .B(n4530), .ZN(n5447) );
  INV_X1 U6983 ( .A(n5447), .ZN(n5445) );
  NAND2_X1 U6984 ( .A1(n5448), .A2(n5447), .ZN(n5450) );
  OAI22_X1 U6985 ( .A1(n9522), .A2(n5493), .B1(n9514), .B2(n8588), .ZN(n8732)
         );
  MUX2_X1 U6986 ( .A(n10114), .B(n6820), .S(n4660), .Z(n5474) );
  XNOR2_X1 U6987 ( .A(n5474), .B(SI_16_), .ZN(n5454) );
  XNOR2_X1 U6988 ( .A(n5476), .B(n5454), .ZN(n6795) );
  NAND2_X1 U6989 ( .A1(n6795), .A2(n4905), .ZN(n5459) );
  NAND2_X1 U6990 ( .A1(n4492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5455) );
  MUX2_X1 U6991 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5455), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5457) );
  NAND2_X1 U6992 ( .A1(n5457), .A2(n5481), .ZN(n7221) );
  AOI22_X1 U6993 ( .A1(n5548), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5547), .B2(
        n7227), .ZN(n5458) );
  NAND2_X1 U6994 ( .A1(n5460), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6995 ( .A1(n5461), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5467) );
  INV_X1 U6996 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6997 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  AND2_X1 U6998 ( .A1(n5487), .A2(n5464), .ZN(n8652) );
  NAND2_X1 U6999 ( .A1(n5631), .A2(n8652), .ZN(n5466) );
  NAND2_X1 U7000 ( .A1(n6497), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5465) );
  AOI22_X1 U7001 ( .A1(n9101), .A2(n8593), .B1(n4402), .B2(n9298), .ZN(n5469)
         );
  XOR2_X1 U7002 ( .A(n4413), .B(n5469), .Z(n5471) );
  INV_X1 U7003 ( .A(n5616), .ZN(n5593) );
  OAI22_X1 U7004 ( .A1(n4668), .A2(n5593), .B1(n8661), .B2(n8588), .ZN(n5470)
         );
  NOR2_X1 U7005 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  AOI21_X1 U7006 ( .B1(n5471), .B2(n5470), .A(n5472), .ZN(n8647) );
  INV_X1 U7007 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U7008 ( .A1(n8645), .A2(n5473), .ZN(n8656) );
  MUX2_X1 U7009 ( .A(n6866), .B(n6863), .S(n5876), .Z(n5478) );
  NAND2_X1 U7010 ( .A1(n5478), .A2(n5477), .ZN(n5502) );
  INV_X1 U7011 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U7012 ( .A1(n5479), .A2(SI_17_), .ZN(n5480) );
  NAND2_X1 U7013 ( .A1(n5502), .A2(n5480), .ZN(n5500) );
  XNOR2_X1 U7014 ( .A(n5501), .B(n5500), .ZN(n6862) );
  NAND2_X1 U7015 ( .A1(n6862), .A2(n4905), .ZN(n5486) );
  NAND2_X1 U7016 ( .A1(n5481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5482) );
  MUX2_X1 U7017 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5482), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n5484) );
  NAND2_X1 U7018 ( .A1(n5484), .A2(n5483), .ZN(n7305) );
  INV_X1 U7019 ( .A(n7305), .ZN(n7296) );
  AOI22_X1 U7020 ( .A1(n5548), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5547), .B2(
        n7296), .ZN(n5485) );
  NAND2_X1 U7021 ( .A1(n6497), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7022 ( .A1(n5657), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5491) );
  AND2_X1 U7023 ( .A1(n5487), .A2(n10081), .ZN(n5488) );
  NOR2_X1 U7024 ( .A1(n5551), .A2(n5488), .ZN(n9290) );
  NAND2_X1 U7025 ( .A1(n5631), .A2(n9290), .ZN(n5490) );
  NAND2_X1 U7026 ( .A1(n5661), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5489) );
  NAND4_X1 U7027 ( .A1(n5492), .A2(n5491), .A3(n5490), .A4(n5489), .ZN(n9483)
         );
  OAI22_X1 U7028 ( .A1(n9509), .A2(n5493), .B1(n9102), .B2(n8588), .ZN(n5497)
         );
  NAND2_X1 U7029 ( .A1(n9292), .A2(n8593), .ZN(n5495) );
  NAND2_X1 U7030 ( .A1(n9483), .A2(n4402), .ZN(n5494) );
  NAND2_X1 U7031 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  XNOR2_X1 U7032 ( .A(n5496), .B(n4413), .ZN(n5498) );
  XOR2_X1 U7033 ( .A(n5497), .B(n5498), .Z(n8657) );
  MUX2_X1 U7034 ( .A(n10172), .B(n6918), .S(n4660), .Z(n5503) );
  XNOR2_X1 U7035 ( .A(n5503), .B(SI_18_), .ZN(n5541) );
  INV_X1 U7036 ( .A(n5541), .ZN(n5506) );
  INV_X1 U7037 ( .A(n5503), .ZN(n5504) );
  NAND2_X1 U7038 ( .A1(n5504), .A2(SI_18_), .ZN(n5505) );
  OAI21_X1 U7039 ( .B1(n5542), .B2(n5506), .A(n5505), .ZN(n5527) );
  MUX2_X1 U7040 ( .A(n7683), .B(n7617), .S(n5876), .Z(n5508) );
  NAND2_X1 U7041 ( .A1(n5508), .A2(n5507), .ZN(n5511) );
  INV_X1 U7042 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7043 ( .A1(n5509), .A2(SI_19_), .ZN(n5510) );
  NAND2_X1 U7044 ( .A1(n5511), .A2(n5510), .ZN(n5526) );
  MUX2_X1 U7045 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4660), .Z(n5576) );
  XNOR2_X1 U7046 ( .A(n5576), .B(n5578), .ZN(n5513) );
  XNOR2_X1 U7047 ( .A(n5579), .B(n5513), .ZN(n7204) );
  NAND2_X1 U7048 ( .A1(n7204), .A2(n4905), .ZN(n5515) );
  INV_X1 U7049 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7203) );
  OR2_X1 U7050 ( .A1(n8823), .A2(n7203), .ZN(n5514) );
  NAND2_X1 U7051 ( .A1(n9377), .A2(n8593), .ZN(n5522) );
  NAND2_X1 U7052 ( .A1(n6497), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7053 ( .A1(n5657), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7054 ( .A1(n5551), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5552) );
  INV_X1 U7055 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7056 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n5530), .ZN(n5585) );
  OAI21_X1 U7057 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5530), .A(n5585), .ZN(
        n5516) );
  INV_X1 U7058 ( .A(n5516), .ZN(n9258) );
  NAND2_X1 U7059 ( .A1(n5631), .A2(n9258), .ZN(n5518) );
  NAND2_X1 U7060 ( .A1(n5661), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5517) );
  NAND4_X1 U7061 ( .A1(n5520), .A2(n5519), .A3(n5518), .A4(n5517), .ZN(n9370)
         );
  NAND2_X1 U7062 ( .A1(n9370), .A2(n4402), .ZN(n5521) );
  NAND2_X1 U7063 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  XNOR2_X1 U7064 ( .A(n5523), .B(n4530), .ZN(n5570) );
  NAND2_X1 U7065 ( .A1(n9377), .A2(n5616), .ZN(n5525) );
  NAND2_X1 U7066 ( .A1(n9370), .A2(n5639), .ZN(n5524) );
  NAND2_X1 U7067 ( .A1(n5525), .A2(n5524), .ZN(n5571) );
  XNOR2_X1 U7068 ( .A(n5527), .B(n5526), .ZN(n7616) );
  NAND2_X1 U7069 ( .A1(n7616), .A2(n4905), .ZN(n5529) );
  AOI22_X1 U7070 ( .A1(n5548), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5547), .B2(
        n9493), .ZN(n5528) );
  NAND2_X1 U7071 ( .A1(n9384), .A2(n8593), .ZN(n5537) );
  AOI21_X1 U7072 ( .B1(n5552), .B2(n5531), .A(n5530), .ZN(n9280) );
  NAND2_X1 U7073 ( .A1(n5631), .A2(n9280), .ZN(n5535) );
  NAND2_X1 U7074 ( .A1(n5661), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7075 ( .A1(n6497), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7076 ( .A1(n5657), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5532) );
  NAND4_X1 U7077 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n9484)
         );
  NAND2_X1 U7078 ( .A1(n9484), .A2(n5616), .ZN(n5536) );
  NAND2_X1 U7079 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  XNOR2_X1 U7080 ( .A(n5538), .B(n4413), .ZN(n5566) );
  NAND2_X1 U7081 ( .A1(n9384), .A2(n5616), .ZN(n5540) );
  NAND2_X1 U7082 ( .A1(n9484), .A2(n5639), .ZN(n5539) );
  NAND2_X1 U7083 ( .A1(n5540), .A2(n5539), .ZN(n8575) );
  NAND2_X1 U7084 ( .A1(n5566), .A2(n8575), .ZN(n8676) );
  XNOR2_X1 U7085 ( .A(n5542), .B(n5541), .ZN(n6916) );
  NAND2_X1 U7086 ( .A1(n6916), .A2(n4905), .ZN(n5550) );
  OR2_X1 U7087 ( .A1(n5544), .A2(n5543), .ZN(n5545) );
  AND2_X1 U7088 ( .A1(n5546), .A2(n5545), .ZN(n7418) );
  AOI22_X1 U7089 ( .A1(n5548), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5547), .B2(
        n7418), .ZN(n5549) );
  NAND2_X1 U7090 ( .A1(n9488), .A2(n8593), .ZN(n5559) );
  NAND2_X1 U7091 ( .A1(n5657), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5557) );
  OR2_X1 U7092 ( .A1(n5551), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7093 ( .A1(n5553), .A2(n5552), .ZN(n9500) );
  INV_X1 U7094 ( .A(n9500), .ZN(n8727) );
  NAND2_X1 U7095 ( .A1(n5631), .A2(n8727), .ZN(n5556) );
  NAND2_X1 U7096 ( .A1(n5661), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7097 ( .A1(n6497), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5554) );
  NAND4_X1 U7098 ( .A1(n5557), .A2(n5556), .A3(n5555), .A4(n5554), .ZN(n9299)
         );
  NAND2_X1 U7099 ( .A1(n9299), .A2(n5616), .ZN(n5558) );
  NAND2_X1 U7100 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  XNOR2_X1 U7101 ( .A(n5560), .B(n4530), .ZN(n8573) );
  NAND2_X1 U7102 ( .A1(n9488), .A2(n4402), .ZN(n5562) );
  NAND2_X1 U7103 ( .A1(n9299), .A2(n5639), .ZN(n5561) );
  NAND2_X1 U7104 ( .A1(n5562), .A2(n5561), .ZN(n8572) );
  NAND2_X1 U7105 ( .A1(n8573), .A2(n8572), .ZN(n5563) );
  NAND2_X1 U7106 ( .A1(n8676), .A2(n5563), .ZN(n5564) );
  INV_X1 U7107 ( .A(n5566), .ZN(n8576) );
  OAI21_X1 U7108 ( .B1(n8573), .B2(n8572), .A(n8575), .ZN(n5568) );
  NOR3_X1 U7109 ( .A1(n8573), .A2(n8575), .A3(n8572), .ZN(n5567) );
  AOI21_X1 U7110 ( .B1(n8576), .B2(n5568), .A(n5567), .ZN(n5569) );
  INV_X1 U7111 ( .A(n5570), .ZN(n5573) );
  INV_X1 U7112 ( .A(n5571), .ZN(n5572) );
  NAND2_X1 U7113 ( .A1(n5573), .A2(n5572), .ZN(n8616) );
  INV_X1 U7114 ( .A(n5576), .ZN(n5577) );
  MUX2_X1 U7115 ( .A(n10110), .B(n7294), .S(n5876), .Z(n5600) );
  XNOR2_X1 U7116 ( .A(n5600), .B(SI_21_), .ZN(n5582) );
  XNOR2_X1 U7117 ( .A(n5604), .B(n5582), .ZN(n7292) );
  NAND2_X1 U7118 ( .A1(n7292), .A2(n4905), .ZN(n5584) );
  OR2_X1 U7119 ( .A1(n8823), .A2(n7294), .ZN(n5583) );
  AND2_X2 U7120 ( .A1(n5584), .A2(n5583), .ZN(n9250) );
  INV_X2 U7121 ( .A(n9250), .ZN(n9371) );
  NAND2_X1 U7122 ( .A1(n6497), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7123 ( .A1(n5657), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5590) );
  OAI21_X1 U7124 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n5586), .A(n5629), .ZN(
        n5587) );
  INV_X1 U7125 ( .A(n5587), .ZN(n9246) );
  NAND2_X1 U7126 ( .A1(n5631), .A2(n9246), .ZN(n5589) );
  NAND2_X1 U7127 ( .A1(n5661), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5588) );
  AOI22_X1 U7128 ( .A1(n9371), .A2(n8593), .B1(n4402), .B2(n9363), .ZN(n5592)
         );
  XNOR2_X1 U7129 ( .A(n5592), .B(n4413), .ZN(n5597) );
  OAI22_X1 U7130 ( .A1(n9250), .A2(n5593), .B1(n9232), .B2(n8588), .ZN(n5595)
         );
  XNOR2_X1 U7131 ( .A(n5597), .B(n5595), .ZN(n8614) );
  INV_X1 U7132 ( .A(n5595), .ZN(n5596) );
  NAND2_X1 U7133 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  INV_X1 U7134 ( .A(SI_21_), .ZN(n5599) );
  AND2_X1 U7135 ( .A1(n5600), .A2(n5599), .ZN(n5603) );
  INV_X1 U7136 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7137 ( .A1(n5601), .A2(SI_21_), .ZN(n5602) );
  MUX2_X1 U7138 ( .A(n7437), .B(n7439), .S(n4660), .Z(n5606) );
  INV_X1 U7139 ( .A(SI_22_), .ZN(n5605) );
  NAND2_X1 U7140 ( .A1(n5606), .A2(n5605), .ZN(n5617) );
  INV_X1 U7141 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U7142 ( .A1(n5607), .A2(SI_22_), .ZN(n5608) );
  NAND2_X1 U7143 ( .A1(n5617), .A2(n5608), .ZN(n5618) );
  XNOR2_X1 U7144 ( .A(n5619), .B(n5618), .ZN(n7436) );
  NAND2_X1 U7145 ( .A1(n7436), .A2(n4905), .ZN(n5610) );
  OR2_X1 U7146 ( .A1(n8823), .A2(n7439), .ZN(n5609) );
  NAND2_X1 U7147 ( .A1(n6497), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7148 ( .A1(n5657), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5613) );
  XNOR2_X1 U7149 ( .A(n5629), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U7150 ( .A1(n5631), .A2(n9230), .ZN(n5612) );
  NAND2_X1 U7151 ( .A1(n5661), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5611) );
  AOI22_X1 U7152 ( .A1(n9364), .A2(n8593), .B1(n4402), .B2(n9242), .ZN(n5615)
         );
  XNOR2_X1 U7153 ( .A(n5615), .B(n4530), .ZN(n5646) );
  OAI22_X1 U7154 ( .A1(n9235), .A2(n5493), .B1(n9356), .B2(n8588), .ZN(n8686)
         );
  MUX2_X1 U7155 ( .A(n7507), .B(n10037), .S(n4660), .Z(n5621) );
  INV_X1 U7156 ( .A(SI_23_), .ZN(n5620) );
  NAND2_X1 U7157 ( .A1(n5621), .A2(n5620), .ZN(n5650) );
  INV_X1 U7158 ( .A(n5621), .ZN(n5622) );
  NAND2_X1 U7159 ( .A1(n5622), .A2(SI_23_), .ZN(n5623) );
  NAND2_X1 U7160 ( .A1(n7509), .A2(n4905), .ZN(n5625) );
  OR2_X1 U7161 ( .A1(n8823), .A2(n10037), .ZN(n5624) );
  NAND2_X1 U7162 ( .A1(n9213), .A2(n8593), .ZN(n5637) );
  NAND2_X1 U7163 ( .A1(n5657), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7164 ( .A1(n6497), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5634) );
  INV_X1 U7165 ( .A(n5629), .ZN(n5627) );
  AND2_X1 U7166 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5626) );
  NAND2_X1 U7167 ( .A1(n5627), .A2(n5626), .ZN(n5659) );
  INV_X1 U7168 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8689) );
  INV_X1 U7169 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5628) );
  OAI21_X1 U7170 ( .B1(n5629), .B2(n8689), .A(n5628), .ZN(n5630) );
  AND2_X1 U7171 ( .A1(n5659), .A2(n5630), .ZN(n9214) );
  NAND2_X1 U7172 ( .A1(n5631), .A2(n9214), .ZN(n5633) );
  NAND2_X1 U7173 ( .A1(n5661), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5632) );
  NAND4_X1 U7174 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n9226)
         );
  NAND2_X1 U7175 ( .A1(n9226), .A2(n5616), .ZN(n5636) );
  NAND2_X1 U7176 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  XNOR2_X1 U7177 ( .A(n5638), .B(n8591), .ZN(n5641) );
  AND2_X1 U7178 ( .A1(n9226), .A2(n5639), .ZN(n5640) );
  AOI21_X1 U7179 ( .B1(n9213), .B2(n5616), .A(n5640), .ZN(n5642) );
  NAND2_X1 U7180 ( .A1(n5641), .A2(n5642), .ZN(n8665) );
  INV_X1 U7181 ( .A(n5641), .ZN(n5644) );
  INV_X1 U7182 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7183 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  INV_X1 U7184 ( .A(n5646), .ZN(n5647) );
  INV_X1 U7185 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7564) );
  INV_X1 U7186 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7566) );
  MUX2_X1 U7187 ( .A(n7564), .B(n7566), .S(n4660), .Z(n5652) );
  INV_X1 U7188 ( .A(SI_24_), .ZN(n5651) );
  NAND2_X1 U7189 ( .A1(n5652), .A2(n5651), .ZN(n5680) );
  INV_X1 U7190 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7191 ( .A1(n5653), .A2(SI_24_), .ZN(n5654) );
  XNOR2_X1 U7192 ( .A(n5679), .B(n5678), .ZN(n7563) );
  NAND2_X1 U7193 ( .A1(n7563), .A2(n4905), .ZN(n5656) );
  OR2_X1 U7194 ( .A1(n8823), .A2(n7566), .ZN(n5655) );
  NAND2_X1 U7195 ( .A1(n5657), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7196 ( .A1(n6497), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5664) );
  INV_X1 U7197 ( .A(n5659), .ZN(n5658) );
  NAND2_X1 U7198 ( .A1(n5658), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5689) );
  INV_X1 U7199 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U7200 ( .A1(n5659), .A2(n10131), .ZN(n5660) );
  AND2_X1 U7201 ( .A1(n5689), .A2(n5660), .ZN(n9205) );
  NAND2_X1 U7202 ( .A1(n5210), .A2(n9205), .ZN(n5663) );
  NAND2_X1 U7203 ( .A1(n5461), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5662) );
  OAI22_X1 U7204 ( .A1(n9208), .A2(n5666), .B1(n9191), .B2(n5493), .ZN(n5667)
         );
  XNOR2_X1 U7205 ( .A(n5667), .B(n8591), .ZN(n5670) );
  OR2_X1 U7206 ( .A1(n9208), .A2(n5493), .ZN(n5669) );
  OR2_X1 U7207 ( .A1(n9191), .A2(n8588), .ZN(n5668) );
  NAND2_X1 U7208 ( .A1(n5670), .A2(n5671), .ZN(n5677) );
  INV_X1 U7209 ( .A(n5670), .ZN(n5673) );
  INV_X1 U7210 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U7211 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  NAND2_X1 U7212 ( .A1(n5679), .A2(n5678), .ZN(n5681) );
  INV_X1 U7213 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7570) );
  INV_X1 U7214 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7572) );
  MUX2_X1 U7215 ( .A(n7570), .B(n7572), .S(n4660), .Z(n5683) );
  INV_X1 U7216 ( .A(SI_25_), .ZN(n5682) );
  NAND2_X1 U7217 ( .A1(n5683), .A2(n5682), .ZN(n5704) );
  INV_X1 U7218 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U7219 ( .A1(n5684), .A2(SI_25_), .ZN(n5685) );
  XNOR2_X1 U7220 ( .A(n5703), .B(n5702), .ZN(n7569) );
  NAND2_X1 U7221 ( .A1(n7569), .A2(n4905), .ZN(n5687) );
  OR2_X1 U7222 ( .A1(n8823), .A2(n7572), .ZN(n5686) );
  NAND2_X1 U7223 ( .A1(n5657), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7224 ( .A1(n6497), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5693) );
  INV_X1 U7225 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7226 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  AND2_X1 U7227 ( .A1(n5711), .A2(n5690), .ZN(n9189) );
  NAND2_X1 U7228 ( .A1(n5210), .A2(n9189), .ZN(n5692) );
  NAND2_X1 U7229 ( .A1(n5661), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5691) );
  NAND4_X1 U7230 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(n9201)
         );
  INV_X1 U7231 ( .A(n9201), .ZN(n8747) );
  OAI22_X1 U7232 ( .A1(n9193), .A2(n5493), .B1(n8747), .B2(n8588), .ZN(n5699)
         );
  NAND2_X1 U7233 ( .A1(n9346), .A2(n8593), .ZN(n5696) );
  NAND2_X1 U7234 ( .A1(n9201), .A2(n4402), .ZN(n5695) );
  NAND2_X1 U7235 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  XNOR2_X1 U7236 ( .A(n5697), .B(n4413), .ZN(n5698) );
  XOR2_X1 U7237 ( .A(n5699), .B(n5698), .Z(n8639) );
  INV_X1 U7238 ( .A(n5698), .ZN(n5701) );
  INV_X1 U7239 ( .A(n5699), .ZN(n5700) );
  NAND2_X1 U7240 ( .A1(n5701), .A2(n5700), .ZN(n5746) );
  INV_X1 U7241 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7576) );
  INV_X1 U7242 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7577) );
  MUX2_X1 U7243 ( .A(n7576), .B(n7577), .S(n4660), .Z(n5706) );
  INV_X1 U7244 ( .A(SI_26_), .ZN(n5705) );
  NAND2_X1 U7245 ( .A1(n5706), .A2(n5705), .ZN(n5824) );
  INV_X1 U7246 ( .A(n5706), .ZN(n5707) );
  NAND2_X1 U7247 ( .A1(n5707), .A2(SI_26_), .ZN(n5708) );
  NAND2_X1 U7248 ( .A1(n7575), .A2(n4905), .ZN(n5710) );
  OR2_X1 U7249 ( .A1(n8823), .A2(n7577), .ZN(n5709) );
  NAND2_X1 U7250 ( .A1(n9339), .A2(n8593), .ZN(n5718) );
  NAND2_X1 U7251 ( .A1(n8598), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7252 ( .A1(n5657), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5715) );
  INV_X1 U7253 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7254 ( .A1(n5711), .A2(n5763), .ZN(n5712) );
  NAND2_X1 U7255 ( .A1(n5210), .A2(n9169), .ZN(n5714) );
  NAND2_X1 U7256 ( .A1(n5461), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5713) );
  OR2_X1 U7257 ( .A1(n9332), .A2(n5593), .ZN(n5717) );
  NAND2_X1 U7258 ( .A1(n5718), .A2(n5717), .ZN(n5720) );
  XNOR2_X1 U7259 ( .A(n5720), .B(n4530), .ZN(n7583) );
  NOR2_X1 U7260 ( .A1(n9332), .A2(n8588), .ZN(n5721) );
  AOI21_X1 U7261 ( .B1(n9339), .B2(n4402), .A(n5721), .ZN(n7584) );
  XNOR2_X1 U7262 ( .A(n7583), .B(n7584), .ZN(n5748) );
  NAND2_X1 U7263 ( .A1(n7574), .A2(P1_B_REG_SCAN_IN), .ZN(n5723) );
  INV_X1 U7264 ( .A(n7568), .ZN(n5722) );
  MUX2_X1 U7265 ( .A(n5723), .B(P1_B_REG_SCAN_IN), .S(n5722), .Z(n5724) );
  NAND2_X1 U7266 ( .A1(n7579), .A2(n7568), .ZN(n9403) );
  INV_X1 U7267 ( .A(n9313), .ZN(n9387) );
  NAND2_X1 U7268 ( .A1(n7579), .A2(n7574), .ZN(n9402) );
  OAI21_X1 U7269 ( .B1(n6950), .B2(P1_D_REG_1__SCAN_IN), .A(n9402), .ZN(n9311)
         );
  INV_X1 U7270 ( .A(n9311), .ZN(n6954) );
  INV_X1 U7271 ( .A(n6950), .ZN(n5735) );
  NOR2_X1 U7272 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n9985) );
  NOR4_X1 U7273 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5728) );
  NOR4_X1 U7274 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5727) );
  NOR4_X1 U7275 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5726) );
  AND4_X1 U7276 ( .A1(n9985), .A2(n5728), .A3(n5727), .A4(n5726), .ZN(n5734)
         );
  NOR4_X1 U7277 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5732) );
  NOR4_X1 U7278 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5731) );
  NOR4_X1 U7279 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n5730) );
  NOR4_X1 U7280 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5729) );
  AND4_X1 U7281 ( .A1(n5732), .A2(n5731), .A3(n5730), .A4(n5729), .ZN(n5733)
         );
  NAND2_X1 U7282 ( .A1(n5734), .A2(n5733), .ZN(n6952) );
  NAND2_X1 U7283 ( .A1(n5735), .A2(n6952), .ZN(n9310) );
  AND3_X1 U7284 ( .A1(n9387), .A2(n6954), .A3(n9310), .ZN(n5767) );
  NAND2_X1 U7285 ( .A1(n8912), .A2(n8835), .ZN(n7002) );
  INV_X1 U7286 ( .A(n7002), .ZN(n9561) );
  OR2_X1 U7287 ( .A1(n9625), .A2(n8904), .ZN(n5751) );
  INV_X1 U7288 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7289 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  NAND2_X1 U7290 ( .A1(n5742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5744) );
  NOR2_X1 U7291 ( .A1(n5751), .A2(n9307), .ZN(n5745) );
  OAI211_X1 U7292 ( .C1(n5749), .C2(n5748), .A(n8722), .B(n7600), .ZN(n5773)
         );
  INV_X1 U7293 ( .A(n5767), .ZN(n5757) );
  INV_X1 U7294 ( .A(n8904), .ZN(n5750) );
  OR2_X1 U7295 ( .A1(n5768), .A2(P1_U3086), .ZN(n7201) );
  NAND3_X1 U7296 ( .A1(n5751), .A2(n7003), .A3(n7201), .ZN(n5752) );
  NAND2_X1 U7297 ( .A1(n5757), .A2(n5752), .ZN(n5753) );
  AND2_X1 U7298 ( .A1(n8904), .A2(n5738), .ZN(n9308) );
  INV_X1 U7299 ( .A(n9308), .ZN(n6953) );
  NAND2_X1 U7300 ( .A1(n5753), .A2(n6953), .ZN(n6695) );
  OAI21_X1 U7301 ( .B1(n6695), .B2(n5754), .A(P1_STATE_REG_SCAN_IN), .ZN(n5755) );
  OR2_X1 U7302 ( .A1(n9307), .A2(n5738), .ZN(n5756) );
  NOR2_X1 U7303 ( .A1(n5757), .A2(n5756), .ZN(n5762) );
  NAND2_X1 U7304 ( .A1(n5657), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7305 ( .A1(n8598), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7306 ( .A(n7604), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U7307 ( .A1(n5210), .A2(n9156), .ZN(n5759) );
  NAND2_X1 U7308 ( .A1(n5461), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5758) );
  NOR2_X1 U7309 ( .A1(n8704), .A2(n9325), .ZN(n5765) );
  OAI22_X1 U7310 ( .A1(n8737), .A2(n8747), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5763), .ZN(n5764) );
  AOI211_X1 U7311 ( .C1(n9169), .C2(n8742), .A(n5765), .B(n5764), .ZN(n5772)
         );
  INV_X1 U7312 ( .A(n9339), .ZN(n9171) );
  OR2_X1 U7313 ( .A1(n7002), .A2(n5768), .ZN(n9492) );
  NOR2_X1 U7314 ( .A1(n9307), .A2(n9492), .ZN(n5766) );
  NAND2_X1 U7315 ( .A1(n5767), .A2(n5766), .ZN(n5769) );
  NAND2_X1 U7316 ( .A1(n9668), .A2(n8835), .ZN(n9309) );
  NAND2_X1 U7317 ( .A1(n9339), .A2(n5770), .ZN(n5771) );
  NAND3_X1 U7318 ( .A1(n5773), .A2(n5772), .A3(n5771), .ZN(P1_U3240) );
  INV_X1 U7319 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7320 ( .A1(n9891), .A2(n5774), .ZN(n5906) );
  INV_X1 U7321 ( .A(n5906), .ZN(n5776) );
  NAND2_X1 U7322 ( .A1(n5776), .A2(n5775), .ZN(n5924) );
  INV_X1 U7323 ( .A(n5934), .ZN(n5778) );
  NAND2_X1 U7324 ( .A1(n5778), .A2(n5777), .ZN(n5947) );
  INV_X1 U7325 ( .A(n5960), .ZN(n5780) );
  INV_X1 U7326 ( .A(n6016), .ZN(n5783) );
  INV_X1 U7327 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U7328 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5785) );
  INV_X1 U7329 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5787) );
  INV_X1 U7330 ( .A(n6117), .ZN(n5790) );
  INV_X1 U7331 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5789) );
  INV_X1 U7332 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5791) );
  INV_X1 U7333 ( .A(n6153), .ZN(n5794) );
  INV_X1 U7334 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5793) );
  INV_X1 U7335 ( .A(n6175), .ZN(n5796) );
  INV_X1 U7336 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7337 ( .A1(n5796), .A2(n5795), .ZN(n6177) );
  NAND2_X1 U7338 ( .A1(n6177), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7339 ( .A1(n8150), .A2(n5797), .ZN(n8169) );
  NOR2_X1 U7340 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5806) );
  NAND4_X1 U7341 ( .A1(n5806), .A2(n5981), .A3(n6202), .A4(n6205), .ZN(n5807)
         );
  INV_X1 U7342 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5813) );
  XNOR2_X2 U7343 ( .A(n5814), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7344 ( .A1(n8169), .A2(n6191), .ZN(n5821) );
  INV_X1 U7345 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U7346 ( .A1(n7894), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7347 ( .A1(n5889), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5817) );
  OAI211_X1 U7348 ( .C1(n8383), .C2(n5870), .A(n5818), .B(n5817), .ZN(n5819)
         );
  INV_X1 U7349 ( .A(n5819), .ZN(n5820) );
  INV_X1 U7350 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10163) );
  INV_X1 U7351 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10186) );
  MUX2_X1 U7352 ( .A(n10163), .B(n10186), .S(n4660), .Z(n5827) );
  INV_X1 U7353 ( .A(SI_27_), .ZN(n5826) );
  NAND2_X1 U7354 ( .A1(n5827), .A2(n5826), .ZN(n5830) );
  INV_X1 U7355 ( .A(n5827), .ZN(n5828) );
  NAND2_X1 U7356 ( .A1(n5828), .A2(SI_27_), .ZN(n5829) );
  INV_X1 U7357 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10065) );
  INV_X1 U7358 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10051) );
  MUX2_X1 U7359 ( .A(n10065), .B(n10051), .S(n4660), .Z(n6189) );
  XNOR2_X1 U7360 ( .A(n6189), .B(SI_28_), .ZN(n6187) );
  INV_X1 U7361 ( .A(n5831), .ZN(n5834) );
  NAND2_X1 U7362 ( .A1(n5837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7363 ( .A1(n5834), .A2(n5833), .ZN(n6239) );
  NAND2_X1 U7364 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5835) );
  AOI22_X1 U7365 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n6200), .B1(n5835), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7366 ( .A1(n8585), .A2(n7890), .ZN(n5840) );
  NAND2_X2 U7367 ( .A1(n5862), .A2(n4660), .ZN(n5864) );
  OR2_X1 U7368 ( .A1(n5864), .A2(n10065), .ZN(n5839) );
  INV_X1 U7369 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10092) );
  OR2_X1 U7370 ( .A1(n5870), .A2(n10092), .ZN(n5844) );
  INV_X1 U7371 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7264) );
  OR2_X1 U7372 ( .A1(n5868), .A2(n7264), .ZN(n5843) );
  NAND2_X1 U7373 ( .A1(n5889), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5842) );
  INV_X1 U7374 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7267) );
  OR2_X1 U7375 ( .A1(n5869), .A2(n7267), .ZN(n5841) );
  OR2_X1 U7376 ( .A1(n5865), .A2(n6471), .ZN(n5883) );
  OR2_X1 U7377 ( .A1(n5864), .A2(n6455), .ZN(n5882) );
  OR2_X1 U7378 ( .A1(n5845), .A2(n6200), .ZN(n5847) );
  XNOR2_X2 U7379 ( .A(n5847), .B(n5846), .ZN(n6454) );
  OR2_X1 U7380 ( .A1(n5896), .A2(n6454), .ZN(n5881) );
  OR2_X1 U7381 ( .A1(n9884), .A2(n7263), .ZN(n7942) );
  NAND2_X1 U7382 ( .A1(n9884), .A2(n7263), .ZN(n7940) );
  NAND2_X1 U7383 ( .A1(n5889), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7384 ( .A1(n5868), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5852) );
  INV_X1 U7385 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5848) );
  OR2_X1 U7386 ( .A1(n5870), .A2(n5848), .ZN(n5851) );
  INV_X1 U7387 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7388 ( .A1(n5869), .A2(n5849), .ZN(n5850) );
  NAND2_X1 U7389 ( .A1(n5854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5856) );
  INV_X1 U7390 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7391 ( .A1(n5865), .A2(n6469), .ZN(n5858) );
  INV_X1 U7392 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6456) );
  OR2_X1 U7393 ( .A1(n5864), .A2(n6456), .ZN(n5857) );
  OAI211_X1 U7394 ( .C1(n5896), .C2(n9724), .A(n5858), .B(n5857), .ZN(n9896)
         );
  NAND2_X1 U7395 ( .A1(n8112), .A2(n9896), .ZN(n5880) );
  AND2_X1 U7396 ( .A1(n9878), .A2(n5880), .ZN(n5888) );
  INV_X1 U7397 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9706) );
  INV_X1 U7398 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7140) );
  NAND2_X1 U7399 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5859) );
  MUX2_X1 U7400 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5859), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5860) );
  INV_X1 U7401 ( .A(n9703), .ZN(n5861) );
  OR2_X1 U7402 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  OAI21_X1 U7403 ( .B1(P1_DATAO_REG_1__SCAN_IN), .B2(n5864), .A(n5863), .ZN(
        n5867) );
  NOR2_X1 U7404 ( .A1(n5865), .A2(n6457), .ZN(n5866) );
  NOR2_X2 U7405 ( .A1(n5867), .A2(n5866), .ZN(n6880) );
  NAND2_X1 U7406 ( .A1(n5889), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5873) );
  INV_X1 U7407 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6811) );
  OR2_X1 U7408 ( .A1(n5868), .A2(n6811), .ZN(n5872) );
  INV_X1 U7409 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7288) );
  OR2_X1 U7410 ( .A1(n5869), .A2(n7288), .ZN(n5871) );
  NAND4_X1 U7411 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n4451), .ZN(n6214)
         );
  INV_X1 U7412 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5874) );
  OAI21_X1 U7413 ( .B1(n5876), .B2(n5875), .A(n5874), .ZN(n5877) );
  AND2_X1 U7414 ( .A1(n5878), .A2(n5877), .ZN(n8551) );
  MUX2_X1 U7415 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8551), .S(n5896), .Z(n6808) );
  NAND2_X1 U7416 ( .A1(n6214), .A2(n6808), .ZN(n6841) );
  OR2_X1 U7417 ( .A1(n6731), .A2(n6880), .ZN(n5879) );
  INV_X1 U7418 ( .A(n5880), .ZN(n5887) );
  NAND3_X1 U7419 ( .A1(n5883), .A2(n5882), .A3(n5881), .ZN(n6805) );
  OR2_X1 U7420 ( .A1(n9884), .A2(n6805), .ZN(n9880) );
  INV_X1 U7421 ( .A(n9880), .ZN(n5885) );
  NOR2_X1 U7422 ( .A1(n8112), .A2(n9896), .ZN(n5884) );
  NOR2_X1 U7423 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  AOI21_X2 U7424 ( .B1(n5888), .B2(n9879), .A(n5034), .ZN(n6929) );
  NAND2_X1 U7425 ( .A1(n7894), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5895) );
  INV_X1 U7426 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5890) );
  OR2_X1 U7427 ( .A1(n6244), .A2(n5890), .ZN(n5894) );
  NAND2_X1 U7428 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5891) );
  AND2_X1 U7429 ( .A1(n5906), .A2(n5891), .ZN(n6909) );
  OR2_X1 U7430 ( .A1(n6109), .A2(n6909), .ZN(n5893) );
  INV_X1 U7431 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6398) );
  OR2_X1 U7432 ( .A1(n5870), .A2(n6398), .ZN(n5892) );
  OR2_X1 U7433 ( .A1(n5865), .A2(n6473), .ZN(n5904) );
  OR2_X1 U7434 ( .A1(n5864), .A2(n6461), .ZN(n5903) );
  INV_X1 U7435 ( .A(n5897), .ZN(n5901) );
  NAND2_X1 U7436 ( .A1(n5898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5899) );
  MUX2_X1 U7437 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5899), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5900) );
  NAND2_X1 U7438 ( .A1(n5901), .A2(n5900), .ZN(n6460) );
  OR2_X1 U7439 ( .A1(n5896), .A2(n6460), .ZN(n5902) );
  NAND2_X1 U7440 ( .A1(n5889), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5912) );
  INV_X1 U7441 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5905) );
  OR2_X1 U7442 ( .A1(n5869), .A2(n5905), .ZN(n5911) );
  NAND2_X1 U7443 ( .A1(n5906), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5907) );
  AND2_X1 U7444 ( .A1(n5924), .A2(n5907), .ZN(n7317) );
  OR2_X1 U7445 ( .A1(n6109), .A2(n7317), .ZN(n5910) );
  INV_X1 U7446 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5908) );
  OR2_X1 U7447 ( .A1(n5870), .A2(n5908), .ZN(n5909) );
  OR2_X1 U7448 ( .A1(n5897), .A2(n6200), .ZN(n5914) );
  XNOR2_X1 U7449 ( .A(n5914), .B(n5913), .ZN(n6462) );
  OR2_X1 U7450 ( .A1(n5865), .A2(n6475), .ZN(n5916) );
  OR2_X1 U7451 ( .A1(n5864), .A2(n6463), .ZN(n5915) );
  OAI211_X1 U7452 ( .C1(n5896), .C2(n6462), .A(n5916), .B(n5915), .ZN(n7052)
         );
  NOR2_X1 U7453 ( .A1(n8111), .A2(n7052), .ZN(n7045) );
  NAND2_X1 U7454 ( .A1(n8111), .A2(n7052), .ZN(n7043) );
  NOR2_X1 U7455 ( .A1(n5917), .A2(n6200), .ZN(n5918) );
  MUX2_X1 U7456 ( .A(n6200), .B(n5918), .S(P2_IR_REG_6__SCAN_IN), .Z(n5921) );
  INV_X1 U7457 ( .A(n5919), .ZN(n5920) );
  OR2_X1 U7458 ( .A1(n5865), .A2(n6467), .ZN(n5923) );
  INV_X1 U7459 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6468) );
  OR2_X1 U7460 ( .A1(n5864), .A2(n6468), .ZN(n5922) );
  OAI211_X1 U7461 ( .C1(n5896), .C2(n9756), .A(n5923), .B(n5922), .ZN(n7137)
         );
  NAND2_X1 U7462 ( .A1(n7129), .A2(n7137), .ZN(n5930) );
  NAND2_X1 U7463 ( .A1(n5889), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5929) );
  INV_X1 U7464 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6304) );
  OR2_X1 U7465 ( .A1(n5870), .A2(n6304), .ZN(n5928) );
  NAND2_X1 U7466 ( .A1(n5924), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5925) );
  AND2_X1 U7467 ( .A1(n5934), .A2(n5925), .ZN(n7135) );
  OR2_X1 U7468 ( .A1(n6109), .A2(n7135), .ZN(n5927) );
  INV_X1 U7469 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7134) );
  OR2_X1 U7470 ( .A1(n5869), .A2(n7134), .ZN(n5926) );
  NAND2_X1 U7471 ( .A1(n5930), .A2(n7273), .ZN(n5932) );
  NAND2_X1 U7472 ( .A1(n5932), .A2(n5931), .ZN(n7271) );
  NAND2_X1 U7473 ( .A1(n7894), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5939) );
  INV_X1 U7474 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5933) );
  OR2_X1 U7475 ( .A1(n6244), .A2(n5933), .ZN(n5938) );
  NAND2_X1 U7476 ( .A1(n5934), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5935) );
  AND2_X1 U7477 ( .A1(n5947), .A2(n5935), .ZN(n7274) );
  OR2_X1 U7478 ( .A1(n6109), .A2(n7274), .ZN(n5937) );
  OR2_X1 U7479 ( .A1(n5870), .A2(n9945), .ZN(n5936) );
  NAND4_X1 U7480 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n8109)
         );
  OR2_X1 U7481 ( .A1(n5865), .A2(n6478), .ZN(n5944) );
  OR2_X1 U7482 ( .A1(n5864), .A2(n10052), .ZN(n5943) );
  NAND2_X1 U7483 ( .A1(n5919), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5941) );
  INV_X1 U7484 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7485 ( .A(n5941), .B(n5940), .ZN(n6890) );
  OR2_X1 U7486 ( .A1(n5896), .A2(n6890), .ZN(n5942) );
  OR2_X1 U7487 ( .A1(n8109), .A2(n7275), .ZN(n7971) );
  NAND2_X1 U7488 ( .A1(n8109), .A2(n7275), .ZN(n7327) );
  NAND2_X1 U7489 ( .A1(n7971), .A2(n7327), .ZN(n7907) );
  INV_X1 U7490 ( .A(n7275), .ZN(n9917) );
  OR2_X1 U7491 ( .A1(n8109), .A2(n9917), .ZN(n5945) );
  NAND2_X1 U7492 ( .A1(n5889), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5953) );
  INV_X1 U7493 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5946) );
  OR2_X1 U7494 ( .A1(n5869), .A2(n5946), .ZN(n5952) );
  NAND2_X1 U7495 ( .A1(n5947), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5948) );
  AND2_X1 U7496 ( .A1(n5960), .A2(n5948), .ZN(n7371) );
  OR2_X1 U7497 ( .A1(n6109), .A2(n7371), .ZN(n5951) );
  INV_X1 U7498 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5949) );
  OR2_X1 U7499 ( .A1(n5870), .A2(n5949), .ZN(n5950) );
  NAND4_X1 U7500 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n8108)
         );
  OR2_X1 U7501 ( .A1(n5864), .A2(n6479), .ZN(n5956) );
  NAND2_X1 U7502 ( .A1(n4441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7503 ( .A(n5954), .B(n5799), .ZN(n9780) );
  OR2_X1 U7504 ( .A1(n5896), .A2(n9780), .ZN(n5955) );
  NAND2_X1 U7505 ( .A1(n8108), .A2(n9919), .ZN(n7979) );
  INV_X1 U7506 ( .A(n7918), .ZN(n5958) );
  INV_X1 U7507 ( .A(n9919), .ZN(n7368) );
  NAND2_X1 U7508 ( .A1(n8108), .A2(n7368), .ZN(n5959) );
  NAND2_X1 U7509 ( .A1(n7324), .A2(n5959), .ZN(n7385) );
  NAND2_X1 U7510 ( .A1(n5889), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5965) );
  INV_X1 U7511 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6303) );
  OR2_X1 U7512 ( .A1(n5869), .A2(n6303), .ZN(n5964) );
  NAND2_X1 U7513 ( .A1(n5960), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5961) );
  AND2_X1 U7514 ( .A1(n5972), .A2(n5961), .ZN(n7484) );
  OR2_X1 U7515 ( .A1(n6109), .A2(n7484), .ZN(n5963) );
  INV_X1 U7516 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6302) );
  OR2_X1 U7517 ( .A1(n5870), .A2(n6302), .ZN(n5962) );
  NAND4_X1 U7518 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n8107)
         );
  NAND2_X1 U7519 ( .A1(n5966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  XNOR2_X1 U7520 ( .A(n5967), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6403) );
  INV_X1 U7521 ( .A(n6403), .ZN(n9790) );
  OR2_X1 U7522 ( .A1(n5865), .A2(n6483), .ZN(n5969) );
  OR2_X1 U7523 ( .A1(n5864), .A2(n6482), .ZN(n5968) );
  OAI211_X1 U7524 ( .C1(n5896), .C2(n9790), .A(n5969), .B(n5968), .ZN(n7481)
         );
  OR2_X1 U7525 ( .A1(n8107), .A2(n7481), .ZN(n5970) );
  NAND2_X1 U7526 ( .A1(n7385), .A2(n5970), .ZN(n7409) );
  NAND2_X1 U7527 ( .A1(n7894), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5978) );
  INV_X1 U7528 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5971) );
  OR2_X1 U7529 ( .A1(n6244), .A2(n5971), .ZN(n5977) );
  NAND2_X1 U7530 ( .A1(n5972), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5973) );
  AND2_X1 U7531 ( .A1(n5988), .A2(n5973), .ZN(n7723) );
  OR2_X1 U7532 ( .A1(n6109), .A2(n7723), .ZN(n5976) );
  INV_X1 U7533 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5974) );
  OR2_X1 U7534 ( .A1(n5870), .A2(n5974), .ZN(n5975) );
  NOR2_X1 U7535 ( .A1(n5982), .A2(n6200), .ZN(n5979) );
  MUX2_X1 U7536 ( .A(n6200), .B(n5979), .S(P2_IR_REG_10__SCAN_IN), .Z(n5980)
         );
  INV_X1 U7537 ( .A(n5980), .ZN(n5983) );
  INV_X1 U7538 ( .A(n5996), .ZN(n6199) );
  NAND2_X1 U7539 ( .A1(n5983), .A2(n6199), .ZN(n7491) );
  INV_X1 U7540 ( .A(n7491), .ZN(n6326) );
  AOI22_X1 U7541 ( .A1(n7889), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6092), .B2(
        n6326), .ZN(n5985) );
  NAND2_X1 U7542 ( .A1(n6485), .A2(n7890), .ZN(n5984) );
  NAND2_X1 U7543 ( .A1(n5985), .A2(n5984), .ZN(n7730) );
  NAND2_X1 U7544 ( .A1(n8106), .A2(n7730), .ZN(n5986) );
  NAND2_X1 U7545 ( .A1(n8107), .A2(n7481), .ZN(n7408) );
  AND2_X1 U7546 ( .A1(n5986), .A2(n7408), .ZN(n5987) );
  AOI21_X2 U7547 ( .B1(n7409), .B2(n5987), .A(n4433), .ZN(n7373) );
  NAND2_X1 U7548 ( .A1(n5889), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5993) );
  INV_X1 U7549 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6301) );
  OR2_X1 U7550 ( .A1(n5869), .A2(n6301), .ZN(n5992) );
  NAND2_X1 U7551 ( .A1(n5988), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5989) );
  AND2_X1 U7552 ( .A1(n6004), .A2(n5989), .ZN(n7378) );
  OR2_X1 U7553 ( .A1(n6109), .A2(n7378), .ZN(n5991) );
  INV_X1 U7554 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6300) );
  OR2_X1 U7555 ( .A1(n5870), .A2(n6300), .ZN(n5990) );
  NAND2_X1 U7556 ( .A1(n6502), .A2(n7890), .ZN(n5999) );
  NOR2_X1 U7557 ( .A1(n5996), .A2(n6200), .ZN(n5994) );
  MUX2_X1 U7558 ( .A(n6200), .B(n5994), .S(P2_IR_REG_11__SCAN_IN), .Z(n5997)
         );
  NOR2_X1 U7559 ( .A1(n5997), .A2(n6013), .ZN(n6377) );
  AOI22_X1 U7560 ( .A1(n7889), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6092), .B2(
        n6377), .ZN(n5998) );
  NAND2_X1 U7561 ( .A1(n5999), .A2(n5998), .ZN(n7377) );
  OR2_X1 U7562 ( .A1(n7728), .A2(n7377), .ZN(n7992) );
  NAND2_X1 U7563 ( .A1(n7728), .A2(n7377), .ZN(n7994) );
  NAND2_X1 U7564 ( .A1(n7992), .A2(n7994), .ZN(n7923) );
  NAND2_X1 U7565 ( .A1(n7373), .A2(n7923), .ZN(n7372) );
  INV_X1 U7566 ( .A(n7728), .ZN(n8369) );
  NAND2_X1 U7567 ( .A1(n7377), .A2(n8369), .ZN(n6000) );
  NAND2_X1 U7568 ( .A1(n7372), .A2(n6000), .ZN(n8368) );
  NAND2_X1 U7569 ( .A1(n6505), .A2(n7890), .ZN(n6003) );
  OR2_X1 U7570 ( .A1(n6013), .A2(n6200), .ZN(n6001) );
  XNOR2_X1 U7571 ( .A(n6001), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7528) );
  AOI22_X1 U7572 ( .A1(n7889), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6092), .B2(
        n7528), .ZN(n6002) );
  NAND2_X1 U7573 ( .A1(n5889), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6009) );
  INV_X1 U7574 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8374) );
  OR2_X1 U7575 ( .A1(n5869), .A2(n8374), .ZN(n6008) );
  NAND2_X1 U7576 ( .A1(n6004), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6005) );
  AND2_X1 U7577 ( .A1(n6016), .A2(n6005), .ZN(n7755) );
  OR2_X1 U7578 ( .A1(n6109), .A2(n7755), .ZN(n6007) );
  INV_X1 U7579 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8431) );
  OR2_X1 U7580 ( .A1(n5870), .A2(n8431), .ZN(n6006) );
  NAND4_X1 U7581 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .ZN(n8105)
         );
  OR2_X1 U7582 ( .A1(n8533), .A2(n8105), .ZN(n6010) );
  NAND2_X1 U7583 ( .A1(n8533), .A2(n8105), .ZN(n6011) );
  NAND2_X1 U7584 ( .A1(n6522), .A2(n7890), .ZN(n6015) );
  NAND2_X1 U7585 ( .A1(n6053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6023) );
  XNOR2_X1 U7586 ( .A(n6023), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U7587 ( .A1(n7889), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6092), .B2(
        n9822), .ZN(n6014) );
  NAND2_X1 U7588 ( .A1(n6015), .A2(n6014), .ZN(n8526) );
  NAND2_X1 U7589 ( .A1(n5889), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6021) );
  INV_X1 U7590 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9821) );
  OR2_X1 U7591 ( .A1(n5870), .A2(n9821), .ZN(n6020) );
  NAND2_X1 U7592 ( .A1(n6016), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6017) );
  AND2_X1 U7593 ( .A1(n6029), .A2(n6017), .ZN(n8356) );
  OR2_X1 U7594 ( .A1(n6109), .A2(n8356), .ZN(n6019) );
  INV_X1 U7595 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8357) );
  OR2_X1 U7596 ( .A1(n5869), .A2(n8357), .ZN(n6018) );
  OR2_X1 U7597 ( .A1(n8526), .A2(n8332), .ZN(n8003) );
  NAND2_X1 U7598 ( .A1(n8526), .A2(n8332), .ZN(n8002) );
  INV_X1 U7599 ( .A(n8526), .ZN(n7816) );
  NAND2_X1 U7600 ( .A1(n7816), .A2(n8332), .ZN(n6022) );
  NAND2_X1 U7601 ( .A1(n8343), .A2(n6022), .ZN(n8328) );
  NAND2_X1 U7602 ( .A1(n6661), .A2(n7890), .ZN(n6028) );
  NAND2_X1 U7603 ( .A1(n6023), .A2(n6051), .ZN(n6024) );
  NAND2_X1 U7604 ( .A1(n6024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7605 ( .A1(n6025), .A2(n6050), .ZN(n6038) );
  OR2_X1 U7606 ( .A1(n6025), .A2(n6050), .ZN(n6026) );
  AOI22_X1 U7607 ( .A1(n7889), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6092), .B2(
        n8119), .ZN(n6027) );
  NAND2_X1 U7608 ( .A1(n5889), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6034) );
  INV_X1 U7609 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6383) );
  OR2_X1 U7610 ( .A1(n5869), .A2(n6383), .ZN(n6033) );
  NAND2_X1 U7611 ( .A1(n6029), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6030) );
  AND2_X1 U7612 ( .A1(n6042), .A2(n6030), .ZN(n8335) );
  OR2_X1 U7613 ( .A1(n6109), .A2(n8335), .ZN(n6032) );
  INV_X1 U7614 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8424) );
  OR2_X1 U7615 ( .A1(n5870), .A2(n8424), .ZN(n6031) );
  NAND4_X1 U7616 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n8104)
         );
  NAND2_X1 U7617 ( .A1(n8520), .A2(n8104), .ZN(n6035) );
  NAND2_X1 U7618 ( .A1(n8328), .A2(n6035), .ZN(n6037) );
  OR2_X1 U7619 ( .A1(n8520), .A2(n8104), .ZN(n6036) );
  NAND2_X1 U7620 ( .A1(n6037), .A2(n6036), .ZN(n8319) );
  NAND2_X1 U7621 ( .A1(n6690), .A2(n7890), .ZN(n6041) );
  NAND2_X1 U7622 ( .A1(n6038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6039) );
  XNOR2_X1 U7623 ( .A(n6039), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6413) );
  AOI22_X1 U7624 ( .A1(n7889), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6413), .B2(
        n6092), .ZN(n6040) );
  NAND2_X1 U7625 ( .A1(n5889), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6047) );
  INV_X1 U7626 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10055) );
  OR2_X1 U7627 ( .A1(n5870), .A2(n10055), .ZN(n6046) );
  NAND2_X1 U7628 ( .A1(n6042), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6043) );
  AND2_X1 U7629 ( .A1(n6058), .A2(n6043), .ZN(n7870) );
  OR2_X1 U7630 ( .A1(n6109), .A2(n7870), .ZN(n6045) );
  INV_X1 U7631 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8322) );
  OR2_X1 U7632 ( .A1(n5869), .A2(n8322), .ZN(n6044) );
  NAND4_X1 U7633 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n8330)
         );
  NOR2_X1 U7634 ( .A1(n8421), .A2(n8330), .ZN(n6048) );
  INV_X1 U7635 ( .A(n8421), .ZN(n8514) );
  NAND2_X1 U7636 ( .A1(n6795), .A2(n7890), .ZN(n6057) );
  NAND3_X1 U7637 ( .A1(n6051), .A2(n6050), .A3(n6049), .ZN(n6052) );
  INV_X1 U7638 ( .A(n6067), .ZN(n6054) );
  NAND2_X1 U7639 ( .A1(n6054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6055) );
  XNOR2_X1 U7640 ( .A(n6055), .B(P2_IR_REG_16__SCAN_IN), .ZN(n6416) );
  AOI22_X1 U7641 ( .A1(n7889), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6092), .B2(
        n6416), .ZN(n6056) );
  NAND2_X1 U7642 ( .A1(n5889), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6063) );
  INV_X1 U7643 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10125) );
  OR2_X1 U7644 ( .A1(n5869), .A2(n10125), .ZN(n6062) );
  NAND2_X1 U7645 ( .A1(n6058), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6059) );
  AND2_X1 U7646 ( .A1(n6080), .A2(n6059), .ZN(n8313) );
  OR2_X1 U7647 ( .A1(n6109), .A2(n8313), .ZN(n6061) );
  INV_X1 U7648 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8417) );
  OR2_X1 U7649 ( .A1(n5870), .A2(n8417), .ZN(n6060) );
  NAND2_X1 U7650 ( .A1(n8508), .A2(n8321), .ZN(n8015) );
  NAND2_X1 U7651 ( .A1(n8018), .A2(n8015), .ZN(n8307) );
  NAND2_X1 U7652 ( .A1(n8306), .A2(n8307), .ZN(n6065) );
  INV_X1 U7653 ( .A(n8321), .ZN(n8103) );
  NAND2_X1 U7654 ( .A1(n8508), .A2(n8103), .ZN(n6064) );
  NAND2_X1 U7655 ( .A1(n6065), .A2(n6064), .ZN(n8296) );
  NAND2_X1 U7656 ( .A1(n6862), .A2(n7890), .ZN(n6070) );
  NAND2_X1 U7657 ( .A1(n6067), .A2(n6066), .ZN(n6077) );
  NAND2_X1 U7658 ( .A1(n6077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6068) );
  XNOR2_X1 U7659 ( .A(n6068), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U7660 ( .A1(n7889), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6092), .B2(
        n9857), .ZN(n6069) );
  NAND2_X1 U7661 ( .A1(n5889), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6074) );
  INV_X1 U7662 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10211) );
  OR2_X1 U7663 ( .A1(n5869), .A2(n10211), .ZN(n6073) );
  INV_X1 U7664 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9877) );
  XNOR2_X1 U7665 ( .A(n6080), .B(n9877), .ZN(n7790) );
  OR2_X1 U7666 ( .A1(n6109), .A2(n7790), .ZN(n6072) );
  INV_X1 U7667 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10128) );
  OR2_X1 U7668 ( .A1(n5870), .A2(n10128), .ZN(n6071) );
  OR2_X1 U7669 ( .A1(n8502), .A2(n8310), .ZN(n8020) );
  NAND2_X1 U7670 ( .A1(n8502), .A2(n8310), .ZN(n8025) );
  NAND2_X1 U7671 ( .A1(n8020), .A2(n8025), .ZN(n7905) );
  NAND2_X1 U7672 ( .A1(n8296), .A2(n7905), .ZN(n6076) );
  NAND2_X1 U7673 ( .A1(n8502), .A2(n8102), .ZN(n6075) );
  NAND2_X1 U7674 ( .A1(n6076), .A2(n6075), .ZN(n8282) );
  NAND2_X1 U7675 ( .A1(n6916), .A2(n7890), .ZN(n6079) );
  XNOR2_X1 U7676 ( .A(n4409), .B(P2_IR_REG_18__SCAN_IN), .ZN(n6420) );
  AOI22_X1 U7677 ( .A1(n7889), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6420), .B2(
        n6092), .ZN(n6078) );
  NAND2_X1 U7678 ( .A1(n5889), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6085) );
  INV_X1 U7679 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8290) );
  OR2_X1 U7680 ( .A1(n5869), .A2(n8290), .ZN(n6084) );
  OAI21_X1 U7681 ( .B1(n6080), .B2(P2_REG3_REG_17__SCAN_IN), .A(
        P2_REG3_REG_18__SCAN_IN), .ZN(n6081) );
  AND2_X1 U7682 ( .A1(n6095), .A2(n6081), .ZN(n8289) );
  OR2_X1 U7683 ( .A1(n6109), .A2(n8289), .ZN(n6083) );
  INV_X1 U7684 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10222) );
  OR2_X1 U7685 ( .A1(n5870), .A2(n10222), .ZN(n6082) );
  NAND4_X1 U7686 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n8298)
         );
  AND2_X1 U7687 ( .A1(n8287), .A2(n8298), .ZN(n6087) );
  OR2_X1 U7688 ( .A1(n8287), .A2(n8298), .ZN(n6086) );
  OAI21_X1 U7689 ( .B1(n8282), .B2(n6087), .A(n6086), .ZN(n8271) );
  INV_X1 U7690 ( .A(n8271), .ZN(n6103) );
  NAND2_X1 U7691 ( .A1(n7616), .A2(n7890), .ZN(n6094) );
  NAND2_X1 U7692 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  AOI22_X1 U7693 ( .A1(n8090), .A2(n6092), .B1(n7889), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6093) );
  INV_X1 U7694 ( .A(n5870), .ZN(n6241) );
  NAND2_X1 U7695 ( .A1(n6241), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6101) );
  INV_X1 U7696 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10040) );
  OR2_X1 U7697 ( .A1(n6244), .A2(n10040), .ZN(n6100) );
  NAND2_X1 U7698 ( .A1(n6095), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6096) );
  AND2_X1 U7699 ( .A1(n6107), .A2(n6096), .ZN(n8277) );
  OR2_X1 U7700 ( .A1(n6109), .A2(n8277), .ZN(n6099) );
  INV_X1 U7701 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6097) );
  OR2_X1 U7702 ( .A1(n5869), .A2(n6097), .ZN(n6098) );
  NAND2_X1 U7703 ( .A1(n8279), .A2(n8284), .ZN(n8031) );
  NAND2_X1 U7704 ( .A1(n6103), .A2(n6102), .ZN(n8273) );
  NAND2_X1 U7705 ( .A1(n8279), .A2(n8262), .ZN(n6104) );
  NAND2_X1 U7706 ( .A1(n7204), .A2(n7890), .ZN(n6106) );
  INV_X1 U7707 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7205) );
  OR2_X1 U7708 ( .A1(n5864), .A2(n7205), .ZN(n6105) );
  NAND2_X1 U7709 ( .A1(n7894), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6113) );
  INV_X1 U7710 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8486) );
  OR2_X1 U7711 ( .A1(n6244), .A2(n8486), .ZN(n6112) );
  NAND2_X1 U7712 ( .A1(n6107), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6108) );
  AND2_X1 U7713 ( .A1(n6117), .A2(n6108), .ZN(n7807) );
  OR2_X1 U7714 ( .A1(n6109), .A2(n7807), .ZN(n6111) );
  INV_X1 U7715 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8406) );
  OR2_X1 U7716 ( .A1(n5870), .A2(n8406), .ZN(n6110) );
  NAND2_X1 U7717 ( .A1(n8487), .A2(n8252), .ZN(n8245) );
  NAND2_X1 U7718 ( .A1(n8035), .A2(n8245), .ZN(n8261) );
  INV_X1 U7719 ( .A(n8252), .ZN(n8274) );
  OR2_X1 U7720 ( .A1(n8487), .A2(n8274), .ZN(n6114) );
  NAND2_X1 U7721 ( .A1(n7292), .A2(n7890), .ZN(n6116) );
  OR2_X1 U7722 ( .A1(n5864), .A2(n10110), .ZN(n6115) );
  NAND2_X1 U7723 ( .A1(n6117), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7724 ( .A1(n6127), .A2(n6118), .ZN(n8253) );
  NAND2_X1 U7725 ( .A1(n6191), .A2(n8253), .ZN(n6122) );
  INV_X1 U7726 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n10083) );
  OR2_X1 U7727 ( .A1(n6244), .A2(n10083), .ZN(n6121) );
  INV_X1 U7728 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8255) );
  OR2_X1 U7729 ( .A1(n5869), .A2(n8255), .ZN(n6120) );
  INV_X1 U7730 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8404) );
  OR2_X1 U7731 ( .A1(n5870), .A2(n8404), .ZN(n6119) );
  NAND2_X1 U7732 ( .A1(n8403), .A2(n8237), .ZN(n8041) );
  NAND2_X1 U7733 ( .A1(n8040), .A2(n8041), .ZN(n8249) );
  OR2_X1 U7734 ( .A1(n8403), .A2(n8263), .ZN(n6123) );
  NAND2_X1 U7735 ( .A1(n6124), .A2(n6123), .ZN(n8233) );
  NAND2_X1 U7736 ( .A1(n7436), .A2(n7890), .ZN(n6126) );
  OR2_X1 U7737 ( .A1(n5864), .A2(n7437), .ZN(n6125) );
  NAND2_X1 U7738 ( .A1(n6127), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7739 ( .A1(n6136), .A2(n6128), .ZN(n8240) );
  NAND2_X1 U7740 ( .A1(n8240), .A2(n6191), .ZN(n6132) );
  NAND2_X1 U7741 ( .A1(n5889), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7742 ( .A1(n6241), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7743 ( .A1(n7894), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7744 ( .A1(n7822), .A2(n8251), .ZN(n8044) );
  NAND2_X1 U7745 ( .A1(n8045), .A2(n8044), .ZN(n8238) );
  INV_X1 U7746 ( .A(n8251), .ZN(n8227) );
  OR2_X1 U7747 ( .A1(n7822), .A2(n8227), .ZN(n6133) );
  NAND2_X1 U7748 ( .A1(n7509), .A2(n7890), .ZN(n6135) );
  OR2_X1 U7749 ( .A1(n5864), .A2(n7507), .ZN(n6134) );
  INV_X1 U7750 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U7751 ( .A1(n6136), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7752 ( .A1(n6146), .A2(n6137), .ZN(n8230) );
  NAND2_X1 U7753 ( .A1(n8230), .A2(n6191), .ZN(n6141) );
  NAND2_X1 U7754 ( .A1(n7894), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7755 ( .A1(n5889), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6138) );
  AND2_X1 U7756 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7757 ( .A1(n8474), .A2(n8215), .ZN(n6142) );
  NAND2_X1 U7758 ( .A1(n6143), .A2(n6142), .ZN(n8212) );
  NAND2_X1 U7759 ( .A1(n7563), .A2(n7890), .ZN(n6145) );
  OR2_X1 U7760 ( .A1(n5864), .A2(n7564), .ZN(n6144) );
  NAND2_X1 U7761 ( .A1(n6146), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7762 ( .A1(n6153), .A2(n6147), .ZN(n8217) );
  NAND2_X1 U7763 ( .A1(n8217), .A2(n6191), .ZN(n6150) );
  AOI22_X1 U7764 ( .A1(n7894), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n5889), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6149) );
  INV_X1 U7765 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8393) );
  OR2_X1 U7766 ( .A1(n5870), .A2(n8393), .ZN(n6148) );
  NAND2_X1 U7767 ( .A1(n8468), .A2(n7764), .ZN(n6227) );
  NAND2_X1 U7768 ( .A1(n8047), .A2(n6227), .ZN(n8210) );
  NAND2_X1 U7769 ( .A1(n7569), .A2(n7890), .ZN(n6152) );
  OR2_X1 U7770 ( .A1(n5864), .A2(n7570), .ZN(n6151) );
  NAND2_X1 U7771 ( .A1(n6153), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7772 ( .A1(n6162), .A2(n6154), .ZN(n8199) );
  NAND2_X1 U7773 ( .A1(n8199), .A2(n6191), .ZN(n6159) );
  INV_X1 U7774 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U7775 ( .A1(n7894), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7776 ( .A1(n5889), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6155) );
  OAI211_X1 U7777 ( .C1(n8390), .C2(n5870), .A(n6156), .B(n6155), .ZN(n6157)
         );
  INV_X1 U7778 ( .A(n6157), .ZN(n6158) );
  NOR2_X1 U7779 ( .A1(n8462), .A2(n8214), .ZN(n7904) );
  NAND2_X1 U7780 ( .A1(n7575), .A2(n7890), .ZN(n6161) );
  OR2_X1 U7781 ( .A1(n5864), .A2(n7576), .ZN(n6160) );
  NAND2_X1 U7782 ( .A1(n6162), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7783 ( .A1(n6175), .A2(n6163), .ZN(n8182) );
  NAND2_X1 U7784 ( .A1(n8182), .A2(n6191), .ZN(n6169) );
  INV_X1 U7785 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U7786 ( .A1(n5889), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6166) );
  INV_X1 U7787 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6164) );
  OR2_X1 U7788 ( .A1(n5869), .A2(n6164), .ZN(n6165) );
  OAI211_X1 U7789 ( .C1(n10130), .C2(n5870), .A(n6166), .B(n6165), .ZN(n6167)
         );
  INV_X1 U7790 ( .A(n6167), .ZN(n6168) );
  INV_X1 U7791 ( .A(n8456), .ZN(n7865) );
  INV_X1 U7792 ( .A(n8172), .ZN(n6184) );
  NAND2_X1 U7793 ( .A1(n7580), .A2(n7890), .ZN(n6174) );
  OR2_X1 U7794 ( .A1(n5864), .A2(n10163), .ZN(n6173) );
  NAND2_X1 U7795 ( .A1(n6175), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7796 ( .A1(n6177), .A2(n6176), .ZN(n8177) );
  NAND2_X1 U7797 ( .A1(n8177), .A2(n6191), .ZN(n6182) );
  INV_X1 U7798 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10224) );
  NAND2_X1 U7799 ( .A1(n5889), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6179) );
  INV_X1 U7800 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8176) );
  OR2_X1 U7801 ( .A1(n5869), .A2(n8176), .ZN(n6178) );
  OAI211_X1 U7802 ( .C1(n10224), .C2(n5870), .A(n6179), .B(n6178), .ZN(n6180)
         );
  INV_X1 U7803 ( .A(n6180), .ZN(n6181) );
  NAND2_X2 U7804 ( .A1(n6182), .A2(n6181), .ZN(n8185) );
  INV_X1 U7805 ( .A(n8450), .ZN(n7707) );
  AOI21_X2 U7806 ( .B1(n6184), .B2(n6183), .A(n5029), .ZN(n8166) );
  OAI21_X1 U7807 ( .B1(n8174), .B2(n8444), .A(n8166), .ZN(n6186) );
  INV_X1 U7808 ( .A(n8174), .ZN(n7703) );
  NAND2_X1 U7809 ( .A1(n8444), .A2(n8174), .ZN(n6185) );
  NAND2_X1 U7810 ( .A1(n6186), .A2(n6185), .ZN(n6197) );
  INV_X1 U7811 ( .A(SI_28_), .ZN(n6188) );
  INV_X1 U7812 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7684) );
  INV_X1 U7813 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8806) );
  MUX2_X1 U7814 ( .A(n7684), .B(n8806), .S(n4660), .Z(n7689) );
  OR2_X1 U7815 ( .A1(n5864), .A2(n7684), .ZN(n6190) );
  INV_X1 U7816 ( .A(n8150), .ZN(n6192) );
  NAND2_X1 U7817 ( .A1(n6192), .A2(n6191), .ZN(n7896) );
  INV_X1 U7818 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U7819 ( .A1(n7894), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7820 ( .A1(n6241), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7821 ( .C1(n6244), .C2(n10093), .A(n6194), .B(n6193), .ZN(n6195)
         );
  INV_X1 U7822 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U7823 ( .A1(n6293), .A2(n8101), .ZN(n7892) );
  XNOR2_X1 U7824 ( .A(n6197), .B(n8073), .ZN(n6213) );
  NAND2_X1 U7825 ( .A1(n6201), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n6204) );
  INV_X1 U7826 ( .A(n6201), .ZN(n6203) );
  INV_X1 U7827 ( .A(n8092), .ZN(n6266) );
  NAND2_X1 U7828 ( .A1(n8090), .A2(n6266), .ZN(n6425) );
  NAND2_X1 U7829 ( .A1(n6208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7830 ( .A1(n4512), .A2(n6729), .ZN(n6211) );
  NAND2_X1 U7831 ( .A1(n6213), .A2(n6212), .ZN(n6250) );
  OR2_X1 U7832 ( .A1(n6214), .A2(n7291), .ZN(n7914) );
  INV_X1 U7833 ( .A(n7914), .ZN(n6215) );
  NAND2_X1 U7834 ( .A1(n6215), .A2(n7912), .ZN(n6837) );
  NAND2_X1 U7835 ( .A1(n6837), .A2(n7945), .ZN(n6897) );
  XNOR2_X1 U7836 ( .A(n8112), .B(n9896), .ZN(n9887) );
  NAND2_X1 U7837 ( .A1(n9888), .A2(n9887), .ZN(n6216) );
  INV_X1 U7838 ( .A(n9896), .ZN(n7939) );
  OR2_X1 U7839 ( .A1(n8112), .A2(n7939), .ZN(n7953) );
  NAND2_X1 U7840 ( .A1(n6216), .A2(n7953), .ZN(n6928) );
  NAND2_X1 U7841 ( .A1(n9885), .A2(n9901), .ZN(n7957) );
  OR2_X1 U7842 ( .A1(n9885), .A2(n9901), .ZN(n7964) );
  INV_X1 U7843 ( .A(n7052), .ZN(n7318) );
  NOR2_X1 U7844 ( .A1(n8111), .A2(n7318), .ZN(n7963) );
  INV_X1 U7845 ( .A(n7963), .ZN(n6217) );
  NAND2_X1 U7846 ( .A1(n8111), .A2(n7318), .ZN(n7954) );
  NAND2_X1 U7847 ( .A1(n6218), .A2(n7954), .ZN(n7128) );
  INV_X1 U7848 ( .A(n7128), .ZN(n6221) );
  INV_X1 U7849 ( .A(n7137), .ZN(n9906) );
  AND2_X1 U7850 ( .A1(n8110), .A2(n9906), .ZN(n7955) );
  OR2_X1 U7851 ( .A1(n8110), .A2(n9906), .ZN(n7959) );
  INV_X1 U7852 ( .A(n7481), .ZN(n9924) );
  OR2_X1 U7853 ( .A1(n8107), .A2(n9924), .ZN(n7985) );
  NAND2_X1 U7854 ( .A1(n8107), .A2(n9924), .ZN(n7980) );
  NAND2_X1 U7855 ( .A1(n8106), .A2(n9929), .ZN(n7991) );
  AND2_X1 U7856 ( .A1(n7980), .A2(n7991), .ZN(n7986) );
  INV_X1 U7857 ( .A(n7923), .ZN(n7638) );
  NAND2_X1 U7858 ( .A1(n8533), .A2(n8350), .ZN(n7998) );
  NAND2_X1 U7859 ( .A1(n7999), .A2(n7998), .ZN(n8362) );
  INV_X1 U7860 ( .A(n7994), .ZN(n8363) );
  NOR2_X1 U7861 ( .A1(n8362), .A2(n8363), .ZN(n6222) );
  NOR2_X1 U7862 ( .A1(n8520), .A2(n8348), .ZN(n8006) );
  NAND2_X1 U7863 ( .A1(n8520), .A2(n8348), .ZN(n7927) );
  OR2_X1 U7864 ( .A1(n8421), .A2(n7926), .ZN(n8011) );
  NAND2_X1 U7865 ( .A1(n8317), .A2(n8011), .ZN(n6223) );
  NAND2_X1 U7866 ( .A1(n8421), .A2(n7926), .ZN(n8013) );
  NAND2_X1 U7867 ( .A1(n6223), .A2(n8013), .ZN(n8305) );
  INV_X1 U7868 ( .A(n8015), .ZN(n8021) );
  NAND2_X1 U7869 ( .A1(n6224), .A2(n8018), .ZN(n8295) );
  NAND2_X1 U7870 ( .A1(n8287), .A2(n7736), .ZN(n8026) );
  NAND2_X1 U7871 ( .A1(n8027), .A2(n8026), .ZN(n8285) );
  NAND2_X1 U7872 ( .A1(n8269), .A2(n8028), .ZN(n6225) );
  AND2_X1 U7873 ( .A1(n8041), .A2(n8245), .ZN(n8036) );
  NAND2_X1 U7874 ( .A1(n8239), .A2(n8044), .ZN(n6226) );
  NAND2_X1 U7875 ( .A1(n6226), .A2(n8045), .ZN(n8206) );
  NAND2_X1 U7876 ( .A1(n8474), .A2(n8236), .ZN(n8208) );
  NAND2_X1 U7877 ( .A1(n8206), .A2(n6228), .ZN(n6231) );
  INV_X1 U7878 ( .A(n6228), .ZN(n8048) );
  NOR2_X1 U7879 ( .A1(n8462), .A2(n8187), .ZN(n6232) );
  NAND2_X1 U7880 ( .A1(n8462), .A2(n8187), .ZN(n6233) );
  NAND2_X1 U7881 ( .A1(n6235), .A2(n8061), .ZN(n8171) );
  NAND2_X1 U7882 ( .A1(n8450), .A2(n7861), .ZN(n7903) );
  NOR2_X1 U7883 ( .A1(n8450), .A2(n7861), .ZN(n8067) );
  NAND2_X1 U7884 ( .A1(n8444), .A2(n7703), .ZN(n6236) );
  INV_X1 U7885 ( .A(n8068), .ZN(n8073) );
  AND2_X1 U7886 ( .A1(n6720), .A2(n9933), .ZN(n7286) );
  OAI21_X1 U7887 ( .B1(n8090), .B2(n8092), .A(n6728), .ZN(n6238) );
  INV_X1 U7888 ( .A(n8544), .ZN(n6352) );
  NAND2_X1 U7889 ( .A1(n6352), .A2(n8548), .ZN(n8095) );
  INV_X1 U7890 ( .A(n8548), .ZN(n9462) );
  NAND2_X1 U7891 ( .A1(n8544), .A2(n9462), .ZN(n6351) );
  INV_X1 U7892 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U7893 ( .A1(n7894), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7894 ( .A1(n6241), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6242) );
  OAI211_X1 U7895 ( .C1(n6244), .C2(n10174), .A(n6243), .B(n6242), .ZN(n6245)
         );
  INV_X1 U7896 ( .A(n6245), .ZN(n6246) );
  AND2_X1 U7897 ( .A1(n7896), .A2(n6246), .ZN(n7900) );
  NAND2_X1 U7898 ( .A1(n5896), .A2(P2_B_REG_SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7899 ( .A1(n8370), .A2(n6247), .ZN(n8148) );
  OAI22_X1 U7900 ( .A1(n7703), .A2(n8351), .B1(n7900), .B2(n8148), .ZN(n6248)
         );
  AOI21_X1 U7901 ( .B1(n8155), .B2(n6927), .A(n6248), .ZN(n6249) );
  NOR2_X1 U7902 ( .A1(n8156), .A2(n6251), .ZN(n6424) );
  NAND2_X1 U7903 ( .A1(n6821), .A2(n7913), .ZN(n6715) );
  MUX2_X1 U7904 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6253), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n6255) );
  NAND2_X1 U7905 ( .A1(n6255), .A2(n6254), .ZN(n7565) );
  XNOR2_X1 U7906 ( .A(n7565), .B(P2_B_REG_SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7907 ( .A1(n6254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6257) );
  NOR2_X1 U7908 ( .A1(n6259), .A2(n5813), .ZN(n6262) );
  INV_X1 U7909 ( .A(n6262), .ZN(n6261) );
  NAND2_X1 U7910 ( .A1(n6261), .A2(n6260), .ZN(n6264) );
  NAND2_X1 U7911 ( .A1(n6262), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6263) );
  INV_X1 U7912 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U7913 ( .A1(n6275), .A2(n10228), .ZN(n6265) );
  NAND2_X1 U7914 ( .A1(n4527), .A2(n7565), .ZN(n6489) );
  NAND2_X1 U7915 ( .A1(n6715), .A2(n6726), .ZN(n6268) );
  NAND3_X1 U7916 ( .A1(n6237), .A2(n6266), .A3(n6729), .ZN(n6267) );
  NAND2_X1 U7917 ( .A1(n6268), .A2(n6922), .ZN(n6292) );
  NAND2_X1 U7918 ( .A1(n6728), .A2(n8083), .ZN(n6704) );
  NAND2_X1 U7919 ( .A1(n7505), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6487) );
  INV_X1 U7920 ( .A(n7565), .ZN(n6273) );
  INV_X1 U7921 ( .A(n7571), .ZN(n6272) );
  INV_X1 U7922 ( .A(n6275), .ZN(n6488) );
  NOR2_X1 U7923 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .ZN(
        n6279) );
  NOR4_X1 U7924 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6278) );
  NOR4_X1 U7925 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6277) );
  NOR4_X1 U7926 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6276) );
  NAND4_X1 U7927 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n6285)
         );
  NOR4_X1 U7928 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6283) );
  NOR4_X1 U7929 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6282) );
  NOR4_X1 U7930 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6281) );
  NOR4_X1 U7931 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6280) );
  NAND4_X1 U7932 ( .A1(n6283), .A2(n6282), .A3(n6281), .A4(n6280), .ZN(n6284)
         );
  NOR2_X1 U7933 ( .A1(n6285), .A2(n6284), .ZN(n6286) );
  NOR2_X1 U7934 ( .A1(n6714), .A2(n6702), .ZN(n6428) );
  AND2_X1 U7935 ( .A1(n6704), .A2(n6428), .ZN(n6926) );
  INV_X1 U7936 ( .A(n6922), .ZN(n6289) );
  INV_X1 U7937 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U7938 ( .A1(n6275), .A2(n6496), .ZN(n6288) );
  NAND2_X1 U7939 ( .A1(n4527), .A2(n7571), .ZN(n6287) );
  AOI21_X1 U7940 ( .B1(n6289), .B2(n6920), .A(n6699), .ZN(n6290) );
  NAND2_X1 U7941 ( .A1(n6296), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6294) );
  INV_X1 U7942 ( .A(n6297), .ZN(n6703) );
  NAND2_X1 U7943 ( .A1(n6703), .A2(n8078), .ZN(n6298) );
  NAND2_X1 U7944 ( .A1(n6298), .A2(n7505), .ZN(n6350) );
  NAND2_X1 U7945 ( .A1(n6350), .A2(n5896), .ZN(n6299) );
  NAND2_X1 U7946 ( .A1(n6299), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  MUX2_X1 U7947 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8548), .Z(n6346) );
  XNOR2_X1 U7948 ( .A(n9857), .B(n6346), .ZN(n9866) );
  MUX2_X1 U7949 ( .A(n10125), .B(n8417), .S(n8548), .Z(n6344) );
  NOR2_X1 U7950 ( .A1(n6344), .A2(n6416), .ZN(n8132) );
  INV_X1 U7951 ( .A(n6413), .ZN(n9840) );
  MUX2_X1 U7952 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8548), .Z(n6341) );
  NOR2_X1 U7953 ( .A1(n9840), .A2(n6341), .ZN(n6343) );
  MUX2_X1 U7954 ( .A(n6383), .B(n8424), .S(n8548), .Z(n6339) );
  AND2_X1 U7955 ( .A1(n6339), .A2(n8119), .ZN(n6340) );
  MUX2_X1 U7956 ( .A(n8357), .B(n9821), .S(n8548), .Z(n6336) );
  AND2_X1 U7957 ( .A1(n6336), .A2(n9822), .ZN(n6337) );
  MUX2_X1 U7958 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8548), .Z(n6331) );
  NAND2_X1 U7959 ( .A1(n6331), .A2(n6507), .ZN(n6334) );
  MUX2_X1 U7960 ( .A(n6301), .B(n6300), .S(n8548), .Z(n6328) );
  NAND2_X1 U7961 ( .A1(n6328), .A2(n6377), .ZN(n6330) );
  INV_X1 U7962 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U7963 ( .A(n10124), .B(n5974), .S(n8548), .Z(n6325) );
  AND2_X1 U7964 ( .A1(n6325), .A2(n6326), .ZN(n6327) );
  MUX2_X1 U7965 ( .A(n6303), .B(n6302), .S(n8548), .Z(n6322) );
  AND2_X1 U7966 ( .A1(n6322), .A2(n6403), .ZN(n6323) );
  MUX2_X1 U7967 ( .A(n5946), .B(n5949), .S(n8548), .Z(n6319) );
  AND2_X1 U7968 ( .A1(n6319), .A2(n4727), .ZN(n6320) );
  MUX2_X1 U7969 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8548), .Z(n6316) );
  XOR2_X1 U7970 ( .A(n6890), .B(n6316), .Z(n6889) );
  MUX2_X1 U7971 ( .A(n7134), .B(n6304), .S(n8548), .Z(n6306) );
  INV_X1 U7972 ( .A(n9756), .ZN(n6305) );
  NAND2_X1 U7973 ( .A1(n6306), .A2(n6305), .ZN(n6315) );
  OAI21_X1 U7974 ( .B1(n6306), .B2(n6305), .A(n6315), .ZN(n9758) );
  MUX2_X1 U7975 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8548), .Z(n6312) );
  INV_X1 U7976 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6393) );
  MUX2_X1 U7977 ( .A(n9706), .B(n6393), .S(n8548), .Z(n6307) );
  XNOR2_X1 U7978 ( .A(n6307), .B(n9703), .ZN(n9713) );
  INV_X1 U7979 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6391) );
  MUX2_X1 U7980 ( .A(n7288), .B(n6391), .S(n8548), .Z(n6525) );
  NAND2_X1 U7981 ( .A1(n6525), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9714) );
  INV_X1 U7982 ( .A(n6307), .ZN(n6308) );
  AOI22_X1 U7983 ( .A1(n9713), .A2(n9714), .B1(n9703), .B2(n6308), .ZN(n6603)
         );
  MUX2_X1 U7984 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8548), .Z(n6309) );
  XNOR2_X1 U7985 ( .A(n6309), .B(n6454), .ZN(n6602) );
  INV_X1 U7986 ( .A(n6454), .ZN(n6611) );
  INV_X1 U7987 ( .A(n6309), .ZN(n6310) );
  OAI22_X1 U7988 ( .A1(n6603), .A2(n6602), .B1(n6611), .B2(n6310), .ZN(n9727)
         );
  MUX2_X1 U7989 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8548), .Z(n6311) );
  XNOR2_X1 U7990 ( .A(n6311), .B(n9724), .ZN(n9728) );
  NOR2_X1 U7991 ( .A1(n6311), .A2(n9724), .ZN(n6749) );
  XNOR2_X1 U7992 ( .A(n6312), .B(n6460), .ZN(n6752) );
  NOR3_X1 U7993 ( .A1(n9726), .A2(n6749), .A3(n6752), .ZN(n6750) );
  AOI21_X1 U7994 ( .B1(n6312), .B2(n6460), .A(n6750), .ZN(n9744) );
  MUX2_X1 U7995 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8548), .Z(n6313) );
  XNOR2_X1 U7996 ( .A(n6313), .B(n6462), .ZN(n9745) );
  INV_X1 U7997 ( .A(n6313), .ZN(n6314) );
  OAI22_X1 U7998 ( .A1(n9744), .A2(n9745), .B1(n4855), .B2(n6314), .ZN(n9759)
         );
  NAND2_X1 U7999 ( .A1(n6889), .A2(n6888), .ZN(n6887) );
  OAI21_X1 U8000 ( .B1(n6316), .B2(n6890), .A(n6887), .ZN(n6317) );
  INV_X1 U8001 ( .A(n6320), .ZN(n6318) );
  OAI21_X1 U8002 ( .B1(n4727), .B2(n6319), .A(n6318), .ZN(n9774) );
  INV_X1 U8003 ( .A(n6323), .ZN(n6321) );
  OAI21_X1 U8004 ( .B1(n6403), .B2(n6322), .A(n6321), .ZN(n9795) );
  NOR2_X1 U8005 ( .A1(n9794), .A2(n9795), .ZN(n9793) );
  NOR2_X1 U8006 ( .A1(n6323), .A2(n9793), .ZN(n7493) );
  INV_X1 U8007 ( .A(n6327), .ZN(n6324) );
  OAI21_X1 U8008 ( .B1(n6326), .B2(n6325), .A(n6324), .ZN(n7494) );
  NOR2_X1 U8009 ( .A1(n6327), .A2(n7492), .ZN(n9810) );
  OAI21_X1 U8010 ( .B1(n6328), .B2(n6377), .A(n6330), .ZN(n9811) );
  NOR2_X1 U8011 ( .A1(n9810), .A2(n9811), .ZN(n9809) );
  INV_X1 U8012 ( .A(n9809), .ZN(n6329) );
  NAND2_X1 U8013 ( .A1(n6330), .A2(n6329), .ZN(n7532) );
  INV_X1 U8014 ( .A(n7532), .ZN(n6332) );
  XNOR2_X1 U8015 ( .A(n6331), .B(n7528), .ZN(n7533) );
  NAND2_X1 U8016 ( .A1(n6332), .A2(n7533), .ZN(n6333) );
  NAND2_X1 U8017 ( .A1(n6334), .A2(n6333), .ZN(n9828) );
  INV_X1 U8018 ( .A(n6337), .ZN(n6335) );
  OAI21_X1 U8019 ( .B1(n9822), .B2(n6336), .A(n6335), .ZN(n9829) );
  NOR2_X1 U8020 ( .A1(n6337), .A2(n9827), .ZN(n8117) );
  INV_X1 U8021 ( .A(n6340), .ZN(n6338) );
  OAI21_X1 U8022 ( .B1(n8119), .B2(n6339), .A(n6338), .ZN(n8118) );
  NOR2_X1 U8023 ( .A1(n6340), .A2(n8116), .ZN(n9845) );
  AOI21_X1 U8024 ( .B1(n6341), .B2(n9840), .A(n6343), .ZN(n6342) );
  INV_X1 U8025 ( .A(n6342), .ZN(n9846) );
  NOR2_X1 U8026 ( .A1(n9845), .A2(n9846), .ZN(n9844) );
  NOR2_X1 U8027 ( .A1(n6343), .A2(n9844), .ZN(n8134) );
  AND2_X1 U8028 ( .A1(n6344), .A2(n6416), .ZN(n8133) );
  INV_X1 U8029 ( .A(n8133), .ZN(n6345) );
  NAND2_X1 U8030 ( .A1(n9866), .A2(n9867), .ZN(n9865) );
  OAI21_X1 U8031 ( .B1(n6864), .B2(n6346), .A(n9865), .ZN(n6348) );
  MUX2_X1 U8032 ( .A(n8290), .B(n10222), .S(n8548), .Z(n6347) );
  NOR2_X1 U8033 ( .A1(n6348), .A2(n6347), .ZN(n9461) );
  NAND2_X1 U8034 ( .A1(n6348), .A2(n6347), .ZN(n9459) );
  INV_X1 U8035 ( .A(n9459), .ZN(n6349) );
  NOR2_X1 U8036 ( .A1(n9461), .A2(n6349), .ZN(n6356) );
  INV_X1 U8037 ( .A(n6356), .ZN(n6355) );
  NAND2_X1 U8038 ( .A1(n6350), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6360) );
  OR2_X1 U8039 ( .A1(n6360), .A2(n6351), .ZN(n6354) );
  NAND2_X1 U8040 ( .A1(P2_U3893), .A2(n6352), .ZN(n6353) );
  OAI21_X1 U8041 ( .B1(n6355), .B2(n8113), .A(n9841), .ZN(n6358) );
  NOR2_X1 U8042 ( .A1(n6356), .A2(n9847), .ZN(n6357) );
  INV_X1 U8043 ( .A(n6420), .ZN(n9460) );
  INV_X1 U8044 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7845) );
  INV_X1 U8045 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9452) );
  NOR2_X1 U8046 ( .A1(n6360), .A2(n8544), .ZN(n6527) );
  INV_X1 U8047 ( .A(n6527), .ZN(n6361) );
  NAND2_X1 U8048 ( .A1(n9756), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6369) );
  NOR2_X1 U8049 ( .A1(n7288), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8050 ( .A1(n5845), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U8051 ( .B1(n9703), .B2(n6362), .A(n6363), .ZN(n9707) );
  NAND2_X1 U8052 ( .A1(n9709), .A2(n6363), .ZN(n6613) );
  XNOR2_X1 U8053 ( .A(n6454), .B(n7267), .ZN(n6614) );
  NAND2_X1 U8054 ( .A1(n6613), .A2(n6614), .ZN(n6612) );
  NAND2_X1 U8055 ( .A1(n6454), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8056 ( .A1(n6612), .A2(n6364), .ZN(n6365) );
  NAND2_X1 U8057 ( .A1(n6365), .A2(n9724), .ZN(n6759) );
  INV_X1 U8058 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10188) );
  MUX2_X1 U8059 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10188), .S(n6460), .Z(n6758)
         );
  NAND2_X1 U8060 ( .A1(n6460), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8061 ( .A1(n6762), .A2(n6366), .ZN(n6367) );
  OAI21_X1 U8062 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9756), .A(n6369), .ZN(
        n9761) );
  INV_X1 U8063 ( .A(n9760), .ZN(n6368) );
  NAND2_X1 U8064 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n9780), .ZN(n6372) );
  OAI21_X1 U8065 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9780), .A(n6372), .ZN(
        n9778) );
  NOR2_X1 U8066 ( .A1(n6403), .A2(n6373), .ZN(n6374) );
  XNOR2_X1 U8067 ( .A(n6373), .B(n6403), .ZN(n9792) );
  NOR2_X1 U8068 ( .A1(n6303), .A2(n9792), .ZN(n9791) );
  NOR2_X1 U8069 ( .A1(n6374), .A2(n9791), .ZN(n7487) );
  NAND2_X1 U8070 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7491), .ZN(n6375) );
  OAI21_X1 U8071 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7491), .A(n6375), .ZN(
        n7486) );
  NOR2_X1 U8072 ( .A1(n7487), .A2(n7486), .ZN(n7485) );
  AND2_X1 U8073 ( .A1(n7491), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6376) );
  INV_X1 U8074 ( .A(n6377), .ZN(n9806) );
  NAND2_X1 U8075 ( .A1(n6379), .A2(n9806), .ZN(n6378) );
  INV_X1 U8076 ( .A(n6378), .ZN(n6380) );
  NOR2_X1 U8077 ( .A1(n6301), .A2(n9808), .ZN(n9807) );
  AOI22_X1 U8078 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7528), .B1(n6507), .B2(
        n8374), .ZN(n7522) );
  NOR2_X1 U8079 ( .A1(n7523), .A2(n7522), .ZN(n7521) );
  NOR2_X1 U8080 ( .A1(n9822), .A2(n6381), .ZN(n6382) );
  AOI22_X1 U8081 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8119), .B1(n6662), .B2(
        n6383), .ZN(n8115) );
  NOR2_X1 U8082 ( .A1(n6413), .A2(n6384), .ZN(n6385) );
  INV_X1 U8083 ( .A(n6416), .ZN(n8138) );
  AOI22_X1 U8084 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n6416), .B1(n8138), .B2(
        n10125), .ZN(n8131) );
  NOR2_X1 U8085 ( .A1(n6416), .A2(n10125), .ZN(n6386) );
  NAND2_X1 U8086 ( .A1(n6388), .A2(n6864), .ZN(n6387) );
  OAI21_X1 U8087 ( .B1(n6388), .B2(n6864), .A(n6387), .ZN(n9861) );
  OR2_X1 U8088 ( .A1(n6420), .A2(n8290), .ZN(n9471) );
  NAND2_X1 U8089 ( .A1(n6420), .A2(n8290), .ZN(n6389) );
  NAND2_X1 U8090 ( .A1(n9471), .A2(n6389), .ZN(n6390) );
  AOI21_X1 U8091 ( .B1(n4479), .B2(n6390), .A(n9470), .ZN(n6423) );
  INV_X1 U8092 ( .A(n6460), .ZN(n6764) );
  NOR2_X1 U8093 ( .A1(n6391), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8094 ( .A1(n5845), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8095 ( .A1(n6395), .A2(n6394), .ZN(n6606) );
  XNOR2_X1 U8096 ( .A(n6454), .B(n10092), .ZN(n6605) );
  NAND2_X1 U8097 ( .A1(n6454), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6396) );
  MUX2_X1 U8098 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6398), .S(n6460), .Z(n6754)
         );
  NAND2_X1 U8099 ( .A1(n9756), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6399) );
  OAI21_X1 U8100 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n9756), .A(n6399), .ZN(
        n9754) );
  INV_X1 U8101 ( .A(n6399), .ZN(n6400) );
  INV_X1 U8102 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9945) );
  NAND2_X1 U8103 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n9780), .ZN(n6402) );
  OAI21_X1 U8104 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n9780), .A(n6402), .ZN(
        n9771) );
  NOR2_X1 U8105 ( .A1(n6403), .A2(n6404), .ZN(n6405) );
  NAND2_X1 U8106 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7491), .ZN(n6406) );
  OAI21_X1 U8107 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7491), .A(n6406), .ZN(
        n7489) );
  AND2_X1 U8108 ( .A1(n7491), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8109 ( .A1(n6409), .A2(n9806), .ZN(n6408) );
  INV_X1 U8110 ( .A(n6408), .ZN(n6410) );
  OAI21_X1 U8111 ( .B1(n6409), .B2(n9806), .A(n6408), .ZN(n9804) );
  AOI22_X1 U8112 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7528), .B1(n6507), .B2(
        n8431), .ZN(n7526) );
  NOR2_X1 U8113 ( .A1(n9822), .A2(n6411), .ZN(n6412) );
  AOI22_X1 U8114 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8119), .B1(n6662), .B2(
        n8424), .ZN(n8124) );
  NOR2_X1 U8115 ( .A1(n6413), .A2(n6414), .ZN(n6415) );
  XNOR2_X1 U8116 ( .A(n6414), .B(n6413), .ZN(n9837) );
  NOR2_X1 U8117 ( .A1(n10055), .A2(n9837), .ZN(n9836) );
  AOI22_X1 U8118 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n6416), .B1(n8138), .B2(
        n8417), .ZN(n8140) );
  INV_X1 U8119 ( .A(n6417), .ZN(n6419) );
  OAI21_X1 U8120 ( .B1(n6418), .B2(n6864), .A(n6417), .ZN(n9860) );
  NOR2_X1 U8121 ( .A1(n6419), .A2(n9859), .ZN(n6422) );
  OR2_X1 U8122 ( .A1(n6420), .A2(n10222), .ZN(n9455) );
  OAI21_X1 U8123 ( .B1(n9460), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9455), .ZN(
        n6421) );
  NOR2_X1 U8124 ( .A1(n6421), .A2(n6422), .ZN(n9457) );
  AND2_X1 U8125 ( .A1(n8078), .A2(n9933), .ZN(n6426) );
  NAND2_X1 U8126 ( .A1(n6741), .A2(n6426), .ZN(n6738) );
  NAND2_X1 U8127 ( .A1(n6738), .A2(n8336), .ZN(n6700) );
  NOR2_X1 U8128 ( .A1(n6726), .A2(n6702), .ZN(n6427) );
  INV_X1 U8129 ( .A(n6714), .ZN(n6709) );
  NAND2_X1 U8130 ( .A1(n6700), .A2(n6743), .ZN(n6431) );
  NAND2_X1 U8131 ( .A1(n6720), .A2(n6741), .ZN(n6429) );
  NAND2_X1 U8132 ( .A1(n6739), .A2(n6429), .ZN(n6430) );
  OAI21_X1 U8133 ( .B1(n6424), .B2(n9941), .A(n5032), .ZN(P2_U3456) );
  NOR2_X1 U8134 ( .A1(n6433), .A2(P1_U3086), .ZN(n6434) );
  NAND2_X1 U8135 ( .A1(n9307), .A2(n8970), .ZN(n6439) );
  INV_X1 U8136 ( .A(n6439), .ZN(n6438) );
  NAND2_X1 U8137 ( .A1(n8904), .A2(n6435), .ZN(n6436) );
  AND2_X1 U8138 ( .A1(n6437), .A2(n6436), .ZN(n6440) );
  INV_X1 U8139 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9417) );
  NOR2_X1 U8140 ( .A1(n9026), .A2(n9417), .ZN(n6453) );
  INV_X1 U8141 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7012) );
  MUX2_X1 U8142 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7012), .S(n6549), .Z(n6443)
         );
  NAND2_X1 U8143 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n8994) );
  INV_X1 U8144 ( .A(n8994), .ZN(n6442) );
  NAND2_X1 U8145 ( .A1(n6440), .A2(n6439), .ZN(n6450) );
  OR2_X1 U8146 ( .A1(n5160), .A2(n8992), .ZN(n6441) );
  OR2_X1 U8147 ( .A1(n6450), .A2(n6441), .ZN(n7300) );
  NAND2_X1 U8148 ( .A1(n6443), .A2(n6442), .ZN(n6533) );
  OAI211_X1 U8149 ( .C1(n6443), .C2(n6442), .A(n9075), .B(n6533), .ZN(n6448)
         );
  AND2_X1 U8150 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6446) );
  INV_X1 U8151 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6444) );
  MUX2_X1 U8152 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6444), .S(n6549), .Z(n6445)
         );
  INV_X1 U8153 ( .A(n6450), .ZN(n6672) );
  NAND2_X1 U8154 ( .A1(n6445), .A2(n6446), .ZN(n6551) );
  OAI211_X1 U8155 ( .C1(n6446), .C2(n6445), .A(n9084), .B(n6551), .ZN(n6447)
         );
  NAND2_X1 U8156 ( .A1(n6448), .A2(n6447), .ZN(n6452) );
  INV_X1 U8157 ( .A(n6549), .ZN(n6458) );
  INV_X1 U8158 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7011) );
  OAI22_X1 U8159 ( .A1(n9070), .A2(n6458), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7011), .ZN(n6451) );
  OR3_X1 U8160 ( .A1(n6453), .A2(n6452), .A3(n6451), .ZN(P1_U3244) );
  XNOR2_X1 U8161 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U8162 ( .A1(n4660), .A2(P2_U3151), .ZN(n8540) );
  NAND2_X1 U8163 ( .A1(n7885), .A2(P2_U3151), .ZN(n8546) );
  OAI222_X1 U8164 ( .A1(n8540), .A2(n6455), .B1(n8546), .B2(n6471), .C1(
        P2_U3151), .C2(n6454), .ZN(P2_U3293) );
  OAI222_X1 U8165 ( .A1(n8540), .A2(n6456), .B1(n8546), .B2(n6469), .C1(
        P2_U3151), .C2(n9724), .ZN(P2_U3292) );
  AND2_X1 U8166 ( .A1(n7885), .A2(P1_U3086), .ZN(n9409) );
  INV_X2 U8167 ( .A(n9409), .ZN(n7618) );
  INV_X1 U8168 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6459) );
  AND2_X1 U8169 ( .A1(n4660), .A2(P1_U3086), .ZN(n7508) );
  INV_X2 U8170 ( .A(n7508), .ZN(n9411) );
  INV_X1 U8171 ( .A(n6457), .ZN(n6464) );
  OAI222_X1 U8172 ( .A1(n7618), .A2(n6459), .B1(n9411), .B2(n6464), .C1(
        P1_U3086), .C2(n6458), .ZN(P1_U3354) );
  OAI222_X1 U8173 ( .A1(n8540), .A2(n6461), .B1(n8546), .B2(n6473), .C1(
        P2_U3151), .C2(n6460), .ZN(P2_U3291) );
  OAI222_X1 U8174 ( .A1(n8540), .A2(n6463), .B1(n8546), .B2(n6475), .C1(
        P2_U3151), .C2(n6462), .ZN(P2_U3290) );
  INV_X1 U8175 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6465) );
  INV_X1 U8176 ( .A(n8546), .ZN(n7504) );
  INV_X1 U8177 ( .A(n7504), .ZN(n8550) );
  OAI222_X1 U8178 ( .A1(n8540), .A2(n6465), .B1(n8550), .B2(n6464), .C1(
        P2_U3151), .C2(n9703), .ZN(P2_U3294) );
  OAI222_X1 U8179 ( .A1(n7618), .A2(n6466), .B1(n9411), .B2(n6467), .C1(
        P1_U3086), .C2(n9061), .ZN(P1_U3349) );
  OAI222_X1 U8180 ( .A1(n8540), .A2(n6468), .B1(n8546), .B2(n6467), .C1(
        P2_U3151), .C2(n9756), .ZN(P2_U3289) );
  OAI222_X1 U8181 ( .A1(n7618), .A2(n6470), .B1(n9411), .B2(n6469), .C1(
        P1_U3086), .C2(n9016), .ZN(P1_U3352) );
  OAI222_X1 U8182 ( .A1(n7618), .A2(n6472), .B1(n9411), .B2(n6471), .C1(
        P1_U3086), .C2(n6547), .ZN(P1_U3353) );
  OAI222_X1 U8183 ( .A1(n7618), .A2(n6474), .B1(n9411), .B2(n6473), .C1(
        P1_U3086), .C2(n9032), .ZN(P1_U3351) );
  OAI222_X1 U8184 ( .A1(n7618), .A2(n6476), .B1(n9411), .B2(n6475), .C1(
        P1_U3086), .C2(n9041), .ZN(P1_U3350) );
  OAI222_X1 U8185 ( .A1(n7618), .A2(n6477), .B1(n9411), .B2(n6478), .C1(
        P1_U3086), .C2(n9069), .ZN(P1_U3348) );
  OAI222_X1 U8186 ( .A1(n8540), .A2(n10052), .B1(n8546), .B2(n6478), .C1(
        P2_U3151), .C2(n6890), .ZN(P2_U3288) );
  OAI222_X1 U8187 ( .A1(n8540), .A2(n6479), .B1(n8546), .B2(n6480), .C1(
        P2_U3151), .C2(n9780), .ZN(P2_U3287) );
  OAI222_X1 U8188 ( .A1(n7618), .A2(n6481), .B1(n9411), .B2(n6480), .C1(
        P1_U3086), .C2(n6582), .ZN(P1_U3347) );
  INV_X1 U8189 ( .A(n8540), .ZN(n6523) );
  INV_X1 U8190 ( .A(n6523), .ZN(n8547) );
  OAI222_X1 U8191 ( .A1(n8550), .A2(n6483), .B1(n9790), .B2(P2_U3151), .C1(
        n6482), .C2(n8547), .ZN(P2_U3286) );
  OAI222_X1 U8192 ( .A1(n7618), .A2(n6484), .B1(n9411), .B2(n6483), .C1(n6595), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8193 ( .A(n6485), .ZN(n6492) );
  INV_X1 U8194 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6486) );
  OAI222_X1 U8195 ( .A1(n8550), .A2(n6492), .B1(n7491), .B2(P2_U3151), .C1(
        n6486), .C2(n8547), .ZN(P2_U3285) );
  INV_X1 U8196 ( .A(n6487), .ZN(n6490) );
  NAND2_X1 U8197 ( .A1(n6490), .A2(n6488), .ZN(n6508) );
  INV_X1 U8198 ( .A(n6489), .ZN(n6491) );
  AOI22_X1 U8199 ( .A1(n6508), .A2(n10228), .B1(n6491), .B2(n6490), .ZN(
        P2_U3376) );
  INV_X1 U8200 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6493) );
  INV_X1 U8201 ( .A(n6579), .ZN(n6627) );
  OAI222_X1 U8202 ( .A1(n7618), .A2(n6493), .B1(n9411), .B2(n6492), .C1(n6627), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U8203 ( .A1(n6709), .A2(n6494), .ZN(n6495) );
  OAI21_X1 U8204 ( .B1(n6709), .B2(n6496), .A(n6495), .ZN(P2_U3377) );
  INV_X1 U8205 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U8206 ( .A1(n6497), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8207 ( .A1(n5461), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U8208 ( .A1(n5657), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6498) );
  AND3_X1 U8209 ( .A1(n6500), .A2(n6499), .A3(n6498), .ZN(n9092) );
  INV_X1 U8210 ( .A(n9092), .ZN(n8828) );
  NAND2_X1 U8211 ( .A1(n8828), .A2(P1_U3973), .ZN(n6501) );
  OAI21_X1 U8212 ( .B1(n10158), .B2(P1_U3973), .A(n6501), .ZN(P1_U3585) );
  INV_X1 U8213 ( .A(n6502), .ZN(n6503) );
  INV_X1 U8214 ( .A(n6578), .ZN(n6637) );
  OAI222_X1 U8215 ( .A1(n7618), .A2(n6530), .B1(n9411), .B2(n6503), .C1(
        P1_U3086), .C2(n6637), .ZN(P1_U3344) );
  OAI222_X1 U8216 ( .A1(n8540), .A2(n6504), .B1(n8546), .B2(n6503), .C1(
        P2_U3151), .C2(n9806), .ZN(P2_U3284) );
  INV_X1 U8217 ( .A(n9026), .ZN(n9073) );
  NOR2_X1 U8218 ( .A1(n9073), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8219 ( .A(n6505), .ZN(n6520) );
  INV_X1 U8220 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6506) );
  OAI222_X1 U8221 ( .A1(n8550), .A2(n6520), .B1(n6507), .B2(P2_U3151), .C1(
        n6506), .C2(n8547), .ZN(P2_U3283) );
  INV_X1 U8222 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U8223 ( .A1(n6674), .A2(n6509), .ZN(P2_U3254) );
  INV_X1 U8224 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6510) );
  NOR2_X1 U8225 ( .A1(n6674), .A2(n6510), .ZN(P2_U3249) );
  INV_X1 U8226 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10194) );
  NOR2_X1 U8227 ( .A1(n6674), .A2(n10194), .ZN(P2_U3257) );
  INV_X1 U8228 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6511) );
  NOR2_X1 U8229 ( .A1(n6674), .A2(n6511), .ZN(P2_U3247) );
  INV_X1 U8230 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U8231 ( .A1(n6674), .A2(n6512), .ZN(P2_U3255) );
  INV_X1 U8232 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U8233 ( .A1(n6674), .A2(n6513), .ZN(P2_U3250) );
  INV_X1 U8234 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6514) );
  NOR2_X1 U8235 ( .A1(n6674), .A2(n6514), .ZN(P2_U3253) );
  INV_X1 U8236 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6515) );
  NOR2_X1 U8237 ( .A1(n6674), .A2(n6515), .ZN(P2_U3251) );
  INV_X1 U8238 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6516) );
  NOR2_X1 U8239 ( .A1(n6674), .A2(n6516), .ZN(P2_U3248) );
  INV_X1 U8240 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6517) );
  NOR2_X1 U8241 ( .A1(n6674), .A2(n6517), .ZN(P2_U3252) );
  INV_X1 U8242 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6518) );
  NOR2_X1 U8243 ( .A1(n6674), .A2(n6518), .ZN(P2_U3246) );
  INV_X1 U8244 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6519) );
  NOR2_X1 U8245 ( .A1(n6674), .A2(n6519), .ZN(P2_U3256) );
  INV_X1 U8246 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6521) );
  OAI222_X1 U8247 ( .A1(n7618), .A2(n6521), .B1(n9411), .B2(n6520), .C1(n6640), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8248 ( .A(n6522), .ZN(n6600) );
  AOI22_X1 U8249 ( .A1(n9822), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6523), .ZN(n6524) );
  OAI21_X1 U8250 ( .B1(n6600), .B2(n8546), .A(n6524), .ZN(P2_U3282) );
  INV_X1 U8251 ( .A(n9841), .ZN(n9858) );
  AOI22_X1 U8252 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n9858), .B1(n9856), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n6529) );
  OAI21_X1 U8253 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6525), .A(n9714), .ZN(n6526) );
  OAI21_X1 U8254 ( .B1(n6527), .B2(n9868), .A(n6526), .ZN(n6528) );
  OAI211_X1 U8255 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6811), .A(n6529), .B(n6528), .ZN(P2_U3182) );
  MUX2_X1 U8256 ( .A(n6530), .B(n7728), .S(P2_U3893), .Z(n6531) );
  INV_X1 U8257 ( .A(n6531), .ZN(P2_U3502) );
  INV_X1 U8258 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7072) );
  MUX2_X1 U8259 ( .A(n7072), .B(P1_REG2_REG_2__SCAN_IN), .S(n6547), .Z(n9007)
         );
  NAND2_X1 U8260 ( .A1(n6549), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8261 ( .A1(n6533), .A2(n6532), .ZN(n9006) );
  NAND2_X1 U8262 ( .A1(n9007), .A2(n9006), .ZN(n9005) );
  INV_X1 U8263 ( .A(n6547), .ZN(n9002) );
  NAND2_X1 U8264 ( .A1(n9002), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8265 ( .A1(n9005), .A2(n6534), .ZN(n9014) );
  INV_X1 U8266 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6535) );
  MUX2_X1 U8267 ( .A(n6535), .B(P1_REG2_REG_3__SCAN_IN), .S(n9016), .Z(n9015)
         );
  NAND2_X1 U8268 ( .A1(n9014), .A2(n9015), .ZN(n9013) );
  INV_X1 U8269 ( .A(n9016), .ZN(n6536) );
  NAND2_X1 U8270 ( .A1(n6536), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8271 ( .A1(n9013), .A2(n6537), .ZN(n9030) );
  XNOR2_X1 U8272 ( .A(n9032), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U8273 ( .A1(n9030), .A2(n9031), .ZN(n9029) );
  INV_X1 U8274 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6538) );
  OR2_X1 U8275 ( .A1(n9032), .A2(n6538), .ZN(n6539) );
  NAND2_X1 U8276 ( .A1(n9029), .A2(n6539), .ZN(n9045) );
  INV_X1 U8277 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10176) );
  MUX2_X1 U8278 ( .A(n10176), .B(P1_REG2_REG_5__SCAN_IN), .S(n9041), .Z(n9046)
         );
  NAND2_X1 U8279 ( .A1(n9045), .A2(n9046), .ZN(n9044) );
  OR2_X1 U8280 ( .A1(n9041), .A2(n10176), .ZN(n6540) );
  NAND2_X1 U8281 ( .A1(n9044), .A2(n6540), .ZN(n9058) );
  INV_X1 U8282 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U8283 ( .A(n10157), .B(P1_REG2_REG_6__SCAN_IN), .S(n9061), .Z(n9059)
         );
  NAND2_X1 U8284 ( .A1(n9058), .A2(n9059), .ZN(n9057) );
  INV_X1 U8285 ( .A(n9061), .ZN(n6561) );
  NAND2_X1 U8286 ( .A1(n6561), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U8287 ( .A1(n9057), .A2(n6541), .ZN(n9076) );
  XNOR2_X1 U8288 ( .A(n9069), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U8289 ( .A1(n9076), .A2(n9077), .ZN(n9074) );
  INV_X1 U8290 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6542) );
  OR2_X1 U8291 ( .A1(n9069), .A2(n6542), .ZN(n6543) );
  NAND2_X1 U8292 ( .A1(n9074), .A2(n6543), .ZN(n6544) );
  INV_X1 U8293 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10230) );
  MUX2_X1 U8294 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10230), .S(n6572), .Z(n6545)
         );
  AND2_X1 U8295 ( .A1(n6544), .A2(n6545), .ZN(n6571) );
  OAI21_X1 U8296 ( .B1(n6545), .B2(n6544), .A(n9075), .ZN(n6569) );
  AND2_X1 U8297 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7444) );
  NOR2_X1 U8298 ( .A1(n9070), .A2(n6582), .ZN(n6546) );
  AOI211_X1 U8299 ( .C1(n9073), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7444), .B(
        n6546), .ZN(n6568) );
  INV_X1 U8300 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6548) );
  MUX2_X1 U8301 ( .A(n6548), .B(P1_REG1_REG_2__SCAN_IN), .S(n6547), .Z(n9004)
         );
  NAND2_X1 U8302 ( .A1(n6549), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8303 ( .A1(n6551), .A2(n6550), .ZN(n9003) );
  NAND2_X1 U8304 ( .A1(n9004), .A2(n9003), .ZN(n9018) );
  NAND2_X1 U8305 ( .A1(n9002), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U8306 ( .A1(n9018), .A2(n9017), .ZN(n6554) );
  INV_X1 U8307 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6552) );
  MUX2_X1 U8308 ( .A(n6552), .B(P1_REG1_REG_3__SCAN_IN), .S(n9016), .Z(n6553)
         );
  NAND2_X1 U8309 ( .A1(n6554), .A2(n6553), .ZN(n9035) );
  OR2_X1 U8310 ( .A1(n9016), .A2(n6552), .ZN(n9034) );
  NAND2_X1 U8311 ( .A1(n9035), .A2(n9034), .ZN(n6557) );
  INV_X1 U8312 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6555) );
  MUX2_X1 U8313 ( .A(n6555), .B(P1_REG1_REG_4__SCAN_IN), .S(n9032), .Z(n6556)
         );
  NAND2_X1 U8314 ( .A1(n6557), .A2(n6556), .ZN(n9050) );
  INV_X1 U8315 ( .A(n9032), .ZN(n6558) );
  NAND2_X1 U8316 ( .A1(n6558), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9049) );
  INV_X1 U8317 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U8318 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9680), .S(n9041), .Z(n9048)
         );
  AOI21_X1 U8319 ( .B1(n9050), .B2(n9049), .A(n9048), .ZN(n9047) );
  NOR2_X1 U8320 ( .A1(n9041), .A2(n9680), .ZN(n9060) );
  INV_X1 U8321 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6559) );
  MUX2_X1 U8322 ( .A(n6559), .B(P1_REG1_REG_6__SCAN_IN), .S(n9061), .Z(n6560)
         );
  OAI21_X1 U8323 ( .B1(n9047), .B2(n9060), .A(n6560), .ZN(n9081) );
  NAND2_X1 U8324 ( .A1(n6561), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9080) );
  INV_X1 U8325 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9683) );
  MUX2_X1 U8326 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9683), .S(n9069), .Z(n9079)
         );
  AOI21_X1 U8327 ( .B1(n9081), .B2(n9080), .A(n9079), .ZN(n9078) );
  NOR2_X1 U8328 ( .A1(n9069), .A2(n9683), .ZN(n6565) );
  INV_X1 U8329 ( .A(n6565), .ZN(n6563) );
  INV_X1 U8330 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9685) );
  MUX2_X1 U8331 ( .A(n9685), .B(P1_REG1_REG_8__SCAN_IN), .S(n6572), .Z(n6562)
         );
  NAND2_X1 U8332 ( .A1(n6563), .A2(n6562), .ZN(n6566) );
  MUX2_X1 U8333 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9685), .S(n6572), .Z(n6564)
         );
  OAI21_X1 U8334 ( .B1(n9078), .B2(n6565), .A(n6564), .ZN(n6581) );
  OAI211_X1 U8335 ( .C1(n9078), .C2(n6566), .A(n9084), .B(n6581), .ZN(n6567)
         );
  OAI211_X1 U8336 ( .C1(n6571), .C2(n6569), .A(n6568), .B(n6567), .ZN(P1_U3251) );
  INV_X1 U8337 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10023) );
  NOR2_X1 U8338 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10023), .ZN(n8700) );
  INV_X1 U8339 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6570) );
  AOI22_X1 U8340 ( .A1(n6579), .A2(n6570), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6627), .ZN(n6621) );
  INV_X1 U8341 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U8342 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6580), .B1(n6595), .B2(
        n10056), .ZN(n6590) );
  AOI21_X1 U8343 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6572), .A(n6571), .ZN(
        n6592) );
  NAND2_X1 U8344 ( .A1(n6590), .A2(n6592), .ZN(n6591) );
  OAI21_X1 U8345 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6580), .A(n6591), .ZN(
        n6620) );
  NOR2_X1 U8346 ( .A1(n6621), .A2(n6620), .ZN(n6619) );
  AOI21_X1 U8347 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6579), .A(n6619), .ZN(
        n6576) );
  NAND2_X1 U8348 ( .A1(n6578), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6632) );
  OR2_X1 U8349 ( .A1(n6578), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6573) );
  NAND2_X1 U8350 ( .A1(n6632), .A2(n6573), .ZN(n6575) );
  OR2_X1 U8351 ( .A1(n6576), .A2(n6575), .ZN(n6633) );
  INV_X1 U8352 ( .A(n6633), .ZN(n6574) );
  AOI211_X1 U8353 ( .C1(n6576), .C2(n6575), .A(n6574), .B(n7300), .ZN(n6577)
         );
  AOI211_X1 U8354 ( .C1(n9073), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8700), .B(
        n6577), .ZN(n6586) );
  MUX2_X1 U8355 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9691), .S(n6578), .Z(n6584)
         );
  INV_X1 U8356 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9689) );
  MUX2_X1 U8357 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9689), .S(n6579), .Z(n6623)
         );
  INV_X1 U8358 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9687) );
  MUX2_X1 U8359 ( .A(n9687), .B(P1_REG1_REG_9__SCAN_IN), .S(n6580), .Z(n6588)
         );
  OAI21_X1 U8360 ( .B1(n9685), .B2(n6582), .A(n6581), .ZN(n6589) );
  NOR2_X1 U8361 ( .A1(n6588), .A2(n6589), .ZN(n6587) );
  AOI21_X1 U8362 ( .B1(n6595), .B2(n9687), .A(n6587), .ZN(n6624) );
  NAND2_X1 U8363 ( .A1(n6623), .A2(n6624), .ZN(n6622) );
  OAI21_X1 U8364 ( .B1(n6627), .B2(n9689), .A(n6622), .ZN(n6583) );
  NAND2_X1 U8365 ( .A1(n6584), .A2(n6583), .ZN(n6636) );
  OAI211_X1 U8366 ( .C1(n6584), .C2(n6583), .A(n9084), .B(n6636), .ZN(n6585)
         );
  OAI211_X1 U8367 ( .C1(n9070), .C2(n6637), .A(n6586), .B(n6585), .ZN(P1_U3254) );
  AOI21_X1 U8368 ( .B1(n6589), .B2(n6588), .A(n6587), .ZN(n6599) );
  AOI221_X1 U8369 ( .B1(n6592), .B2(n6591), .C1(n6590), .C2(n6591), .A(n7300), 
        .ZN(n6593) );
  INV_X1 U8370 ( .A(n6593), .ZN(n6598) );
  NOR2_X1 U8371 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6594), .ZN(n7400) );
  NOR2_X1 U8372 ( .A1(n9070), .A2(n6595), .ZN(n6596) );
  AOI211_X1 U8373 ( .C1(n9073), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7400), .B(
        n6596), .ZN(n6597) );
  OAI211_X1 U8374 ( .C1(n6599), .C2(n7429), .A(n6598), .B(n6597), .ZN(P1_U3252) );
  INV_X1 U8375 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6601) );
  INV_X1 U8376 ( .A(n6777), .ZN(n6646) );
  OAI222_X1 U8377 ( .A1(n7618), .A2(n6601), .B1(n9411), .B2(n6600), .C1(
        P1_U3086), .C2(n6646), .ZN(P1_U3342) );
  XNOR2_X1 U8378 ( .A(n6603), .B(n6602), .ZN(n6618) );
  OAI21_X1 U8379 ( .B1(n6606), .B2(n6605), .A(n6604), .ZN(n6607) );
  INV_X1 U8380 ( .A(n6607), .ZN(n6608) );
  NOR2_X1 U8381 ( .A1(n6608), .A2(n9872), .ZN(n6610) );
  NOR2_X1 U8382 ( .A1(n7264), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6609) );
  AOI211_X1 U8383 ( .C1(n9858), .C2(n6611), .A(n6610), .B(n6609), .ZN(n6617)
         );
  OAI21_X1 U8384 ( .B1(n6614), .B2(n6613), .A(n6612), .ZN(n6615) );
  AOI22_X1 U8385 ( .A1(n9863), .A2(n6615), .B1(n9856), .B2(
        P2_ADDR_REG_2__SCAN_IN), .ZN(n6616) );
  OAI211_X1 U8386 ( .C1(n9847), .C2(n6618), .A(n6617), .B(n6616), .ZN(P2_U3184) );
  AOI211_X1 U8387 ( .C1(n6621), .C2(n6620), .A(n6619), .B(n7300), .ZN(n6629)
         );
  OAI211_X1 U8388 ( .C1(n6624), .C2(n6623), .A(n9084), .B(n6622), .ZN(n6626)
         );
  INV_X1 U8389 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U8390 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10213), .ZN(n7542) );
  AOI21_X1 U8391 ( .B1(n9073), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7542), .ZN(
        n6625) );
  OAI211_X1 U8392 ( .C1(n9070), .C2(n6627), .A(n6626), .B(n6625), .ZN(n6628)
         );
  OR2_X1 U8393 ( .A1(n6629), .A2(n6628), .ZN(P1_U3253) );
  INV_X1 U8394 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6630) );
  AOI22_X1 U8395 ( .A1(n6777), .A2(n6630), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n6646), .ZN(n6635) );
  NOR2_X1 U8396 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6659), .ZN(n6631) );
  AOI21_X1 U8397 ( .B1(n6659), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6631), .ZN(
        n6654) );
  AND2_X1 U8398 ( .A1(n6633), .A2(n6632), .ZN(n6656) );
  NAND2_X1 U8399 ( .A1(n6654), .A2(n6656), .ZN(n6655) );
  OAI21_X1 U8400 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6659), .A(n6655), .ZN(
        n6634) );
  NOR2_X1 U8401 ( .A1(n6635), .A2(n6634), .ZN(n6770) );
  AOI211_X1 U8402 ( .C1(n6635), .C2(n6634), .A(n6770), .B(n7300), .ZN(n6648)
         );
  INV_X1 U8403 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9693) );
  INV_X1 U8404 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9691) );
  OAI21_X1 U8405 ( .B1(n9691), .B2(n6637), .A(n6636), .ZN(n6650) );
  NAND2_X1 U8406 ( .A1(n6640), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6638) );
  OAI21_X1 U8407 ( .B1(n6640), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6638), .ZN(
        n6639) );
  INV_X1 U8408 ( .A(n6639), .ZN(n6651) );
  NOR2_X1 U8409 ( .A1(n6650), .A2(n6651), .ZN(n6649) );
  AOI21_X1 U8410 ( .B1(n9693), .B2(n6640), .A(n6649), .ZN(n6643) );
  NOR2_X1 U8411 ( .A1(n6777), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6641) );
  AOI21_X1 U8412 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6777), .A(n6641), .ZN(
        n6642) );
  NAND2_X1 U8413 ( .A1(n6642), .A2(n6643), .ZN(n6781) );
  OAI211_X1 U8414 ( .C1(n6643), .C2(n6642), .A(n9084), .B(n6781), .ZN(n6645)
         );
  NOR2_X1 U8415 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10195), .ZN(n7629) );
  AOI21_X1 U8416 ( .B1(n9073), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7629), .ZN(
        n6644) );
  OAI211_X1 U8417 ( .C1(n9070), .C2(n6646), .A(n6645), .B(n6644), .ZN(n6647)
         );
  OR2_X1 U8418 ( .A1(n6648), .A2(n6647), .ZN(P1_U3256) );
  INV_X1 U8419 ( .A(n9070), .ZN(n9001) );
  AOI21_X1 U8420 ( .B1(n6651), .B2(n6650), .A(n6649), .ZN(n6653) );
  AND2_X1 U8421 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8631) );
  AOI21_X1 U8422 ( .B1(n9073), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8631), .ZN(
        n6652) );
  OAI21_X1 U8423 ( .B1(n7429), .B2(n6653), .A(n6652), .ZN(n6658) );
  AOI221_X1 U8424 ( .B1(n6656), .B2(n6655), .C1(n6654), .C2(n6655), .A(n7300), 
        .ZN(n6657) );
  AOI211_X1 U8425 ( .C1(n9001), .C2(n6659), .A(n6658), .B(n6657), .ZN(n6660)
         );
  INV_X1 U8426 ( .A(n6660), .ZN(P1_U3255) );
  INV_X1 U8427 ( .A(n6661), .ZN(n6663) );
  INV_X1 U8428 ( .A(n6780), .ZN(n6868) );
  OAI222_X1 U8429 ( .A1(n7618), .A2(n10206), .B1(n9411), .B2(n6663), .C1(
        P1_U3086), .C2(n6868), .ZN(P1_U3341) );
  OAI222_X1 U8430 ( .A1(n8540), .A2(n6664), .B1(n8546), .B2(n6663), .C1(
        P2_U3151), .C2(n6662), .ZN(P2_U3281) );
  NOR2_X1 U8431 ( .A1(n8992), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6665) );
  OR2_X1 U8432 ( .A1(n5160), .A2(n6665), .ZN(n8995) );
  INV_X1 U8433 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9674) );
  AOI21_X1 U8434 ( .B1(n8992), .B2(n9674), .A(n8995), .ZN(n6666) );
  MUX2_X1 U8435 ( .A(n8995), .B(n6666), .S(n4710), .Z(n6671) );
  INV_X1 U8436 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6668) );
  INV_X1 U8437 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6667) );
  OAI22_X1 U8438 ( .A1(n9026), .A2(n6668), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6667), .ZN(n6670) );
  NOR3_X1 U8439 ( .A1(n7429), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n4710), .ZN(
        n6669) );
  AOI211_X1 U8440 ( .C1(n6672), .C2(n6671), .A(n6670), .B(n6669), .ZN(n6673)
         );
  INV_X1 U8441 ( .A(n6673), .ZN(P1_U3243) );
  INV_X1 U8442 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6675) );
  NOR2_X1 U8443 ( .A1(n6674), .A2(n6675), .ZN(P2_U3261) );
  INV_X1 U8444 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10251) );
  NOR2_X1 U8445 ( .A1(n6674), .A2(n10251), .ZN(P2_U3258) );
  INV_X1 U8446 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U8447 ( .A1(n6674), .A2(n6676), .ZN(P2_U3260) );
  INV_X1 U8448 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6677) );
  NOR2_X1 U8449 ( .A1(n6674), .A2(n6677), .ZN(P2_U3259) );
  INV_X1 U8450 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6678) );
  NOR2_X1 U8451 ( .A1(n6674), .A2(n6678), .ZN(P2_U3263) );
  INV_X1 U8452 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6679) );
  NOR2_X1 U8453 ( .A1(n6674), .A2(n6679), .ZN(P2_U3237) );
  INV_X1 U8454 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6680) );
  NOR2_X1 U8455 ( .A1(n6674), .A2(n6680), .ZN(P2_U3245) );
  INV_X1 U8456 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6681) );
  NOR2_X1 U8457 ( .A1(n6674), .A2(n6681), .ZN(P2_U3243) );
  INV_X1 U8458 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U8459 ( .A1(n6674), .A2(n6682), .ZN(P2_U3242) );
  INV_X1 U8460 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10242) );
  NOR2_X1 U8461 ( .A1(n6674), .A2(n10242), .ZN(P2_U3241) );
  INV_X1 U8462 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6683) );
  NOR2_X1 U8463 ( .A1(n6674), .A2(n6683), .ZN(P2_U3240) );
  INV_X1 U8464 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U8465 ( .A1(n6674), .A2(n10035), .ZN(P2_U3239) );
  INV_X1 U8466 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U8467 ( .A1(n6674), .A2(n6684), .ZN(P2_U3238) );
  INV_X1 U8468 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U8469 ( .A1(n6674), .A2(n6685), .ZN(P2_U3262) );
  INV_X1 U8470 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U8471 ( .A1(n6674), .A2(n6686), .ZN(P2_U3244) );
  INV_X1 U8472 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U8473 ( .A1(n6674), .A2(n6687), .ZN(P2_U3236) );
  INV_X1 U8474 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6688) );
  NOR2_X1 U8475 ( .A1(n6674), .A2(n6688), .ZN(P2_U3235) );
  INV_X1 U8476 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U8477 ( .A1(n6674), .A2(n6689), .ZN(P2_U3234) );
  INV_X1 U8478 ( .A(n6690), .ZN(n6692) );
  OAI222_X1 U8479 ( .A1(n8550), .A2(n6692), .B1(n9840), .B2(P2_U3151), .C1(
        n6691), .C2(n8547), .ZN(P2_U3280) );
  INV_X1 U8480 ( .A(n6962), .ZN(n6969) );
  OAI222_X1 U8481 ( .A1(n7618), .A2(n10143), .B1(n9411), .B2(n6692), .C1(n6969), .C2(P1_U3086), .ZN(P1_U3340) );
  XOR2_X1 U8482 ( .A(n6693), .B(n4403), .Z(n8993) );
  INV_X1 U8483 ( .A(n8993), .ZN(n6698) );
  OR2_X1 U8484 ( .A1(n6695), .A2(n9307), .ZN(n8715) );
  INV_X1 U8485 ( .A(n9569), .ZN(n8920) );
  OAI22_X1 U8486 ( .A1(n8920), .A2(n8704), .B1(n8739), .B2(n6947), .ZN(n6696)
         );
  AOI21_X1 U8487 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8715), .A(n6696), .ZN(
        n6697) );
  OAI21_X1 U8488 ( .B1(n6698), .B2(n8745), .A(n6697), .ZN(P1_U3232) );
  INV_X1 U8489 ( .A(n6699), .ZN(n6701) );
  OAI21_X1 U8490 ( .B1(n6702), .B2(n6701), .A(n6700), .ZN(n6708) );
  AND2_X1 U8491 ( .A1(n6703), .A2(n7505), .ZN(n6705) );
  OAI211_X1 U8492 ( .C1(n6741), .C2(n6711), .A(n6705), .B(n6704), .ZN(n6706)
         );
  INV_X1 U8493 ( .A(n6706), .ZN(n6707) );
  AOI21_X1 U8494 ( .B1(n6708), .B2(n6707), .A(P2_U3151), .ZN(n6713) );
  INV_X1 U8495 ( .A(n6720), .ZN(n6710) );
  NAND2_X1 U8496 ( .A1(n6710), .A2(n6709), .ZN(n8096) );
  NOR2_X1 U8497 ( .A1(n8096), .A2(n6711), .ZN(n6712) );
  NOR2_X1 U8498 ( .A1(n7875), .A2(P2_U3151), .ZN(n6812) );
  NAND2_X1 U8499 ( .A1(n6739), .A2(n9918), .ZN(n6716) );
  NOR2_X1 U8500 ( .A1(n6720), .A2(n6717), .ZN(n6718) );
  INV_X1 U8501 ( .A(n7858), .ZN(n7873) );
  INV_X1 U8502 ( .A(n6214), .ZN(n6722) );
  INV_X1 U8503 ( .A(n9884), .ZN(n6796) );
  NOR2_X1 U8504 ( .A1(n6720), .A2(n6719), .ZN(n6721) );
  OAI22_X1 U8505 ( .A1(n7873), .A2(n6722), .B1(n6796), .B2(n7860), .ZN(n6723)
         );
  AOI21_X1 U8506 ( .B1(n6880), .B2(n7850), .A(n6723), .ZN(n6748) );
  INV_X1 U8507 ( .A(n6724), .ZN(n6725) );
  NAND2_X1 U8508 ( .A1(n6726), .A2(n6725), .ZN(n6727) );
  INV_X1 U8509 ( .A(n6732), .ZN(n6730) );
  NAND2_X1 U8510 ( .A1(n6730), .A2(n6731), .ZN(n6733) );
  INV_X1 U8511 ( .A(n6731), .ZN(n6802) );
  NAND2_X1 U8512 ( .A1(n6802), .A2(n6732), .ZN(n6797) );
  OR2_X1 U8513 ( .A1(n7118), .A2(n6808), .ZN(n6735) );
  NAND2_X1 U8514 ( .A1(n7914), .A2(n6735), .ZN(n6737) );
  OAI21_X1 U8515 ( .B1(n6736), .B2(n6737), .A(n6798), .ZN(n6746) );
  INV_X1 U8516 ( .A(n6738), .ZN(n6740) );
  NAND2_X1 U8517 ( .A1(n6740), .A2(n6739), .ZN(n6745) );
  INV_X1 U8518 ( .A(n6741), .ZN(n6742) );
  NAND2_X1 U8519 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  NAND2_X1 U8520 ( .A1(n6746), .A2(n7866), .ZN(n6747) );
  OAI211_X1 U8521 ( .C1(n6812), .C2(n7140), .A(n6748), .B(n6747), .ZN(P2_U3162) );
  OR2_X1 U8522 ( .A1(n9726), .A2(n6749), .ZN(n6751) );
  AOI211_X1 U8523 ( .C1(n6752), .C2(n6751), .A(n9847), .B(n6750), .ZN(n6769)
         );
  NOR2_X1 U8524 ( .A1(n4834), .A2(n6754), .ZN(n6755) );
  NAND2_X1 U8525 ( .A1(n9730), .A2(n6755), .ZN(n6756) );
  AND2_X1 U8526 ( .A1(n6757), .A2(n6756), .ZN(n6767) );
  INV_X1 U8527 ( .A(n6758), .ZN(n6760) );
  NAND3_X1 U8528 ( .A1(n9720), .A2(n6760), .A3(n6759), .ZN(n6761) );
  AOI21_X1 U8529 ( .B1(n6762), .B2(n6761), .A(n9849), .ZN(n6763) );
  AOI21_X1 U8530 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(n9856), .A(n6763), .ZN(
        n6766) );
  AND2_X1 U8531 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6911) );
  AOI21_X1 U8532 ( .B1(n9858), .B2(n6764), .A(n6911), .ZN(n6765) );
  OAI211_X1 U8533 ( .C1(n6767), .C2(n9872), .A(n6766), .B(n6765), .ZN(n6768)
         );
  OR2_X1 U8534 ( .A1(n6769), .A2(n6768), .ZN(P2_U3186) );
  NAND2_X1 U8535 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8556) );
  INV_X1 U8536 ( .A(n8556), .ZN(n6776) );
  AOI21_X1 U8537 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n6777), .A(n6770), .ZN(
        n6774) );
  NAND2_X1 U8538 ( .A1(n6780), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6872) );
  OR2_X1 U8539 ( .A1(n6780), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U8540 ( .A1(n6872), .A2(n6771), .ZN(n6773) );
  INV_X1 U8541 ( .A(n6873), .ZN(n6772) );
  AOI211_X1 U8542 ( .C1(n6774), .C2(n6773), .A(n6772), .B(n7300), .ZN(n6775)
         );
  AOI211_X1 U8543 ( .C1(n9073), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n6776), .B(
        n6775), .ZN(n6787) );
  NAND2_X1 U8544 ( .A1(n6780), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8545 ( .A1(n6777), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8546 ( .A1(n6783), .A2(n6781), .ZN(n6778) );
  OAI211_X1 U8547 ( .C1(n6780), .C2(P1_REG1_REG_14__SCAN_IN), .A(n6779), .B(
        n6778), .ZN(n6867) );
  INV_X1 U8548 ( .A(n6781), .ZN(n6782) );
  AOI21_X1 U8549 ( .B1(n6868), .B2(P1_REG1_REG_14__SCAN_IN), .A(n6782), .ZN(
        n6784) );
  OAI211_X1 U8550 ( .C1(P1_REG1_REG_14__SCAN_IN), .C2(n6868), .A(n6784), .B(
        n6783), .ZN(n6785) );
  NAND3_X1 U8551 ( .A1(n9084), .A2(n6867), .A3(n6785), .ZN(n6786) );
  OAI211_X1 U8552 ( .C1(n9070), .C2(n6868), .A(n6787), .B(n6786), .ZN(P1_U3257) );
  AOI21_X1 U8553 ( .B1(n6789), .B2(n6788), .A(n6828), .ZN(n6794) );
  NOR2_X1 U8554 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6791), .ZN(n9012) );
  INV_X1 U8555 ( .A(n8990), .ZN(n9580) );
  OAI22_X1 U8556 ( .A1(n9580), .A2(n8737), .B1(n8704), .B2(n7086), .ZN(n6790)
         );
  AOI211_X1 U8557 ( .C1(n7060), .C2(n5770), .A(n9012), .B(n6790), .ZN(n6793)
         );
  NAND2_X1 U8558 ( .A1(n8742), .A2(n6791), .ZN(n6792) );
  OAI211_X1 U8559 ( .C1(n6794), .C2(n8745), .A(n6793), .B(n6792), .ZN(P1_U3218) );
  INV_X1 U8560 ( .A(n6795), .ZN(n6819) );
  OAI222_X1 U8561 ( .A1(n8550), .A2(n6819), .B1(n8138), .B2(P2_U3151), .C1(
        n10114), .C2(n8547), .ZN(P2_U3279) );
  XNOR2_X1 U8562 ( .A(n6846), .B(n6796), .ZN(n6800) );
  NAND2_X1 U8563 ( .A1(n6798), .A2(n6797), .ZN(n6799) );
  NAND2_X1 U8564 ( .A1(n6799), .A2(n6800), .ZN(n6848) );
  OAI21_X1 U8565 ( .B1(n6800), .B2(n6799), .A(n6848), .ZN(n6801) );
  NAND2_X1 U8566 ( .A1(n6801), .A2(n7866), .ZN(n6807) );
  INV_X1 U8567 ( .A(n8112), .ZN(n6803) );
  OAI22_X1 U8568 ( .A1(n7873), .A2(n6802), .B1(n6803), .B2(n7860), .ZN(n6804)
         );
  AOI21_X1 U8569 ( .B1(n6805), .B2(n7850), .A(n6804), .ZN(n6806) );
  OAI211_X1 U8570 ( .C1(n6812), .C2(n7264), .A(n6807), .B(n6806), .ZN(P2_U3177) );
  NAND2_X1 U8571 ( .A1(n6214), .A2(n7291), .ZN(n7911) );
  NAND2_X1 U8572 ( .A1(n7914), .A2(n7911), .ZN(n7285) );
  INV_X1 U8573 ( .A(n7860), .ZN(n7871) );
  AOI22_X1 U8574 ( .A1(n7866), .A2(n7285), .B1(n7871), .B2(n6731), .ZN(n6810)
         );
  NAND2_X1 U8575 ( .A1(n7850), .A2(n6808), .ZN(n6809) );
  OAI211_X1 U8576 ( .C1(n6812), .C2(n6811), .A(n6810), .B(n6809), .ZN(P2_U3172) );
  INV_X1 U8577 ( .A(n8711), .ZN(n6814) );
  AOI21_X1 U8578 ( .B1(n6815), .B2(n6813), .A(n6814), .ZN(n6818) );
  INV_X1 U8579 ( .A(n8737), .ZN(n8714) );
  AOI22_X1 U8580 ( .A1(n8714), .A2(n8991), .B1(n5770), .B2(n8919), .ZN(n6817)
         );
  INV_X1 U8581 ( .A(n8704), .ZN(n8734) );
  AOI22_X1 U8582 ( .A1(n8734), .A2(n8990), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8715), .ZN(n6816) );
  OAI211_X1 U8583 ( .C1(n6818), .C2(n8745), .A(n6817), .B(n6816), .ZN(P1_U3222) );
  OAI222_X1 U8584 ( .A1(n7618), .A2(n6820), .B1(n9411), .B2(n6819), .C1(n7221), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8585 ( .A(n6927), .ZN(n7389) );
  INV_X1 U8586 ( .A(n6821), .ZN(n9925) );
  OAI21_X1 U8587 ( .B1(n9938), .B2(n6212), .A(n7285), .ZN(n6822) );
  NAND2_X1 U8588 ( .A1(n6731), .A2(n8370), .ZN(n7283) );
  NAND2_X1 U8589 ( .A1(n6822), .A2(n7283), .ZN(n6860) );
  INV_X1 U8590 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6823) );
  OAI22_X1 U8591 ( .A1(n7291), .A2(n8513), .B1(n9939), .B2(n6823), .ZN(n6824)
         );
  AOI21_X1 U8592 ( .B1(n9939), .B2(n6860), .A(n6824), .ZN(n6825) );
  INV_X1 U8593 ( .A(n6825), .ZN(P2_U3390) );
  INV_X1 U8594 ( .A(n8742), .ZN(n7453) );
  INV_X1 U8595 ( .A(n7063), .ZN(n6835) );
  OAI21_X1 U8596 ( .B1(n6828), .B2(n6827), .A(n6826), .ZN(n6829) );
  NAND3_X1 U8597 ( .A1(n6830), .A2(n8722), .A3(n6829), .ZN(n6834) );
  INV_X1 U8598 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6831) );
  NOR2_X1 U8599 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6831), .ZN(n9024) );
  INV_X1 U8600 ( .A(n9586), .ZN(n7079) );
  OAI22_X1 U8601 ( .A1(n7079), .A2(n8737), .B1(n8704), .B2(n9605), .ZN(n6832)
         );
  AOI211_X1 U8602 ( .C1(n9585), .C2(n5770), .A(n9024), .B(n6832), .ZN(n6833)
         );
  OAI211_X1 U8603 ( .C1(n7453), .C2(n6835), .A(n6834), .B(n6833), .ZN(P1_U3230) );
  NAND2_X1 U8604 ( .A1(n8113), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6836) );
  OAI21_X1 U8605 ( .B1(n7900), .B2(n8113), .A(n6836), .ZN(P2_U3521) );
  INV_X1 U8606 ( .A(n9938), .ZN(n9912) );
  INV_X1 U8607 ( .A(n6837), .ZN(n6839) );
  AOI22_X1 U8608 ( .A1(n6839), .A2(n7945), .B1(n7914), .B2(n6838), .ZN(n7146)
         );
  OAI21_X1 U8609 ( .B1(n6838), .B2(n6841), .A(n6840), .ZN(n6842) );
  AOI222_X1 U8610 ( .A1(n6212), .A2(n6842), .B1(n9884), .B2(n8370), .C1(n6214), 
        .C2(n9883), .ZN(n7142) );
  OAI21_X1 U8611 ( .B1(n9912), .B2(n7146), .A(n7142), .ZN(n6879) );
  INV_X1 U8612 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6843) );
  OAI22_X1 U8613 ( .A1(n7141), .A2(n8513), .B1(n9939), .B2(n6843), .ZN(n6844)
         );
  AOI21_X1 U8614 ( .B1(n6879), .B2(n9939), .A(n6844), .ZN(n6845) );
  INV_X1 U8615 ( .A(n6845), .ZN(P2_U3393) );
  INV_X1 U8616 ( .A(n7875), .ZN(n7848) );
  OR2_X1 U8617 ( .A1(n6846), .A2(n9884), .ZN(n6847) );
  NAND2_X1 U8618 ( .A1(n6848), .A2(n6847), .ZN(n6849) );
  XNOR2_X1 U8619 ( .A(n6904), .B(n8112), .ZN(n6850) );
  AOI21_X1 U8620 ( .B1(n6849), .B2(n6850), .A(n7852), .ZN(n6853) );
  INV_X1 U8621 ( .A(n6849), .ZN(n6852) );
  INV_X1 U8622 ( .A(n6850), .ZN(n6851) );
  NAND2_X1 U8623 ( .A1(n6853), .A2(n6906), .ZN(n6858) );
  NAND2_X1 U8624 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9736) );
  INV_X1 U8625 ( .A(n9736), .ZN(n6854) );
  AOI21_X1 U8626 ( .B1(n7858), .B2(n9884), .A(n6854), .ZN(n6855) );
  OAI21_X1 U8627 ( .B1(n4753), .B2(n7860), .A(n6855), .ZN(n6856) );
  AOI21_X1 U8628 ( .B1(n9896), .B2(n7850), .A(n6856), .ZN(n6857) );
  OAI211_X1 U8629 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7848), .A(n6858), .B(
        n6857), .ZN(P2_U3158) );
  OAI22_X1 U8630 ( .A1(n8414), .A2(n7291), .B1(n9951), .B2(n6391), .ZN(n6859)
         );
  AOI21_X1 U8631 ( .B1(n9951), .B2(n6860), .A(n6859), .ZN(n6861) );
  INV_X1 U8632 ( .A(n6861), .ZN(P2_U3459) );
  INV_X1 U8633 ( .A(n6862), .ZN(n6865) );
  OAI222_X1 U8634 ( .A1(n7618), .A2(n6863), .B1(n9411), .B2(n6865), .C1(
        P1_U3086), .C2(n7305), .ZN(P1_U3338) );
  OAI222_X1 U8635 ( .A1(n8547), .A2(n6866), .B1(n8546), .B2(n6865), .C1(
        P2_U3151), .C2(n6864), .ZN(P2_U3278) );
  INV_X1 U8636 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6871) );
  INV_X1 U8637 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9698) );
  OAI21_X1 U8638 ( .B1(n9698), .B2(n6868), .A(n6867), .ZN(n6961) );
  XNOR2_X1 U8639 ( .A(n6961), .B(n6969), .ZN(n6869) );
  NAND2_X1 U8640 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n6869), .ZN(n6963) );
  OAI211_X1 U8641 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n6869), .A(n9084), .B(
        n6963), .ZN(n6870) );
  NAND2_X1 U8642 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8735) );
  OAI211_X1 U8643 ( .C1(n9026), .C2(n6871), .A(n6870), .B(n8735), .ZN(n6877)
         );
  INV_X1 U8644 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6875) );
  XOR2_X1 U8645 ( .A(n6970), .B(n6962), .Z(n6874) );
  NOR2_X1 U8646 ( .A1(n6875), .A2(n6874), .ZN(n6971) );
  AOI211_X1 U8647 ( .C1(n6875), .C2(n6874), .A(n6971), .B(n7300), .ZN(n6876)
         );
  AOI211_X1 U8648 ( .C1(n9001), .C2(n6962), .A(n6877), .B(n6876), .ZN(n6878)
         );
  INV_X1 U8649 ( .A(n6878), .ZN(P1_U3258) );
  INV_X1 U8650 ( .A(n6879), .ZN(n6882) );
  AOI22_X1 U8651 ( .A1(n8432), .A2(n6880), .B1(n6296), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n6881) );
  OAI21_X1 U8652 ( .B1(n6882), .B2(n6296), .A(n6881), .ZN(P2_U3460) );
  AOI21_X1 U8653 ( .B1(n9945), .B2(n6884), .A(n6883), .ZN(n6895) );
  OAI21_X1 U8654 ( .B1(n4502), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6885), .ZN(
        n6886) );
  AOI22_X1 U8655 ( .A1(n9863), .A2(n6886), .B1(n9856), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n6894) );
  OAI21_X1 U8656 ( .B1(n6889), .B2(n6888), .A(n6887), .ZN(n6892) );
  AND2_X1 U8657 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7241) );
  NOR2_X1 U8658 ( .A1(n9841), .A2(n6890), .ZN(n6891) );
  AOI211_X1 U8659 ( .C1(n9868), .C2(n6892), .A(n7241), .B(n6891), .ZN(n6893)
         );
  OAI211_X1 U8660 ( .C1(n6895), .C2(n9872), .A(n6894), .B(n6893), .ZN(P2_U3189) );
  XNOR2_X1 U8661 ( .A(n9879), .B(n6896), .ZN(n6900) );
  XNOR2_X1 U8662 ( .A(n6897), .B(n6896), .ZN(n6901) );
  NAND2_X1 U8663 ( .A1(n6901), .A2(n6927), .ZN(n6899) );
  AOI22_X1 U8664 ( .A1(n9883), .A2(n6731), .B1(n8112), .B2(n8370), .ZN(n6898)
         );
  OAI211_X1 U8665 ( .C1(n6900), .C2(n8347), .A(n6899), .B(n6898), .ZN(n7266)
         );
  INV_X1 U8666 ( .A(n6901), .ZN(n7270) );
  OAI22_X1 U8667 ( .A1(n7270), .A2(n9925), .B1(n7263), .B2(n9933), .ZN(n6902)
         );
  NOR2_X1 U8668 ( .A1(n7266), .A2(n6902), .ZN(n9894) );
  MUX2_X1 U8669 ( .A(n10092), .B(n9894), .S(n9951), .Z(n6903) );
  INV_X1 U8670 ( .A(n6903), .ZN(P2_U3461) );
  NAND2_X1 U8671 ( .A1(n6904), .A2(n8112), .ZN(n6905) );
  XNOR2_X1 U8672 ( .A(n7118), .B(n9901), .ZN(n6907) );
  NAND2_X1 U8673 ( .A1(n6907), .A2(n9885), .ZN(n6908) );
  NAND2_X1 U8674 ( .A1(n6987), .A2(n6908), .ZN(n6986) );
  NOR2_X1 U8675 ( .A1(n6984), .A2(n6986), .ZN(n6983) );
  AOI21_X1 U8676 ( .B1(n6984), .B2(n6986), .A(n6983), .ZN(n6915) );
  INV_X1 U8677 ( .A(n6909), .ZN(n6933) );
  INV_X1 U8678 ( .A(n8111), .ZN(n7114) );
  NOR2_X1 U8679 ( .A1(n7860), .A2(n7114), .ZN(n6910) );
  AOI211_X1 U8680 ( .C1(n7858), .C2(n8112), .A(n6911), .B(n6910), .ZN(n6912)
         );
  OAI21_X1 U8681 ( .B1(n9901), .B2(n7878), .A(n6912), .ZN(n6913) );
  AOI21_X1 U8682 ( .B1(n6933), .B2(n7875), .A(n6913), .ZN(n6914) );
  OAI21_X1 U8683 ( .B1(n6915), .B2(n7852), .A(n6914), .ZN(P2_U3170) );
  INV_X1 U8684 ( .A(n6916), .ZN(n6917) );
  OAI222_X1 U8685 ( .A1(n8550), .A2(n6917), .B1(n9460), .B2(P2_U3151), .C1(
        n10172), .C2(n8547), .ZN(P2_U3277) );
  OAI222_X1 U8686 ( .A1(n7618), .A2(n6918), .B1(n9411), .B2(n6917), .C1(n7315), 
        .C2(P1_U3086), .ZN(P1_U3337) );
  AND2_X1 U8687 ( .A1(n6919), .A2(n4512), .ZN(n7262) );
  OR2_X1 U8688 ( .A1(n6922), .A2(n6920), .ZN(n6925) );
  INV_X1 U8689 ( .A(n6726), .ZN(n6921) );
  NAND2_X1 U8690 ( .A1(n6921), .A2(n6920), .ZN(n6924) );
  NAND2_X1 U8691 ( .A1(n6922), .A2(n6726), .ZN(n6923) );
  NAND4_X1 U8692 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n6931)
         );
  INV_X1 U8693 ( .A(n7950), .ZN(n7916) );
  XNOR2_X1 U8694 ( .A(n6928), .B(n7916), .ZN(n9902) );
  XNOR2_X1 U8695 ( .A(n6929), .B(n7950), .ZN(n6930) );
  AOI222_X1 U8696 ( .A1(n6212), .A2(n6930), .B1(n8111), .B2(n8370), .C1(n8112), 
        .C2(n9883), .ZN(n9900) );
  MUX2_X1 U8697 ( .A(n10188), .B(n9900), .S(n8373), .Z(n6936) );
  INV_X1 U8698 ( .A(n6931), .ZN(n6932) );
  INV_X1 U8699 ( .A(n8336), .ZN(n8352) );
  INV_X1 U8700 ( .A(n9901), .ZN(n6934) );
  AOI22_X1 U8701 ( .A1(n9889), .A2(n6934), .B1(n9890), .B2(n6933), .ZN(n6935)
         );
  OAI211_X1 U8702 ( .C1(n8378), .C2(n9902), .A(n6936), .B(n6935), .ZN(P2_U3229) );
  NAND2_X1 U8703 ( .A1(n6938), .A2(n6937), .ZN(n6940) );
  XNOR2_X1 U8704 ( .A(n6940), .B(n6939), .ZN(n6946) );
  INV_X1 U8705 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6941) );
  NOR2_X1 U8706 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6941), .ZN(n9043) );
  OAI22_X1 U8707 ( .A1(n7086), .A2(n8737), .B1(n8704), .B2(n7162), .ZN(n6942)
         );
  AOI211_X1 U8708 ( .C1(n9594), .C2(n5770), .A(n9043), .B(n6942), .ZN(n6945)
         );
  NAND2_X1 U8709 ( .A1(n8742), .A2(n6943), .ZN(n6944) );
  OAI211_X1 U8710 ( .C1(n6946), .C2(n8745), .A(n6945), .B(n6944), .ZN(P1_U3227) );
  INV_X1 U8711 ( .A(n9535), .ZN(n9277) );
  NOR2_X1 U8712 ( .A1(n8920), .A2(n9277), .ZN(n9559) );
  NOR2_X1 U8713 ( .A1(n8991), .A2(n6947), .ZN(n7004) );
  AND2_X1 U8714 ( .A1(n6947), .A2(n8991), .ZN(n8916) );
  NOR2_X1 U8715 ( .A1(n7004), .A2(n8916), .ZN(n9556) );
  INV_X1 U8716 ( .A(n7003), .ZN(n6948) );
  NOR3_X1 U8717 ( .A1(n9556), .A2(n6948), .A3(n9561), .ZN(n6949) );
  AOI211_X1 U8718 ( .C1(n9541), .C2(P1_REG3_REG_0__SCAN_IN), .A(n9559), .B(
        n6949), .ZN(n6960) );
  INV_X1 U8719 ( .A(n9307), .ZN(n6951) );
  OAI21_X1 U8720 ( .B1(n6952), .B2(n9307), .A(n9555), .ZN(n6955) );
  NAND4_X1 U8721 ( .A1(n6955), .A2(n6954), .A3(n9313), .A4(n6953), .ZN(n6956)
         );
  NAND2_X1 U8722 ( .A1(n9301), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6959) );
  NOR2_X1 U8723 ( .A1(n9295), .A2(n9487), .ZN(n9179) );
  OAI21_X1 U8724 ( .B1(n9179), .B2(n9291), .A(n9560), .ZN(n6958) );
  OAI211_X1 U8725 ( .C1(n6960), .C2(n9553), .A(n6959), .B(n6958), .ZN(P1_U3293) );
  NAND2_X1 U8726 ( .A1(n6962), .A2(n6961), .ZN(n6964) );
  NAND2_X1 U8727 ( .A1(n6964), .A2(n6963), .ZN(n6968) );
  NAND2_X1 U8728 ( .A1(n7221), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6965) );
  OAI21_X1 U8729 ( .B1(n7221), .B2(P1_REG1_REG_16__SCAN_IN), .A(n6965), .ZN(
        n6966) );
  INV_X1 U8730 ( .A(n6966), .ZN(n6967) );
  NOR2_X1 U8731 ( .A1(n6967), .A2(n6968), .ZN(n7220) );
  AOI21_X1 U8732 ( .B1(n6968), .B2(n6967), .A(n7220), .ZN(n6981) );
  NOR2_X1 U8733 ( .A1(n6970), .A2(n6969), .ZN(n6972) );
  NOR2_X1 U8734 ( .A1(n6972), .A2(n6971), .ZN(n6975) );
  NAND2_X1 U8735 ( .A1(n7227), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6973) );
  OAI21_X1 U8736 ( .B1(n7227), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6973), .ZN(
        n6974) );
  NOR2_X1 U8737 ( .A1(n6975), .A2(n6974), .ZN(n7226) );
  AOI211_X1 U8738 ( .C1(n6975), .C2(n6974), .A(n7226), .B(n7300), .ZN(n6976)
         );
  INV_X1 U8739 ( .A(n6976), .ZN(n6980) );
  INV_X1 U8740 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8741 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8649) );
  OAI21_X1 U8742 ( .B1(n9026), .B2(n6977), .A(n8649), .ZN(n6978) );
  AOI21_X1 U8743 ( .B1(n7227), .B2(n9001), .A(n6978), .ZN(n6979) );
  OAI211_X1 U8744 ( .C1(n6981), .C2(n7429), .A(n6980), .B(n6979), .ZN(P1_U3259) );
  INV_X1 U8745 ( .A(n6987), .ZN(n6982) );
  XNOR2_X1 U8746 ( .A(n7118), .B(n7052), .ZN(n7115) );
  XNOR2_X1 U8747 ( .A(n7115), .B(n8111), .ZN(n6985) );
  NOR3_X1 U8748 ( .A1(n6983), .A2(n6982), .A3(n6985), .ZN(n6993) );
  INV_X1 U8749 ( .A(n6984), .ZN(n6991) );
  INV_X1 U8750 ( .A(n6985), .ZN(n6988) );
  NOR2_X1 U8751 ( .A1(n6986), .A2(n6988), .ZN(n6990) );
  INV_X1 U8752 ( .A(n7117), .ZN(n6992) );
  OAI21_X1 U8753 ( .B1(n6993), .B2(n6992), .A(n7866), .ZN(n6998) );
  NAND2_X1 U8754 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9751) );
  INV_X1 U8755 ( .A(n9751), .ZN(n6994) );
  AOI21_X1 U8756 ( .B1(n7858), .B2(n9885), .A(n6994), .ZN(n6995) );
  OAI21_X1 U8757 ( .B1(n7273), .B2(n7860), .A(n6995), .ZN(n6996) );
  AOI21_X1 U8758 ( .B1(n7052), .B2(n7850), .A(n6996), .ZN(n6997) );
  OAI211_X1 U8759 ( .C1(n7317), .C2(n7848), .A(n6998), .B(n6997), .ZN(P2_U3167) );
  NAND2_X1 U8760 ( .A1(n8991), .A2(n9560), .ZN(n7019) );
  XNOR2_X1 U8761 ( .A(n9569), .B(n9565), .ZN(n8844) );
  INV_X1 U8762 ( .A(n8844), .ZN(n7005) );
  XNOR2_X1 U8763 ( .A(n7019), .B(n7005), .ZN(n9563) );
  OR2_X1 U8764 ( .A1(n6999), .A2(n8972), .ZN(n7017) );
  NOR2_X1 U8765 ( .A1(n9553), .A2(n7017), .ZN(n9550) );
  INV_X1 U8766 ( .A(n9550), .ZN(n7180) );
  NAND2_X1 U8767 ( .A1(n7000), .A2(n5738), .ZN(n7001) );
  NAND3_X1 U8768 ( .A1(n7003), .A2(n7002), .A3(n7001), .ZN(n9318) );
  AOI22_X1 U8769 ( .A1(n9535), .A2(n8990), .B1(n8991), .B2(n9626), .ZN(n7009)
         );
  NAND2_X1 U8770 ( .A1(n7004), .A2(n7005), .ZN(n7025) );
  OAI21_X1 U8771 ( .B1(n7005), .B2(n7004), .A(n7025), .ZN(n7007) );
  NAND2_X1 U8772 ( .A1(n5737), .A2(n9493), .ZN(n7006) );
  NAND2_X1 U8773 ( .A1(n7007), .A2(n9486), .ZN(n7008) );
  OAI211_X1 U8774 ( .C1(n9563), .C2(n9318), .A(n7009), .B(n7008), .ZN(n9566)
         );
  NAND2_X1 U8775 ( .A1(n9566), .A2(n9494), .ZN(n7016) );
  XNOR2_X1 U8776 ( .A(n9560), .B(n9565), .ZN(n7010) );
  NAND2_X1 U8777 ( .A1(n7010), .A2(n9546), .ZN(n9564) );
  NOR2_X1 U8778 ( .A1(n9295), .A2(n9564), .ZN(n7014) );
  OAI22_X1 U8779 ( .A1(n9494), .A2(n7012), .B1(n7011), .B2(n9499), .ZN(n7013)
         );
  AOI211_X1 U8780 ( .C1(n9291), .C2(n8919), .A(n7014), .B(n7013), .ZN(n7015)
         );
  OAI211_X1 U8781 ( .C1(n9563), .C2(n7180), .A(n7016), .B(n7015), .ZN(P1_U3292) );
  AND2_X1 U8782 ( .A1(n9318), .A2(n7017), .ZN(n7018) );
  NAND2_X1 U8783 ( .A1(n8844), .A2(n7019), .ZN(n7021) );
  NAND2_X1 U8784 ( .A1(n8920), .A2(n9565), .ZN(n7020) );
  NAND2_X1 U8785 ( .A1(n7021), .A2(n7020), .ZN(n7071) );
  XNOR2_X1 U8786 ( .A(n7026), .B(n8990), .ZN(n7077) );
  NAND2_X1 U8787 ( .A1(n7071), .A2(n7077), .ZN(n7023) );
  NAND2_X1 U8788 ( .A1(n9580), .A2(n7026), .ZN(n7022) );
  NAND2_X1 U8789 ( .A1(n7023), .A2(n7022), .ZN(n7055) );
  XNOR2_X1 U8790 ( .A(n9579), .B(n9586), .ZN(n8845) );
  INV_X1 U8791 ( .A(n8845), .ZN(n7058) );
  XNOR2_X1 U8792 ( .A(n7055), .B(n7058), .ZN(n9578) );
  NAND2_X1 U8793 ( .A1(n8920), .A2(n8919), .ZN(n7024) );
  NAND2_X1 U8794 ( .A1(n7025), .A2(n7024), .ZN(n7078) );
  NAND2_X1 U8795 ( .A1(n7026), .A2(n8990), .ZN(n8922) );
  NAND2_X1 U8796 ( .A1(n7078), .A2(n8922), .ZN(n7028) );
  NAND2_X1 U8797 ( .A1(n9580), .A2(n9570), .ZN(n7027) );
  NAND2_X1 U8798 ( .A1(n7028), .A2(n7027), .ZN(n7059) );
  XNOR2_X1 U8799 ( .A(n7059), .B(n7058), .ZN(n7029) );
  AOI22_X1 U8800 ( .A1(n7029), .A2(n9486), .B1(n9535), .B2(n9595), .ZN(n9577)
         );
  MUX2_X1 U8801 ( .A(n6535), .B(n9577), .S(n9494), .Z(n7033) );
  AOI211_X1 U8802 ( .C1(n7060), .C2(n7073), .A(n9487), .B(n7066), .ZN(n9582)
         );
  NOR2_X1 U8803 ( .A1(n9248), .A2(n9580), .ZN(n7031) );
  OAI22_X1 U8804 ( .A1(n9544), .A2(n9579), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9499), .ZN(n7030) );
  AOI211_X1 U8805 ( .C1(n9582), .C2(n9549), .A(n7031), .B(n7030), .ZN(n7032)
         );
  OAI211_X1 U8806 ( .C1(n9286), .C2(n9578), .A(n7033), .B(n7032), .ZN(P1_U3290) );
  INV_X1 U8807 ( .A(n7034), .ZN(n7036) );
  NAND2_X1 U8808 ( .A1(n7036), .A2(n7035), .ZN(n7037) );
  XNOR2_X1 U8809 ( .A(n7038), .B(n7037), .ZN(n7042) );
  AND2_X1 U8810 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9056) );
  OAI22_X1 U8811 ( .A1(n9605), .A2(n8737), .B1(n8704), .B2(n7443), .ZN(n7039)
         );
  AOI211_X1 U8812 ( .C1(n7155), .C2(n5770), .A(n9056), .B(n7039), .ZN(n7041)
         );
  NAND2_X1 U8813 ( .A1(n8742), .A2(n7154), .ZN(n7040) );
  OAI211_X1 U8814 ( .C1(n7042), .C2(n8745), .A(n7041), .B(n7040), .ZN(P1_U3239) );
  INV_X1 U8815 ( .A(n7043), .ZN(n7044) );
  OR2_X1 U8816 ( .A1(n7045), .A2(n7044), .ZN(n7906) );
  XNOR2_X1 U8817 ( .A(n7046), .B(n7906), .ZN(n7321) );
  XNOR2_X1 U8818 ( .A(n7047), .B(n7906), .ZN(n7048) );
  OAI222_X1 U8819 ( .A1(n8349), .A2(n7273), .B1(n8351), .B2(n4753), .C1(n7048), 
        .C2(n8347), .ZN(n7316) );
  AOI21_X1 U8820 ( .B1(n9938), .B2(n7321), .A(n7316), .ZN(n7054) );
  INV_X1 U8821 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7049) );
  OAI22_X1 U8822 ( .A1(n7318), .A2(n8513), .B1(n9939), .B2(n7049), .ZN(n7050)
         );
  INV_X1 U8823 ( .A(n7050), .ZN(n7051) );
  OAI21_X1 U8824 ( .B1(n7054), .B2(n9941), .A(n7051), .ZN(P2_U3405) );
  AOI22_X1 U8825 ( .A1(n8432), .A2(n7052), .B1(n6296), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7053) );
  OAI21_X1 U8826 ( .B1(n7054), .B2(n6296), .A(n7053), .ZN(P2_U3464) );
  NAND2_X1 U8827 ( .A1(n7055), .A2(n8845), .ZN(n7057) );
  NAND2_X1 U8828 ( .A1(n7079), .A2(n9579), .ZN(n7056) );
  NAND2_X1 U8829 ( .A1(n7057), .A2(n7056), .ZN(n7084) );
  NAND2_X1 U8830 ( .A1(n7086), .A2(n9585), .ZN(n7090) );
  NAND2_X1 U8831 ( .A1(n7090), .A2(n8923), .ZN(n7083) );
  INV_X1 U8832 ( .A(n7083), .ZN(n8843) );
  XNOR2_X1 U8833 ( .A(n7084), .B(n8843), .ZN(n9589) );
  XNOR2_X1 U8834 ( .A(n7092), .B(n7083), .ZN(n7062) );
  OAI22_X1 U8835 ( .A1(n7062), .A2(n9557), .B1(n9605), .B2(n9277), .ZN(n9591)
         );
  NAND2_X1 U8836 ( .A1(n9591), .A2(n9494), .ZN(n7070) );
  INV_X1 U8837 ( .A(n9248), .ZN(n7102) );
  AOI22_X1 U8838 ( .A1(n9553), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7063), .B2(
        n9541), .ZN(n7064) );
  OAI21_X1 U8839 ( .B1(n9544), .B2(n7085), .A(n7064), .ZN(n7068) );
  AND2_X1 U8840 ( .A1(n7066), .A2(n7085), .ZN(n7099) );
  INV_X1 U8841 ( .A(n7099), .ZN(n7065) );
  OAI211_X1 U8842 ( .C1(n7085), .C2(n7066), .A(n7065), .B(n9546), .ZN(n9587)
         );
  NOR2_X1 U8843 ( .A1(n9587), .A2(n9295), .ZN(n7067) );
  AOI211_X1 U8844 ( .C1(n7102), .C2(n9586), .A(n7068), .B(n7067), .ZN(n7069)
         );
  OAI211_X1 U8845 ( .C1(n9589), .C2(n9286), .A(n7070), .B(n7069), .ZN(P1_U3289) );
  INV_X1 U8846 ( .A(n7077), .ZN(n8846) );
  XNOR2_X1 U8847 ( .A(n7071), .B(n8846), .ZN(n9573) );
  INV_X1 U8848 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8998) );
  OAI22_X1 U8849 ( .A1(n9494), .A2(n7072), .B1(n8998), .B2(n9499), .ZN(n7076)
         );
  OAI21_X1 U8850 ( .B1(n9560), .B2(n8919), .A(n9570), .ZN(n7074) );
  NAND3_X1 U8851 ( .A1(n7074), .A2(n9546), .A3(n7073), .ZN(n9571) );
  OAI22_X1 U8852 ( .A1(n9571), .A2(n9295), .B1(n9248), .B2(n8920), .ZN(n7075)
         );
  AOI211_X1 U8853 ( .C1(n9291), .C2(n9570), .A(n7076), .B(n7075), .ZN(n7082)
         );
  XNOR2_X1 U8854 ( .A(n7078), .B(n7077), .ZN(n7080) );
  OAI22_X1 U8855 ( .A1(n7080), .A2(n9557), .B1(n7079), .B2(n9277), .ZN(n9575)
         );
  NAND2_X1 U8856 ( .A1(n9575), .A2(n9494), .ZN(n7081) );
  OAI211_X1 U8857 ( .C1(n9573), .C2(n9286), .A(n7082), .B(n7081), .ZN(P1_U3291) );
  NAND2_X1 U8858 ( .A1(n7084), .A2(n7083), .ZN(n7088) );
  NAND2_X1 U8859 ( .A1(n7086), .A2(n7085), .ZN(n7087) );
  NAND2_X1 U8860 ( .A1(n7088), .A2(n7087), .ZN(n7147) );
  NAND2_X1 U8861 ( .A1(n9605), .A2(n9594), .ZN(n7089) );
  NAND2_X1 U8862 ( .A1(n7148), .A2(n8989), .ZN(n8924) );
  NAND2_X1 U8863 ( .A1(n7089), .A2(n8924), .ZN(n8840) );
  INV_X1 U8864 ( .A(n8840), .ZN(n7094) );
  XNOR2_X1 U8865 ( .A(n7147), .B(n7094), .ZN(n9593) );
  INV_X1 U8866 ( .A(n7090), .ZN(n7091) );
  NAND2_X1 U8867 ( .A1(n7093), .A2(n7094), .ZN(n7151) );
  NOR2_X1 U8868 ( .A1(n7094), .A2(n4689), .ZN(n7095) );
  AOI21_X1 U8869 ( .B1(n7096), .B2(n7095), .A(n9557), .ZN(n7097) );
  INV_X1 U8870 ( .A(n7162), .ZN(n9536) );
  AOI22_X1 U8871 ( .A1(n7151), .A2(n7097), .B1(n9535), .B2(n9536), .ZN(n9598)
         );
  MUX2_X1 U8872 ( .A(n10176), .B(n9598), .S(n9494), .Z(n7104) );
  OAI22_X1 U8873 ( .A1(n9544), .A2(n7148), .B1(n7098), .B2(n9499), .ZN(n7101)
         );
  OAI211_X1 U8874 ( .C1(n7099), .C2(n7148), .A(n9546), .B(n7153), .ZN(n9596)
         );
  NOR2_X1 U8875 ( .A1(n9596), .A2(n9295), .ZN(n7100) );
  AOI211_X1 U8876 ( .C1(n7102), .C2(n9595), .A(n7101), .B(n7100), .ZN(n7103)
         );
  OAI211_X1 U8877 ( .C1(n9593), .C2(n9286), .A(n7104), .B(n7103), .ZN(P1_U3288) );
  INV_X1 U8878 ( .A(n7105), .ZN(n7106) );
  XNOR2_X1 U8879 ( .A(n7107), .B(n7106), .ZN(n7108) );
  XNOR2_X1 U8880 ( .A(n4515), .B(n7108), .ZN(n7113) );
  INV_X1 U8881 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U8882 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10231), .ZN(n9072) );
  OAI22_X1 U8883 ( .A1(n7162), .A2(n8737), .B1(n8704), .B2(n7254), .ZN(n7110)
         );
  AOI211_X1 U8884 ( .C1(n7165), .C2(n5770), .A(n9072), .B(n7110), .ZN(n7112)
         );
  NAND2_X1 U8885 ( .A1(n8742), .A2(n9542), .ZN(n7111) );
  OAI211_X1 U8886 ( .C1(n7113), .C2(n8745), .A(n7112), .B(n7111), .ZN(P1_U3213) );
  NAND2_X1 U8887 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  NAND2_X1 U8888 ( .A1(n7117), .A2(n7116), .ZN(n7119) );
  CLKBUF_X3 U8889 ( .A(n7118), .Z(n7664) );
  XNOR2_X1 U8890 ( .A(n7664), .B(n9906), .ZN(n7234) );
  XNOR2_X1 U8891 ( .A(n7234), .B(n8110), .ZN(n7120) );
  AOI21_X1 U8892 ( .B1(n7119), .B2(n7120), .A(n7852), .ZN(n7122) );
  NAND2_X1 U8893 ( .A1(n7122), .A2(n7236), .ZN(n7127) );
  INV_X1 U8894 ( .A(n8109), .ZN(n7237) );
  NAND2_X1 U8895 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9767) );
  INV_X1 U8896 ( .A(n9767), .ZN(n7123) );
  AOI21_X1 U8897 ( .B1(n7858), .B2(n8111), .A(n7123), .ZN(n7124) );
  OAI21_X1 U8898 ( .B1(n7237), .B2(n7860), .A(n7124), .ZN(n7125) );
  AOI21_X1 U8899 ( .B1(n7137), .B2(n7850), .A(n7125), .ZN(n7126) );
  OAI211_X1 U8900 ( .C1(n7135), .C2(n7848), .A(n7127), .B(n7126), .ZN(P2_U3179) );
  NAND2_X1 U8901 ( .A1(n6220), .A2(n7959), .ZN(n7909) );
  XOR2_X1 U8902 ( .A(n7909), .B(n7128), .Z(n9907) );
  INV_X1 U8903 ( .A(n7909), .ZN(n7130) );
  XNOR2_X1 U8904 ( .A(n7129), .B(n7130), .ZN(n7131) );
  NAND2_X1 U8905 ( .A1(n7131), .A2(n6212), .ZN(n7133) );
  AOI22_X1 U8906 ( .A1(n9883), .A2(n8111), .B1(n8109), .B2(n8370), .ZN(n7132)
         );
  AND2_X1 U8907 ( .A1(n7133), .A2(n7132), .ZN(n9905) );
  MUX2_X1 U8908 ( .A(n7134), .B(n9905), .S(n8373), .Z(n7139) );
  INV_X1 U8909 ( .A(n7135), .ZN(n7136) );
  AOI22_X1 U8910 ( .A1(n9889), .A2(n7137), .B1(n9890), .B2(n7136), .ZN(n7138)
         );
  OAI211_X1 U8911 ( .C1(n9907), .C2(n8378), .A(n7139), .B(n7138), .ZN(P2_U3227) );
  OAI22_X1 U8912 ( .A1(n8288), .A2(n7141), .B1(n7140), .B2(n8355), .ZN(n7144)
         );
  NOR2_X1 U8913 ( .A1(n7142), .A2(n8340), .ZN(n7143) );
  AOI211_X1 U8914 ( .C1(n8340), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7144), .B(
        n7143), .ZN(n7145) );
  OAI21_X1 U8915 ( .B1(n8378), .B2(n7146), .A(n7145), .ZN(P2_U3232) );
  NAND2_X1 U8916 ( .A1(n7147), .A2(n8840), .ZN(n7150) );
  NAND2_X1 U8917 ( .A1(n9605), .A2(n7148), .ZN(n7149) );
  NAND2_X1 U8918 ( .A1(n7150), .A2(n7149), .ZN(n7161) );
  NAND2_X1 U8919 ( .A1(n7162), .A2(n7155), .ZN(n7168) );
  INV_X1 U8920 ( .A(n7155), .ZN(n9604) );
  NAND2_X1 U8921 ( .A1(n9604), .A2(n9536), .ZN(n7186) );
  NAND2_X1 U8922 ( .A1(n7168), .A2(n7186), .ZN(n7160) );
  INV_X1 U8923 ( .A(n7160), .ZN(n8841) );
  XNOR2_X1 U8924 ( .A(n7161), .B(n8841), .ZN(n9603) );
  XNOR2_X1 U8925 ( .A(n7169), .B(n7160), .ZN(n7152) );
  AOI22_X1 U8926 ( .A1(n7152), .A2(n9486), .B1(n9535), .B2(n8988), .ZN(n9602)
         );
  MUX2_X1 U8927 ( .A(n10157), .B(n9602), .S(n9494), .Z(n7159) );
  AOI211_X1 U8928 ( .C1(n7155), .C2(n7153), .A(n9487), .B(n4496), .ZN(n9607)
         );
  AOI22_X1 U8929 ( .A1(n9291), .A2(n7155), .B1(n7154), .B2(n9541), .ZN(n7156)
         );
  OAI21_X1 U8930 ( .B1(n9605), .B2(n9248), .A(n7156), .ZN(n7157) );
  AOI21_X1 U8931 ( .B1(n9607), .B2(n9549), .A(n7157), .ZN(n7158) );
  OAI211_X1 U8932 ( .C1(n9603), .C2(n9286), .A(n7159), .B(n7158), .ZN(P1_U3287) );
  NAND2_X1 U8933 ( .A1(n7254), .A2(n7177), .ZN(n7247) );
  NAND2_X1 U8934 ( .A1(n7247), .A2(n7249), .ZN(n7191) );
  NAND2_X1 U8935 ( .A1(n7161), .A2(n7160), .ZN(n7164) );
  NAND2_X1 U8936 ( .A1(n7162), .A2(n9604), .ZN(n7163) );
  NAND2_X1 U8937 ( .A1(n7164), .A2(n7163), .ZN(n9531) );
  NAND2_X1 U8938 ( .A1(n7443), .A2(n7165), .ZN(n7181) );
  NAND2_X1 U8939 ( .A1(n9612), .A2(n8988), .ZN(n7184) );
  NAND2_X1 U8940 ( .A1(n7181), .A2(n7184), .ZN(n9532) );
  NAND2_X1 U8941 ( .A1(n9531), .A2(n9532), .ZN(n7167) );
  NAND2_X1 U8942 ( .A1(n7443), .A2(n9612), .ZN(n7166) );
  XOR2_X1 U8943 ( .A(n7191), .B(n7192), .Z(n9617) );
  XOR2_X1 U8944 ( .A(n7191), .B(n7248), .Z(n7171) );
  OAI22_X1 U8945 ( .A1(n7443), .A2(n9656), .B1(n7447), .B2(n9277), .ZN(n7170)
         );
  AOI21_X1 U8946 ( .B1(n7171), .B2(n9486), .A(n7170), .ZN(n7172) );
  OAI21_X1 U8947 ( .B1(n9617), .B2(n9318), .A(n7172), .ZN(n9620) );
  NAND2_X1 U8948 ( .A1(n9620), .A2(n9494), .ZN(n7179) );
  INV_X1 U8949 ( .A(n7173), .ZN(n7452) );
  OAI22_X1 U8950 ( .A1(n9494), .A2(n10230), .B1(n7452), .B2(n9499), .ZN(n7176)
         );
  INV_X1 U8951 ( .A(n9547), .ZN(n7174) );
  OAI211_X1 U8952 ( .C1(n7174), .C2(n9619), .A(n9546), .B(n7255), .ZN(n9618)
         );
  NOR2_X1 U8953 ( .A1(n9618), .A2(n9295), .ZN(n7175) );
  AOI211_X1 U8954 ( .C1(n9291), .C2(n7177), .A(n7176), .B(n7175), .ZN(n7178)
         );
  OAI211_X1 U8955 ( .C1(n9617), .C2(n7180), .A(n7179), .B(n7178), .ZN(P1_U3285) );
  NAND2_X1 U8956 ( .A1(n7447), .A2(n9624), .ZN(n8757) );
  NAND2_X1 U8957 ( .A1(n8757), .A2(n7247), .ZN(n8753) );
  INV_X1 U8958 ( .A(n7181), .ZN(n7182) );
  INV_X1 U8959 ( .A(n7447), .ZN(n8987) );
  NAND2_X1 U8960 ( .A1(n8765), .A2(n7249), .ZN(n8749) );
  NAND2_X1 U8961 ( .A1(n8749), .A2(n8757), .ZN(n7183) );
  NAND2_X1 U8962 ( .A1(n7249), .A2(n7184), .ZN(n8752) );
  INV_X1 U8963 ( .A(n8765), .ZN(n7185) );
  NAND2_X1 U8964 ( .A1(n9636), .A2(n8986), .ZN(n8929) );
  NAND2_X1 U8965 ( .A1(n7404), .A2(n7548), .ZN(n8764) );
  NAND2_X1 U8966 ( .A1(n8929), .A2(n8764), .ZN(n8851) );
  NAND2_X1 U8967 ( .A1(n7187), .A2(n8851), .ZN(n7188) );
  NAND2_X1 U8968 ( .A1(n7210), .A2(n7188), .ZN(n7190) );
  OAI22_X1 U8969 ( .A1(n7447), .A2(n9656), .B1(n7546), .B2(n9277), .ZN(n7189)
         );
  AOI21_X1 U8970 ( .B1(n7190), .B2(n9486), .A(n7189), .ZN(n9635) );
  NAND2_X1 U8971 ( .A1(n7254), .A2(n9619), .ZN(n7193) );
  NAND2_X1 U8972 ( .A1(n8757), .A2(n8765), .ZN(n7251) );
  XNOR2_X1 U8973 ( .A(n7207), .B(n8851), .ZN(n9638) );
  NAND2_X1 U8974 ( .A1(n9638), .A2(n9480), .ZN(n7200) );
  OAI22_X1 U8975 ( .A1(n9494), .A2(n6570), .B1(n7195), .B2(n9499), .ZN(n7198)
         );
  OR2_X1 U8976 ( .A1(n7255), .A2(n9624), .ZN(n7256) );
  XNOR2_X1 U8977 ( .A(n7256), .B(n9636), .ZN(n7196) );
  NAND2_X1 U8978 ( .A1(n7196), .A2(n9546), .ZN(n9634) );
  NOR2_X1 U8979 ( .A1(n9634), .A2(n9295), .ZN(n7197) );
  AOI211_X1 U8980 ( .C1(n9291), .C2(n7548), .A(n7198), .B(n7197), .ZN(n7199)
         );
  OAI211_X1 U8981 ( .C1(n9301), .C2(n9635), .A(n7200), .B(n7199), .ZN(P1_U3283) );
  NAND2_X1 U8982 ( .A1(n7204), .A2(n7508), .ZN(n7202) );
  OAI211_X1 U8983 ( .C1(n7203), .C2(n7618), .A(n7202), .B(n7201), .ZN(P1_U3335) );
  INV_X1 U8984 ( .A(n7204), .ZN(n7206) );
  OAI222_X1 U8985 ( .A1(n8550), .A2(n7206), .B1(P2_U3151), .B2(n8088), .C1(
        n7205), .C2(n8547), .ZN(P2_U3275) );
  NAND2_X1 U8986 ( .A1(n7207), .A2(n8851), .ZN(n7209) );
  NAND2_X1 U8987 ( .A1(n9636), .A2(n7404), .ZN(n7208) );
  NAND2_X1 U8988 ( .A1(n7209), .A2(n7208), .ZN(n7333) );
  OR2_X1 U8989 ( .A1(n8706), .A2(n7546), .ZN(n8767) );
  NAND2_X1 U8990 ( .A1(n8706), .A2(n7546), .ZN(n8768) );
  NAND2_X1 U8991 ( .A1(n8767), .A2(n8768), .ZN(n8852) );
  XNOR2_X1 U8992 ( .A(n7333), .B(n8852), .ZN(n9643) );
  INV_X1 U8993 ( .A(n9318), .ZN(n9540) );
  NAND2_X1 U8994 ( .A1(n7210), .A2(n8764), .ZN(n7338) );
  XNOR2_X1 U8995 ( .A(n7338), .B(n8852), .ZN(n7212) );
  INV_X1 U8996 ( .A(n9657), .ZN(n8984) );
  AOI22_X1 U8997 ( .A1(n8984), .A2(n9535), .B1(n9626), .B2(n8986), .ZN(n7211)
         );
  OAI21_X1 U8998 ( .B1(n7212), .B2(n9557), .A(n7211), .ZN(n7213) );
  AOI21_X1 U8999 ( .B1(n9643), .B2(n9540), .A(n7213), .ZN(n9645) );
  INV_X1 U9000 ( .A(n8706), .ZN(n9641) );
  NAND2_X1 U9001 ( .A1(n7214), .A2(n9641), .ZN(n7351) );
  OAI211_X1 U9002 ( .C1(n7214), .C2(n9641), .A(n9546), .B(n7351), .ZN(n9640)
         );
  AOI22_X1 U9003 ( .A1(n9301), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8701), .B2(
        n9541), .ZN(n7216) );
  NAND2_X1 U9004 ( .A1(n9291), .A2(n8706), .ZN(n7215) );
  OAI211_X1 U9005 ( .C1(n9640), .C2(n9295), .A(n7216), .B(n7215), .ZN(n7217)
         );
  AOI21_X1 U9006 ( .B1(n9643), .B2(n9550), .A(n7217), .ZN(n7218) );
  OAI21_X1 U9007 ( .B1(n9645), .B2(n9301), .A(n7218), .ZN(P1_U3282) );
  NOR2_X1 U9008 ( .A1(n7305), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7219) );
  AOI21_X1 U9009 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n7305), .A(n7219), .ZN(
        n7223) );
  INV_X1 U9010 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9519) );
  AOI21_X1 U9011 ( .B1(n7221), .B2(n9519), .A(n7220), .ZN(n7222) );
  NOR2_X1 U9012 ( .A1(n7222), .A2(n7223), .ZN(n7306) );
  AOI21_X1 U9013 ( .B1(n7223), .B2(n7222), .A(n7306), .ZN(n7225) );
  NAND2_X1 U9014 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U9015 ( .A1(n9073), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n7224) );
  OAI211_X1 U9016 ( .C1(n7429), .C2(n7225), .A(n8659), .B(n7224), .ZN(n7232)
         );
  AOI21_X1 U9017 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n7227), .A(n7226), .ZN(
        n7230) );
  NOR2_X1 U9018 ( .A1(n7296), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7228) );
  AOI21_X1 U9019 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n7296), .A(n7228), .ZN(
        n7229) );
  NAND2_X1 U9020 ( .A1(n7229), .A2(n7230), .ZN(n7295) );
  AOI221_X1 U9021 ( .B1(n7230), .B2(n7295), .C1(n7229), .C2(n7295), .A(n7300), 
        .ZN(n7231) );
  AOI211_X1 U9022 ( .C1(n9001), .C2(n7296), .A(n7232), .B(n7231), .ZN(n7233)
         );
  INV_X1 U9023 ( .A(n7233), .ZN(P1_U3260) );
  NAND2_X1 U9024 ( .A1(n7234), .A2(n8110), .ZN(n7235) );
  XNOR2_X1 U9025 ( .A(n7664), .B(n7275), .ZN(n7360) );
  XNOR2_X1 U9026 ( .A(n7360), .B(n7237), .ZN(n7238) );
  OAI21_X1 U9027 ( .B1(n7239), .B2(n7238), .A(n7361), .ZN(n7240) );
  NAND2_X1 U9028 ( .A1(n7240), .A2(n7866), .ZN(n7245) );
  INV_X1 U9029 ( .A(n8108), .ZN(n7363) );
  AOI21_X1 U9030 ( .B1(n7858), .B2(n8110), .A(n7241), .ZN(n7242) );
  OAI21_X1 U9031 ( .B1(n7363), .B2(n7860), .A(n7242), .ZN(n7243) );
  AOI21_X1 U9032 ( .B1(n9917), .B2(n7850), .A(n7243), .ZN(n7244) );
  OAI211_X1 U9033 ( .C1(n7274), .C2(n7848), .A(n7245), .B(n7244), .ZN(P2_U3153) );
  XOR2_X1 U9034 ( .A(n7251), .B(n7246), .Z(n9630) );
  NAND2_X1 U9035 ( .A1(n8751), .A2(n7249), .ZN(n7250) );
  XOR2_X1 U9036 ( .A(n7251), .B(n7250), .Z(n7252) );
  NOR2_X1 U9037 ( .A1(n7252), .A2(n9557), .ZN(n9632) );
  NAND2_X1 U9038 ( .A1(n9632), .A2(n9494), .ZN(n7261) );
  AOI22_X1 U9039 ( .A1(n9301), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7401), .B2(
        n9541), .ZN(n7253) );
  OAI21_X1 U9040 ( .B1(n9248), .B2(n7254), .A(n7253), .ZN(n7259) );
  AOI21_X1 U9041 ( .B1(n7255), .B2(n9624), .A(n9487), .ZN(n7257) );
  AOI22_X1 U9042 ( .A1(n7257), .A2(n7256), .B1(n9535), .B2(n8986), .ZN(n9629)
         );
  NOR2_X1 U9043 ( .A1(n9629), .A2(n9295), .ZN(n7258) );
  AOI211_X1 U9044 ( .C1(n9291), .C2(n9624), .A(n7259), .B(n7258), .ZN(n7260)
         );
  OAI211_X1 U9045 ( .C1(n9630), .C2(n9286), .A(n7261), .B(n7260), .ZN(P1_U3284) );
  NAND2_X1 U9046 ( .A1(n8373), .A2(n7262), .ZN(n8162) );
  OAI22_X1 U9047 ( .A1(n8355), .A2(n7264), .B1(n7263), .B2(n8336), .ZN(n7265)
         );
  NOR2_X1 U9048 ( .A1(n7266), .A2(n7265), .ZN(n7268) );
  MUX2_X1 U9049 ( .A(n7268), .B(n7267), .S(n8340), .Z(n7269) );
  OAI21_X1 U9050 ( .B1(n7270), .B2(n8162), .A(n7269), .ZN(P2_U3231) );
  XNOR2_X1 U9051 ( .A(n7271), .B(n7976), .ZN(n7272) );
  OAI222_X1 U9052 ( .A1(n8351), .A2(n7273), .B1(n8349), .B2(n7363), .C1(n8347), 
        .C2(n7272), .ZN(n9915) );
  INV_X1 U9053 ( .A(n9915), .ZN(n7282) );
  OAI22_X1 U9054 ( .A1(n8288), .A2(n7275), .B1(n7274), .B2(n8355), .ZN(n7277)
         );
  NOR2_X1 U9055 ( .A1(n8373), .A2(n4726), .ZN(n7276) );
  NOR2_X1 U9056 ( .A1(n7277), .A2(n7276), .ZN(n7281) );
  NOR2_X1 U9057 ( .A1(n7278), .A2(n7976), .ZN(n9914) );
  INV_X1 U9058 ( .A(n9914), .ZN(n7279) );
  NAND3_X1 U9059 ( .A1(n7279), .A2(n9892), .A3(n9911), .ZN(n7280) );
  OAI211_X1 U9060 ( .C1(n7282), .C2(n8340), .A(n7281), .B(n7280), .ZN(P2_U3226) );
  INV_X1 U9061 ( .A(n7283), .ZN(n7284) );
  AOI21_X1 U9062 ( .B1(n7286), .B2(n7285), .A(n7284), .ZN(n7287) );
  MUX2_X1 U9063 ( .A(n7288), .B(n7287), .S(n8373), .Z(n7290) );
  NAND2_X1 U9064 ( .A1(n9890), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7289) );
  OAI211_X1 U9065 ( .C1(n8288), .C2(n7291), .A(n7290), .B(n7289), .ZN(P2_U3233) );
  INV_X1 U9066 ( .A(n7292), .ZN(n7293) );
  OAI222_X1 U9067 ( .A1(n8550), .A2(n7293), .B1(P2_U3151), .B2(n7913), .C1(
        n10110), .C2(n8547), .ZN(P2_U3274) );
  OAI222_X1 U9068 ( .A1(n7618), .A2(n7294), .B1(n9411), .B2(n7293), .C1(n8835), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U9069 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8724) );
  INV_X1 U9070 ( .A(n8724), .ZN(n7304) );
  OAI21_X1 U9071 ( .B1(n7296), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7295), .ZN(
        n7302) );
  NAND2_X1 U9072 ( .A1(n7315), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7299) );
  INV_X1 U9073 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U9074 ( .A1(n7418), .A2(n7297), .ZN(n7298) );
  AND2_X1 U9075 ( .A1(n7299), .A2(n7298), .ZN(n7301) );
  NOR2_X1 U9076 ( .A1(n7302), .A2(n7301), .ZN(n7420) );
  AOI211_X1 U9077 ( .C1(n7302), .C2(n7301), .A(n7420), .B(n7300), .ZN(n7303)
         );
  AOI211_X1 U9078 ( .C1(n9073), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n7304), .B(
        n7303), .ZN(n7314) );
  INV_X1 U9079 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U9080 ( .A1(n7315), .A2(n9506), .ZN(n7307) );
  INV_X1 U9081 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U9082 ( .A1(n7305), .A2(n10221), .ZN(n7309) );
  NAND2_X1 U9083 ( .A1(n7418), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7423) );
  INV_X1 U9084 ( .A(n7306), .ZN(n7308) );
  NAND4_X1 U9085 ( .A1(n7307), .A2(n7309), .A3(n7423), .A4(n7308), .ZN(n7424)
         );
  NAND2_X1 U9086 ( .A1(n7315), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U9087 ( .A1(n7309), .A2(n7308), .ZN(n7310) );
  OAI211_X1 U9088 ( .C1(n7315), .C2(P1_REG1_REG_18__SCAN_IN), .A(n7311), .B(
        n7310), .ZN(n7312) );
  NAND3_X1 U9089 ( .A1(n9084), .A2(n7424), .A3(n7312), .ZN(n7313) );
  OAI211_X1 U9090 ( .C1(n9070), .C2(n7315), .A(n7314), .B(n7313), .ZN(P1_U3261) );
  INV_X1 U9091 ( .A(n7316), .ZN(n7323) );
  NOR2_X1 U9092 ( .A1(n8373), .A2(n5905), .ZN(n7320) );
  OAI22_X1 U9093 ( .A1(n8288), .A2(n7318), .B1(n7317), .B2(n8355), .ZN(n7319)
         );
  AOI211_X1 U9094 ( .C1(n7321), .C2(n9892), .A(n7320), .B(n7319), .ZN(n7322)
         );
  OAI21_X1 U9095 ( .B1(n7323), .B2(n8340), .A(n7322), .ZN(P2_U3228) );
  OAI211_X1 U9096 ( .C1(n4498), .C2(n5958), .A(n6212), .B(n7324), .ZN(n7326)
         );
  AOI22_X1 U9097 ( .A1(n9883), .A2(n8109), .B1(n8107), .B2(n8370), .ZN(n7325)
         );
  NAND2_X1 U9098 ( .A1(n7326), .A2(n7325), .ZN(n9920) );
  INV_X1 U9099 ( .A(n9920), .ZN(n7332) );
  NAND2_X1 U9100 ( .A1(n9911), .A2(n7327), .ZN(n7328) );
  XOR2_X1 U9101 ( .A(n7918), .B(n7328), .Z(n9922) );
  NOR2_X1 U9102 ( .A1(n8373), .A2(n5946), .ZN(n7330) );
  OAI22_X1 U9103 ( .A1(n8288), .A2(n9919), .B1(n7371), .B2(n8355), .ZN(n7329)
         );
  AOI211_X1 U9104 ( .C1(n9922), .C2(n9892), .A(n7330), .B(n7329), .ZN(n7331)
         );
  OAI21_X1 U9105 ( .B1(n7332), .B2(n8340), .A(n7331), .ZN(P2_U3225) );
  NAND2_X1 U9106 ( .A1(n7333), .A2(n8852), .ZN(n7335) );
  OR2_X1 U9107 ( .A1(n8706), .A2(n8985), .ZN(n7334) );
  NAND2_X1 U9108 ( .A1(n7335), .A2(n7334), .ZN(n7346) );
  OR2_X1 U9109 ( .A1(n7354), .A2(n9657), .ZN(n8770) );
  NAND2_X1 U9110 ( .A1(n7354), .A2(n9657), .ZN(n8936) );
  NAND2_X1 U9111 ( .A1(n8770), .A2(n8936), .ZN(n8854) );
  NAND2_X1 U9112 ( .A1(n7346), .A2(n8854), .ZN(n7337) );
  OR2_X1 U9113 ( .A1(n7354), .A2(n8984), .ZN(n7336) );
  OR2_X1 U9114 ( .A1(n7621), .A2(n8633), .ZN(n8939) );
  NAND2_X1 U9115 ( .A1(n7621), .A2(n8633), .ZN(n8937) );
  NAND2_X1 U9116 ( .A1(n8939), .A2(n8937), .ZN(n7455) );
  INV_X1 U9117 ( .A(n7455), .ZN(n8855) );
  XNOR2_X1 U9118 ( .A(n7456), .B(n8855), .ZN(n9655) );
  NAND3_X1 U9119 ( .A1(n7347), .A2(n8936), .A3(n7455), .ZN(n7339) );
  AND2_X1 U9120 ( .A1(n7457), .A2(n7339), .ZN(n7340) );
  OAI22_X1 U9121 ( .A1(n7340), .A2(n9557), .B1(n8738), .B2(n9277), .ZN(n9661)
         );
  NAND2_X1 U9122 ( .A1(n9661), .A2(n9494), .ZN(n7345) );
  AOI211_X1 U9123 ( .C1(n7621), .C2(n7352), .A(n9487), .B(n7463), .ZN(n9660)
         );
  NAND2_X1 U9124 ( .A1(n7621), .A2(n9291), .ZN(n7342) );
  AOI22_X1 U9125 ( .A1(n9301), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7632), .B2(
        n9541), .ZN(n7341) );
  OAI211_X1 U9126 ( .C1(n9657), .C2(n9248), .A(n7342), .B(n7341), .ZN(n7343)
         );
  AOI21_X1 U9127 ( .B1(n9660), .B2(n9549), .A(n7343), .ZN(n7344) );
  OAI211_X1 U9128 ( .C1(n9655), .C2(n9286), .A(n7345), .B(n7344), .ZN(P1_U3280) );
  XNOR2_X1 U9129 ( .A(n7346), .B(n8854), .ZN(n9651) );
  INV_X1 U9130 ( .A(n9651), .ZN(n7359) );
  INV_X1 U9131 ( .A(n7347), .ZN(n7348) );
  AOI21_X1 U9132 ( .B1(n8854), .B2(n7349), .A(n7348), .ZN(n7350) );
  OAI222_X1 U9133 ( .A1(n9277), .A2(n8633), .B1(n9656), .B2(n7546), .C1(n9557), 
        .C2(n7350), .ZN(n9649) );
  INV_X1 U9134 ( .A(n7351), .ZN(n7353) );
  INV_X1 U9135 ( .A(n7354), .ZN(n9648) );
  OAI211_X1 U9136 ( .C1(n7353), .C2(n9648), .A(n9546), .B(n7352), .ZN(n9647)
         );
  AOI22_X1 U9137 ( .A1(n9553), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8635), .B2(
        n9541), .ZN(n7356) );
  NAND2_X1 U9138 ( .A1(n7354), .A2(n9291), .ZN(n7355) );
  OAI211_X1 U9139 ( .C1(n9647), .C2(n9295), .A(n7356), .B(n7355), .ZN(n7357)
         );
  AOI21_X1 U9140 ( .B1(n9649), .B2(n9494), .A(n7357), .ZN(n7358) );
  OAI21_X1 U9141 ( .B1(n7359), .B2(n9286), .A(n7358), .ZN(P1_U3281) );
  XNOR2_X1 U9142 ( .A(n7664), .B(n9919), .ZN(n7470) );
  OAI21_X1 U9143 ( .B1(n7363), .B2(n7362), .A(n7473), .ZN(n7364) );
  NAND2_X1 U9144 ( .A1(n7364), .A2(n7866), .ZN(n7370) );
  INV_X1 U9145 ( .A(n8107), .ZN(n7412) );
  NAND2_X1 U9146 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9784) );
  INV_X1 U9147 ( .A(n9784), .ZN(n7365) );
  AOI21_X1 U9148 ( .B1(n7858), .B2(n8109), .A(n7365), .ZN(n7366) );
  OAI21_X1 U9149 ( .B1(n7412), .B2(n7860), .A(n7366), .ZN(n7367) );
  AOI21_X1 U9150 ( .B1(n7368), .B2(n7850), .A(n7367), .ZN(n7369) );
  OAI211_X1 U9151 ( .C1(n7371), .C2(n7848), .A(n7370), .B(n7369), .ZN(P2_U3161) );
  OAI211_X1 U9152 ( .C1(n7373), .C2(n7923), .A(n7372), .B(n6212), .ZN(n7375)
         );
  AOI22_X1 U9153 ( .A1(n9883), .A2(n8106), .B1(n8105), .B2(n8370), .ZN(n7374)
         );
  NAND2_X1 U9154 ( .A1(n7375), .A2(n7374), .ZN(n9935) );
  INV_X1 U9155 ( .A(n9935), .ZN(n7382) );
  OAI21_X1 U9156 ( .B1(n7376), .B2(n7638), .A(n8361), .ZN(n9937) );
  INV_X1 U9157 ( .A(n7377), .ZN(n9934) );
  INV_X1 U9158 ( .A(n7378), .ZN(n7840) );
  AOI22_X1 U9159 ( .A1(n8340), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n9890), .B2(
        n7840), .ZN(n7379) );
  OAI21_X1 U9160 ( .B1(n9934), .B2(n8288), .A(n7379), .ZN(n7380) );
  AOI21_X1 U9161 ( .B1(n9937), .B2(n9892), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9162 ( .B1(n7382), .B2(n8340), .A(n7381), .ZN(P2_U3222) );
  OAI21_X1 U9163 ( .B1(n7384), .B2(n7920), .A(n7383), .ZN(n9926) );
  XNOR2_X1 U9164 ( .A(n7385), .B(n7920), .ZN(n7386) );
  NAND2_X1 U9165 ( .A1(n7386), .A2(n6212), .ZN(n7388) );
  AOI22_X1 U9166 ( .A1(n8370), .A2(n8106), .B1(n8108), .B2(n9883), .ZN(n7387)
         );
  OAI211_X1 U9167 ( .C1(n7389), .C2(n9926), .A(n7388), .B(n7387), .ZN(n9928)
         );
  NAND2_X1 U9168 ( .A1(n9928), .A2(n8373), .ZN(n7392) );
  OAI22_X1 U9169 ( .A1(n8373), .A2(n6303), .B1(n7484), .B2(n8355), .ZN(n7390)
         );
  AOI21_X1 U9170 ( .B1(n9889), .B2(n7481), .A(n7390), .ZN(n7391) );
  OAI211_X1 U9171 ( .C1(n9926), .C2(n8162), .A(n7392), .B(n7391), .ZN(P2_U3224) );
  NOR2_X1 U9172 ( .A1(n7394), .A2(n7393), .ZN(n7396) );
  AOI21_X1 U9173 ( .B1(n7394), .B2(n7393), .A(n7396), .ZN(n7441) );
  NAND2_X1 U9174 ( .A1(n7441), .A2(n5299), .ZN(n7440) );
  NOR2_X1 U9175 ( .A1(n7396), .A2(n7395), .ZN(n7399) );
  INV_X1 U9176 ( .A(n7397), .ZN(n7398) );
  AOI21_X1 U9177 ( .B1(n7440), .B2(n7399), .A(n7398), .ZN(n7407) );
  AOI21_X1 U9178 ( .B1(n8714), .B2(n9627), .A(n7400), .ZN(n7403) );
  NAND2_X1 U9179 ( .A1(n8742), .A2(n7401), .ZN(n7402) );
  OAI211_X1 U9180 ( .C1(n7404), .C2(n8704), .A(n7403), .B(n7402), .ZN(n7405)
         );
  AOI21_X1 U9181 ( .B1(n9624), .B2(n5770), .A(n7405), .ZN(n7406) );
  OAI21_X1 U9182 ( .B1(n7407), .B2(n8745), .A(n7406), .ZN(P1_U3231) );
  NAND2_X1 U9183 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  NAND2_X1 U9184 ( .A1(n7989), .A2(n7991), .ZN(n7921) );
  XNOR2_X1 U9185 ( .A(n7410), .B(n7921), .ZN(n7411) );
  OAI222_X1 U9186 ( .A1(n8351), .A2(n7412), .B1(n8349), .B2(n7728), .C1(n7411), 
        .C2(n8347), .ZN(n9930) );
  INV_X1 U9187 ( .A(n9930), .ZN(n7417) );
  NAND2_X1 U9188 ( .A1(n7383), .A2(n7980), .ZN(n7413) );
  XNOR2_X1 U9189 ( .A(n7413), .B(n7921), .ZN(n9932) );
  NOR2_X1 U9190 ( .A1(n8288), .A2(n9929), .ZN(n7415) );
  OAI22_X1 U9191 ( .A1(n8373), .A2(n10124), .B1(n7723), .B2(n8355), .ZN(n7414)
         );
  AOI211_X1 U9192 ( .C1(n9932), .C2(n9892), .A(n7415), .B(n7414), .ZN(n7416)
         );
  OAI21_X1 U9193 ( .B1(n7417), .B2(n8340), .A(n7416), .ZN(P2_U3223) );
  INV_X1 U9194 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7435) );
  AND2_X1 U9195 ( .A1(n7418), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7419) );
  OR2_X1 U9196 ( .A1(n7420), .A2(n7419), .ZN(n7422) );
  INV_X1 U9197 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7421) );
  XNOR2_X1 U9198 ( .A(n7422), .B(n7421), .ZN(n7427) );
  NAND2_X1 U9199 ( .A1(n7424), .A2(n7423), .ZN(n7426) );
  INV_X1 U9200 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7425) );
  XNOR2_X1 U9201 ( .A(n7426), .B(n7425), .ZN(n7428) );
  AOI22_X1 U9202 ( .A1(n7427), .A2(n9075), .B1(n9084), .B2(n7428), .ZN(n7433)
         );
  INV_X1 U9203 ( .A(n7427), .ZN(n7431) );
  OAI21_X1 U9204 ( .B1(n7429), .B2(n7428), .A(n9070), .ZN(n7430) );
  AOI21_X1 U9205 ( .B1(n7431), .B2(n9075), .A(n7430), .ZN(n7432) );
  MUX2_X1 U9206 ( .A(n7433), .B(n7432), .S(n9493), .Z(n7434) );
  NAND2_X1 U9207 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8580) );
  OAI211_X1 U9208 ( .C1(n7435), .C2(n9026), .A(n7434), .B(n8580), .ZN(P1_U3262) );
  INV_X1 U9209 ( .A(n7436), .ZN(n7438) );
  OAI222_X1 U9210 ( .A1(n8547), .A2(n7437), .B1(n8550), .B2(n7438), .C1(n8092), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9211 ( .A1(n7618), .A2(n7439), .B1(n9411), .B2(n7438), .C1(
        P1_U3086), .C2(n8912), .ZN(P1_U3333) );
  OAI21_X1 U9212 ( .B1(n5299), .B2(n7441), .A(n7440), .ZN(n7442) );
  NAND2_X1 U9213 ( .A1(n7442), .A2(n8722), .ZN(n7451) );
  OR2_X1 U9214 ( .A1(n8737), .A2(n7443), .ZN(n7446) );
  INV_X1 U9215 ( .A(n7444), .ZN(n7445) );
  OAI211_X1 U9216 ( .C1(n8704), .C2(n7447), .A(n7446), .B(n7445), .ZN(n7449)
         );
  NOR2_X1 U9217 ( .A1(n8739), .A2(n9619), .ZN(n7448) );
  NOR2_X1 U9218 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  OAI211_X1 U9219 ( .C1(n7453), .C2(n7452), .A(n7451), .B(n7450), .ZN(P1_U3221) );
  NOR2_X1 U9220 ( .A1(n7621), .A2(n8983), .ZN(n7454) );
  OR2_X1 U9221 ( .A1(n7517), .A2(n8738), .ZN(n8938) );
  NAND2_X1 U9222 ( .A1(n7517), .A2(n8738), .ZN(n8761) );
  NAND2_X1 U9223 ( .A1(n8938), .A2(n8761), .ZN(n8857) );
  INV_X1 U9224 ( .A(n8857), .ZN(n8772) );
  XNOR2_X1 U9225 ( .A(n7518), .B(n8772), .ZN(n9669) );
  AND3_X1 U9226 ( .A1(n7457), .A2(n8937), .A3(n8857), .ZN(n7458) );
  OAI21_X1 U9227 ( .B1(n7511), .B2(n7458), .A(n9486), .ZN(n7461) );
  OAI22_X1 U9228 ( .A1(n8633), .A2(n9656), .B1(n9514), .B2(n9277), .ZN(n7459)
         );
  INV_X1 U9229 ( .A(n7459), .ZN(n7460) );
  NAND2_X1 U9230 ( .A1(n7461), .A2(n7460), .ZN(n7462) );
  AOI21_X1 U9231 ( .B1(n9669), .B2(n9540), .A(n7462), .ZN(n9671) );
  OAI21_X1 U9232 ( .B1(n7463), .B2(n9666), .A(n9546), .ZN(n7464) );
  OR2_X1 U9233 ( .A1(n7464), .A2(n7513), .ZN(n9664) );
  AOI22_X1 U9234 ( .A1(n9301), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8560), .B2(
        n9541), .ZN(n7466) );
  NAND2_X1 U9235 ( .A1(n7517), .A2(n9291), .ZN(n7465) );
  OAI211_X1 U9236 ( .C1(n9664), .C2(n9295), .A(n7466), .B(n7465), .ZN(n7467)
         );
  AOI21_X1 U9237 ( .B1(n9669), .B2(n9550), .A(n7467), .ZN(n7468) );
  OAI21_X1 U9238 ( .B1(n9671), .B2(n9553), .A(n7468), .ZN(P1_U3279) );
  INV_X1 U9239 ( .A(n7470), .ZN(n7471) );
  NAND2_X1 U9240 ( .A1(n7469), .A2(n7471), .ZN(n7472) );
  NAND2_X1 U9241 ( .A1(n7473), .A2(n7472), .ZN(n7474) );
  XNOR2_X1 U9242 ( .A(n7664), .B(n9924), .ZN(n7635) );
  XNOR2_X1 U9243 ( .A(n7635), .B(n8107), .ZN(n7475) );
  AOI21_X1 U9244 ( .B1(n7474), .B2(n7475), .A(n7852), .ZN(n7477) );
  NAND2_X1 U9245 ( .A1(n7477), .A2(n7637), .ZN(n7483) );
  INV_X1 U9246 ( .A(n8106), .ZN(n7479) );
  NOR2_X1 U9247 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5779), .ZN(n9800) );
  AOI21_X1 U9248 ( .B1(n7858), .B2(n8108), .A(n9800), .ZN(n7478) );
  OAI21_X1 U9249 ( .B1(n7479), .B2(n7860), .A(n7478), .ZN(n7480) );
  AOI21_X1 U9250 ( .B1(n7481), .B2(n7850), .A(n7480), .ZN(n7482) );
  OAI211_X1 U9251 ( .C1(n7484), .C2(n7848), .A(n7483), .B(n7482), .ZN(P2_U3171) );
  AOI21_X1 U9252 ( .B1(n7487), .B2(n7486), .A(n7485), .ZN(n7503) );
  AOI21_X1 U9253 ( .B1(n4499), .B2(n7489), .A(n7488), .ZN(n7490) );
  NOR2_X1 U9254 ( .A1(n7490), .A2(n9872), .ZN(n7501) );
  INV_X1 U9255 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U9256 ( .A1(n9839), .A2(n10103), .ZN(n7500) );
  NOR2_X1 U9257 ( .A1(n9841), .A2(n7491), .ZN(n7499) );
  AOI21_X1 U9258 ( .B1(n7494), .B2(n7493), .A(n7492), .ZN(n7497) );
  INV_X1 U9259 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7495) );
  NOR2_X1 U9260 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7495), .ZN(n7725) );
  INV_X1 U9261 ( .A(n7725), .ZN(n7496) );
  OAI21_X1 U9262 ( .B1(n9847), .B2(n7497), .A(n7496), .ZN(n7498) );
  NOR4_X1 U9263 ( .A1(n7501), .A2(n7500), .A3(n7499), .A4(n7498), .ZN(n7502)
         );
  OAI21_X1 U9264 ( .B1(n7503), .B2(n9849), .A(n7502), .ZN(P2_U3192) );
  NAND2_X1 U9265 ( .A1(n7509), .A2(n7504), .ZN(n7506) );
  NOR2_X1 U9266 ( .A1(n7505), .A2(P2_U3151), .ZN(n8093) );
  INV_X1 U9267 ( .A(n8093), .ZN(n8098) );
  OAI211_X1 U9268 ( .C1(n7507), .C2(n8540), .A(n7506), .B(n8098), .ZN(P2_U3272) );
  NAND2_X1 U9269 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  OAI211_X1 U9270 ( .C1(n10037), .C2(n7618), .A(n7510), .B(n8970), .ZN(
        P1_U3332) );
  XNOR2_X1 U9271 ( .A(n7558), .B(n8981), .ZN(n8859) );
  INV_X1 U9272 ( .A(n8761), .ZN(n8775) );
  XOR2_X1 U9273 ( .A(n8859), .B(n4483), .Z(n7512) );
  AOI222_X1 U9274 ( .A1(n9486), .A2(n7512), .B1(n9298), .B2(n9535), .C1(n8982), 
        .C2(n9626), .ZN(n9521) );
  OAI211_X1 U9275 ( .C1(n7513), .C2(n9522), .A(n9546), .B(n7552), .ZN(n9520)
         );
  INV_X1 U9276 ( .A(n9520), .ZN(n7516) );
  AOI22_X1 U9277 ( .A1(n9301), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8743), .B2(
        n9541), .ZN(n7514) );
  OAI21_X1 U9278 ( .B1(n9522), .B2(n9544), .A(n7514), .ZN(n7515) );
  AOI21_X1 U9279 ( .B1(n7516), .B2(n9549), .A(n7515), .ZN(n7520) );
  XOR2_X1 U9280 ( .A(n8859), .B(n7557), .Z(n9524) );
  NAND2_X1 U9281 ( .A1(n9524), .A2(n9480), .ZN(n7519) );
  OAI211_X1 U9282 ( .C1(n9521), .C2(n9553), .A(n7520), .B(n7519), .ZN(P1_U3278) );
  AOI21_X1 U9283 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7537) );
  NOR2_X1 U9284 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7524), .ZN(n7756) );
  AOI21_X1 U9285 ( .B1(n7527), .B2(n7526), .A(n7525), .ZN(n7530) );
  AOI22_X1 U9286 ( .A1(n9858), .A2(n7528), .B1(n9856), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n7529) );
  OAI21_X1 U9287 ( .B1(n9872), .B2(n7530), .A(n7529), .ZN(n7531) );
  NOR2_X1 U9288 ( .A1(n7756), .A2(n7531), .ZN(n7536) );
  XNOR2_X1 U9289 ( .A(n7533), .B(n7532), .ZN(n7534) );
  NAND2_X1 U9290 ( .A1(n9868), .A2(n7534), .ZN(n7535) );
  OAI211_X1 U9291 ( .C1(n7537), .C2(n9849), .A(n7536), .B(n7535), .ZN(P2_U3194) );
  INV_X1 U9292 ( .A(n8698), .ZN(n7539) );
  AOI21_X1 U9293 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7550) );
  AOI21_X1 U9294 ( .B1(n8714), .B2(n8987), .A(n7542), .ZN(n7545) );
  NAND2_X1 U9295 ( .A1(n8742), .A2(n7543), .ZN(n7544) );
  OAI211_X1 U9296 ( .C1(n7546), .C2(n8704), .A(n7545), .B(n7544), .ZN(n7547)
         );
  AOI21_X1 U9297 ( .B1(n7548), .B2(n5770), .A(n7547), .ZN(n7549) );
  OAI21_X1 U9298 ( .B1(n7550), .B2(n8745), .A(n7549), .ZN(P1_U3217) );
  NAND2_X1 U9299 ( .A1(n9101), .A2(n8661), .ZN(n8942) );
  INV_X1 U9300 ( .A(n8861), .ZN(n8892) );
  XNOR2_X1 U9301 ( .A(n4484), .B(n8892), .ZN(n7551) );
  OAI22_X1 U9302 ( .A1(n7551), .A2(n9557), .B1(n9102), .B2(n9277), .ZN(n9517)
         );
  INV_X1 U9303 ( .A(n9517), .ZN(n7562) );
  AOI21_X1 U9304 ( .B1(n7552), .B2(n9101), .A(n9487), .ZN(n7553) );
  NAND2_X1 U9305 ( .A1(n9101), .A2(n9291), .ZN(n7555) );
  AOI22_X1 U9306 ( .A1(n9301), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8652), .B2(
        n9541), .ZN(n7554) );
  OAI211_X1 U9307 ( .C1(n9514), .C2(n9248), .A(n7555), .B(n7554), .ZN(n7556)
         );
  AOI21_X1 U9308 ( .B1(n9516), .B2(n9549), .A(n7556), .ZN(n7561) );
  AND2_X1 U9309 ( .A1(n7559), .A2(n8861), .ZN(n9512) );
  OR3_X1 U9310 ( .A1(n9513), .A2(n9512), .A3(n9286), .ZN(n7560) );
  OAI211_X1 U9311 ( .C1(n7562), .C2(n9553), .A(n7561), .B(n7560), .ZN(P1_U3277) );
  INV_X1 U9312 ( .A(n7563), .ZN(n7567) );
  OAI222_X1 U9313 ( .A1(n8550), .A2(n7567), .B1(P2_U3151), .B2(n7565), .C1(
        n7564), .C2(n8547), .ZN(P2_U3271) );
  OAI222_X1 U9314 ( .A1(n7568), .A2(P1_U3086), .B1(n9411), .B2(n7567), .C1(
        n7566), .C2(n7618), .ZN(P1_U3331) );
  INV_X1 U9315 ( .A(n7569), .ZN(n7573) );
  OAI222_X1 U9316 ( .A1(n8550), .A2(n7573), .B1(P2_U3151), .B2(n7571), .C1(
        n7570), .C2(n8547), .ZN(P2_U3270) );
  OAI222_X1 U9317 ( .A1(n7574), .A2(P1_U3086), .B1(n9411), .B2(n7573), .C1(
        n7572), .C2(n7618), .ZN(P1_U3330) );
  INV_X1 U9318 ( .A(n7575), .ZN(n7578) );
  OAI222_X1 U9319 ( .A1(n8546), .A2(n7578), .B1(P2_U3151), .B2(n4527), .C1(
        n7576), .C2(n8547), .ZN(P2_U3269) );
  OAI222_X1 U9320 ( .A1(n7579), .A2(P1_U3086), .B1(n9411), .B2(n7578), .C1(
        n7577), .C2(n7618), .ZN(P1_U3329) );
  NAND2_X1 U9321 ( .A1(n7580), .A2(n4905), .ZN(n7582) );
  OR2_X1 U9322 ( .A1(n8823), .A2(n10186), .ZN(n7581) );
  INV_X1 U9323 ( .A(n9335), .ZN(n7615) );
  INV_X1 U9324 ( .A(n7583), .ZN(n7585) );
  OR2_X1 U9325 ( .A1(n7585), .A2(n7584), .ZN(n7596) );
  NAND2_X1 U9326 ( .A1(n9335), .A2(n8593), .ZN(n7587) );
  OR2_X1 U9327 ( .A1(n9325), .A2(n5593), .ZN(n7586) );
  NAND2_X1 U9328 ( .A1(n7587), .A2(n7586), .ZN(n7588) );
  XNOR2_X1 U9329 ( .A(n7588), .B(n8591), .ZN(n7592) );
  INV_X1 U9330 ( .A(n7592), .ZN(n7594) );
  NOR2_X1 U9331 ( .A1(n9325), .A2(n8588), .ZN(n7590) );
  AOI21_X1 U9332 ( .B1(n9335), .B2(n5616), .A(n7590), .ZN(n7591) );
  INV_X1 U9333 ( .A(n7591), .ZN(n7593) );
  AOI21_X1 U9334 ( .B1(n7594), .B2(n7593), .A(n8607), .ZN(n7595) );
  AOI21_X1 U9335 ( .B1(n7600), .B2(n7596), .A(n7595), .ZN(n7601) );
  INV_X1 U9336 ( .A(n7595), .ZN(n7598) );
  INV_X1 U9337 ( .A(n7596), .ZN(n7597) );
  NOR2_X1 U9338 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  AND2_X2 U9339 ( .A1(n7600), .A2(n7599), .ZN(n8597) );
  OAI21_X1 U9340 ( .B1(n7601), .B2(n8597), .A(n8722), .ZN(n7614) );
  NAND2_X1 U9341 ( .A1(n8598), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9342 ( .A1(n5657), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7608) );
  NAND2_X1 U9343 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7602) );
  INV_X1 U9344 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7610) );
  INV_X1 U9345 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7603) );
  OAI21_X1 U9346 ( .B1(n7604), .B2(n7610), .A(n7603), .ZN(n7605) );
  NAND2_X1 U9347 ( .A1(n5210), .A2(n9144), .ZN(n7607) );
  NAND2_X1 U9348 ( .A1(n5461), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7606) );
  NOR2_X1 U9349 ( .A1(n8704), .A2(n9116), .ZN(n7612) );
  OAI22_X1 U9350 ( .A1(n8737), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7610), .ZN(n7611) );
  AOI211_X1 U9351 ( .C1(n9156), .C2(n8742), .A(n7612), .B(n7611), .ZN(n7613)
         );
  OAI211_X1 U9352 ( .C1(n7615), .C2(n8739), .A(n7614), .B(n7613), .ZN(P1_U3214) );
  INV_X1 U9353 ( .A(n7616), .ZN(n7682) );
  OAI222_X1 U9354 ( .A1(n7618), .A2(n7617), .B1(n9411), .B2(n7682), .C1(
        P1_U3086), .C2(n8972), .ZN(P1_U3336) );
  INV_X1 U9355 ( .A(n7619), .ZN(n7686) );
  OAI222_X1 U9356 ( .A1(n7618), .A2(n8806), .B1(P1_U3086), .B2(n7620), .C1(
        n7686), .C2(n9411), .ZN(P1_U3326) );
  INV_X1 U9357 ( .A(n7621), .ZN(n9658) );
  NAND2_X1 U9358 ( .A1(n8624), .A2(n7622), .ZN(n8629) );
  NAND2_X1 U9359 ( .A1(n8629), .A2(n7623), .ZN(n7626) );
  OAI21_X1 U9360 ( .B1(n7627), .B2(n7626), .A(n7625), .ZN(n7628) );
  NAND2_X1 U9361 ( .A1(n7628), .A2(n8722), .ZN(n7634) );
  AOI21_X1 U9362 ( .B1(n8714), .B2(n8984), .A(n7629), .ZN(n7630) );
  OAI21_X1 U9363 ( .B1(n8738), .B2(n8704), .A(n7630), .ZN(n7631) );
  AOI21_X1 U9364 ( .B1(n7632), .B2(n8742), .A(n7631), .ZN(n7633) );
  OAI211_X1 U9365 ( .C1(n9658), .C2(n8739), .A(n7634), .B(n7633), .ZN(P1_U3234) );
  XNOR2_X1 U9366 ( .A(n7822), .B(n7664), .ZN(n7659) );
  XNOR2_X1 U9367 ( .A(n8279), .B(n7664), .ZN(n7655) );
  XNOR2_X1 U9368 ( .A(n8502), .B(n7664), .ZN(n7652) );
  INV_X1 U9369 ( .A(n7652), .ZN(n7653) );
  XNOR2_X1 U9370 ( .A(n8421), .B(n7664), .ZN(n7649) );
  XNOR2_X1 U9371 ( .A(n9929), .B(n7664), .ZN(n7722) );
  XNOR2_X1 U9372 ( .A(n7923), .B(n7664), .ZN(n7832) );
  NAND2_X1 U9373 ( .A1(n7635), .A2(n8107), .ZN(n7636) );
  NOR3_X1 U9374 ( .A1(n8106), .A2(n7664), .A3(n7730), .ZN(n7639) );
  AOI211_X1 U9375 ( .C1(n7728), .C2(n7664), .A(n7639), .B(n7638), .ZN(n7642)
         );
  NOR3_X1 U9376 ( .A1(n7667), .A2(n9929), .A3(n8106), .ZN(n7640) );
  AOI211_X1 U9377 ( .C1(n7728), .C2(n7667), .A(n7923), .B(n7640), .ZN(n7641)
         );
  XNOR2_X1 U9378 ( .A(n8533), .B(n7664), .ZN(n7643) );
  NAND2_X1 U9379 ( .A1(n7643), .A2(n8350), .ZN(n7751) );
  OAI21_X1 U9380 ( .B1(n7642), .B2(n7641), .A(n7751), .ZN(n7645) );
  INV_X1 U9381 ( .A(n7643), .ZN(n7644) );
  NAND2_X1 U9382 ( .A1(n7644), .A2(n8105), .ZN(n7752) );
  XNOR2_X1 U9383 ( .A(n8526), .B(n7664), .ZN(n7646) );
  XNOR2_X1 U9384 ( .A(n7646), .B(n8332), .ZN(n7813) );
  INV_X1 U9385 ( .A(n7646), .ZN(n7647) );
  INV_X1 U9386 ( .A(n8332), .ZN(n8371) );
  XNOR2_X1 U9387 ( .A(n8520), .B(n7664), .ZN(n7648) );
  XNOR2_X1 U9388 ( .A(n7648), .B(n8104), .ZN(n7709) );
  XNOR2_X1 U9389 ( .A(n7649), .B(n8330), .ZN(n7868) );
  XNOR2_X1 U9390 ( .A(n8508), .B(n7664), .ZN(n7650) );
  XNOR2_X1 U9391 ( .A(n7650), .B(n8321), .ZN(n7778) );
  INV_X1 U9392 ( .A(n7650), .ZN(n7651) );
  NOR2_X1 U9393 ( .A1(n7651), .A2(n8103), .ZN(n7786) );
  XNOR2_X1 U9394 ( .A(n7652), .B(n8102), .ZN(n7785) );
  XNOR2_X1 U9395 ( .A(n8287), .B(n7664), .ZN(n7654) );
  XNOR2_X1 U9396 ( .A(n7654), .B(n8298), .ZN(n7844) );
  XNOR2_X1 U9397 ( .A(n7655), .B(n8262), .ZN(n7734) );
  XNOR2_X1 U9398 ( .A(n8487), .B(n7664), .ZN(n7656) );
  NOR2_X1 U9399 ( .A1(n7656), .A2(n8252), .ZN(n7804) );
  XNOR2_X1 U9400 ( .A(n8403), .B(n7667), .ZN(n7657) );
  NOR2_X1 U9401 ( .A1(n7657), .A2(n8263), .ZN(n7658) );
  AOI21_X1 U9402 ( .B1(n7657), .B2(n8263), .A(n7658), .ZN(n7743) );
  INV_X1 U9403 ( .A(n7658), .ZN(n7823) );
  XNOR2_X1 U9404 ( .A(n7659), .B(n8251), .ZN(n7824) );
  XNOR2_X1 U9405 ( .A(n8474), .B(n7664), .ZN(n7765) );
  XNOR2_X1 U9406 ( .A(n8468), .B(n7667), .ZN(n7660) );
  NAND2_X1 U9407 ( .A1(n7660), .A2(n8226), .ZN(n7769) );
  OAI21_X1 U9408 ( .B1(n8236), .B2(n7765), .A(n7769), .ZN(n7663) );
  NAND3_X1 U9409 ( .A1(n7769), .A2(n8236), .A3(n7765), .ZN(n7662) );
  INV_X1 U9410 ( .A(n7660), .ZN(n7661) );
  NAND2_X1 U9411 ( .A1(n7661), .A2(n7764), .ZN(n7771) );
  XNOR2_X1 U9412 ( .A(n8462), .B(n7664), .ZN(n7665) );
  XNOR2_X1 U9413 ( .A(n7665), .B(n8214), .ZN(n7770) );
  NAND2_X1 U9414 ( .A1(n7665), .A2(n8187), .ZN(n7666) );
  XNOR2_X1 U9415 ( .A(n8456), .B(n7667), .ZN(n7669) );
  INV_X1 U9416 ( .A(n7669), .ZN(n7670) );
  NAND2_X1 U9417 ( .A1(n7668), .A2(n7670), .ZN(n7671) );
  XNOR2_X1 U9418 ( .A(n8450), .B(n7664), .ZN(n7672) );
  XNOR2_X1 U9419 ( .A(n7672), .B(n7861), .ZN(n7699) );
  INV_X1 U9420 ( .A(n7672), .ZN(n7673) );
  NAND2_X1 U9421 ( .A1(n7673), .A2(n8185), .ZN(n7674) );
  NAND2_X1 U9422 ( .A1(n7700), .A2(n7674), .ZN(n7676) );
  XNOR2_X1 U9423 ( .A(n7676), .B(n7675), .ZN(n7681) );
  AOI22_X1 U9424 ( .A1(n8185), .A2(n7858), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7678) );
  NAND2_X1 U9425 ( .A1(n8169), .A2(n7875), .ZN(n7677) );
  OAI211_X1 U9426 ( .C1(n8101), .C2(n7860), .A(n7678), .B(n7677), .ZN(n7679)
         );
  AOI21_X1 U9427 ( .B1(n8444), .B2(n7850), .A(n7679), .ZN(n7680) );
  OAI21_X1 U9428 ( .B1(n7681), .B2(n7852), .A(n7680), .ZN(P2_U3160) );
  OAI222_X1 U9429 ( .A1(n8540), .A2(n7683), .B1(n8550), .B2(n7682), .C1(n6237), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U9430 ( .A(n7580), .ZN(n8549) );
  OAI222_X1 U9431 ( .A1(n7618), .A2(n10186), .B1(n9411), .B2(n8549), .C1(n8992), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U9432 ( .A1(n8550), .A2(n7686), .B1(n7685), .B2(P2_U3151), .C1(
        n7684), .C2(n8547), .ZN(P2_U3266) );
  INV_X1 U9433 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7879) );
  INV_X1 U9434 ( .A(SI_29_), .ZN(n7687) );
  INV_X1 U9435 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8822) );
  MUX2_X1 U9436 ( .A(n8822), .B(n7879), .S(n7885), .Z(n7694) );
  INV_X1 U9437 ( .A(SI_30_), .ZN(n7693) );
  NAND2_X1 U9438 ( .A1(n7694), .A2(n7693), .ZN(n7882) );
  INV_X1 U9439 ( .A(n7694), .ZN(n7695) );
  NAND2_X1 U9440 ( .A1(n7695), .A2(SI_30_), .ZN(n7696) );
  NAND2_X1 U9441 ( .A1(n7882), .A2(n7696), .ZN(n7883) );
  INV_X1 U9442 ( .A(n8821), .ZN(n7698) );
  OAI222_X1 U9443 ( .A1(n8540), .A2(n7879), .B1(n8546), .B2(n7698), .C1(
        P2_U3151), .C2(n5815), .ZN(P2_U3265) );
  INV_X1 U9444 ( .A(n8585), .ZN(n8545) );
  OAI222_X1 U9445 ( .A1(n7618), .A2(n10051), .B1(n9411), .B2(n8545), .C1(n5160), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U9446 ( .A1(n7618), .A2(n8822), .B1(n9411), .B2(n7698), .C1(n7697), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  NAND2_X1 U9447 ( .A1(n7701), .A2(n7700), .ZN(n7706) );
  AOI22_X1 U9448 ( .A1(n8197), .A2(n7858), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7702) );
  OAI21_X1 U9449 ( .B1(n7703), .B2(n7860), .A(n7702), .ZN(n7704) );
  AOI21_X1 U9450 ( .B1(n8177), .B2(n7875), .A(n7704), .ZN(n7705) );
  OAI211_X1 U9451 ( .C1(n7707), .C2(n7878), .A(n7706), .B(n7705), .ZN(P2_U3154) );
  XOR2_X1 U9452 ( .A(n7709), .B(n4411), .Z(n7715) );
  INV_X1 U9453 ( .A(n8335), .ZN(n7713) );
  NAND2_X1 U9454 ( .A1(n7858), .A2(n8371), .ZN(n7710) );
  NAND2_X1 U9455 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8120) );
  OAI211_X1 U9456 ( .C1(n7926), .C2(n7860), .A(n7710), .B(n8120), .ZN(n7712)
         );
  INV_X1 U9457 ( .A(n8520), .ZN(n8337) );
  NOR2_X1 U9458 ( .A1(n8337), .A2(n7878), .ZN(n7711) );
  AOI211_X1 U9459 ( .C1(n7713), .C2(n7875), .A(n7712), .B(n7711), .ZN(n7714)
         );
  OAI21_X1 U9460 ( .B1(n7715), .B2(n7852), .A(n7714), .ZN(P2_U3155) );
  XNOR2_X1 U9461 ( .A(n7767), .B(n7765), .ZN(n7768) );
  XNOR2_X1 U9462 ( .A(n7768), .B(n8215), .ZN(n7720) );
  AOI22_X1 U9463 ( .A1(n8226), .A2(n7871), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7717) );
  NAND2_X1 U9464 ( .A1(n7875), .A2(n8230), .ZN(n7716) );
  OAI211_X1 U9465 ( .C1(n8251), .C2(n7873), .A(n7717), .B(n7716), .ZN(n7718)
         );
  AOI21_X1 U9466 ( .B1(n8474), .B2(n7850), .A(n7718), .ZN(n7719) );
  OAI21_X1 U9467 ( .B1(n7720), .B2(n7852), .A(n7719), .ZN(P2_U3156) );
  XNOR2_X1 U9468 ( .A(n7750), .B(n8106), .ZN(n7721) );
  NOR2_X1 U9469 ( .A1(n7721), .A2(n7722), .ZN(n7834) );
  AOI21_X1 U9470 ( .B1(n7722), .B2(n7721), .A(n7834), .ZN(n7732) );
  INV_X1 U9471 ( .A(n7723), .ZN(n7724) );
  NAND2_X1 U9472 ( .A1(n7875), .A2(n7724), .ZN(n7727) );
  AOI21_X1 U9473 ( .B1(n7858), .B2(n8107), .A(n7725), .ZN(n7726) );
  OAI211_X1 U9474 ( .C1(n7728), .C2(n7860), .A(n7727), .B(n7726), .ZN(n7729)
         );
  AOI21_X1 U9475 ( .B1(n7730), .B2(n7850), .A(n7729), .ZN(n7731) );
  OAI21_X1 U9476 ( .B1(n7732), .B2(n7852), .A(n7731), .ZN(P2_U3157) );
  INV_X1 U9477 ( .A(n8279), .ZN(n8492) );
  OAI211_X1 U9478 ( .C1(n7735), .C2(n7734), .A(n7733), .B(n7866), .ZN(n7740)
         );
  NAND2_X1 U9479 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9466) );
  OAI21_X1 U9480 ( .B1(n7873), .B2(n7736), .A(n9466), .ZN(n7738) );
  NOR2_X1 U9481 ( .A1(n7848), .A2(n8277), .ZN(n7737) );
  AOI211_X1 U9482 ( .C1(n7871), .C2(n8274), .A(n7738), .B(n7737), .ZN(n7739)
         );
  OAI211_X1 U9483 ( .C1(n8492), .C2(n7878), .A(n7740), .B(n7739), .ZN(P2_U3159) );
  INV_X1 U9484 ( .A(n8403), .ZN(n7749) );
  OAI21_X1 U9485 ( .B1(n7743), .B2(n7741), .A(n4407), .ZN(n7744) );
  NAND2_X1 U9486 ( .A1(n7744), .A2(n7866), .ZN(n7748) );
  AOI22_X1 U9487 ( .A1(n7871), .A2(n8227), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7745) );
  OAI21_X1 U9488 ( .B1(n8252), .B2(n7873), .A(n7745), .ZN(n7746) );
  AOI21_X1 U9489 ( .B1(n8253), .B2(n7875), .A(n7746), .ZN(n7747) );
  OAI211_X1 U9490 ( .C1(n7749), .C2(n7878), .A(n7748), .B(n7747), .ZN(P2_U3163) );
  NOR2_X1 U9491 ( .A1(n7750), .A2(n8106), .ZN(n7833) );
  NOR3_X1 U9492 ( .A1(n7834), .A2(n7833), .A3(n7832), .ZN(n7831) );
  AOI21_X1 U9493 ( .B1(n8369), .B2(n7832), .A(n7831), .ZN(n7754) );
  NAND2_X1 U9494 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  XNOR2_X1 U9495 ( .A(n7754), .B(n7753), .ZN(n7761) );
  INV_X1 U9496 ( .A(n7755), .ZN(n8375) );
  NAND2_X1 U9497 ( .A1(n7875), .A2(n8375), .ZN(n7758) );
  AOI21_X1 U9498 ( .B1(n7858), .B2(n8369), .A(n7756), .ZN(n7757) );
  OAI211_X1 U9499 ( .C1(n8332), .C2(n7860), .A(n7758), .B(n7757), .ZN(n7759)
         );
  AOI21_X1 U9500 ( .B1(n8533), .B2(n7850), .A(n7759), .ZN(n7760) );
  OAI21_X1 U9501 ( .B1(n7761), .B2(n7852), .A(n7760), .ZN(P2_U3164) );
  AOI22_X1 U9502 ( .A1(n8197), .A2(n7871), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7763) );
  NAND2_X1 U9503 ( .A1(n7875), .A2(n8199), .ZN(n7762) );
  OAI211_X1 U9504 ( .C1(n7764), .C2(n7873), .A(n7763), .B(n7762), .ZN(n7776)
         );
  INV_X1 U9505 ( .A(n7765), .ZN(n7766) );
  AOI22_X1 U9506 ( .A1(n7768), .A2(n8215), .B1(n7767), .B2(n7766), .ZN(n7797)
         );
  AND2_X1 U9507 ( .A1(n7769), .A2(n7771), .ZN(n7798) );
  NAND2_X1 U9508 ( .A1(n7797), .A2(n7798), .ZN(n7796) );
  INV_X1 U9509 ( .A(n7770), .ZN(n7772) );
  NAND3_X1 U9510 ( .A1(n7796), .A2(n7772), .A3(n7771), .ZN(n7774) );
  AOI21_X1 U9511 ( .B1(n7774), .B2(n7773), .A(n7852), .ZN(n7775) );
  AOI21_X1 U9512 ( .B1(n7778), .B2(n7777), .A(n7787), .ZN(n7783) );
  NAND2_X1 U9513 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8136) );
  OAI21_X1 U9514 ( .B1(n7860), .B2(n8310), .A(n8136), .ZN(n7779) );
  AOI21_X1 U9515 ( .B1(n7858), .B2(n8330), .A(n7779), .ZN(n7780) );
  OAI21_X1 U9516 ( .B1(n7848), .B2(n8313), .A(n7780), .ZN(n7781) );
  AOI21_X1 U9517 ( .B1(n8508), .B2(n7850), .A(n7781), .ZN(n7782) );
  OAI21_X1 U9518 ( .B1(n7783), .B2(n7852), .A(n7782), .ZN(P2_U3166) );
  INV_X1 U9519 ( .A(n8502), .ZN(n7795) );
  INV_X1 U9520 ( .A(n4410), .ZN(n7789) );
  NOR3_X1 U9521 ( .A1(n7787), .A2(n7786), .A3(n7785), .ZN(n7788) );
  OAI21_X1 U9522 ( .B1(n7789), .B2(n7788), .A(n7866), .ZN(n7794) );
  INV_X1 U9523 ( .A(n7790), .ZN(n8302) );
  AOI22_X1 U9524 ( .A1(n7871), .A2(n8298), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n7791) );
  OAI21_X1 U9525 ( .B1(n8321), .B2(n7873), .A(n7791), .ZN(n7792) );
  AOI21_X1 U9526 ( .B1(n8302), .B2(n7875), .A(n7792), .ZN(n7793) );
  OAI211_X1 U9527 ( .C1(n7795), .C2(n7878), .A(n7794), .B(n7793), .ZN(P2_U3168) );
  INV_X1 U9528 ( .A(n8468), .ZN(n8219) );
  OAI21_X1 U9529 ( .B1(n7798), .B2(n7797), .A(n7796), .ZN(n7799) );
  NAND2_X1 U9530 ( .A1(n7799), .A2(n7866), .ZN(n7803) );
  AOI22_X1 U9531 ( .A1(n8214), .A2(n7871), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7800) );
  OAI21_X1 U9532 ( .B1(n8236), .B2(n7873), .A(n7800), .ZN(n7801) );
  AOI21_X1 U9533 ( .B1(n8217), .B2(n7875), .A(n7801), .ZN(n7802) );
  OAI211_X1 U9534 ( .C1(n8219), .C2(n7878), .A(n7803), .B(n7802), .ZN(P2_U3169) );
  NOR2_X1 U9535 ( .A1(n7804), .A2(n4485), .ZN(n7805) );
  XNOR2_X1 U9536 ( .A(n7806), .B(n7805), .ZN(n7812) );
  INV_X1 U9537 ( .A(n7807), .ZN(n8266) );
  NAND2_X1 U9538 ( .A1(n7875), .A2(n8266), .ZN(n7809) );
  AOI22_X1 U9539 ( .A1(n7858), .A2(n8262), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7808) );
  OAI211_X1 U9540 ( .C1(n8237), .C2(n7860), .A(n7809), .B(n7808), .ZN(n7810)
         );
  AOI21_X1 U9541 ( .B1(n8487), .B2(n7850), .A(n7810), .ZN(n7811) );
  OAI21_X1 U9542 ( .B1(n7812), .B2(n7852), .A(n7811), .ZN(P2_U3173) );
  XOR2_X1 U9543 ( .A(n7814), .B(n7813), .Z(n7821) );
  INV_X1 U9544 ( .A(n8356), .ZN(n7819) );
  NAND2_X1 U9545 ( .A1(n7858), .A2(n8105), .ZN(n7815) );
  NAND2_X1 U9546 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9823) );
  OAI211_X1 U9547 ( .C1(n8348), .C2(n7860), .A(n7815), .B(n9823), .ZN(n7818)
         );
  NOR2_X1 U9548 ( .A1(n7816), .A2(n7878), .ZN(n7817) );
  AOI211_X1 U9549 ( .C1(n7819), .C2(n7875), .A(n7818), .B(n7817), .ZN(n7820)
         );
  OAI21_X1 U9550 ( .B1(n7821), .B2(n7852), .A(n7820), .ZN(P2_U3174) );
  AND3_X1 U9551 ( .A1(n4407), .A2(n7824), .A3(n7823), .ZN(n7825) );
  OAI21_X1 U9552 ( .B1(n7826), .B2(n7825), .A(n7866), .ZN(n7830) );
  AOI22_X1 U9553 ( .A1(n7858), .A2(n8263), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7827) );
  OAI21_X1 U9554 ( .B1(n8236), .B2(n7860), .A(n7827), .ZN(n7828) );
  AOI21_X1 U9555 ( .B1(n8240), .B2(n7875), .A(n7828), .ZN(n7829) );
  OAI211_X1 U9556 ( .C1(n8481), .C2(n7878), .A(n7830), .B(n7829), .ZN(P2_U3175) );
  INV_X1 U9557 ( .A(n7831), .ZN(n7836) );
  OAI21_X1 U9558 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n7835) );
  NAND3_X1 U9559 ( .A1(n7836), .A2(n7866), .A3(n7835), .ZN(n7842) );
  NAND2_X1 U9560 ( .A1(n7858), .A2(n8106), .ZN(n7838) );
  AND2_X1 U9561 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9816) );
  INV_X1 U9562 ( .A(n9816), .ZN(n7837) );
  OAI211_X1 U9563 ( .C1(n8350), .C2(n7860), .A(n7838), .B(n7837), .ZN(n7839)
         );
  AOI21_X1 U9564 ( .B1(n7875), .B2(n7840), .A(n7839), .ZN(n7841) );
  OAI211_X1 U9565 ( .C1(n9934), .C2(n7878), .A(n7842), .B(n7841), .ZN(P2_U3176) );
  XOR2_X1 U9566 ( .A(n7844), .B(n7843), .Z(n7853) );
  OAI22_X1 U9567 ( .A1(n7860), .A2(n8284), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7845), .ZN(n7846) );
  AOI21_X1 U9568 ( .B1(n7858), .B2(n8102), .A(n7846), .ZN(n7847) );
  OAI21_X1 U9569 ( .B1(n7848), .B2(n8289), .A(n7847), .ZN(n7849) );
  AOI21_X1 U9570 ( .B1(n8287), .B2(n7850), .A(n7849), .ZN(n7851) );
  OAI21_X1 U9571 ( .B1(n7853), .B2(n7852), .A(n7851), .ZN(P2_U3178) );
  OAI21_X1 U9572 ( .B1(n7856), .B2(n7855), .A(n7854), .ZN(n7857) );
  NAND2_X1 U9573 ( .A1(n7857), .A2(n7866), .ZN(n7864) );
  AOI22_X1 U9574 ( .A1(n8214), .A2(n7858), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7859) );
  OAI21_X1 U9575 ( .B1(n7861), .B2(n7860), .A(n7859), .ZN(n7862) );
  AOI21_X1 U9576 ( .B1(n8182), .B2(n7875), .A(n7862), .ZN(n7863) );
  OAI211_X1 U9577 ( .C1(n7865), .C2(n7878), .A(n7864), .B(n7863), .ZN(P2_U3180) );
  OAI211_X1 U9578 ( .C1(n7869), .C2(n7868), .A(n7867), .B(n7866), .ZN(n7877)
         );
  INV_X1 U9579 ( .A(n7870), .ZN(n8323) );
  NOR2_X1 U9580 ( .A1(n10237), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9853) );
  AOI21_X1 U9581 ( .B1(n7871), .B2(n8103), .A(n9853), .ZN(n7872) );
  OAI21_X1 U9582 ( .B1(n8348), .B2(n7873), .A(n7872), .ZN(n7874) );
  AOI21_X1 U9583 ( .B1(n8323), .B2(n7875), .A(n7874), .ZN(n7876) );
  OAI211_X1 U9584 ( .C1(n8514), .C2(n7878), .A(n7877), .B(n7876), .ZN(P2_U3181) );
  NAND2_X1 U9585 ( .A1(n8821), .A2(n7890), .ZN(n7881) );
  OR2_X1 U9586 ( .A1(n5864), .A2(n7879), .ZN(n7880) );
  INV_X1 U9587 ( .A(n8439), .ZN(n8154) );
  OAI21_X1 U9588 ( .B1(n7884), .B2(n7883), .A(n7882), .ZN(n7888) );
  INV_X1 U9589 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8814) );
  MUX2_X1 U9590 ( .A(n8814), .B(n10158), .S(n7885), .Z(n7886) );
  XNOR2_X1 U9591 ( .A(n7886), .B(SI_31_), .ZN(n7887) );
  XNOR2_X1 U9592 ( .A(n7888), .B(n7887), .ZN(n8813) );
  AOI22_X1 U9593 ( .A1(n8813), .A2(n7890), .B1(n7889), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8438) );
  INV_X1 U9594 ( .A(n8438), .ZN(n8379) );
  NAND2_X1 U9595 ( .A1(n8439), .A2(n7900), .ZN(n8076) );
  NAND2_X1 U9596 ( .A1(n8076), .A2(n7892), .ZN(n8081) );
  INV_X1 U9597 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7897) );
  AOI22_X1 U9598 ( .A1(n7894), .A2(P2_REG2_REG_31__SCAN_IN), .B1(n5889), .B2(
        P2_REG0_REG_31__SCAN_IN), .ZN(n7895) );
  OAI211_X1 U9599 ( .C1(n5870), .C2(n7897), .A(n7896), .B(n7895), .ZN(n8100)
         );
  INV_X1 U9600 ( .A(n8100), .ZN(n8149) );
  NOR2_X1 U9601 ( .A1(n8379), .A2(n8149), .ZN(n8087) );
  INV_X1 U9602 ( .A(n8087), .ZN(n7898) );
  OAI211_X1 U9603 ( .C1(n8154), .C2(n8379), .A(n7899), .B(n7898), .ZN(n7938)
         );
  OR2_X1 U9604 ( .A1(n8439), .A2(n7900), .ZN(n8077) );
  INV_X1 U9605 ( .A(n8077), .ZN(n7901) );
  NOR2_X1 U9606 ( .A1(n8438), .A2(n8100), .ZN(n8085) );
  AOI211_X1 U9607 ( .C1(n7901), .C2(n8379), .A(n7913), .B(n8085), .ZN(n7937)
         );
  INV_X1 U9608 ( .A(n8062), .ZN(n7902) );
  INV_X1 U9609 ( .A(n7903), .ZN(n8066) );
  INV_X1 U9610 ( .A(n8210), .ZN(n8213) );
  INV_X1 U9611 ( .A(n8285), .ZN(n7930) );
  INV_X1 U9612 ( .A(n7906), .ZN(n7910) );
  INV_X1 U9613 ( .A(n7945), .ZN(n7908) );
  NOR4_X1 U9614 ( .A1(n7910), .A2(n7909), .A3(n7908), .A4(n7907), .ZN(n7919)
         );
  NAND2_X1 U9615 ( .A1(n7912), .A2(n7911), .ZN(n7946) );
  AND2_X1 U9616 ( .A1(n7914), .A2(n7913), .ZN(n7947) );
  INV_X1 U9617 ( .A(n7947), .ZN(n7915) );
  NOR4_X1 U9618 ( .A1(n9878), .A2(n7946), .A3(n7916), .A4(n7915), .ZN(n7917)
         );
  NAND4_X1 U9619 ( .A1(n7919), .A2(n7918), .A3(n7917), .A4(n9887), .ZN(n7924)
         );
  INV_X1 U9620 ( .A(n7920), .ZN(n7922) );
  NOR4_X1 U9621 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n7925)
         );
  INV_X1 U9622 ( .A(n8362), .ZN(n8367) );
  NAND3_X1 U9623 ( .A1(n7925), .A2(n8367), .A3(n8353), .ZN(n7928) );
  XNOR2_X1 U9624 ( .A(n8421), .B(n7926), .ZN(n8318) );
  INV_X1 U9625 ( .A(n7927), .ZN(n8007) );
  NOR4_X1 U9626 ( .A1(n8307), .A2(n7928), .A3(n8318), .A4(n8329), .ZN(n7929)
         );
  NAND4_X1 U9627 ( .A1(n8270), .A2(n8297), .A3(n7930), .A4(n7929), .ZN(n7931)
         );
  NOR4_X1 U9628 ( .A1(n8238), .A2(n8249), .A3(n8261), .A4(n7931), .ZN(n7932)
         );
  NAND4_X1 U9629 ( .A1(n8196), .A2(n8213), .A3(n8225), .A4(n7932), .ZN(n7933)
         );
  NOR3_X1 U9630 ( .A1(n8180), .A2(n8173), .A3(n7933), .ZN(n7934) );
  NAND4_X1 U9631 ( .A1(n8077), .A2(n7934), .A3(n8165), .A4(n7891), .ZN(n7935)
         );
  NOR4_X1 U9632 ( .A1(n8085), .A2(n8087), .A3(n8081), .A4(n7935), .ZN(n7936)
         );
  NAND2_X1 U9633 ( .A1(n7946), .A2(n7945), .ZN(n7941) );
  NAND2_X1 U9634 ( .A1(n8112), .A2(n7939), .ZN(n7962) );
  OAI211_X1 U9635 ( .C1(n7941), .C2(n9878), .A(n7940), .B(n7962), .ZN(n7944)
         );
  NAND2_X1 U9636 ( .A1(n7942), .A2(n7953), .ZN(n7943) );
  MUX2_X1 U9637 ( .A(n7944), .B(n7943), .S(n8078), .Z(n7952) );
  OAI21_X1 U9638 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n7949) );
  NOR2_X1 U9639 ( .A1(n9878), .A2(n8083), .ZN(n7948) );
  AND2_X1 U9640 ( .A1(n7949), .A2(n7948), .ZN(n7951) );
  OAI21_X1 U9641 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n7966) );
  INV_X1 U9642 ( .A(n7953), .ZN(n7958) );
  INV_X1 U9643 ( .A(n7954), .ZN(n7956) );
  NOR2_X1 U9644 ( .A1(n7956), .A2(n7955), .ZN(n7967) );
  OAI211_X1 U9645 ( .C1(n7966), .C2(n7958), .A(n7967), .B(n7957), .ZN(n7961)
         );
  AOI21_X1 U9646 ( .B1(n7963), .B2(n6220), .A(n6219), .ZN(n7960) );
  NAND2_X1 U9647 ( .A1(n7961), .A2(n7960), .ZN(n7970) );
  INV_X1 U9648 ( .A(n7962), .ZN(n7965) );
  OAI211_X1 U9649 ( .C1(n7966), .C2(n7965), .A(n6217), .B(n7964), .ZN(n7968)
         );
  AOI21_X1 U9650 ( .B1(n7968), .B2(n7967), .A(n6219), .ZN(n7969) );
  NAND2_X1 U9651 ( .A1(n7978), .A2(n7971), .ZN(n7974) );
  INV_X1 U9652 ( .A(n7972), .ZN(n7973) );
  MUX2_X1 U9653 ( .A(n7974), .B(n7973), .S(n8078), .Z(n7975) );
  AOI21_X1 U9654 ( .B1(n7977), .B2(n7976), .A(n7975), .ZN(n7984) );
  NAND2_X1 U9655 ( .A1(n7978), .A2(n7985), .ZN(n7982) );
  NAND2_X1 U9656 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  MUX2_X1 U9657 ( .A(n7982), .B(n7981), .S(n8083), .Z(n7983) );
  AND2_X1 U9658 ( .A1(n7989), .A2(n7985), .ZN(n7987) );
  MUX2_X1 U9659 ( .A(n7987), .B(n7986), .S(n8078), .Z(n7988) );
  NAND3_X1 U9660 ( .A1(n7993), .A2(n7994), .A3(n7989), .ZN(n7990) );
  NAND2_X1 U9661 ( .A1(n7990), .A2(n7992), .ZN(n7997) );
  NAND3_X1 U9662 ( .A1(n7993), .A2(n7992), .A3(n7991), .ZN(n7995) );
  NAND2_X1 U9663 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  MUX2_X1 U9664 ( .A(n7997), .B(n7996), .S(n8083), .Z(n8001) );
  MUX2_X1 U9665 ( .A(n7999), .B(n7998), .S(n8078), .Z(n8000) );
  OAI211_X1 U9666 ( .C1(n8001), .C2(n8362), .A(n8353), .B(n8000), .ZN(n8005)
         );
  INV_X1 U9667 ( .A(n8329), .ZN(n8326) );
  MUX2_X1 U9668 ( .A(n8003), .B(n8002), .S(n8083), .Z(n8004) );
  NAND3_X1 U9669 ( .A1(n8005), .A2(n8326), .A3(n8004), .ZN(n8010) );
  MUX2_X1 U9670 ( .A(n8007), .B(n8006), .S(n8083), .Z(n8008) );
  NOR2_X1 U9671 ( .A1(n8318), .A2(n8008), .ZN(n8009) );
  NAND2_X1 U9672 ( .A1(n8010), .A2(n8009), .ZN(n8016) );
  AND2_X1 U9673 ( .A1(n8018), .A2(n8011), .ZN(n8012) );
  MUX2_X1 U9674 ( .A(n8013), .B(n8012), .S(n8078), .Z(n8014) );
  NAND3_X1 U9675 ( .A1(n8016), .A2(n8015), .A3(n8014), .ZN(n8017) );
  NAND2_X1 U9676 ( .A1(n8017), .A2(n8297), .ZN(n8022) );
  INV_X1 U9677 ( .A(n8018), .ZN(n8019) );
  NOR2_X1 U9678 ( .A1(n8022), .A2(n8019), .ZN(n8023) );
  NAND3_X1 U9679 ( .A1(n8030), .A2(n8031), .A3(n8026), .ZN(n8024) );
  NAND3_X1 U9680 ( .A1(n8024), .A2(n8035), .A3(n8028), .ZN(n8034) );
  NAND2_X1 U9681 ( .A1(n8026), .A2(n8025), .ZN(n8029) );
  OAI211_X1 U9682 ( .C1(n8030), .C2(n8029), .A(n8028), .B(n8027), .ZN(n8032)
         );
  NAND2_X1 U9683 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  INV_X1 U9684 ( .A(n8245), .ZN(n8039) );
  AND2_X1 U9685 ( .A1(n8040), .A2(n8035), .ZN(n8037) );
  MUX2_X1 U9686 ( .A(n8037), .B(n8036), .S(n8078), .Z(n8038) );
  INV_X1 U9687 ( .A(n8238), .ZN(n8234) );
  MUX2_X1 U9688 ( .A(n8041), .B(n8040), .S(n8078), .Z(n8042) );
  NAND3_X1 U9689 ( .A1(n8043), .A2(n8234), .A3(n8042), .ZN(n8052) );
  AND2_X1 U9690 ( .A1(n8208), .A2(n8044), .ZN(n8046) );
  MUX2_X1 U9691 ( .A(n8046), .B(n8045), .S(n8083), .Z(n8051) );
  NAND2_X1 U9692 ( .A1(n8047), .A2(n8207), .ZN(n8049) );
  MUX2_X1 U9693 ( .A(n8049), .B(n8048), .S(n8083), .Z(n8050) );
  AOI21_X1 U9694 ( .B1(n8052), .B2(n8051), .A(n8050), .ZN(n8056) );
  INV_X1 U9695 ( .A(n6227), .ZN(n8053) );
  MUX2_X1 U9696 ( .A(n8054), .B(n8053), .S(n8078), .Z(n8055) );
  OAI21_X1 U9697 ( .B1(n8056), .B2(n8055), .A(n8196), .ZN(n8060) );
  NAND2_X1 U9698 ( .A1(n8214), .A2(n8083), .ZN(n8058) );
  NAND2_X1 U9699 ( .A1(n8187), .A2(n8078), .ZN(n8057) );
  MUX2_X1 U9700 ( .A(n8058), .B(n8057), .S(n8462), .Z(n8059) );
  INV_X1 U9701 ( .A(n8061), .ZN(n8063) );
  MUX2_X1 U9702 ( .A(n8063), .B(n8062), .S(n8078), .Z(n8064) );
  MUX2_X1 U9703 ( .A(n8067), .B(n8066), .S(n8083), .Z(n8069) );
  MUX2_X1 U9704 ( .A(n8174), .B(n8444), .S(n8078), .Z(n8072) );
  INV_X1 U9705 ( .A(n8082), .ZN(n8075) );
  INV_X1 U9706 ( .A(n8076), .ZN(n8079) );
  OAI21_X1 U9707 ( .B1(n8079), .B2(n8078), .A(n8077), .ZN(n8086) );
  NOR2_X1 U9708 ( .A1(n8080), .A2(n8174), .ZN(n8084) );
  XNOR2_X1 U9709 ( .A(n8091), .B(n8090), .ZN(n8099) );
  NAND2_X1 U9710 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  OAI211_X1 U9711 ( .C1(n8096), .C2(n8095), .A(P2_B_REG_SCAN_IN), .B(n8094), 
        .ZN(n8097) );
  OAI21_X1 U9712 ( .B1(n8099), .B2(n8098), .A(n8097), .ZN(P2_U3296) );
  MUX2_X1 U9713 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8100), .S(P2_U3893), .Z(
        P2_U3522) );
  INV_X1 U9714 ( .A(n8101), .ZN(n8167) );
  MUX2_X1 U9715 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8167), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9716 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8174), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9717 ( .A(n8185), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8113), .Z(
        P2_U3518) );
  MUX2_X1 U9718 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8197), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9719 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8214), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9720 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8226), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9721 ( .A(n8215), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8113), .Z(
        P2_U3514) );
  MUX2_X1 U9722 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8227), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9723 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8263), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9724 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8274), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9725 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8262), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9726 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8298), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9727 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8102), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9728 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8103), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9729 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8330), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9730 ( .A(n8104), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8113), .Z(
        P2_U3505) );
  MUX2_X1 U9731 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8371), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9732 ( .A(n8105), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8113), .Z(
        P2_U3503) );
  MUX2_X1 U9733 ( .A(n8106), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8113), .Z(
        P2_U3501) );
  MUX2_X1 U9734 ( .A(n8107), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8113), .Z(
        P2_U3500) );
  MUX2_X1 U9735 ( .A(n8108), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8113), .Z(
        P2_U3499) );
  MUX2_X1 U9736 ( .A(n8109), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8113), .Z(
        P2_U3498) );
  MUX2_X1 U9737 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8110), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9738 ( .A(n8111), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8113), .Z(
        P2_U3496) );
  MUX2_X1 U9739 ( .A(n9885), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8113), .Z(
        P2_U3495) );
  MUX2_X1 U9740 ( .A(n8112), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8113), .Z(
        P2_U3494) );
  MUX2_X1 U9741 ( .A(n9884), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8113), .Z(
        P2_U3493) );
  MUX2_X1 U9742 ( .A(n6731), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8113), .Z(
        P2_U3492) );
  MUX2_X1 U9743 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6214), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U9744 ( .B1(n4486), .B2(n8115), .A(n8114), .ZN(n8129) );
  AOI21_X1 U9745 ( .B1(n8118), .B2(n8117), .A(n8116), .ZN(n8122) );
  NAND2_X1 U9746 ( .A1(n9858), .A2(n8119), .ZN(n8121) );
  OAI211_X1 U9747 ( .C1(n8122), .C2(n9847), .A(n8121), .B(n8120), .ZN(n8127)
         );
  AOI21_X1 U9748 ( .B1(n4491), .B2(n8124), .A(n8123), .ZN(n8125) );
  NOR2_X1 U9749 ( .A1(n8125), .A2(n9872), .ZN(n8126) );
  AOI211_X1 U9750 ( .C1(n9856), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8127), .B(
        n8126), .ZN(n8128) );
  OAI21_X1 U9751 ( .B1(n8129), .B2(n9849), .A(n8128), .ZN(P2_U3196) );
  AOI21_X1 U9752 ( .B1(n4487), .B2(n8131), .A(n8130), .ZN(n8147) );
  NOR2_X1 U9753 ( .A1(n8133), .A2(n8132), .ZN(n8135) );
  XOR2_X1 U9754 ( .A(n8135), .B(n8134), .Z(n8145) );
  NAND2_X1 U9755 ( .A1(n9856), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8137) );
  OAI211_X1 U9756 ( .C1(n9841), .C2(n8138), .A(n8137), .B(n8136), .ZN(n8144)
         );
  AOI21_X1 U9757 ( .B1(n8141), .B2(n8140), .A(n8139), .ZN(n8142) );
  NOR2_X1 U9758 ( .A1(n8142), .A2(n9872), .ZN(n8143) );
  AOI211_X1 U9759 ( .C1(n9868), .C2(n8145), .A(n8144), .B(n8143), .ZN(n8146)
         );
  OAI21_X1 U9760 ( .B1(n8147), .B2(n9849), .A(n8146), .ZN(P2_U3198) );
  NOR2_X1 U9761 ( .A1(n8149), .A2(n8148), .ZN(n8436) );
  NOR2_X1 U9762 ( .A1(n8150), .A2(n8355), .ZN(n8159) );
  AOI21_X1 U9763 ( .B1(n8436), .B2(n8373), .A(n8159), .ZN(n8153) );
  NAND2_X1 U9764 ( .A1(n8340), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8151) );
  OAI211_X1 U9765 ( .C1(n8438), .C2(n8288), .A(n8153), .B(n8151), .ZN(P2_U3202) );
  NAND2_X1 U9766 ( .A1(n8340), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8152) );
  OAI211_X1 U9767 ( .C1(n8154), .C2(n8288), .A(n8153), .B(n8152), .ZN(P2_U3203) );
  INV_X1 U9768 ( .A(n8155), .ZN(n8163) );
  NAND2_X1 U9769 ( .A1(n8156), .A2(n8373), .ZN(n8161) );
  NOR2_X1 U9770 ( .A1(n8157), .A2(n8288), .ZN(n8158) );
  AOI211_X1 U9771 ( .C1(n8340), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8159), .B(
        n8158), .ZN(n8160) );
  OAI211_X1 U9772 ( .C1(n8163), .C2(n8162), .A(n8161), .B(n8160), .ZN(P2_U3204) );
  XOR2_X1 U9773 ( .A(n8165), .B(n8164), .Z(n8447) );
  INV_X1 U9774 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8168) );
  AOI22_X1 U9775 ( .A1(n8444), .A2(n9889), .B1(n9890), .B2(n8169), .ZN(n8170)
         );
  XOR2_X1 U9776 ( .A(n8173), .B(n8171), .Z(n8453) );
  XOR2_X1 U9777 ( .A(n8173), .B(n8172), .Z(n8175) );
  AOI222_X1 U9778 ( .A1(n6212), .A2(n8175), .B1(n8197), .B2(n9883), .C1(n8174), 
        .C2(n8370), .ZN(n8448) );
  MUX2_X1 U9779 ( .A(n8176), .B(n8448), .S(n8373), .Z(n8179) );
  AOI22_X1 U9780 ( .A1(n8450), .A2(n9889), .B1(n9890), .B2(n8177), .ZN(n8178)
         );
  OAI211_X1 U9781 ( .C1(n8453), .C2(n8378), .A(n8179), .B(n8178), .ZN(P2_U3206) );
  XNOR2_X1 U9782 ( .A(n8181), .B(n8180), .ZN(n8459) );
  INV_X1 U9783 ( .A(n8182), .ZN(n8190) );
  XNOR2_X1 U9784 ( .A(n8184), .B(n8183), .ZN(n8189) );
  NAND2_X1 U9785 ( .A1(n8185), .A2(n8370), .ZN(n8186) );
  OAI21_X1 U9786 ( .B1(n8187), .B2(n8351), .A(n8186), .ZN(n8188) );
  AOI21_X1 U9787 ( .B1(n8189), .B2(n6212), .A(n8188), .ZN(n8454) );
  OAI21_X1 U9788 ( .B1(n8190), .B2(n8355), .A(n8454), .ZN(n8191) );
  NAND2_X1 U9789 ( .A1(n8191), .A2(n8373), .ZN(n8193) );
  AOI22_X1 U9790 ( .A1(n8456), .A2(n9889), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8340), .ZN(n8192) );
  OAI211_X1 U9791 ( .C1(n8459), .C2(n8378), .A(n8193), .B(n8192), .ZN(P2_U3207) );
  XNOR2_X1 U9792 ( .A(n8194), .B(n8196), .ZN(n8465) );
  XOR2_X1 U9793 ( .A(n8196), .B(n8195), .Z(n8198) );
  AOI222_X1 U9794 ( .A1(n6212), .A2(n8198), .B1(n8197), .B2(n8370), .C1(n8226), 
        .C2(n9883), .ZN(n8460) );
  INV_X1 U9795 ( .A(n8460), .ZN(n8203) );
  INV_X1 U9796 ( .A(n8462), .ZN(n8201) );
  INV_X1 U9797 ( .A(n8199), .ZN(n8200) );
  OAI22_X1 U9798 ( .A1(n8201), .A2(n8336), .B1(n8200), .B2(n8355), .ZN(n8202)
         );
  OAI21_X1 U9799 ( .B1(n8203), .B2(n8202), .A(n8373), .ZN(n8205) );
  NAND2_X1 U9800 ( .A1(n8340), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8204) );
  OAI211_X1 U9801 ( .C1(n8465), .C2(n8378), .A(n8205), .B(n8204), .ZN(P2_U3208) );
  INV_X1 U9802 ( .A(n8207), .ZN(n8209) );
  OAI21_X1 U9803 ( .B1(n8206), .B2(n8209), .A(n8208), .ZN(n8211) );
  XNOR2_X1 U9804 ( .A(n8211), .B(n8210), .ZN(n8471) );
  XNOR2_X1 U9805 ( .A(n8212), .B(n8213), .ZN(n8216) );
  AOI222_X1 U9806 ( .A1(n6212), .A2(n8216), .B1(n8215), .B2(n9883), .C1(n8214), 
        .C2(n8370), .ZN(n8466) );
  INV_X1 U9807 ( .A(n8466), .ZN(n8221) );
  INV_X1 U9808 ( .A(n8217), .ZN(n8218) );
  OAI22_X1 U9809 ( .A1(n8219), .A2(n8336), .B1(n8218), .B2(n8355), .ZN(n8220)
         );
  OAI21_X1 U9810 ( .B1(n8221), .B2(n8220), .A(n8373), .ZN(n8223) );
  NAND2_X1 U9811 ( .A1(n8340), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8222) );
  OAI211_X1 U9812 ( .C1(n8471), .C2(n8378), .A(n8223), .B(n8222), .ZN(P2_U3209) );
  XNOR2_X1 U9813 ( .A(n8206), .B(n8225), .ZN(n8477) );
  INV_X1 U9814 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8229) );
  XOR2_X1 U9815 ( .A(n8224), .B(n8225), .Z(n8228) );
  AOI222_X1 U9816 ( .A1(n6212), .A2(n8228), .B1(n8227), .B2(n9883), .C1(n8226), 
        .C2(n8370), .ZN(n8472) );
  MUX2_X1 U9817 ( .A(n8229), .B(n8472), .S(n8373), .Z(n8232) );
  AOI22_X1 U9818 ( .A1(n8474), .A2(n9889), .B1(n9890), .B2(n8230), .ZN(n8231)
         );
  OAI211_X1 U9819 ( .C1(n8477), .C2(n8378), .A(n8232), .B(n8231), .ZN(P2_U3210) );
  XNOR2_X1 U9820 ( .A(n8233), .B(n8234), .ZN(n8235) );
  OAI222_X1 U9821 ( .A1(n8351), .A2(n8237), .B1(n8349), .B2(n8236), .C1(n8347), 
        .C2(n8235), .ZN(n8398) );
  INV_X1 U9822 ( .A(n8398), .ZN(n8244) );
  XNOR2_X1 U9823 ( .A(n8239), .B(n8238), .ZN(n8399) );
  AOI22_X1 U9824 ( .A1(n8340), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9890), .B2(
        n8240), .ZN(n8241) );
  OAI21_X1 U9825 ( .B1(n8481), .B2(n8288), .A(n8241), .ZN(n8242) );
  AOI21_X1 U9826 ( .B1(n8399), .B2(n9892), .A(n8242), .ZN(n8243) );
  OAI21_X1 U9827 ( .B1(n8244), .B2(n8340), .A(n8243), .ZN(P2_U3211) );
  NAND2_X1 U9828 ( .A1(n8246), .A2(n8245), .ZN(n8247) );
  XNOR2_X1 U9829 ( .A(n8247), .B(n8249), .ZN(n8484) );
  XOR2_X1 U9830 ( .A(n8249), .B(n8248), .Z(n8250) );
  OAI222_X1 U9831 ( .A1(n8351), .A2(n8252), .B1(n8349), .B2(n8251), .C1(n8347), 
        .C2(n8250), .ZN(n8402) );
  NAND2_X1 U9832 ( .A1(n8402), .A2(n8373), .ZN(n8258) );
  INV_X1 U9833 ( .A(n8253), .ZN(n8254) );
  OAI22_X1 U9834 ( .A1(n8373), .A2(n8255), .B1(n8254), .B2(n8355), .ZN(n8256)
         );
  AOI21_X1 U9835 ( .B1(n8403), .B2(n9889), .A(n8256), .ZN(n8257) );
  OAI211_X1 U9836 ( .C1(n8484), .C2(n8378), .A(n8258), .B(n8257), .ZN(P2_U3212) );
  XNOR2_X1 U9837 ( .A(n8259), .B(n8261), .ZN(n8490) );
  INV_X1 U9838 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8265) );
  OAI21_X1 U9839 ( .B1(n4471), .B2(n8261), .A(n8260), .ZN(n8264) );
  AOI222_X1 U9840 ( .A1(n6212), .A2(n8264), .B1(n8263), .B2(n8370), .C1(n8262), 
        .C2(n9883), .ZN(n8485) );
  MUX2_X1 U9841 ( .A(n8265), .B(n8485), .S(n8373), .Z(n8268) );
  AOI22_X1 U9842 ( .A1(n8487), .A2(n9889), .B1(n9890), .B2(n8266), .ZN(n8267)
         );
  OAI211_X1 U9843 ( .C1(n8490), .C2(n8378), .A(n8268), .B(n8267), .ZN(P2_U3213) );
  XOR2_X1 U9844 ( .A(n8270), .B(n8269), .Z(n8493) );
  NAND2_X1 U9845 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  NAND3_X1 U9846 ( .A1(n8273), .A2(n6212), .A3(n8272), .ZN(n8276) );
  AOI22_X1 U9847 ( .A1(n8274), .A2(n8370), .B1(n9883), .B2(n8298), .ZN(n8275)
         );
  NAND2_X1 U9848 ( .A1(n8276), .A2(n8275), .ZN(n8491) );
  NOR2_X1 U9849 ( .A1(n8355), .A2(n8277), .ZN(n8278) );
  OAI21_X1 U9850 ( .B1(n8491), .B2(n8278), .A(n8373), .ZN(n8281) );
  AOI22_X1 U9851 ( .A1(n8279), .A2(n9889), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n8340), .ZN(n8280) );
  OAI211_X1 U9852 ( .C1(n8493), .C2(n8378), .A(n8281), .B(n8280), .ZN(P2_U3214) );
  XNOR2_X1 U9853 ( .A(n8282), .B(n8285), .ZN(n8283) );
  OAI222_X1 U9854 ( .A1(n8349), .A2(n8284), .B1(n8351), .B2(n8310), .C1(n8283), 
        .C2(n8347), .ZN(n8411) );
  INV_X1 U9855 ( .A(n8411), .ZN(n8294) );
  AOI21_X1 U9856 ( .B1(n8286), .B2(n8285), .A(n4489), .ZN(n8412) );
  INV_X1 U9857 ( .A(n8287), .ZN(n8499) );
  NOR2_X1 U9858 ( .A1(n8499), .A2(n8288), .ZN(n8292) );
  OAI22_X1 U9859 ( .A1(n8373), .A2(n8290), .B1(n8289), .B2(n8355), .ZN(n8291)
         );
  AOI211_X1 U9860 ( .C1(n8412), .C2(n9892), .A(n8292), .B(n8291), .ZN(n8293)
         );
  OAI21_X1 U9861 ( .B1(n8294), .B2(n8340), .A(n8293), .ZN(P2_U3215) );
  XNOR2_X1 U9862 ( .A(n8295), .B(n8297), .ZN(n8505) );
  XNOR2_X1 U9863 ( .A(n8296), .B(n8297), .ZN(n8301) );
  NAND2_X1 U9864 ( .A1(n8298), .A2(n8370), .ZN(n8299) );
  OAI21_X1 U9865 ( .B1(n8321), .B2(n8351), .A(n8299), .ZN(n8300) );
  AOI21_X1 U9866 ( .B1(n8301), .B2(n6212), .A(n8300), .ZN(n8500) );
  MUX2_X1 U9867 ( .A(n10211), .B(n8500), .S(n8373), .Z(n8304) );
  AOI22_X1 U9868 ( .A1(n8502), .A2(n9889), .B1(n8302), .B2(n9890), .ZN(n8303)
         );
  OAI211_X1 U9869 ( .C1(n8505), .C2(n8378), .A(n8304), .B(n8303), .ZN(P2_U3216) );
  XNOR2_X1 U9870 ( .A(n8305), .B(n8307), .ZN(n8511) );
  INV_X1 U9871 ( .A(n8307), .ZN(n8308) );
  XNOR2_X1 U9872 ( .A(n8306), .B(n8308), .ZN(n8312) );
  NAND2_X1 U9873 ( .A1(n8330), .A2(n9883), .ZN(n8309) );
  OAI21_X1 U9874 ( .B1(n8310), .B2(n8349), .A(n8309), .ZN(n8311) );
  AOI21_X1 U9875 ( .B1(n8312), .B2(n6212), .A(n8311), .ZN(n8506) );
  MUX2_X1 U9876 ( .A(n10125), .B(n8506), .S(n8373), .Z(n8316) );
  INV_X1 U9877 ( .A(n8313), .ZN(n8314) );
  AOI22_X1 U9878 ( .A1(n8508), .A2(n9889), .B1(n9890), .B2(n8314), .ZN(n8315)
         );
  OAI211_X1 U9879 ( .C1(n8511), .C2(n8378), .A(n8316), .B(n8315), .ZN(P2_U3217) );
  XNOR2_X1 U9880 ( .A(n8317), .B(n8318), .ZN(n8515) );
  XOR2_X1 U9881 ( .A(n8319), .B(n8318), .Z(n8320) );
  OAI222_X1 U9882 ( .A1(n8349), .A2(n8321), .B1(n8351), .B2(n8348), .C1(n8320), 
        .C2(n8347), .ZN(n8512) );
  INV_X1 U9883 ( .A(n8512), .ZN(n8420) );
  MUX2_X1 U9884 ( .A(n8322), .B(n8420), .S(n8373), .Z(n8325) );
  AOI22_X1 U9885 ( .A1(n8421), .A2(n9889), .B1(n9890), .B2(n8323), .ZN(n8324)
         );
  OAI211_X1 U9886 ( .C1(n8515), .C2(n8378), .A(n8325), .B(n8324), .ZN(P2_U3218) );
  XNOR2_X1 U9887 ( .A(n8327), .B(n8326), .ZN(n8523) );
  XNOR2_X1 U9888 ( .A(n8328), .B(n8329), .ZN(n8334) );
  NAND2_X1 U9889 ( .A1(n8330), .A2(n8370), .ZN(n8331) );
  OAI21_X1 U9890 ( .B1(n8332), .B2(n8351), .A(n8331), .ZN(n8333) );
  AOI21_X1 U9891 ( .B1(n8334), .B2(n6212), .A(n8333), .ZN(n8519) );
  INV_X1 U9892 ( .A(n8519), .ZN(n8339) );
  OAI22_X1 U9893 ( .A1(n8337), .A2(n8336), .B1(n8335), .B2(n8355), .ZN(n8338)
         );
  OAI21_X1 U9894 ( .B1(n8339), .B2(n8338), .A(n8373), .ZN(n8342) );
  NAND2_X1 U9895 ( .A1(n8340), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8341) );
  OAI211_X1 U9896 ( .C1(n8523), .C2(n8378), .A(n8342), .B(n8341), .ZN(P2_U3219) );
  INV_X1 U9897 ( .A(n8343), .ZN(n8344) );
  AOI21_X1 U9898 ( .B1(n8353), .B2(n8345), .A(n8344), .ZN(n8346) );
  OAI222_X1 U9899 ( .A1(n8351), .A2(n8350), .B1(n8349), .B2(n8348), .C1(n8347), 
        .C2(n8346), .ZN(n8427) );
  AOI21_X1 U9900 ( .B1(n8352), .B2(n8526), .A(n8427), .ZN(n8360) );
  XOR2_X1 U9901 ( .A(n8354), .B(n8353), .Z(n8528) );
  OAI22_X1 U9902 ( .A1(n8373), .A2(n8357), .B1(n8356), .B2(n8355), .ZN(n8358)
         );
  AOI21_X1 U9903 ( .B1(n8528), .B2(n9892), .A(n8358), .ZN(n8359) );
  OAI21_X1 U9904 ( .B1(n8360), .B2(n8340), .A(n8359), .ZN(P2_U3220) );
  INV_X1 U9905 ( .A(n8361), .ZN(n8364) );
  OAI21_X1 U9906 ( .B1(n8364), .B2(n8363), .A(n8362), .ZN(n8366) );
  NAND2_X1 U9907 ( .A1(n8366), .A2(n8365), .ZN(n8538) );
  XNOR2_X1 U9908 ( .A(n8368), .B(n8367), .ZN(n8372) );
  AOI222_X1 U9909 ( .A1(n6212), .A2(n8372), .B1(n8371), .B2(n8370), .C1(n8369), 
        .C2(n9883), .ZN(n8531) );
  MUX2_X1 U9910 ( .A(n8374), .B(n8531), .S(n8373), .Z(n8377) );
  AOI22_X1 U9911 ( .A1(n9889), .A2(n8533), .B1(n9890), .B2(n8375), .ZN(n8376)
         );
  OAI211_X1 U9912 ( .C1(n8538), .C2(n8378), .A(n8377), .B(n8376), .ZN(P2_U3221) );
  NAND2_X1 U9913 ( .A1(n8379), .A2(n8432), .ZN(n8380) );
  NAND2_X1 U9914 ( .A1(n8436), .A2(n9951), .ZN(n8381) );
  OAI211_X1 U9915 ( .C1(n9951), .C2(n7897), .A(n8380), .B(n8381), .ZN(P2_U3490) );
  INV_X1 U9916 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U9917 ( .A1(n8439), .A2(n8432), .ZN(n8382) );
  OAI211_X1 U9918 ( .C1(n9951), .C2(n10024), .A(n8382), .B(n8381), .ZN(
        P2_U3489) );
  MUX2_X1 U9919 ( .A(n8383), .B(n8442), .S(n9951), .Z(n8385) );
  NAND2_X1 U9920 ( .A1(n8444), .A2(n8432), .ZN(n8384) );
  OAI211_X1 U9921 ( .C1(n8447), .C2(n8435), .A(n8385), .B(n8384), .ZN(P2_U3487) );
  MUX2_X1 U9922 ( .A(n10224), .B(n8448), .S(n9951), .Z(n8387) );
  NAND2_X1 U9923 ( .A1(n8450), .A2(n8432), .ZN(n8386) );
  OAI211_X1 U9924 ( .C1(n8453), .C2(n8435), .A(n8387), .B(n8386), .ZN(P2_U3486) );
  MUX2_X1 U9925 ( .A(n10130), .B(n8454), .S(n9951), .Z(n8389) );
  NAND2_X1 U9926 ( .A1(n8456), .A2(n8432), .ZN(n8388) );
  OAI211_X1 U9927 ( .C1(n8435), .C2(n8459), .A(n8389), .B(n8388), .ZN(P2_U3485) );
  MUX2_X1 U9928 ( .A(n8390), .B(n8460), .S(n9951), .Z(n8392) );
  NAND2_X1 U9929 ( .A1(n8462), .A2(n8432), .ZN(n8391) );
  OAI211_X1 U9930 ( .C1(n8435), .C2(n8465), .A(n8392), .B(n8391), .ZN(P2_U3484) );
  MUX2_X1 U9931 ( .A(n8393), .B(n8466), .S(n9951), .Z(n8395) );
  NAND2_X1 U9932 ( .A1(n8468), .A2(n8432), .ZN(n8394) );
  OAI211_X1 U9933 ( .C1(n8435), .C2(n8471), .A(n8395), .B(n8394), .ZN(P2_U3483) );
  MUX2_X1 U9934 ( .A(n10240), .B(n8472), .S(n9951), .Z(n8397) );
  NAND2_X1 U9935 ( .A1(n8474), .A2(n8432), .ZN(n8396) );
  OAI211_X1 U9936 ( .C1(n8477), .C2(n8435), .A(n8397), .B(n8396), .ZN(P2_U3482) );
  INV_X1 U9937 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8400) );
  AOI21_X1 U9938 ( .B1(n9938), .B2(n8399), .A(n8398), .ZN(n8478) );
  MUX2_X1 U9939 ( .A(n8400), .B(n8478), .S(n9951), .Z(n8401) );
  OAI21_X1 U9940 ( .B1(n8481), .B2(n8414), .A(n8401), .ZN(P2_U3481) );
  AOI21_X1 U9941 ( .B1(n9918), .B2(n8403), .A(n8402), .ZN(n8482) );
  MUX2_X1 U9942 ( .A(n8404), .B(n8482), .S(n9951), .Z(n8405) );
  OAI21_X1 U9943 ( .B1(n8435), .B2(n8484), .A(n8405), .ZN(P2_U3480) );
  MUX2_X1 U9944 ( .A(n8406), .B(n8485), .S(n9951), .Z(n8408) );
  NAND2_X1 U9945 ( .A1(n8487), .A2(n8432), .ZN(n8407) );
  OAI211_X1 U9946 ( .C1(n8435), .C2(n8490), .A(n8408), .B(n8407), .ZN(P2_U3479) );
  MUX2_X1 U9947 ( .A(n8491), .B(P2_REG1_REG_19__SCAN_IN), .S(n6296), .Z(n8410)
         );
  OAI22_X1 U9948 ( .A1(n8493), .A2(n8435), .B1(n8492), .B2(n8414), .ZN(n8409)
         );
  OR2_X1 U9949 ( .A1(n8410), .A2(n8409), .ZN(P2_U3478) );
  AOI21_X1 U9950 ( .B1(n8412), .B2(n9938), .A(n8411), .ZN(n8496) );
  MUX2_X1 U9951 ( .A(n10222), .B(n8496), .S(n9951), .Z(n8413) );
  OAI21_X1 U9952 ( .B1(n8499), .B2(n8414), .A(n8413), .ZN(P2_U3477) );
  MUX2_X1 U9953 ( .A(n10128), .B(n8500), .S(n9951), .Z(n8416) );
  NAND2_X1 U9954 ( .A1(n8502), .A2(n8432), .ZN(n8415) );
  OAI211_X1 U9955 ( .C1(n8505), .C2(n8435), .A(n8416), .B(n8415), .ZN(P2_U3476) );
  MUX2_X1 U9956 ( .A(n8417), .B(n8506), .S(n9951), .Z(n8419) );
  NAND2_X1 U9957 ( .A1(n8508), .A2(n8432), .ZN(n8418) );
  OAI211_X1 U9958 ( .C1(n8435), .C2(n8511), .A(n8419), .B(n8418), .ZN(P2_U3475) );
  MUX2_X1 U9959 ( .A(n10055), .B(n8420), .S(n9951), .Z(n8423) );
  NAND2_X1 U9960 ( .A1(n8421), .A2(n8432), .ZN(n8422) );
  OAI211_X1 U9961 ( .C1(n8515), .C2(n8435), .A(n8423), .B(n8422), .ZN(P2_U3474) );
  MUX2_X1 U9962 ( .A(n8519), .B(n8424), .S(n6296), .Z(n8426) );
  NAND2_X1 U9963 ( .A1(n8520), .A2(n8432), .ZN(n8425) );
  OAI211_X1 U9964 ( .C1(n8523), .C2(n8435), .A(n8426), .B(n8425), .ZN(P2_U3473) );
  INV_X1 U9965 ( .A(n8427), .ZN(n8524) );
  MUX2_X1 U9966 ( .A(n9821), .B(n8524), .S(n9951), .Z(n8430) );
  INV_X1 U9967 ( .A(n8435), .ZN(n8428) );
  AOI22_X1 U9968 ( .A1(n8528), .A2(n8428), .B1(n8432), .B2(n8526), .ZN(n8429)
         );
  NAND2_X1 U9969 ( .A1(n8430), .A2(n8429), .ZN(P2_U3472) );
  MUX2_X1 U9970 ( .A(n8431), .B(n8531), .S(n9951), .Z(n8434) );
  NAND2_X1 U9971 ( .A1(n8432), .A2(n8533), .ZN(n8433) );
  OAI211_X1 U9972 ( .C1(n8435), .C2(n8538), .A(n8434), .B(n8433), .ZN(P2_U3471) );
  NAND2_X1 U9973 ( .A1(n9941), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U9974 ( .A1(n8436), .A2(n9939), .ZN(n8440) );
  OAI211_X1 U9975 ( .C1(n8438), .C2(n8513), .A(n8437), .B(n8440), .ZN(P2_U3458) );
  NAND2_X1 U9976 ( .A1(n8439), .A2(n8534), .ZN(n8441) );
  OAI211_X1 U9977 ( .C1(n9939), .C2(n10174), .A(n8441), .B(n8440), .ZN(
        P2_U3457) );
  INV_X1 U9978 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8443) );
  MUX2_X1 U9979 ( .A(n8443), .B(n8442), .S(n9939), .Z(n8446) );
  NAND2_X1 U9980 ( .A1(n8444), .A2(n8534), .ZN(n8445) );
  OAI211_X1 U9981 ( .C1(n8447), .C2(n8537), .A(n8446), .B(n8445), .ZN(P2_U3455) );
  INV_X1 U9982 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8449) );
  MUX2_X1 U9983 ( .A(n8449), .B(n8448), .S(n9939), .Z(n8452) );
  NAND2_X1 U9984 ( .A1(n8450), .A2(n8534), .ZN(n8451) );
  OAI211_X1 U9985 ( .C1(n8453), .C2(n8537), .A(n8452), .B(n8451), .ZN(P2_U3454) );
  INV_X1 U9986 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8455) );
  MUX2_X1 U9987 ( .A(n8455), .B(n8454), .S(n9939), .Z(n8458) );
  NAND2_X1 U9988 ( .A1(n8456), .A2(n8534), .ZN(n8457) );
  OAI211_X1 U9989 ( .C1(n8459), .C2(n8537), .A(n8458), .B(n8457), .ZN(P2_U3453) );
  INV_X1 U9990 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8461) );
  MUX2_X1 U9991 ( .A(n8461), .B(n8460), .S(n9939), .Z(n8464) );
  NAND2_X1 U9992 ( .A1(n8462), .A2(n8534), .ZN(n8463) );
  OAI211_X1 U9993 ( .C1(n8465), .C2(n8537), .A(n8464), .B(n8463), .ZN(P2_U3452) );
  INV_X1 U9994 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8467) );
  MUX2_X1 U9995 ( .A(n8467), .B(n8466), .S(n9939), .Z(n8470) );
  NAND2_X1 U9996 ( .A1(n8468), .A2(n8534), .ZN(n8469) );
  OAI211_X1 U9997 ( .C1(n8471), .C2(n8537), .A(n8470), .B(n8469), .ZN(P2_U3451) );
  INV_X1 U9998 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U9999 ( .A(n8473), .B(n8472), .S(n9939), .Z(n8476) );
  NAND2_X1 U10000 ( .A1(n8474), .A2(n8534), .ZN(n8475) );
  OAI211_X1 U10001 ( .C1(n8477), .C2(n8537), .A(n8476), .B(n8475), .ZN(
        P2_U3450) );
  INV_X1 U10002 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8479) );
  MUX2_X1 U10003 ( .A(n8479), .B(n8478), .S(n9939), .Z(n8480) );
  OAI21_X1 U10004 ( .B1(n8481), .B2(n8513), .A(n8480), .ZN(P2_U3449) );
  MUX2_X1 U10005 ( .A(n10083), .B(n8482), .S(n9939), .Z(n8483) );
  OAI21_X1 U10006 ( .B1(n8484), .B2(n8537), .A(n8483), .ZN(P2_U3448) );
  MUX2_X1 U10007 ( .A(n8486), .B(n8485), .S(n9939), .Z(n8489) );
  NAND2_X1 U10008 ( .A1(n8487), .A2(n8534), .ZN(n8488) );
  OAI211_X1 U10009 ( .C1(n8490), .C2(n8537), .A(n8489), .B(n8488), .ZN(
        P2_U3447) );
  MUX2_X1 U10010 ( .A(n8491), .B(P2_REG0_REG_19__SCAN_IN), .S(n9941), .Z(n8495) );
  OAI22_X1 U10011 ( .A1(n8493), .A2(n8537), .B1(n8492), .B2(n8513), .ZN(n8494)
         );
  OR2_X1 U10012 ( .A1(n8495), .A2(n8494), .ZN(P2_U3446) );
  INV_X1 U10013 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8497) );
  MUX2_X1 U10014 ( .A(n8497), .B(n8496), .S(n9939), .Z(n8498) );
  OAI21_X1 U10015 ( .B1(n8499), .B2(n8513), .A(n8498), .ZN(P2_U3444) );
  INV_X1 U10016 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8501) );
  MUX2_X1 U10017 ( .A(n8501), .B(n8500), .S(n9939), .Z(n8504) );
  NAND2_X1 U10018 ( .A1(n8502), .A2(n8534), .ZN(n8503) );
  OAI211_X1 U10019 ( .C1(n8505), .C2(n8537), .A(n8504), .B(n8503), .ZN(
        P2_U3441) );
  INV_X1 U10020 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8507) );
  MUX2_X1 U10021 ( .A(n8507), .B(n8506), .S(n9939), .Z(n8510) );
  NAND2_X1 U10022 ( .A1(n8508), .A2(n8534), .ZN(n8509) );
  OAI211_X1 U10023 ( .C1(n8511), .C2(n8537), .A(n8510), .B(n8509), .ZN(
        P2_U3438) );
  MUX2_X1 U10024 ( .A(n8512), .B(P2_REG0_REG_15__SCAN_IN), .S(n9941), .Z(n8517) );
  OAI22_X1 U10025 ( .A1(n8515), .A2(n8537), .B1(n8514), .B2(n8513), .ZN(n8516)
         );
  OR2_X1 U10026 ( .A1(n8517), .A2(n8516), .ZN(P2_U3435) );
  INV_X1 U10027 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8518) );
  MUX2_X1 U10028 ( .A(n8519), .B(n8518), .S(n9941), .Z(n8522) );
  NAND2_X1 U10029 ( .A1(n8520), .A2(n8534), .ZN(n8521) );
  OAI211_X1 U10030 ( .C1(n8523), .C2(n8537), .A(n8522), .B(n8521), .ZN(
        P2_U3432) );
  INV_X1 U10031 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8525) );
  MUX2_X1 U10032 ( .A(n8525), .B(n8524), .S(n9939), .Z(n8530) );
  INV_X1 U10033 ( .A(n8537), .ZN(n8527) );
  AOI22_X1 U10034 ( .A1(n8528), .A2(n8527), .B1(n8534), .B2(n8526), .ZN(n8529)
         );
  NAND2_X1 U10035 ( .A1(n8530), .A2(n8529), .ZN(P2_U3429) );
  INV_X1 U10036 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10037 ( .A(n8532), .B(n8531), .S(n9939), .Z(n8536) );
  NAND2_X1 U10038 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  OAI211_X1 U10039 ( .C1(n8538), .C2(n8537), .A(n8536), .B(n8535), .ZN(
        P2_U3426) );
  INV_X1 U10040 ( .A(n8813), .ZN(n9412) );
  NAND3_X1 U10041 ( .A1(n5811), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8541) );
  OAI22_X1 U10042 ( .A1(n8539), .A2(n8541), .B1(n10158), .B2(n8540), .ZN(n8542) );
  INV_X1 U10043 ( .A(n8542), .ZN(n8543) );
  OAI21_X1 U10044 ( .B1(n9412), .B2(n8546), .A(n8543), .ZN(P2_U3264) );
  OAI222_X1 U10045 ( .A1(n8546), .A2(n8545), .B1(n8544), .B2(P2_U3151), .C1(
        n10065), .C2(n8547), .ZN(P2_U3267) );
  OAI222_X1 U10046 ( .A1(n8550), .A2(n8549), .B1(n8548), .B2(P2_U3151), .C1(
        n10163), .C2(n8547), .ZN(P2_U3268) );
  MUX2_X1 U10047 ( .A(n8551), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10048 ( .A(n8552), .ZN(n8553) );
  AOI21_X1 U10049 ( .B1(n8555), .B2(n8554), .A(n8553), .ZN(n8562) );
  NAND2_X1 U10050 ( .A1(n8734), .A2(n8981), .ZN(n8557) );
  OAI211_X1 U10051 ( .C1(n8633), .C2(n8737), .A(n8557), .B(n8556), .ZN(n8559)
         );
  NOR2_X1 U10052 ( .A1(n9666), .A2(n8739), .ZN(n8558) );
  AOI211_X1 U10053 ( .C1(n8560), .C2(n8742), .A(n8559), .B(n8558), .ZN(n8561)
         );
  OAI21_X1 U10054 ( .B1(n8562), .B2(n8745), .A(n8561), .ZN(P1_U3215) );
  INV_X1 U10055 ( .A(n8563), .ZN(n8668) );
  AOI21_X1 U10056 ( .B1(n8565), .B2(n8685), .A(n8564), .ZN(n8566) );
  OAI21_X1 U10057 ( .B1(n8668), .B2(n8566), .A(n8722), .ZN(n8570) );
  AOI22_X1 U10058 ( .A1(n8734), .A2(n9345), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8567) );
  OAI21_X1 U10059 ( .B1(n9356), .B2(n8737), .A(n8567), .ZN(n8568) );
  AOI21_X1 U10060 ( .B1(n9214), .B2(n8742), .A(n8568), .ZN(n8569) );
  OAI211_X1 U10061 ( .C1(n4671), .C2(n8739), .A(n8570), .B(n8569), .ZN(
        P1_U3216) );
  XNOR2_X1 U10062 ( .A(n8571), .B(n8573), .ZN(n8720) );
  INV_X1 U10063 ( .A(n8572), .ZN(n8721) );
  NAND2_X1 U10064 ( .A1(n8720), .A2(n8721), .ZN(n8719) );
  INV_X1 U10065 ( .A(n8573), .ZN(n8574) );
  NAND2_X1 U10066 ( .A1(n8571), .A2(n8574), .ZN(n8577) );
  AND2_X1 U10067 ( .A1(n8719), .A2(n8577), .ZN(n8579) );
  XNOR2_X1 U10068 ( .A(n8576), .B(n8575), .ZN(n8578) );
  NAND3_X1 U10069 ( .A1(n8719), .A2(n8578), .A3(n8577), .ZN(n8677) );
  OAI211_X1 U10070 ( .C1(n8579), .C2(n8578), .A(n8722), .B(n8677), .ZN(n8584)
         );
  NAND2_X1 U10071 ( .A1(n8734), .A2(n9370), .ZN(n8581) );
  OAI211_X1 U10072 ( .C1(n9275), .C2(n8737), .A(n8581), .B(n8580), .ZN(n8582)
         );
  AOI21_X1 U10073 ( .B1(n9280), .B2(n8742), .A(n8582), .ZN(n8583) );
  OAI211_X1 U10074 ( .C1(n9283), .C2(n8739), .A(n8584), .B(n8583), .ZN(
        P1_U3219) );
  OR2_X1 U10075 ( .A1(n8823), .A2(n10051), .ZN(n8586) );
  NAND2_X1 U10076 ( .A1(n9328), .A2(n4402), .ZN(n8590) );
  OR2_X1 U10077 ( .A1(n9116), .A2(n8588), .ZN(n8589) );
  NAND2_X1 U10078 ( .A1(n8590), .A2(n8589), .ZN(n8592) );
  XNOR2_X1 U10079 ( .A(n8592), .B(n8591), .ZN(n8596) );
  NAND2_X1 U10080 ( .A1(n9328), .A2(n8593), .ZN(n8594) );
  OAI21_X1 U10081 ( .B1(n9116), .B2(n5593), .A(n8594), .ZN(n8595) );
  XNOR2_X1 U10082 ( .A(n8596), .B(n8595), .ZN(n8608) );
  OR4_X2 U10083 ( .A1(n8597), .A2(n8607), .A3(n8608), .A4(n8745), .ZN(n8612)
         );
  NAND3_X1 U10084 ( .A1(n8597), .A2(n8722), .A3(n8608), .ZN(n8611) );
  NAND2_X1 U10085 ( .A1(n8598), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U10086 ( .A1(n5657), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8602) );
  INV_X1 U10087 ( .A(n8599), .ZN(n9134) );
  NAND2_X1 U10088 ( .A1(n5210), .A2(n9134), .ZN(n8601) );
  NAND2_X1 U10089 ( .A1(n5461), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8600) );
  INV_X1 U10090 ( .A(n8809), .ZN(n9149) );
  AOI22_X1 U10091 ( .A1(n8734), .A2(n9149), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8604) );
  OAI21_X1 U10092 ( .B1(n9325), .B2(n8737), .A(n8604), .ZN(n8606) );
  NOR2_X1 U10093 ( .A1(n9115), .A2(n8739), .ZN(n8605) );
  AOI211_X1 U10094 ( .C1(n9144), .C2(n8742), .A(n8606), .B(n8605), .ZN(n8610)
         );
  NAND3_X1 U10095 ( .A1(n8608), .A2(n8722), .A3(n8607), .ZN(n8609) );
  NAND4_X1 U10096 ( .A1(n8612), .A2(n8611), .A3(n8610), .A4(n8609), .ZN(
        P1_U3220) );
  INV_X1 U10097 ( .A(n8616), .ZN(n8613) );
  NOR2_X1 U10098 ( .A1(n5039), .A2(n8613), .ZN(n8675) );
  NAND3_X1 U10099 ( .A1(n8677), .A2(n8675), .A3(n8676), .ZN(n8674) );
  INV_X1 U10100 ( .A(n8614), .ZN(n8615) );
  AND3_X1 U10101 ( .A1(n8674), .A2(n8616), .A3(n8615), .ZN(n8619) );
  INV_X1 U10102 ( .A(n8617), .ZN(n8618) );
  OAI21_X1 U10103 ( .B1(n8619), .B2(n8618), .A(n8722), .ZN(n8623) );
  NOR2_X1 U10104 ( .A1(n8704), .A2(n9356), .ZN(n8621) );
  INV_X1 U10105 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10039) );
  OAI22_X1 U10106 ( .A1(n8737), .A2(n9276), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10039), .ZN(n8620) );
  AOI211_X1 U10107 ( .C1(n9246), .C2(n8742), .A(n8621), .B(n8620), .ZN(n8622)
         );
  OAI211_X1 U10108 ( .C1(n9250), .C2(n8739), .A(n8623), .B(n8622), .ZN(
        P1_U3223) );
  AND2_X1 U10109 ( .A1(n8624), .A2(n8695), .ZN(n8697) );
  INV_X1 U10110 ( .A(n8625), .ZN(n8627) );
  NOR3_X1 U10111 ( .A1(n8697), .A2(n8627), .A3(n8626), .ZN(n8630) );
  OAI21_X1 U10112 ( .B1(n8630), .B2(n4493), .A(n8722), .ZN(n8637) );
  AOI21_X1 U10113 ( .B1(n8714), .B2(n8985), .A(n8631), .ZN(n8632) );
  OAI21_X1 U10114 ( .B1(n8633), .B2(n8704), .A(n8632), .ZN(n8634) );
  AOI21_X1 U10115 ( .B1(n8635), .B2(n8742), .A(n8634), .ZN(n8636) );
  OAI211_X1 U10116 ( .C1(n9648), .C2(n8739), .A(n8637), .B(n8636), .ZN(
        P1_U3224) );
  OAI21_X1 U10117 ( .B1(n8639), .B2(n8638), .A(n5747), .ZN(n8640) );
  NAND2_X1 U10118 ( .A1(n8640), .A2(n8722), .ZN(n8644) );
  INV_X1 U10119 ( .A(n9332), .ZN(n9185) );
  AOI22_X1 U10120 ( .A1(n8734), .A2(n9185), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8641) );
  OAI21_X1 U10121 ( .B1(n9191), .B2(n8737), .A(n8641), .ZN(n8642) );
  AOI21_X1 U10122 ( .B1(n9189), .B2(n8742), .A(n8642), .ZN(n8643) );
  OAI211_X1 U10123 ( .C1(n9193), .C2(n8739), .A(n8644), .B(n8643), .ZN(
        P1_U3225) );
  OAI21_X1 U10124 ( .B1(n8647), .B2(n8646), .A(n8645), .ZN(n8648) );
  NAND2_X1 U10125 ( .A1(n8648), .A2(n8722), .ZN(n8654) );
  NAND2_X1 U10126 ( .A1(n8734), .A2(n9483), .ZN(n8650) );
  OAI211_X1 U10127 ( .C1(n9514), .C2(n8737), .A(n8650), .B(n8649), .ZN(n8651)
         );
  AOI21_X1 U10128 ( .B1(n8652), .B2(n8742), .A(n8651), .ZN(n8653) );
  OAI211_X1 U10129 ( .C1(n4668), .C2(n8739), .A(n8654), .B(n8653), .ZN(
        P1_U3226) );
  OAI21_X1 U10130 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8658) );
  NAND2_X1 U10131 ( .A1(n8658), .A2(n8722), .ZN(n8664) );
  NAND2_X1 U10132 ( .A1(n8734), .A2(n9299), .ZN(n8660) );
  OAI211_X1 U10133 ( .C1(n8661), .C2(n8737), .A(n8660), .B(n8659), .ZN(n8662)
         );
  AOI21_X1 U10134 ( .B1(n9290), .B2(n8742), .A(n8662), .ZN(n8663) );
  OAI211_X1 U10135 ( .C1(n9509), .C2(n8739), .A(n8664), .B(n8663), .ZN(
        P1_U3228) );
  INV_X1 U10136 ( .A(n8665), .ZN(n8667) );
  NOR3_X1 U10137 ( .A1(n8668), .A2(n8667), .A3(n8666), .ZN(n8669) );
  OAI21_X1 U10138 ( .B1(n8669), .B2(n5676), .A(n8722), .ZN(n8673) );
  INV_X1 U10139 ( .A(n9226), .ZN(n8789) );
  AOI22_X1 U10140 ( .A1(n8734), .A2(n9201), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8670) );
  OAI21_X1 U10141 ( .B1(n8789), .B2(n8737), .A(n8670), .ZN(n8671) );
  AOI21_X1 U10142 ( .B1(n9205), .B2(n8742), .A(n8671), .ZN(n8672) );
  OAI211_X1 U10143 ( .C1(n9208), .C2(n8739), .A(n8673), .B(n8672), .ZN(
        P1_U3229) );
  INV_X1 U10144 ( .A(n8674), .ZN(n8679) );
  AOI21_X1 U10145 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8678) );
  OAI21_X1 U10146 ( .B1(n8679), .B2(n8678), .A(n8722), .ZN(n8683) );
  INV_X1 U10147 ( .A(n9484), .ZN(n9105) );
  AOI22_X1 U10148 ( .A1(n8734), .A2(n9363), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8680) );
  OAI21_X1 U10149 ( .B1(n9105), .B2(n8737), .A(n8680), .ZN(n8681) );
  AOI21_X1 U10150 ( .B1(n9258), .B2(n8742), .A(n8681), .ZN(n8682) );
  OAI211_X1 U10151 ( .C1(n9260), .C2(n8739), .A(n8683), .B(n8682), .ZN(
        P1_U3233) );
  NAND2_X1 U10152 ( .A1(n8685), .A2(n8684), .ZN(n8687) );
  XNOR2_X1 U10153 ( .A(n8687), .B(n8686), .ZN(n8688) );
  NAND2_X1 U10154 ( .A1(n8688), .A2(n8722), .ZN(n8693) );
  NOR2_X1 U10155 ( .A1(n8704), .A2(n8789), .ZN(n8691) );
  OAI22_X1 U10156 ( .A1(n8737), .A2(n9232), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8689), .ZN(n8690) );
  AOI211_X1 U10157 ( .C1(n9230), .C2(n8742), .A(n8691), .B(n8690), .ZN(n8692)
         );
  OAI211_X1 U10158 ( .C1(n9235), .C2(n8739), .A(n8693), .B(n8692), .ZN(
        P1_U3235) );
  INV_X1 U10159 ( .A(n8694), .ZN(n8696) );
  NOR2_X1 U10160 ( .A1(n8696), .A2(n8695), .ZN(n8699) );
  AOI21_X1 U10161 ( .B1(n8699), .B2(n8698), .A(n8697), .ZN(n8708) );
  AOI21_X1 U10162 ( .B1(n8714), .B2(n8986), .A(n8700), .ZN(n8703) );
  NAND2_X1 U10163 ( .A1(n8742), .A2(n8701), .ZN(n8702) );
  OAI211_X1 U10164 ( .C1(n9657), .C2(n8704), .A(n8703), .B(n8702), .ZN(n8705)
         );
  AOI21_X1 U10165 ( .B1(n8706), .B2(n5770), .A(n8705), .ZN(n8707) );
  OAI21_X1 U10166 ( .B1(n8708), .B2(n8745), .A(n8707), .ZN(P1_U3236) );
  AND3_X1 U10167 ( .A1(n8711), .A2(n8710), .A3(n8709), .ZN(n8712) );
  OAI21_X1 U10168 ( .B1(n8713), .B2(n8712), .A(n8722), .ZN(n8718) );
  AOI22_X1 U10169 ( .A1(n8714), .A2(n9569), .B1(n5770), .B2(n9570), .ZN(n8717)
         );
  AOI22_X1 U10170 ( .A1(n8734), .A2(n9586), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8715), .ZN(n8716) );
  NAND3_X1 U10171 ( .A1(n8718), .A2(n8717), .A3(n8716), .ZN(P1_U3237) );
  OAI21_X1 U10172 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8723) );
  NAND2_X1 U10173 ( .A1(n8723), .A2(n8722), .ZN(n8729) );
  NAND2_X1 U10174 ( .A1(n8734), .A2(n9484), .ZN(n8725) );
  OAI211_X1 U10175 ( .C1(n9102), .C2(n8737), .A(n8725), .B(n8724), .ZN(n8726)
         );
  AOI21_X1 U10176 ( .B1(n8727), .B2(n8742), .A(n8726), .ZN(n8728) );
  OAI211_X1 U10177 ( .C1(n9503), .C2(n8739), .A(n8729), .B(n8728), .ZN(
        P1_U3238) );
  NOR2_X1 U10178 ( .A1(n8733), .A2(n8732), .ZN(n8731) );
  AOI21_X1 U10179 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8746) );
  NAND2_X1 U10180 ( .A1(n8734), .A2(n9298), .ZN(n8736) );
  OAI211_X1 U10181 ( .C1(n8738), .C2(n8737), .A(n8736), .B(n8735), .ZN(n8741)
         );
  NOR2_X1 U10182 ( .A1(n9522), .A2(n8739), .ZN(n8740) );
  AOI211_X1 U10183 ( .C1(n8743), .C2(n8742), .A(n8741), .B(n8740), .ZN(n8744)
         );
  OAI21_X1 U10184 ( .B1(n8746), .B2(n8745), .A(n8744), .ZN(P1_U3241) );
  NAND2_X1 U10185 ( .A1(n9339), .A2(n9332), .ZN(n9126) );
  NAND2_X1 U10186 ( .A1(n9346), .A2(n8747), .ZN(n9125) );
  NAND3_X1 U10187 ( .A1(n9126), .A2(n8826), .A3(n9125), .ZN(n8797) );
  OR2_X1 U10188 ( .A1(n9339), .A2(n9332), .ZN(n8873) );
  OR2_X1 U10189 ( .A1(n9346), .A2(n8747), .ZN(n8836) );
  AND2_X1 U10190 ( .A1(n8873), .A2(n8836), .ZN(n8877) );
  INV_X1 U10191 ( .A(n8826), .ZN(n8831) );
  NAND3_X1 U10192 ( .A1(n8952), .A2(n8877), .A3(n8831), .ZN(n8796) );
  NAND2_X1 U10193 ( .A1(n9371), .A2(n9232), .ZN(n9122) );
  AND2_X1 U10194 ( .A1(n9377), .A2(n9276), .ZN(n9120) );
  INV_X1 U10195 ( .A(n9120), .ZN(n8748) );
  AND2_X1 U10196 ( .A1(n9122), .A2(n8748), .ZN(n8881) );
  INV_X1 U10197 ( .A(n8749), .ZN(n8750) );
  NAND2_X1 U10198 ( .A1(n8751), .A2(n8750), .ZN(n8756) );
  INV_X1 U10199 ( .A(n9532), .ZN(n9533) );
  AOI21_X1 U10200 ( .B1(n9534), .B2(n9533), .A(n8752), .ZN(n8754) );
  OR2_X1 U10201 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  NAND2_X1 U10202 ( .A1(n8766), .A2(n8757), .ZN(n8758) );
  NAND2_X1 U10203 ( .A1(n8768), .A2(n8764), .ZN(n8932) );
  AOI21_X1 U10204 ( .B1(n8758), .B2(n8929), .A(n8932), .ZN(n8759) );
  NAND2_X1 U10205 ( .A1(n8770), .A2(n8767), .ZN(n8933) );
  OAI21_X1 U10206 ( .B1(n8759), .B2(n8933), .A(n8936), .ZN(n8760) );
  NAND2_X1 U10207 ( .A1(n8760), .A2(n8939), .ZN(n8762) );
  NAND3_X1 U10208 ( .A1(n8762), .A2(n8937), .A3(n8761), .ZN(n8763) );
  NAND2_X1 U10209 ( .A1(n8767), .A2(n8929), .ZN(n8769) );
  NAND2_X1 U10210 ( .A1(n8771), .A2(n8937), .ZN(n8773) );
  NAND3_X1 U10211 ( .A1(n8773), .A2(n8772), .A3(n8939), .ZN(n8776) );
  OR2_X1 U10212 ( .A1(n9522), .A2(n8981), .ZN(n8774) );
  NAND2_X1 U10213 ( .A1(n8942), .A2(n8774), .ZN(n8777) );
  NOR2_X1 U10214 ( .A1(n8777), .A2(n8775), .ZN(n8943) );
  AOI22_X1 U10215 ( .A1(n8777), .A2(n8891), .B1(n8826), .B2(n9522), .ZN(n8779)
         );
  AOI21_X1 U10216 ( .B1(n8942), .B2(n8981), .A(n8831), .ZN(n8778) );
  OR2_X1 U10217 ( .A1(n9292), .A2(n9102), .ZN(n8893) );
  NAND2_X1 U10218 ( .A1(n9292), .A2(n9102), .ZN(n8780) );
  OR2_X1 U10219 ( .A1(n9384), .A2(n9105), .ZN(n8838) );
  OR2_X1 U10220 ( .A1(n9488), .A2(n9275), .ZN(n8839) );
  AND2_X1 U10221 ( .A1(n8838), .A2(n8839), .ZN(n8781) );
  INV_X1 U10222 ( .A(n8781), .ZN(n8949) );
  NAND2_X1 U10223 ( .A1(n9488), .A2(n9275), .ZN(n9269) );
  NAND2_X1 U10224 ( .A1(n9269), .A2(n8780), .ZN(n8945) );
  NAND2_X1 U10225 ( .A1(n9384), .A2(n9105), .ZN(n8948) );
  INV_X1 U10226 ( .A(n8948), .ZN(n8896) );
  AOI211_X1 U10227 ( .C1(n8781), .C2(n8945), .A(n8896), .B(n9120), .ZN(n8782)
         );
  OAI21_X1 U10228 ( .B1(n8783), .B2(n8949), .A(n8782), .ZN(n8787) );
  NAND2_X1 U10229 ( .A1(n8839), .A2(n8893), .ZN(n8915) );
  OAI211_X1 U10230 ( .C1(n8784), .C2(n8915), .A(n8948), .B(n9269), .ZN(n8785)
         );
  NAND3_X1 U10231 ( .A1(n8785), .A2(n4428), .A3(n8838), .ZN(n8786) );
  MUX2_X1 U10232 ( .A(n8787), .B(n8786), .S(n8826), .Z(n8788) );
  NAND2_X1 U10233 ( .A1(n9250), .A2(n9363), .ZN(n8897) );
  NAND2_X1 U10234 ( .A1(n8897), .A2(n4428), .ZN(n8914) );
  OR2_X1 U10235 ( .A1(n9364), .A2(n9356), .ZN(n8790) );
  NAND2_X1 U10236 ( .A1(n9364), .A2(n9356), .ZN(n9123) );
  INV_X1 U10237 ( .A(n9225), .ZN(n9229) );
  NAND2_X1 U10238 ( .A1(n9213), .A2(n8789), .ZN(n8875) );
  NAND2_X1 U10239 ( .A1(n8875), .A2(n9123), .ZN(n8880) );
  OR2_X1 U10240 ( .A1(n9213), .A2(n8789), .ZN(n8837) );
  NAND2_X1 U10241 ( .A1(n8837), .A2(n8790), .ZN(n8874) );
  MUX2_X1 U10242 ( .A(n8880), .B(n8874), .S(n8826), .Z(n8792) );
  NAND2_X1 U10243 ( .A1(n9353), .A2(n9191), .ZN(n8885) );
  MUX2_X1 U10244 ( .A(n8837), .B(n8875), .S(n8826), .Z(n8791) );
  OAI211_X1 U10245 ( .C1(n8793), .C2(n8792), .A(n9199), .B(n8791), .ZN(n8795)
         );
  MUX2_X1 U10246 ( .A(n8885), .B(n9182), .S(n8826), .Z(n8794) );
  OR2_X1 U10247 ( .A1(n9328), .A2(n9116), .ZN(n8898) );
  INV_X1 U10248 ( .A(n8898), .ZN(n8805) );
  NAND2_X1 U10249 ( .A1(n8952), .A2(n8831), .ZN(n8799) );
  INV_X1 U10250 ( .A(n9126), .ZN(n8798) );
  NOR2_X1 U10251 ( .A1(n8877), .A2(n8798), .ZN(n8800) );
  AOI211_X1 U10252 ( .C1(n8877), .C2(n9125), .A(n8799), .B(n8800), .ZN(n8803)
         );
  INV_X1 U10253 ( .A(n8800), .ZN(n8801) );
  AOI21_X1 U10254 ( .B1(n8801), .B2(n8952), .A(n8831), .ZN(n8802) );
  NOR2_X1 U10255 ( .A1(n8805), .A2(n8831), .ZN(n8804) );
  NAND2_X1 U10256 ( .A1(n9328), .A2(n9116), .ZN(n9128) );
  NAND2_X1 U10257 ( .A1(n9335), .A2(n9325), .ZN(n9127) );
  NAND2_X1 U10258 ( .A1(n9128), .A2(n9127), .ZN(n8889) );
  NAND2_X1 U10259 ( .A1(n7619), .A2(n4905), .ZN(n8808) );
  OR2_X1 U10260 ( .A1(n8823), .A2(n8806), .ZN(n8807) );
  NAND2_X1 U10261 ( .A1(n9322), .A2(n8809), .ZN(n8871) );
  MUX2_X1 U10262 ( .A(n8899), .B(n8871), .S(n8826), .Z(n8811) );
  NAND2_X1 U10263 ( .A1(n8813), .A2(n4905), .ZN(n8816) );
  OR2_X1 U10264 ( .A1(n8823), .A2(n8814), .ZN(n8815) );
  INV_X1 U10265 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U10266 ( .A1(n5461), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U10267 ( .A1(n5657), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8817) );
  OAI211_X1 U10268 ( .C1(n8820), .C2(n8819), .A(n8818), .B(n8817), .ZN(n9130)
         );
  NAND2_X1 U10269 ( .A1(n8821), .A2(n4905), .ZN(n8825) );
  OR2_X1 U10270 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  OR2_X1 U10271 ( .A1(n8829), .A2(n9092), .ZN(n8973) );
  INV_X1 U10272 ( .A(n8832), .ZN(n8834) );
  NAND2_X1 U10273 ( .A1(n8829), .A2(n9092), .ZN(n8903) );
  INV_X1 U10274 ( .A(n9130), .ZN(n8868) );
  OR2_X1 U10275 ( .A1(n9098), .A2(n8868), .ZN(n8830) );
  NAND2_X1 U10276 ( .A1(n8903), .A2(n8830), .ZN(n8960) );
  AOI22_X1 U10277 ( .A1(n8832), .A2(n8903), .B1(n8831), .B2(n8960), .ZN(n8833)
         );
  AOI21_X1 U10278 ( .B1(n8968), .B2(n5737), .A(n8835), .ZN(n8980) );
  INV_X1 U10279 ( .A(n8973), .ZN(n8905) );
  NAND2_X1 U10280 ( .A1(n8952), .A2(n9127), .ZN(n9114) );
  NAND2_X1 U10281 ( .A1(n8873), .A2(n9126), .ZN(n9166) );
  XNOR2_X1 U10282 ( .A(n9377), .B(n9276), .ZN(n9261) );
  NAND2_X1 U10283 ( .A1(n8838), .A2(n8948), .ZN(n9267) );
  NOR2_X1 U10284 ( .A1(n8840), .A2(n8918), .ZN(n8842) );
  AND4_X1 U10285 ( .A1(n9556), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n8849)
         );
  NOR2_X1 U10286 ( .A1(n8845), .A2(n8844), .ZN(n8848) );
  NAND4_X1 U10287 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), .ZN(n8853)
         );
  NOR4_X1 U10288 ( .A1(n8853), .A2(n8852), .A3(n8851), .A4(n8850), .ZN(n8856)
         );
  NAND3_X1 U10289 ( .A1(n8856), .A2(n8855), .A3(n4886), .ZN(n8858) );
  NOR2_X1 U10290 ( .A1(n8858), .A2(n8857), .ZN(n8860) );
  AND4_X1 U10291 ( .A1(n8895), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(n8862)
         );
  NAND3_X1 U10292 ( .A1(n4548), .A2(n9482), .A3(n8862), .ZN(n8863) );
  NOR2_X1 U10293 ( .A1(n9261), .A2(n8863), .ZN(n8864) );
  XNOR2_X1 U10294 ( .A(n9371), .B(n9232), .ZN(n9240) );
  INV_X1 U10295 ( .A(n9240), .ZN(n9244) );
  AND4_X1 U10296 ( .A1(n9217), .A2(n9225), .A3(n8864), .A4(n9244), .ZN(n8865)
         );
  NAND3_X1 U10297 ( .A1(n9188), .A2(n9199), .A3(n8865), .ZN(n8866) );
  NOR2_X1 U10298 ( .A1(n9166), .A2(n8866), .ZN(n8867) );
  NAND4_X1 U10299 ( .A1(n9118), .A2(n4843), .A3(n9159), .A4(n8867), .ZN(n8870)
         );
  NAND2_X1 U10300 ( .A1(n9098), .A2(n8868), .ZN(n8872) );
  INV_X1 U10301 ( .A(n8872), .ZN(n8869) );
  INV_X1 U10302 ( .A(n8970), .ZN(n8913) );
  NAND4_X1 U10303 ( .A1(n8908), .A2(n9493), .A3(n8913), .A4(n6957), .ZN(n8979)
         );
  NAND2_X1 U10304 ( .A1(n8872), .A2(n8871), .ZN(n8958) );
  INV_X1 U10305 ( .A(n8873), .ZN(n8888) );
  INV_X1 U10306 ( .A(n8874), .ZN(n8876) );
  INV_X1 U10307 ( .A(n8875), .ZN(n9124) );
  OAI21_X1 U10308 ( .B1(n8876), .B2(n9124), .A(n9182), .ZN(n8879) );
  INV_X1 U10309 ( .A(n8877), .ZN(n8878) );
  AOI21_X1 U10310 ( .B1(n8885), .B2(n8879), .A(n8878), .ZN(n8954) );
  INV_X1 U10311 ( .A(n8880), .ZN(n8884) );
  INV_X1 U10312 ( .A(n8881), .ZN(n8882) );
  NAND2_X1 U10313 ( .A1(n8882), .A2(n8897), .ZN(n8883) );
  NAND3_X1 U10314 ( .A1(n8885), .A2(n8884), .A3(n8883), .ZN(n8886) );
  NAND2_X1 U10315 ( .A1(n8954), .A2(n8886), .ZN(n8887) );
  OAI211_X1 U10316 ( .C1(n8888), .C2(n9125), .A(n8887), .B(n9126), .ZN(n8890)
         );
  AOI21_X1 U10317 ( .B1(n8890), .B2(n8952), .A(n8889), .ZN(n8957) );
  INV_X1 U10318 ( .A(n8893), .ZN(n8894) );
  AOI21_X1 U10319 ( .B1(n9297), .B2(n8895), .A(n8894), .ZN(n9481) );
  NAND2_X1 U10320 ( .A1(n9481), .A2(n9482), .ZN(n9271) );
  NAND4_X1 U10321 ( .A1(n9121), .A2(n8954), .A3(n8897), .A4(n8952), .ZN(n8900)
         );
  NAND2_X1 U10322 ( .A1(n8899), .A2(n8898), .ZN(n8955) );
  AOI21_X1 U10323 ( .B1(n8957), .B2(n8900), .A(n8955), .ZN(n8901) );
  AOI211_X1 U10324 ( .C1(n9092), .C2(n9098), .A(n8958), .B(n8901), .ZN(n8902)
         );
  AOI21_X1 U10325 ( .B1(n4504), .B2(n9316), .A(n8902), .ZN(n8906) );
  OAI211_X1 U10326 ( .C1(n8906), .C2(n8905), .A(n8904), .B(n8903), .ZN(n8909)
         );
  NAND2_X1 U10327 ( .A1(n6957), .A2(n8972), .ZN(n8907) );
  AOI211_X1 U10328 ( .C1(n8909), .C2(n8908), .A(n8970), .B(n8907), .ZN(n8967)
         );
  INV_X1 U10329 ( .A(P1_B_REG_SCAN_IN), .ZN(n8911) );
  NOR4_X1 U10330 ( .A1(n9656), .A2(n9307), .A3(n8992), .A4(n5738), .ZN(n8910)
         );
  AOI211_X1 U10331 ( .C1(n8913), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8966)
         );
  INV_X1 U10332 ( .A(n8914), .ZN(n8953) );
  INV_X1 U10333 ( .A(n8915), .ZN(n8947) );
  INV_X1 U10334 ( .A(n8916), .ZN(n8917) );
  OAI211_X1 U10335 ( .C1(n8920), .C2(n8919), .A(n8918), .B(n8917), .ZN(n8927)
         );
  NAND2_X1 U10336 ( .A1(n9579), .A2(n9586), .ZN(n8921) );
  NAND4_X1 U10337 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n8926)
         );
  OAI21_X1 U10338 ( .B1(n8927), .B2(n8926), .A(n8925), .ZN(n8930) );
  OAI211_X1 U10339 ( .C1(n8931), .C2(n8930), .A(n8929), .B(n8928), .ZN(n8935)
         );
  INV_X1 U10340 ( .A(n8932), .ZN(n8934) );
  AOI21_X1 U10341 ( .B1(n8935), .B2(n8934), .A(n8933), .ZN(n8941) );
  NAND2_X1 U10342 ( .A1(n8937), .A2(n8936), .ZN(n8940) );
  OAI211_X1 U10343 ( .C1(n8941), .C2(n8940), .A(n8939), .B(n8938), .ZN(n8944)
         );
  AOI22_X1 U10344 ( .A1(n8944), .A2(n8943), .B1(n8942), .B2(n4490), .ZN(n8946)
         );
  AOI21_X1 U10345 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8950) );
  OAI21_X1 U10346 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8951) );
  NAND4_X1 U10347 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(n8956)
         );
  AOI21_X1 U10348 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(n8959) );
  NOR2_X1 U10349 ( .A1(n8959), .A2(n8958), .ZN(n8961) );
  OAI21_X1 U10350 ( .B1(n8961), .B2(n8960), .A(n8973), .ZN(n8963) );
  INV_X1 U10351 ( .A(n8963), .ZN(n8962) );
  NOR3_X1 U10352 ( .A1(n8962), .A2(n5738), .A3(n8970), .ZN(n8965) );
  NOR4_X1 U10353 ( .A1(n8963), .A2(n6957), .A3(n8970), .A4(n8972), .ZN(n8964)
         );
  NOR4_X1 U10354 ( .A1(n8967), .A2(n8966), .A3(n8965), .A4(n8964), .ZN(n8978)
         );
  INV_X1 U10355 ( .A(n8968), .ZN(n8976) );
  NOR3_X1 U10356 ( .A1(n8970), .A2(n5737), .A3(n8969), .ZN(n8971) );
  INV_X1 U10357 ( .A(n8974), .ZN(n8975) );
  OAI211_X1 U10358 ( .C1(n8980), .C2(n8979), .A(n8978), .B(n8977), .ZN(
        P1_U3242) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9130), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9149), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9117), .S(P1_U3973), .Z(
        P1_U3582) );
  INV_X1 U10362 ( .A(n9325), .ZN(n9175) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9175), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9185), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9201), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9345), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9226), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9242), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9363), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9370), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9484), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9299), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9483), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9298), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8981), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8982), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8983), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8984), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8985), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8986), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8987), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9627), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8988), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9536), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8989), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9595), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9586), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8990), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9569), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8991), .S(P1_U3973), .Z(
        P1_U3554) );
  MUX2_X1 U10391 ( .A(n8994), .B(n8993), .S(n8992), .Z(n8997) );
  NAND2_X1 U10392 ( .A1(n8995), .A2(n4710), .ZN(n8996) );
  OAI211_X1 U10393 ( .C1(n8997), .C2(n5160), .A(P1_U3973), .B(n8996), .ZN(
        n9040) );
  INV_X1 U10394 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8999) );
  OAI22_X1 U10395 ( .A1(n9026), .A2(n8999), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8998), .ZN(n9000) );
  AOI21_X1 U10396 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9010) );
  OAI211_X1 U10397 ( .C1(n9004), .C2(n9003), .A(n9084), .B(n9018), .ZN(n9009)
         );
  OAI211_X1 U10398 ( .C1(n9007), .C2(n9006), .A(n9075), .B(n9005), .ZN(n9008)
         );
  NAND4_X1 U10399 ( .A1(n9040), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(
        P1_U3245) );
  NOR2_X1 U10400 ( .A1(n9070), .A2(n9016), .ZN(n9011) );
  AOI211_X1 U10401 ( .C1(n9073), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9012), .B(
        n9011), .ZN(n9023) );
  OAI211_X1 U10402 ( .C1(n9015), .C2(n9014), .A(n9075), .B(n9013), .ZN(n9022)
         );
  MUX2_X1 U10403 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6552), .S(n9016), .Z(n9019)
         );
  NAND3_X1 U10404 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(n9020) );
  NAND3_X1 U10405 ( .A1(n9084), .A2(n9035), .A3(n9020), .ZN(n9021) );
  NAND3_X1 U10406 ( .A1(n9023), .A2(n9022), .A3(n9021), .ZN(P1_U3246) );
  NOR2_X1 U10407 ( .A1(n9070), .A2(n9032), .ZN(n9028) );
  INV_X1 U10408 ( .A(n9024), .ZN(n9025) );
  OAI21_X1 U10409 ( .B1(n9026), .B2(n10145), .A(n9025), .ZN(n9027) );
  NOR2_X1 U10410 ( .A1(n9028), .A2(n9027), .ZN(n9039) );
  OAI211_X1 U10411 ( .C1(n9031), .C2(n9030), .A(n9075), .B(n9029), .ZN(n9038)
         );
  MUX2_X1 U10412 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6555), .S(n9032), .Z(n9033)
         );
  NAND3_X1 U10413 ( .A1(n9035), .A2(n9034), .A3(n9033), .ZN(n9036) );
  NAND3_X1 U10414 ( .A1(n9084), .A2(n9050), .A3(n9036), .ZN(n9037) );
  NAND4_X1 U10415 ( .A1(n9040), .A2(n9039), .A3(n9038), .A4(n9037), .ZN(
        P1_U3247) );
  NOR2_X1 U10416 ( .A1(n9070), .A2(n9041), .ZN(n9042) );
  AOI211_X1 U10417 ( .C1(n9073), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9043), .B(
        n9042), .ZN(n9054) );
  OAI211_X1 U10418 ( .C1(n9046), .C2(n9045), .A(n9075), .B(n9044), .ZN(n9053)
         );
  INV_X1 U10419 ( .A(n9047), .ZN(n9064) );
  NAND3_X1 U10420 ( .A1(n9050), .A2(n9049), .A3(n9048), .ZN(n9051) );
  NAND3_X1 U10421 ( .A1(n9084), .A2(n9064), .A3(n9051), .ZN(n9052) );
  NAND3_X1 U10422 ( .A1(n9054), .A2(n9053), .A3(n9052), .ZN(P1_U3248) );
  NOR2_X1 U10423 ( .A1(n9070), .A2(n9061), .ZN(n9055) );
  AOI211_X1 U10424 ( .C1(n9073), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9056), .B(
        n9055), .ZN(n9068) );
  OAI211_X1 U10425 ( .C1(n9059), .C2(n9058), .A(n9075), .B(n9057), .ZN(n9067)
         );
  INV_X1 U10426 ( .A(n9060), .ZN(n9063) );
  MUX2_X1 U10427 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6559), .S(n9061), .Z(n9062)
         );
  NAND3_X1 U10428 ( .A1(n9064), .A2(n9063), .A3(n9062), .ZN(n9065) );
  NAND3_X1 U10429 ( .A1(n9084), .A2(n9081), .A3(n9065), .ZN(n9066) );
  NAND3_X1 U10430 ( .A1(n9068), .A2(n9067), .A3(n9066), .ZN(P1_U3249) );
  NOR2_X1 U10431 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  AOI211_X1 U10432 ( .C1(n9073), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n9072), .B(
        n9071), .ZN(n9087) );
  OAI211_X1 U10433 ( .C1(n9077), .C2(n9076), .A(n9075), .B(n9074), .ZN(n9086)
         );
  INV_X1 U10434 ( .A(n9078), .ZN(n9083) );
  NAND3_X1 U10435 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n9082) );
  NAND3_X1 U10436 ( .A1(n9084), .A2(n9083), .A3(n9082), .ZN(n9085) );
  NAND3_X1 U10437 ( .A1(n9087), .A2(n9086), .A3(n9085), .ZN(P1_U3250) );
  INV_X1 U10438 ( .A(n9322), .ZN(n9137) );
  NAND2_X1 U10439 ( .A1(n9204), .A2(n9193), .ZN(n9192) );
  NAND2_X1 U10440 ( .A1(n9316), .A2(n9132), .ZN(n9095) );
  XNOR2_X1 U10441 ( .A(n9306), .B(n9095), .ZN(n9088) );
  NAND2_X1 U10442 ( .A1(n9088), .A2(n9546), .ZN(n9305) );
  NAND2_X1 U10443 ( .A1(n9089), .A2(P1_B_REG_SCAN_IN), .ZN(n9090) );
  AND2_X1 U10444 ( .A1(n9535), .A2(n9090), .ZN(n9129) );
  INV_X1 U10445 ( .A(n9129), .ZN(n9091) );
  OR2_X1 U10446 ( .A1(n9092), .A2(n9091), .ZN(n9314) );
  NOR2_X1 U10447 ( .A1(n9553), .A2(n9314), .ZN(n9097) );
  NOR2_X1 U10448 ( .A1(n9306), .A2(n9544), .ZN(n9093) );
  AOI211_X1 U10449 ( .C1(n9301), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9097), .B(
        n9093), .ZN(n9094) );
  OAI21_X1 U10450 ( .B1(n9295), .B2(n9305), .A(n9094), .ZN(P1_U3263) );
  OAI211_X1 U10451 ( .C1(n9316), .C2(n9132), .A(n9546), .B(n9095), .ZN(n9315)
         );
  AND2_X1 U10452 ( .A1(n9553), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9096) );
  NOR2_X1 U10453 ( .A1(n9097), .A2(n9096), .ZN(n9100) );
  NAND2_X1 U10454 ( .A1(n9098), .A2(n9291), .ZN(n9099) );
  OAI211_X1 U10455 ( .C1(n9315), .C2(n9295), .A(n9100), .B(n9099), .ZN(
        P1_U3264) );
  NOR2_X1 U10456 ( .A1(n9292), .A2(n9483), .ZN(n9103) );
  NAND2_X1 U10457 ( .A1(n9268), .A2(n9104), .ZN(n9106) );
  NOR2_X1 U10458 ( .A1(n9346), .A2(n9201), .ZN(n9111) );
  NAND2_X1 U10459 ( .A1(n9346), .A2(n9201), .ZN(n9112) );
  NAND2_X1 U10460 ( .A1(n9113), .A2(n9112), .ZN(n9165) );
  XNOR2_X1 U10461 ( .A(n9119), .B(n9118), .ZN(n9319) );
  INV_X1 U10462 ( .A(n9319), .ZN(n9140) );
  NAND2_X1 U10463 ( .A1(n9223), .A2(n9123), .ZN(n9218) );
  AOI21_X1 U10464 ( .B1(n9218), .B2(n9217), .A(n9124), .ZN(n9200) );
  NAND2_X1 U10465 ( .A1(n9200), .A2(n9199), .ZN(n9181) );
  NAND3_X1 U10466 ( .A1(n9181), .A2(n9188), .A3(n9182), .ZN(n9183) );
  NAND2_X1 U10467 ( .A1(n9183), .A2(n9125), .ZN(n9173) );
  INV_X1 U10468 ( .A(n9166), .ZN(n9174) );
  AOI22_X1 U10469 ( .A1(n9117), .A2(n9626), .B1(n9130), .B2(n9129), .ZN(n9131)
         );
  INV_X1 U10470 ( .A(n9142), .ZN(n9133) );
  AOI211_X1 U10471 ( .C1(n9322), .C2(n9133), .A(n9487), .B(n9132), .ZN(n9321)
         );
  NAND2_X1 U10472 ( .A1(n9321), .A2(n9549), .ZN(n9136) );
  AOI22_X1 U10473 ( .A1(n9553), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9134), .B2(
        n9541), .ZN(n9135) );
  OAI211_X1 U10474 ( .C1(n9137), .C2(n9544), .A(n9136), .B(n9135), .ZN(n9138)
         );
  AOI21_X1 U10475 ( .B1(n9320), .B2(n9494), .A(n9138), .ZN(n9139) );
  OAI21_X1 U10476 ( .B1(n9140), .B2(n9286), .A(n9139), .ZN(P1_U3356) );
  INV_X1 U10477 ( .A(n9155), .ZN(n9143) );
  AOI211_X1 U10478 ( .C1(n9328), .C2(n9143), .A(n9487), .B(n9142), .ZN(n9326)
         );
  NAND2_X1 U10479 ( .A1(n9328), .A2(n9291), .ZN(n9146) );
  AOI22_X1 U10480 ( .A1(n9301), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9144), .B2(
        n9541), .ZN(n9145) );
  OAI211_X1 U10481 ( .C1(n9325), .C2(n9248), .A(n9146), .B(n9145), .ZN(n9152)
         );
  XNOR2_X1 U10482 ( .A(n9148), .B(n9147), .ZN(n9150) );
  AOI22_X1 U10483 ( .A1(n9150), .A2(n9486), .B1(n9535), .B2(n9149), .ZN(n9330)
         );
  NOR2_X1 U10484 ( .A1(n9330), .A2(n9301), .ZN(n9151) );
  AOI211_X1 U10485 ( .C1(n9326), .C2(n9549), .A(n9152), .B(n9151), .ZN(n9153)
         );
  OAI21_X1 U10486 ( .B1(n9331), .B2(n9286), .A(n9153), .ZN(P1_U3265) );
  XNOR2_X1 U10487 ( .A(n9154), .B(n9159), .ZN(n9338) );
  AOI211_X1 U10488 ( .C1(n9335), .C2(n9167), .A(n9487), .B(n9155), .ZN(n9333)
         );
  NAND2_X1 U10489 ( .A1(n9335), .A2(n9291), .ZN(n9158) );
  AOI22_X1 U10490 ( .A1(n9301), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9156), .B2(
        n9541), .ZN(n9157) );
  OAI211_X1 U10491 ( .C1(n9332), .C2(n9248), .A(n9158), .B(n9157), .ZN(n9163)
         );
  XNOR2_X1 U10492 ( .A(n9160), .B(n9159), .ZN(n9161) );
  AOI22_X1 U10493 ( .A1(n9161), .A2(n9486), .B1(n9535), .B2(n9117), .ZN(n9337)
         );
  NOR2_X1 U10494 ( .A1(n9337), .A2(n9553), .ZN(n9162) );
  AOI211_X1 U10495 ( .C1(n9549), .C2(n9333), .A(n9163), .B(n9162), .ZN(n9164)
         );
  OAI21_X1 U10496 ( .B1(n9338), .B2(n9286), .A(n9164), .ZN(P1_U3266) );
  XNOR2_X1 U10497 ( .A(n9165), .B(n9166), .ZN(n9343) );
  INV_X1 U10498 ( .A(n9167), .ZN(n9168) );
  AOI21_X1 U10499 ( .B1(n9339), .B2(n9192), .A(n9168), .ZN(n9340) );
  AOI22_X1 U10500 ( .A1(n9553), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9169), .B2(
        n9541), .ZN(n9170) );
  OAI21_X1 U10501 ( .B1(n9171), .B2(n9544), .A(n9170), .ZN(n9178) );
  OAI21_X1 U10502 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9176) );
  AOI222_X1 U10503 ( .A1(n9486), .A2(n9176), .B1(n9201), .B2(n9626), .C1(n9175), .C2(n9535), .ZN(n9342) );
  NOR2_X1 U10504 ( .A1(n9342), .A2(n9553), .ZN(n9177) );
  AOI211_X1 U10505 ( .C1(n9340), .C2(n9179), .A(n9178), .B(n9177), .ZN(n9180)
         );
  OAI21_X1 U10506 ( .B1(n9286), .B2(n9343), .A(n9180), .ZN(P1_U3267) );
  AND2_X1 U10507 ( .A1(n9181), .A2(n9182), .ZN(n9184) );
  OAI21_X1 U10508 ( .B1(n9184), .B2(n9188), .A(n9183), .ZN(n9186) );
  AOI22_X1 U10509 ( .A1(n9186), .A2(n9486), .B1(n9535), .B2(n9185), .ZN(n9349)
         );
  XOR2_X1 U10510 ( .A(n9188), .B(n9187), .Z(n9344) );
  NAND2_X1 U10511 ( .A1(n9344), .A2(n9480), .ZN(n9197) );
  AOI22_X1 U10512 ( .A1(n9301), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9189), .B2(
        n9541), .ZN(n9190) );
  OAI21_X1 U10513 ( .B1(n9248), .B2(n9191), .A(n9190), .ZN(n9195) );
  OAI211_X1 U10514 ( .C1(n9204), .C2(n9193), .A(n9546), .B(n9192), .ZN(n9347)
         );
  NOR2_X1 U10515 ( .A1(n9347), .A2(n9295), .ZN(n9194) );
  AOI211_X1 U10516 ( .C1(n9291), .C2(n9346), .A(n9195), .B(n9194), .ZN(n9196)
         );
  OAI211_X1 U10517 ( .C1(n9553), .C2(n9349), .A(n9197), .B(n9196), .ZN(
        P1_U3268) );
  XOR2_X1 U10518 ( .A(n9199), .B(n9198), .Z(n9355) );
  OAI211_X1 U10519 ( .C1(n9200), .C2(n9199), .A(n9181), .B(n9486), .ZN(n9203)
         );
  AOI22_X1 U10520 ( .A1(n9535), .A2(n9201), .B1(n9226), .B2(n9626), .ZN(n9202)
         );
  NAND2_X1 U10521 ( .A1(n9203), .A2(n9202), .ZN(n9351) );
  AOI211_X1 U10522 ( .C1(n9353), .C2(n4673), .A(n9487), .B(n9204), .ZN(n9352)
         );
  NAND2_X1 U10523 ( .A1(n9352), .A2(n9549), .ZN(n9207) );
  AOI22_X1 U10524 ( .A1(n9301), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9205), .B2(
        n9541), .ZN(n9206) );
  OAI211_X1 U10525 ( .C1(n9208), .C2(n9544), .A(n9207), .B(n9206), .ZN(n9209)
         );
  AOI21_X1 U10526 ( .B1(n9351), .B2(n9494), .A(n9209), .ZN(n9210) );
  OAI21_X1 U10527 ( .B1(n9355), .B2(n9286), .A(n9210), .ZN(P1_U3269) );
  XNOR2_X1 U10528 ( .A(n9211), .B(n9217), .ZN(n9361) );
  AOI211_X1 U10529 ( .C1(n9213), .C2(n9233), .A(n9487), .B(n9212), .ZN(n9358)
         );
  NAND2_X1 U10530 ( .A1(n9213), .A2(n9291), .ZN(n9216) );
  AOI22_X1 U10531 ( .A1(n9301), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9214), .B2(
        n9541), .ZN(n9215) );
  OAI211_X1 U10532 ( .C1(n9356), .C2(n9248), .A(n9216), .B(n9215), .ZN(n9221)
         );
  XNOR2_X1 U10533 ( .A(n9218), .B(n9217), .ZN(n9219) );
  AOI22_X1 U10534 ( .A1(n9219), .A2(n9486), .B1(n9535), .B2(n9345), .ZN(n9360)
         );
  NOR2_X1 U10535 ( .A1(n9360), .A2(n9553), .ZN(n9220) );
  AOI211_X1 U10536 ( .C1(n9358), .C2(n9549), .A(n9221), .B(n9220), .ZN(n9222)
         );
  OAI21_X1 U10537 ( .B1(n9361), .B2(n9286), .A(n9222), .ZN(P1_U3270) );
  OAI21_X1 U10538 ( .B1(n9225), .B2(n9224), .A(n9223), .ZN(n9227) );
  AOI22_X1 U10539 ( .A1(n9227), .A2(n9486), .B1(n9535), .B2(n9226), .ZN(n9367)
         );
  XNOR2_X1 U10540 ( .A(n4829), .B(n9229), .ZN(n9362) );
  NAND2_X1 U10541 ( .A1(n9362), .A2(n9480), .ZN(n9239) );
  AOI22_X1 U10542 ( .A1(n9301), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9230), .B2(
        n9541), .ZN(n9231) );
  OAI21_X1 U10543 ( .B1(n9248), .B2(n9232), .A(n9231), .ZN(n9237) );
  INV_X1 U10544 ( .A(n9249), .ZN(n9234) );
  OAI211_X1 U10545 ( .C1(n9235), .C2(n9234), .A(n9233), .B(n9546), .ZN(n9365)
         );
  NOR2_X1 U10546 ( .A1(n9365), .A2(n9295), .ZN(n9236) );
  AOI211_X1 U10547 ( .C1(n9291), .C2(n9364), .A(n9237), .B(n9236), .ZN(n9238)
         );
  OAI211_X1 U10548 ( .C1(n9301), .C2(n9367), .A(n9239), .B(n9238), .ZN(
        P1_U3271) );
  XNOR2_X1 U10549 ( .A(n9241), .B(n9240), .ZN(n9243) );
  AOI22_X1 U10550 ( .A1(n9243), .A2(n9486), .B1(n9535), .B2(n9242), .ZN(n9374)
         );
  XNOR2_X1 U10551 ( .A(n9245), .B(n9244), .ZN(n9369) );
  NAND2_X1 U10552 ( .A1(n9369), .A2(n9480), .ZN(n9254) );
  AOI22_X1 U10553 ( .A1(n9301), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9246), .B2(
        n9541), .ZN(n9247) );
  OAI21_X1 U10554 ( .B1(n9248), .B2(n9276), .A(n9247), .ZN(n9252) );
  OAI211_X1 U10555 ( .C1(n9256), .C2(n9250), .A(n9546), .B(n9249), .ZN(n9372)
         );
  NOR2_X1 U10556 ( .A1(n9372), .A2(n9295), .ZN(n9251) );
  AOI211_X1 U10557 ( .C1(n9291), .C2(n9371), .A(n9252), .B(n9251), .ZN(n9253)
         );
  OAI211_X1 U10558 ( .C1(n9553), .C2(n9374), .A(n9254), .B(n9253), .ZN(
        P1_U3272) );
  XNOR2_X1 U10559 ( .A(n9255), .B(n9261), .ZN(n9380) );
  INV_X1 U10560 ( .A(n9279), .ZN(n9257) );
  AOI211_X1 U10561 ( .C1(n9377), .C2(n9257), .A(n9487), .B(n9256), .ZN(n9376)
         );
  AOI22_X1 U10562 ( .A1(n9301), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9258), .B2(
        n9541), .ZN(n9259) );
  OAI21_X1 U10563 ( .B1(n9260), .B2(n9544), .A(n9259), .ZN(n9265) );
  XNOR2_X1 U10564 ( .A(n9262), .B(n9261), .ZN(n9263) );
  AOI222_X1 U10565 ( .A1(n9486), .A2(n9263), .B1(n9363), .B2(n9535), .C1(n9484), .C2(n9626), .ZN(n9379) );
  NOR2_X1 U10566 ( .A1(n9379), .A2(n9301), .ZN(n9264) );
  AOI211_X1 U10567 ( .C1(n9376), .C2(n9549), .A(n9265), .B(n9264), .ZN(n9266)
         );
  OAI21_X1 U10568 ( .B1(n9380), .B2(n9286), .A(n9266), .ZN(P1_U3273) );
  XNOR2_X1 U10569 ( .A(n9268), .B(n9267), .ZN(n9386) );
  INV_X1 U10570 ( .A(n9269), .ZN(n9270) );
  NOR2_X1 U10571 ( .A1(n4548), .A2(n9270), .ZN(n9273) );
  AOI21_X1 U10572 ( .B1(n9273), .B2(n9271), .A(n9272), .ZN(n9274) );
  OAI222_X1 U10573 ( .A1(n9277), .A2(n9276), .B1(n9656), .B2(n9275), .C1(n9557), .C2(n9274), .ZN(n9382) );
  INV_X1 U10574 ( .A(n9278), .ZN(n9491) );
  AOI211_X1 U10575 ( .C1(n9384), .C2(n9491), .A(n9487), .B(n9279), .ZN(n9383)
         );
  NAND2_X1 U10576 ( .A1(n9383), .A2(n9549), .ZN(n9282) );
  AOI22_X1 U10577 ( .A1(n9553), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9280), .B2(
        n9541), .ZN(n9281) );
  OAI211_X1 U10578 ( .C1(n9283), .C2(n9544), .A(n9282), .B(n9281), .ZN(n9284)
         );
  AOI21_X1 U10579 ( .B1(n9382), .B2(n9494), .A(n9284), .ZN(n9285) );
  OAI21_X1 U10580 ( .B1(n9386), .B2(n9286), .A(n9285), .ZN(P1_U3274) );
  XNOR2_X1 U10581 ( .A(n9287), .B(n9296), .ZN(n9511) );
  AOI21_X1 U10582 ( .B1(n9288), .B2(n9292), .A(n9487), .ZN(n9289) );
  NAND2_X1 U10583 ( .A1(n9289), .A2(n9489), .ZN(n9507) );
  AOI22_X1 U10584 ( .A1(n9301), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9290), .B2(
        n9541), .ZN(n9294) );
  NAND2_X1 U10585 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  OAI211_X1 U10586 ( .C1(n9507), .C2(n9295), .A(n9294), .B(n9293), .ZN(n9303)
         );
  XNOR2_X1 U10587 ( .A(n9297), .B(n9296), .ZN(n9300) );
  AOI222_X1 U10588 ( .A1(n9486), .A2(n9300), .B1(n9299), .B2(n9535), .C1(n9298), .C2(n9626), .ZN(n9508) );
  NOR2_X1 U10589 ( .A1(n9508), .A2(n9301), .ZN(n9302) );
  AOI211_X1 U10590 ( .C1(n9511), .C2(n9480), .A(n9303), .B(n9302), .ZN(n9304)
         );
  INV_X1 U10591 ( .A(n9304), .ZN(P1_U3276) );
  OAI211_X1 U10592 ( .C1(n9306), .C2(n9665), .A(n9305), .B(n9314), .ZN(n9389)
         );
  NOR2_X1 U10593 ( .A1(n9308), .A2(n9307), .ZN(n9312) );
  NAND4_X1 U10594 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n9388)
         );
  MUX2_X1 U10595 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9389), .S(n9381), .Z(
        P1_U3553) );
  OAI211_X1 U10596 ( .C1(n9316), .C2(n9665), .A(n9315), .B(n9314), .ZN(n9390)
         );
  MUX2_X1 U10597 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9390), .S(n9381), .Z(
        P1_U3552) );
  INV_X1 U10598 ( .A(n9668), .ZN(n9317) );
  NAND2_X1 U10599 ( .A1(n9319), .A2(n9652), .ZN(n9324) );
  NAND2_X1 U10600 ( .A1(n9324), .A2(n9323), .ZN(n9391) );
  MUX2_X1 U10601 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9391), .S(n9381), .Z(
        P1_U3551) );
  NOR2_X1 U10602 ( .A1(n9325), .A2(n9656), .ZN(n9327) );
  AOI211_X1 U10603 ( .C1(n9625), .C2(n9328), .A(n9327), .B(n9326), .ZN(n9329)
         );
  OAI211_X1 U10604 ( .C1(n9331), .C2(n9654), .A(n9330), .B(n9329), .ZN(n9392)
         );
  MUX2_X1 U10605 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9392), .S(n9381), .Z(
        P1_U3550) );
  NOR2_X1 U10606 ( .A1(n9332), .A2(n9656), .ZN(n9334) );
  AOI211_X1 U10607 ( .C1(n9625), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9336)
         );
  OAI211_X1 U10608 ( .C1(n9338), .C2(n9654), .A(n9337), .B(n9336), .ZN(n9393)
         );
  MUX2_X1 U10609 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9393), .S(n9381), .Z(
        P1_U3549) );
  AOI22_X1 U10610 ( .A1(n9340), .A2(n9546), .B1(n9625), .B2(n9339), .ZN(n9341)
         );
  OAI211_X1 U10611 ( .C1(n9343), .C2(n9654), .A(n9342), .B(n9341), .ZN(n9394)
         );
  MUX2_X1 U10612 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9394), .S(n9381), .Z(
        P1_U3548) );
  NAND2_X1 U10613 ( .A1(n9344), .A2(n9652), .ZN(n9350) );
  AOI22_X1 U10614 ( .A1(n9346), .A2(n9625), .B1(n9626), .B2(n9345), .ZN(n9348)
         );
  NAND4_X1 U10615 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n9395)
         );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9395), .S(n9381), .Z(
        P1_U3547) );
  AOI211_X1 U10617 ( .C1(n9625), .C2(n9353), .A(n9352), .B(n9351), .ZN(n9354)
         );
  OAI21_X1 U10618 ( .B1(n9355), .B2(n9654), .A(n9354), .ZN(n9396) );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9396), .S(n9381), .Z(
        P1_U3546) );
  OAI22_X1 U10620 ( .A1(n4671), .A2(n9665), .B1(n9356), .B2(n9656), .ZN(n9357)
         );
  NOR2_X1 U10621 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  OAI211_X1 U10622 ( .C1(n9361), .C2(n9654), .A(n9360), .B(n9359), .ZN(n9397)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9397), .S(n9381), .Z(
        P1_U3545) );
  NAND2_X1 U10624 ( .A1(n9362), .A2(n9652), .ZN(n9368) );
  AOI22_X1 U10625 ( .A1(n9364), .A2(n9625), .B1(n9626), .B2(n9363), .ZN(n9366)
         );
  NAND4_X1 U10626 ( .A1(n9368), .A2(n9367), .A3(n9366), .A4(n9365), .ZN(n9398)
         );
  MUX2_X1 U10627 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9398), .S(n9381), .Z(
        P1_U3544) );
  NAND2_X1 U10628 ( .A1(n9369), .A2(n9652), .ZN(n9375) );
  AOI22_X1 U10629 ( .A1(n9371), .A2(n9625), .B1(n9626), .B2(n9370), .ZN(n9373)
         );
  NAND4_X1 U10630 ( .A1(n9375), .A2(n9374), .A3(n9373), .A4(n9372), .ZN(n9399)
         );
  MUX2_X1 U10631 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9399), .S(n9381), .Z(
        P1_U3543) );
  AOI21_X1 U10632 ( .B1(n9625), .B2(n9377), .A(n9376), .ZN(n9378) );
  OAI211_X1 U10633 ( .C1(n9380), .C2(n9654), .A(n9379), .B(n9378), .ZN(n9400)
         );
  MUX2_X1 U10634 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9400), .S(n9381), .Z(
        P1_U3542) );
  AOI211_X1 U10635 ( .C1(n9625), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9385)
         );
  OAI21_X1 U10636 ( .B1(n9654), .B2(n9386), .A(n9385), .ZN(n9401) );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9401), .S(n9700), .Z(
        P1_U3541) );
  MUX2_X1 U10638 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9389), .S(n4404), .Z(
        P1_U3521) );
  MUX2_X1 U10639 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9390), .S(n4404), .Z(
        P1_U3520) );
  MUX2_X1 U10640 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9391), .S(n4404), .Z(
        P1_U3519) );
  MUX2_X1 U10641 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9392), .S(n4404), .Z(
        P1_U3518) );
  MUX2_X1 U10642 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9393), .S(n4404), .Z(
        P1_U3517) );
  MUX2_X1 U10643 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9394), .S(n4404), .Z(
        P1_U3516) );
  MUX2_X1 U10644 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9395), .S(n4404), .Z(
        P1_U3515) );
  MUX2_X1 U10645 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9396), .S(n4404), .Z(
        P1_U3514) );
  MUX2_X1 U10646 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9397), .S(n4404), .Z(
        P1_U3513) );
  MUX2_X1 U10647 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9398), .S(n4404), .Z(
        P1_U3512) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9399), .S(n4404), .Z(
        P1_U3511) );
  MUX2_X1 U10649 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9400), .S(n4404), .Z(
        P1_U3510) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9401), .S(n4404), .Z(
        P1_U3509) );
  MUX2_X1 U10651 ( .A(n9402), .B(P1_D_REG_1__SCAN_IN), .S(n9555), .Z(P1_U3440)
         );
  MUX2_X1 U10652 ( .A(n9403), .B(P1_D_REG_0__SCAN_IN), .S(n9555), .Z(P1_U3439)
         );
  INV_X1 U10653 ( .A(n9404), .ZN(n9407) );
  NOR4_X1 U10654 ( .A1(n9407), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9406), .A4(
        P1_U3086), .ZN(n9408) );
  AOI21_X1 U10655 ( .B1(n9409), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9408), .ZN(
        n9410) );
  OAI21_X1 U10656 ( .B1(n9412), .B2(n9411), .A(n9410), .ZN(P1_U3324) );
  MUX2_X1 U10657 ( .A(n9413), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U10658 ( .A1(n9415), .A2(n9414), .ZN(n9454) );
  NOR2_X1 U10659 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9450) );
  NOR2_X1 U10660 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9448) );
  NOR2_X1 U10661 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9446) );
  NOR2_X1 U10662 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9444) );
  NOR2_X1 U10663 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9442) );
  NOR2_X1 U10664 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9440) );
  NOR2_X1 U10665 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9438) );
  NOR2_X1 U10666 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9434) );
  NOR2_X1 U10667 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9431) );
  NOR2_X1 U10668 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9429) );
  NOR2_X1 U10669 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9427) );
  NOR2_X1 U10670 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9425) );
  NOR2_X1 U10671 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9424) );
  NAND2_X1 U10672 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9422) );
  XOR2_X1 U10673 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10289) );
  NAND2_X1 U10674 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9420) );
  AOI21_X1 U10675 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U10676 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9416) );
  NOR2_X1 U10677 ( .A1(n9417), .A2(n9416), .ZN(n9952) );
  NOR2_X1 U10678 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9952), .ZN(n9418) );
  NOR2_X1 U10679 ( .A1(n9953), .A2(n9418), .ZN(n10287) );
  XNOR2_X1 U10680 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n10185), .ZN(n10286) );
  NAND2_X1 U10681 ( .A1(n10287), .A2(n10286), .ZN(n9419) );
  NAND2_X1 U10682 ( .A1(n9420), .A2(n9419), .ZN(n10288) );
  NAND2_X1 U10683 ( .A1(n10289), .A2(n10288), .ZN(n9421) );
  NAND2_X1 U10684 ( .A1(n9422), .A2(n9421), .ZN(n10291) );
  XOR2_X1 U10685 ( .A(n10145), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10290) );
  NOR2_X1 U10686 ( .A1(n10291), .A2(n10290), .ZN(n9423) );
  NOR2_X1 U10687 ( .A1(n9424), .A2(n9423), .ZN(n10275) );
  XNOR2_X1 U10688 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10274) );
  NOR2_X1 U10689 ( .A1(n10275), .A2(n10274), .ZN(n10273) );
  NOR2_X1 U10690 ( .A1(n9425), .A2(n10273), .ZN(n9975) );
  XNOR2_X1 U10691 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9974) );
  NOR2_X1 U10692 ( .A1(n9975), .A2(n9974), .ZN(n9426) );
  NOR2_X1 U10693 ( .A1(n9427), .A2(n9426), .ZN(n10285) );
  XNOR2_X1 U10694 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10284) );
  NOR2_X1 U10695 ( .A1(n10285), .A2(n10284), .ZN(n9428) );
  NOR2_X1 U10696 ( .A1(n9429), .A2(n9428), .ZN(n10283) );
  XNOR2_X1 U10697 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10282) );
  NOR2_X1 U10698 ( .A1(n10283), .A2(n10282), .ZN(n9430) );
  NOR2_X1 U10699 ( .A1(n9431), .A2(n9430), .ZN(n10281) );
  INV_X1 U10700 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9432) );
  INV_X1 U10701 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9789) );
  AOI22_X1 U10702 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9432), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n9789), .ZN(n10280) );
  NOR2_X1 U10703 ( .A1(n10281), .A2(n10280), .ZN(n9433) );
  NOR2_X1 U10704 ( .A1(n9434), .A2(n9433), .ZN(n9973) );
  AOI22_X1 U10705 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10238), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10103), .ZN(n9972) );
  NOR2_X1 U10706 ( .A1(n9973), .A2(n9972), .ZN(n9435) );
  AOI21_X1 U10707 ( .B1(n10103), .B2(n10238), .A(n9435), .ZN(n9971) );
  INV_X1 U10708 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9436) );
  INV_X1 U10709 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U10710 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9436), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n9805), .ZN(n9970) );
  NOR2_X1 U10711 ( .A1(n9971), .A2(n9970), .ZN(n9437) );
  NOR2_X1 U10712 ( .A1(n9438), .A2(n9437), .ZN(n9969) );
  XNOR2_X1 U10713 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9968) );
  NOR2_X1 U10714 ( .A1(n9969), .A2(n9968), .ZN(n9439) );
  NOR2_X1 U10715 ( .A1(n9440), .A2(n9439), .ZN(n9967) );
  INV_X1 U10716 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10258) );
  XOR2_X1 U10717 ( .A(n10258), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n9966) );
  NOR2_X1 U10718 ( .A1(n9967), .A2(n9966), .ZN(n9441) );
  NOR2_X1 U10719 ( .A1(n9442), .A2(n9441), .ZN(n9965) );
  INV_X1 U10720 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10171) );
  XOR2_X1 U10721 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n10171), .Z(n9964) );
  NOR2_X1 U10722 ( .A1(n9965), .A2(n9964), .ZN(n9443) );
  NOR2_X1 U10723 ( .A1(n9444), .A2(n9443), .ZN(n9963) );
  INV_X1 U10724 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U10725 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n6871), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n9838), .ZN(n9962) );
  NOR2_X1 U10726 ( .A1(n9963), .A2(n9962), .ZN(n9445) );
  NOR2_X1 U10727 ( .A1(n9446), .A2(n9445), .ZN(n9961) );
  XOR2_X1 U10728 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n6977), .Z(n9960) );
  NOR2_X1 U10729 ( .A1(n9961), .A2(n9960), .ZN(n9447) );
  NOR2_X1 U10730 ( .A1(n9448), .A2(n9447), .ZN(n9959) );
  INV_X1 U10731 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10034) );
  INV_X1 U10732 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U10733 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10034), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10254), .ZN(n9958) );
  NOR2_X1 U10734 ( .A1(n9959), .A2(n9958), .ZN(n9449) );
  NOR2_X1 U10735 ( .A1(n9450), .A2(n9449), .ZN(n9956) );
  NAND2_X1 U10736 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9956), .ZN(n9451) );
  NOR2_X1 U10737 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9956), .ZN(n9955) );
  AOI21_X1 U10738 ( .B1(n9452), .B2(n9451), .A(n9955), .ZN(n9453) );
  XOR2_X1 U10739 ( .A(n9454), .B(n9453), .Z(ADD_1068_U4) );
  INV_X1 U10740 ( .A(n9455), .ZN(n9456) );
  NOR2_X1 U10741 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  XNOR2_X1 U10742 ( .A(n8090), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U10743 ( .A(n9458), .B(n9463), .ZN(n9478) );
  OAI21_X1 U10744 ( .B1(n9461), .B2(n9460), .A(n9459), .ZN(n9465) );
  XNOR2_X1 U10745 ( .A(n8090), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9473) );
  MUX2_X1 U10746 ( .A(n9463), .B(n9473), .S(n9462), .Z(n9464) );
  XNOR2_X1 U10747 ( .A(n9465), .B(n9464), .ZN(n9469) );
  INV_X1 U10748 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U10749 ( .A1(n9858), .A2(n8090), .ZN(n9467) );
  OAI211_X1 U10750 ( .C1(n10041), .C2(n9839), .A(n9467), .B(n9466), .ZN(n9468)
         );
  AOI21_X1 U10751 ( .B1(n9868), .B2(n9469), .A(n9468), .ZN(n9477) );
  NAND2_X1 U10752 ( .A1(n9472), .A2(n9471), .ZN(n9474) );
  XNOR2_X1 U10753 ( .A(n9474), .B(n9473), .ZN(n9475) );
  NAND2_X1 U10754 ( .A1(n9475), .A2(n9863), .ZN(n9476) );
  OAI211_X1 U10755 ( .C1(n9478), .C2(n9872), .A(n9477), .B(n9476), .ZN(
        P2_U3201) );
  XNOR2_X1 U10756 ( .A(n9479), .B(n9482), .ZN(n9505) );
  AOI22_X1 U10757 ( .A1(n9505), .A2(n9480), .B1(P1_REG2_REG_18__SCAN_IN), .B2(
        n9553), .ZN(n9498) );
  OAI21_X1 U10758 ( .B1(n9482), .B2(n9481), .A(n9271), .ZN(n9485) );
  AOI222_X1 U10759 ( .A1(n9486), .A2(n9485), .B1(n9484), .B2(n9535), .C1(n9483), .C2(n9626), .ZN(n9502) );
  INV_X1 U10760 ( .A(n9502), .ZN(n9496) );
  AOI21_X1 U10761 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9490) );
  NAND2_X1 U10762 ( .A1(n9491), .A2(n9490), .ZN(n9501) );
  OAI22_X1 U10763 ( .A1(n9501), .A2(n9493), .B1(n9503), .B2(n9492), .ZN(n9495)
         );
  OAI21_X1 U10764 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9497) );
  OAI211_X1 U10765 ( .C1(n9500), .C2(n9499), .A(n9498), .B(n9497), .ZN(
        P1_U3275) );
  OAI211_X1 U10766 ( .C1(n9503), .C2(n9665), .A(n9502), .B(n9501), .ZN(n9504)
         );
  AOI21_X1 U10767 ( .B1(n9505), .B2(n9652), .A(n9504), .ZN(n9526) );
  AOI22_X1 U10768 ( .A1(n9381), .A2(n9526), .B1(n9506), .B2(n9697), .ZN(
        P1_U3540) );
  OAI211_X1 U10769 ( .C1(n9509), .C2(n9665), .A(n9508), .B(n9507), .ZN(n9510)
         );
  AOI21_X1 U10770 ( .B1(n9511), .B2(n9652), .A(n9510), .ZN(n9528) );
  AOI22_X1 U10771 ( .A1(n9381), .A2(n9528), .B1(n10221), .B2(n9697), .ZN(
        P1_U3539) );
  NOR3_X1 U10772 ( .A1(n9513), .A2(n9512), .A3(n9654), .ZN(n9518) );
  OAI22_X1 U10773 ( .A1(n4668), .A2(n9665), .B1(n9514), .B2(n9656), .ZN(n9515)
         );
  NOR4_X1 U10774 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n9529)
         );
  AOI22_X1 U10775 ( .A1(n9381), .A2(n9529), .B1(n9519), .B2(n9697), .ZN(
        P1_U3538) );
  OAI211_X1 U10776 ( .C1(n9522), .C2(n9665), .A(n9521), .B(n9520), .ZN(n9523)
         );
  AOI21_X1 U10777 ( .B1(n9652), .B2(n9524), .A(n9523), .ZN(n9530) );
  INV_X1 U10778 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9525) );
  AOI22_X1 U10779 ( .A1(n9381), .A2(n9530), .B1(n9525), .B2(n9697), .ZN(
        P1_U3537) );
  INV_X1 U10780 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U10781 ( .A1(n4404), .A2(n9526), .B1(n10208), .B2(n9672), .ZN(
        P1_U3507) );
  INV_X1 U10782 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U10783 ( .A1(n4404), .A2(n9528), .B1(n9527), .B2(n9672), .ZN(
        P1_U3504) );
  INV_X1 U10784 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U10785 ( .A1(n4404), .A2(n9529), .B1(n10189), .B2(n9672), .ZN(
        P1_U3501) );
  INV_X1 U10786 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U10787 ( .A1(n4404), .A2(n9530), .B1(n10257), .B2(n9672), .ZN(
        P1_U3498) );
  XNOR2_X1 U10788 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10789 ( .A(n9531), .B(n9532), .ZN(n9616) );
  XNOR2_X1 U10790 ( .A(n9534), .B(n9533), .ZN(n9538) );
  AOI22_X1 U10791 ( .A1(n9626), .A2(n9536), .B1(n9627), .B2(n9535), .ZN(n9537)
         );
  OAI21_X1 U10792 ( .B1(n9538), .B2(n9557), .A(n9537), .ZN(n9539) );
  AOI21_X1 U10793 ( .B1(n9540), .B2(n9616), .A(n9539), .ZN(n9613) );
  AOI22_X1 U10794 ( .A1(n9553), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n9542), .B2(
        n9541), .ZN(n9543) );
  OAI21_X1 U10795 ( .B1(n9544), .B2(n9612), .A(n9543), .ZN(n9545) );
  INV_X1 U10796 ( .A(n9545), .ZN(n9552) );
  OAI211_X1 U10797 ( .C1(n4496), .C2(n9612), .A(n9547), .B(n9546), .ZN(n9611)
         );
  INV_X1 U10798 ( .A(n9611), .ZN(n9548) );
  AOI22_X1 U10799 ( .A1(n9616), .A2(n9550), .B1(n9549), .B2(n9548), .ZN(n9551)
         );
  OAI211_X1 U10800 ( .C1(n9553), .C2(n9613), .A(n9552), .B(n9551), .ZN(
        P1_U3286) );
  INV_X1 U10801 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10205) );
  NOR2_X1 U10802 ( .A1(n9554), .A2(n10205), .ZN(P1_U3294) );
  AND2_X1 U10803 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9555), .ZN(P1_U3295) );
  AND2_X1 U10804 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9555), .ZN(P1_U3296) );
  INV_X1 U10805 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U10806 ( .A1(n9554), .A2(n10049), .ZN(P1_U3297) );
  AND2_X1 U10807 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9555), .ZN(P1_U3298) );
  AND2_X1 U10808 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9555), .ZN(P1_U3299) );
  AND2_X1 U10809 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9555), .ZN(P1_U3300) );
  AND2_X1 U10810 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9555), .ZN(P1_U3301) );
  INV_X1 U10811 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U10812 ( .A1(n9554), .A2(n10225), .ZN(P1_U3302) );
  AND2_X1 U10813 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9555), .ZN(P1_U3303) );
  AND2_X1 U10814 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9555), .ZN(P1_U3304) );
  AND2_X1 U10815 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9555), .ZN(P1_U3305) );
  INV_X1 U10816 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U10817 ( .A1(n9554), .A2(n10191), .ZN(P1_U3306) );
  INV_X1 U10818 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U10819 ( .A1(n9554), .A2(n10066), .ZN(P1_U3307) );
  AND2_X1 U10820 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9555), .ZN(P1_U3308) );
  AND2_X1 U10821 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9555), .ZN(P1_U3309) );
  INV_X1 U10822 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U10823 ( .A1(n9554), .A2(n10252), .ZN(P1_U3310) );
  AND2_X1 U10824 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9555), .ZN(P1_U3311) );
  AND2_X1 U10825 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9555), .ZN(P1_U3312) );
  AND2_X1 U10826 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9555), .ZN(P1_U3313) );
  AND2_X1 U10827 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9555), .ZN(P1_U3314) );
  AND2_X1 U10828 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9555), .ZN(P1_U3315) );
  AND2_X1 U10829 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9555), .ZN(P1_U3316) );
  INV_X1 U10830 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10104) );
  NOR2_X1 U10831 ( .A1(n9554), .A2(n10104), .ZN(P1_U3317) );
  AND2_X1 U10832 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9555), .ZN(P1_U3318) );
  AND2_X1 U10833 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9555), .ZN(P1_U3319) );
  AND2_X1 U10834 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9555), .ZN(P1_U3320) );
  AND2_X1 U10835 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9555), .ZN(P1_U3321) );
  AND2_X1 U10836 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9555), .ZN(P1_U3322) );
  AND2_X1 U10837 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9555), .ZN(P1_U3323) );
  AOI21_X1 U10838 ( .B1(n9654), .B2(n9557), .A(n9556), .ZN(n9558) );
  AOI211_X1 U10839 ( .C1(n9561), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9675)
         );
  INV_X1 U10840 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9562) );
  AOI22_X1 U10841 ( .A1(n4404), .A2(n9675), .B1(n9562), .B2(n9672), .ZN(
        P1_U3453) );
  INV_X1 U10842 ( .A(n9563), .ZN(n9568) );
  OAI21_X1 U10843 ( .B1(n9565), .B2(n9665), .A(n9564), .ZN(n9567) );
  AOI211_X1 U10844 ( .C1(n9668), .C2(n9568), .A(n9567), .B(n9566), .ZN(n9676)
         );
  INV_X1 U10845 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U10846 ( .A1(n4404), .A2(n9676), .B1(n10209), .B2(n9672), .ZN(
        P1_U3456) );
  AOI22_X1 U10847 ( .A1(n9570), .A2(n9625), .B1(n9626), .B2(n9569), .ZN(n9572)
         );
  OAI211_X1 U10848 ( .C1(n9573), .C2(n9654), .A(n9572), .B(n9571), .ZN(n9574)
         );
  NOR2_X1 U10849 ( .A1(n9575), .A2(n9574), .ZN(n9677) );
  INV_X1 U10850 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9576) );
  AOI22_X1 U10851 ( .A1(n4404), .A2(n9677), .B1(n9576), .B2(n9672), .ZN(
        P1_U3459) );
  INV_X1 U10852 ( .A(n9577), .ZN(n9584) );
  NOR2_X1 U10853 ( .A1(n9578), .A2(n9654), .ZN(n9583) );
  OAI22_X1 U10854 ( .A1(n9580), .A2(n9656), .B1(n9579), .B2(n9665), .ZN(n9581)
         );
  NOR4_X1 U10855 ( .A1(n9584), .A2(n9583), .A3(n9582), .A4(n9581), .ZN(n9678)
         );
  INV_X1 U10856 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U10857 ( .A1(n4404), .A2(n9678), .B1(n10102), .B2(n9672), .ZN(
        P1_U3462) );
  AOI22_X1 U10858 ( .A1(n9586), .A2(n9626), .B1(n9585), .B2(n9625), .ZN(n9588)
         );
  OAI211_X1 U10859 ( .C1(n9589), .C2(n9654), .A(n9588), .B(n9587), .ZN(n9590)
         );
  NOR2_X1 U10860 ( .A1(n9591), .A2(n9590), .ZN(n9679) );
  INV_X1 U10861 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9592) );
  AOI22_X1 U10862 ( .A1(n4404), .A2(n9679), .B1(n9592), .B2(n9672), .ZN(
        P1_U3465) );
  INV_X1 U10863 ( .A(n9593), .ZN(n9600) );
  AOI22_X1 U10864 ( .A1(n9595), .A2(n9626), .B1(n9625), .B2(n9594), .ZN(n9597)
         );
  NAND3_X1 U10865 ( .A1(n9598), .A2(n9597), .A3(n9596), .ZN(n9599) );
  AOI21_X1 U10866 ( .B1(n9652), .B2(n9600), .A(n9599), .ZN(n9681) );
  INV_X1 U10867 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9601) );
  AOI22_X1 U10868 ( .A1(n4404), .A2(n9681), .B1(n9601), .B2(n9672), .ZN(
        P1_U3468) );
  INV_X1 U10869 ( .A(n9602), .ZN(n9609) );
  NOR2_X1 U10870 ( .A1(n9603), .A2(n9654), .ZN(n9608) );
  OAI22_X1 U10871 ( .A1(n9605), .A2(n9656), .B1(n9604), .B2(n9665), .ZN(n9606)
         );
  NOR4_X1 U10872 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n9682)
         );
  INV_X1 U10873 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9610) );
  AOI22_X1 U10874 ( .A1(n4404), .A2(n9682), .B1(n9610), .B2(n9672), .ZN(
        P1_U3471) );
  OAI21_X1 U10875 ( .B1(n9612), .B2(n9665), .A(n9611), .ZN(n9615) );
  INV_X1 U10876 ( .A(n9613), .ZN(n9614) );
  AOI211_X1 U10877 ( .C1(n9668), .C2(n9616), .A(n9615), .B(n9614), .ZN(n9684)
         );
  INV_X1 U10878 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U10879 ( .A1(n4404), .A2(n9684), .B1(n10127), .B2(n9672), .ZN(
        P1_U3474) );
  INV_X1 U10880 ( .A(n9617), .ZN(n9622) );
  OAI21_X1 U10881 ( .B1(n9619), .B2(n9665), .A(n9618), .ZN(n9621) );
  AOI211_X1 U10882 ( .C1(n9668), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9686)
         );
  INV_X1 U10883 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9623) );
  AOI22_X1 U10884 ( .A1(n4404), .A2(n9686), .B1(n9623), .B2(n9672), .ZN(
        P1_U3477) );
  AOI22_X1 U10885 ( .A1(n9627), .A2(n9626), .B1(n9625), .B2(n9624), .ZN(n9628)
         );
  OAI211_X1 U10886 ( .C1(n9630), .C2(n9654), .A(n9629), .B(n9628), .ZN(n9631)
         );
  NOR2_X1 U10887 ( .A1(n9632), .A2(n9631), .ZN(n9688) );
  INV_X1 U10888 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9633) );
  AOI22_X1 U10889 ( .A1(n4404), .A2(n9688), .B1(n9633), .B2(n9672), .ZN(
        P1_U3480) );
  OAI211_X1 U10890 ( .C1(n9636), .C2(n9665), .A(n9635), .B(n9634), .ZN(n9637)
         );
  AOI21_X1 U10891 ( .B1(n9652), .B2(n9638), .A(n9637), .ZN(n9690) );
  INV_X1 U10892 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9639) );
  AOI22_X1 U10893 ( .A1(n4404), .A2(n9690), .B1(n9639), .B2(n9672), .ZN(
        P1_U3483) );
  OAI21_X1 U10894 ( .B1(n9641), .B2(n9665), .A(n9640), .ZN(n9642) );
  AOI21_X1 U10895 ( .B1(n9643), .B2(n9668), .A(n9642), .ZN(n9644) );
  AND2_X1 U10896 ( .A1(n9645), .A2(n9644), .ZN(n9692) );
  INV_X1 U10897 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9646) );
  AOI22_X1 U10898 ( .A1(n4404), .A2(n9692), .B1(n9646), .B2(n9672), .ZN(
        P1_U3486) );
  OAI21_X1 U10899 ( .B1(n9648), .B2(n9665), .A(n9647), .ZN(n9650) );
  AOI211_X1 U10900 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9694)
         );
  INV_X1 U10901 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9653) );
  AOI22_X1 U10902 ( .A1(n4404), .A2(n9694), .B1(n9653), .B2(n9672), .ZN(
        P1_U3489) );
  NOR2_X1 U10903 ( .A1(n9655), .A2(n9654), .ZN(n9662) );
  OAI22_X1 U10904 ( .A1(n9658), .A2(n9665), .B1(n9657), .B2(n9656), .ZN(n9659)
         );
  NOR4_X1 U10905 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9696)
         );
  INV_X1 U10906 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U10907 ( .A1(n4404), .A2(n9696), .B1(n9663), .B2(n9672), .ZN(
        P1_U3492) );
  OAI21_X1 U10908 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9667) );
  AOI21_X1 U10909 ( .B1(n9669), .B2(n9668), .A(n9667), .ZN(n9670) );
  AND2_X1 U10910 ( .A1(n9671), .A2(n9670), .ZN(n9699) );
  INV_X1 U10911 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9673) );
  AOI22_X1 U10912 ( .A1(n4404), .A2(n9699), .B1(n9673), .B2(n9672), .ZN(
        P1_U3495) );
  AOI22_X1 U10913 ( .A1(n9381), .A2(n9675), .B1(n9674), .B2(n9697), .ZN(
        P1_U3522) );
  AOI22_X1 U10914 ( .A1(n9381), .A2(n9676), .B1(n6444), .B2(n9697), .ZN(
        P1_U3523) );
  AOI22_X1 U10915 ( .A1(n9381), .A2(n9677), .B1(n6548), .B2(n9697), .ZN(
        P1_U3524) );
  AOI22_X1 U10916 ( .A1(n9700), .A2(n9678), .B1(n6552), .B2(n9697), .ZN(
        P1_U3525) );
  AOI22_X1 U10917 ( .A1(n9700), .A2(n9679), .B1(n6555), .B2(n9697), .ZN(
        P1_U3526) );
  AOI22_X1 U10918 ( .A1(n9700), .A2(n9681), .B1(n9680), .B2(n9697), .ZN(
        P1_U3527) );
  AOI22_X1 U10919 ( .A1(n9700), .A2(n9682), .B1(n6559), .B2(n9697), .ZN(
        P1_U3528) );
  AOI22_X1 U10920 ( .A1(n9700), .A2(n9684), .B1(n9683), .B2(n9697), .ZN(
        P1_U3529) );
  AOI22_X1 U10921 ( .A1(n9700), .A2(n9686), .B1(n9685), .B2(n9697), .ZN(
        P1_U3530) );
  AOI22_X1 U10922 ( .A1(n9700), .A2(n9688), .B1(n9687), .B2(n9697), .ZN(
        P1_U3531) );
  AOI22_X1 U10923 ( .A1(n9700), .A2(n9690), .B1(n9689), .B2(n9697), .ZN(
        P1_U3532) );
  AOI22_X1 U10924 ( .A1(n9700), .A2(n9692), .B1(n9691), .B2(n9697), .ZN(
        P1_U3533) );
  AOI22_X1 U10925 ( .A1(n9700), .A2(n9694), .B1(n9693), .B2(n9697), .ZN(
        P1_U3534) );
  INV_X1 U10926 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10927 ( .A1(n9700), .A2(n9696), .B1(n9695), .B2(n9697), .ZN(
        P1_U3535) );
  AOI22_X1 U10928 ( .A1(n9700), .A2(n9699), .B1(n9698), .B2(n9697), .ZN(
        P1_U3536) );
  XNOR2_X1 U10929 ( .A(n9701), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9702) );
  NOR2_X1 U10930 ( .A1(n9872), .A2(n9702), .ZN(n9705) );
  OAI22_X1 U10931 ( .A1(n9841), .A2(n9703), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7140), .ZN(n9704) );
  NOR2_X1 U10932 ( .A1(n9705), .A2(n9704), .ZN(n9712) );
  NAND2_X1 U10933 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  NAND2_X1 U10934 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  AOI22_X1 U10935 ( .A1(n9863), .A2(n9710), .B1(n9856), .B2(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n9711) );
  AND2_X1 U10936 ( .A1(n9712), .A2(n9711), .ZN(n9717) );
  XOR2_X1 U10937 ( .A(n9713), .B(n9714), .Z(n9715) );
  NAND2_X1 U10938 ( .A1(n9715), .A2(n9868), .ZN(n9716) );
  NAND2_X1 U10939 ( .A1(n9717), .A2(n9716), .ZN(P2_U3183) );
  NAND2_X1 U10940 ( .A1(n9718), .A2(n5849), .ZN(n9719) );
  NAND2_X1 U10941 ( .A1(n9720), .A2(n9719), .ZN(n9721) );
  NAND2_X1 U10942 ( .A1(n9863), .A2(n9721), .ZN(n9723) );
  NAND2_X1 U10943 ( .A1(n9856), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n9722) );
  OAI211_X1 U10944 ( .C1(n9841), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9725)
         );
  INV_X1 U10945 ( .A(n9725), .ZN(n9737) );
  AOI21_X1 U10946 ( .B1(n9728), .B2(n9727), .A(n9726), .ZN(n9729) );
  OR2_X1 U10947 ( .A1(n9729), .A2(n9847), .ZN(n9735) );
  INV_X1 U10948 ( .A(n9730), .ZN(n9733) );
  AND2_X1 U10949 ( .A1(n9731), .A2(n5848), .ZN(n9732) );
  OAI21_X1 U10950 ( .B1(n9733), .B2(n9732), .A(n4902), .ZN(n9734) );
  NAND4_X1 U10951 ( .A1(n9737), .A2(n9736), .A3(n9735), .A4(n9734), .ZN(
        P2_U3185) );
  NOR2_X1 U10952 ( .A1(n9738), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9739) );
  OAI21_X1 U10953 ( .B1(n9740), .B2(n9739), .A(n9863), .ZN(n9743) );
  NAND2_X1 U10954 ( .A1(n9858), .A2(n4855), .ZN(n9742) );
  NAND2_X1 U10955 ( .A1(n9856), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n9741) );
  AND3_X1 U10956 ( .A1(n9743), .A2(n9742), .A3(n9741), .ZN(n9752) );
  XOR2_X1 U10957 ( .A(n9745), .B(n9744), .Z(n9746) );
  NAND2_X1 U10958 ( .A1(n9746), .A2(n9868), .ZN(n9750) );
  NOR2_X1 U10959 ( .A1(n4506), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9747) );
  OAI21_X1 U10960 ( .B1(n9748), .B2(n9747), .A(n4902), .ZN(n9749) );
  NAND4_X1 U10961 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(
        P2_U3187) );
  AOI21_X1 U10962 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(n9769) );
  NOR2_X1 U10963 ( .A1(n9841), .A2(n9756), .ZN(n9766) );
  AOI21_X1 U10964 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9764) );
  AOI21_X1 U10965 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(n9763) );
  OAI22_X1 U10966 ( .A1(n9764), .A2(n9847), .B1(n9763), .B2(n9849), .ZN(n9765)
         );
  AOI211_X1 U10967 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9856), .A(n9766), .B(
        n9765), .ZN(n9768) );
  OAI211_X1 U10968 ( .C1(n9769), .C2(n9872), .A(n9768), .B(n9767), .ZN(
        P2_U3188) );
  AOI21_X1 U10969 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9786) );
  AOI21_X1 U10970 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(n9776) );
  NOR2_X1 U10971 ( .A1(n9776), .A2(n9847), .ZN(n9783) );
  AOI21_X1 U10972 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9781) );
  OAI22_X1 U10973 ( .A1(n9849), .A2(n9781), .B1(n9841), .B2(n9780), .ZN(n9782)
         );
  AOI211_X1 U10974 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9856), .A(n9783), .B(
        n9782), .ZN(n9785) );
  OAI211_X1 U10975 ( .C1(n9786), .C2(n9872), .A(n9785), .B(n9784), .ZN(
        P2_U3190) );
  AOI21_X1 U10976 ( .B1(n6302), .B2(n9788), .A(n9787), .ZN(n9802) );
  OAI22_X1 U10977 ( .A1(n9841), .A2(n9790), .B1(n9839), .B2(n9789), .ZN(n9799)
         );
  AOI21_X1 U10978 ( .B1(n6303), .B2(n9792), .A(n9791), .ZN(n9797) );
  AOI21_X1 U10979 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n9796) );
  OAI22_X1 U10980 ( .A1(n9797), .A2(n9849), .B1(n9796), .B2(n9847), .ZN(n9798)
         );
  NOR3_X1 U10981 ( .A1(n9800), .A2(n9799), .A3(n9798), .ZN(n9801) );
  OAI21_X1 U10982 ( .B1(n9802), .B2(n9872), .A(n9801), .ZN(P2_U3191) );
  AOI21_X1 U10983 ( .B1(n6300), .B2(n9804), .A(n9803), .ZN(n9818) );
  OAI22_X1 U10984 ( .A1(n9841), .A2(n9806), .B1(n9839), .B2(n9805), .ZN(n9815)
         );
  AOI21_X1 U10985 ( .B1(n9808), .B2(n6301), .A(n9807), .ZN(n9813) );
  AOI21_X1 U10986 ( .B1(n9811), .B2(n9810), .A(n9809), .ZN(n9812) );
  OAI22_X1 U10987 ( .A1(n9813), .A2(n9849), .B1(n9812), .B2(n9847), .ZN(n9814)
         );
  NOR3_X1 U10988 ( .A1(n9816), .A2(n9815), .A3(n9814), .ZN(n9817) );
  OAI21_X1 U10989 ( .B1(n9818), .B2(n9872), .A(n9817), .ZN(P2_U3193) );
  AOI21_X1 U10990 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9835) );
  INV_X1 U10991 ( .A(n9822), .ZN(n9824) );
  OAI21_X1 U10992 ( .B1(n9841), .B2(n9824), .A(n9823), .ZN(n9833) );
  AOI21_X1 U10993 ( .B1(n8357), .B2(n9826), .A(n9825), .ZN(n9831) );
  AOI21_X1 U10994 ( .B1(n9829), .B2(n9828), .A(n9827), .ZN(n9830) );
  OAI22_X1 U10995 ( .A1(n9831), .A2(n9849), .B1(n9830), .B2(n9847), .ZN(n9832)
         );
  AOI211_X1 U10996 ( .C1(n9856), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n9833), .B(
        n9832), .ZN(n9834) );
  OAI21_X1 U10997 ( .B1(n9835), .B2(n9872), .A(n9834), .ZN(P2_U3195) );
  AOI21_X1 U10998 ( .B1(n10055), .B2(n9837), .A(n9836), .ZN(n9855) );
  OAI22_X1 U10999 ( .A1(n9841), .A2(n9840), .B1(n9839), .B2(n9838), .ZN(n9852)
         );
  AOI21_X1 U11000 ( .B1(n8322), .B2(n9843), .A(n9842), .ZN(n9850) );
  AOI21_X1 U11001 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9848) );
  OAI22_X1 U11002 ( .A1(n9850), .A2(n9849), .B1(n9848), .B2(n9847), .ZN(n9851)
         );
  NOR3_X1 U11003 ( .A1(n9853), .A2(n9852), .A3(n9851), .ZN(n9854) );
  OAI21_X1 U11004 ( .B1(n9855), .B2(n9872), .A(n9854), .ZN(P2_U3197) );
  AOI22_X1 U11005 ( .A1(n9858), .A2(n9857), .B1(n9856), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9876) );
  AOI21_X1 U11006 ( .B1(n9860), .B2(n10128), .A(n9859), .ZN(n9873) );
  NAND2_X1 U11007 ( .A1(n9861), .A2(n10211), .ZN(n9862) );
  NAND2_X1 U11008 ( .A1(n9862), .A2(n4716), .ZN(n9864) );
  NAND2_X1 U11009 ( .A1(n9864), .A2(n9863), .ZN(n9871) );
  OAI21_X1 U11010 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(n9869) );
  NAND2_X1 U11011 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  OAI211_X1 U11012 ( .C1(n9873), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9874)
         );
  INV_X1 U11013 ( .A(n9874), .ZN(n9875) );
  OAI211_X1 U11014 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9877), .A(n9876), .B(
        n9875), .ZN(P2_U3199) );
  NAND2_X1 U11015 ( .A1(n9879), .A2(n9878), .ZN(n9881) );
  NAND2_X1 U11016 ( .A1(n9881), .A2(n9880), .ZN(n9882) );
  XOR2_X1 U11017 ( .A(n9887), .B(n9882), .Z(n9886) );
  AOI222_X1 U11018 ( .A1(n6212), .A2(n9886), .B1(n9885), .B2(n8370), .C1(n9884), .C2(n9883), .ZN(n9899) );
  XNOR2_X1 U11019 ( .A(n9888), .B(n9887), .ZN(n9897) );
  AOI222_X1 U11020 ( .A1(n9897), .A2(n9892), .B1(n9891), .B2(n9890), .C1(n9896), .C2(n9889), .ZN(n9893) );
  OAI221_X1 U11021 ( .B1(n8340), .B2(n9899), .C1(n8373), .C2(n5849), .A(n9893), 
        .ZN(P2_U3230) );
  INV_X1 U11022 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U11023 ( .A1(n9941), .A2(n9895), .B1(n9894), .B2(n9939), .ZN(
        P2_U3396) );
  INV_X1 U11024 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U11025 ( .A1(n9897), .A2(n9938), .B1(n9918), .B2(n9896), .ZN(n9898)
         );
  AND2_X1 U11026 ( .A1(n9899), .A2(n9898), .ZN(n9942) );
  AOI22_X1 U11027 ( .A1(n9941), .A2(n10115), .B1(n9942), .B2(n9939), .ZN(
        P2_U3399) );
  INV_X1 U11028 ( .A(n9900), .ZN(n9904) );
  OAI22_X1 U11029 ( .A1(n9902), .A2(n9912), .B1(n9901), .B2(n9933), .ZN(n9903)
         );
  NOR2_X1 U11030 ( .A1(n9904), .A2(n9903), .ZN(n9943) );
  AOI22_X1 U11031 ( .A1(n9941), .A2(n5890), .B1(n9943), .B2(n9939), .ZN(
        P2_U3402) );
  INV_X1 U11032 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9910) );
  INV_X1 U11033 ( .A(n9905), .ZN(n9909) );
  OAI22_X1 U11034 ( .A1(n9907), .A2(n9912), .B1(n9906), .B2(n9933), .ZN(n9908)
         );
  NOR2_X1 U11035 ( .A1(n9909), .A2(n9908), .ZN(n9944) );
  AOI22_X1 U11036 ( .A1(n9941), .A2(n9910), .B1(n9944), .B2(n9939), .ZN(
        P2_U3408) );
  INV_X1 U11037 ( .A(n9911), .ZN(n9913) );
  NOR3_X1 U11038 ( .A1(n9914), .A2(n9913), .A3(n9912), .ZN(n9916) );
  AOI211_X1 U11039 ( .C1(n9918), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9946)
         );
  AOI22_X1 U11040 ( .A1(n9941), .A2(n5933), .B1(n9946), .B2(n9939), .ZN(
        P2_U3411) );
  INV_X1 U11041 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9923) );
  NOR2_X1 U11042 ( .A1(n9919), .A2(n9933), .ZN(n9921) );
  AOI211_X1 U11043 ( .C1(n9938), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9947)
         );
  AOI22_X1 U11044 ( .A1(n9941), .A2(n9923), .B1(n9947), .B2(n9939), .ZN(
        P2_U3414) );
  INV_X1 U11045 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10022) );
  OAI22_X1 U11046 ( .A1(n9926), .A2(n9925), .B1(n9924), .B2(n9933), .ZN(n9927)
         );
  NOR2_X1 U11047 ( .A1(n9928), .A2(n9927), .ZN(n9948) );
  AOI22_X1 U11048 ( .A1(n9941), .A2(n10022), .B1(n9948), .B2(n9939), .ZN(
        P2_U3417) );
  NOR2_X1 U11049 ( .A1(n9929), .A2(n9933), .ZN(n9931) );
  AOI211_X1 U11050 ( .C1(n9938), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9949)
         );
  AOI22_X1 U11051 ( .A1(n9941), .A2(n5971), .B1(n9949), .B2(n9939), .ZN(
        P2_U3420) );
  INV_X1 U11052 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U11053 ( .A1(n9934), .A2(n9933), .ZN(n9936) );
  AOI211_X1 U11054 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9950)
         );
  AOI22_X1 U11055 ( .A1(n9941), .A2(n9940), .B1(n9950), .B2(n9939), .ZN(
        P2_U3423) );
  AOI22_X1 U11056 ( .A1(n9951), .A2(n9942), .B1(n5848), .B2(n6296), .ZN(
        P2_U3462) );
  AOI22_X1 U11057 ( .A1(n9951), .A2(n9943), .B1(n6398), .B2(n6296), .ZN(
        P2_U3463) );
  AOI22_X1 U11058 ( .A1(n9951), .A2(n9944), .B1(n6304), .B2(n6296), .ZN(
        P2_U3465) );
  AOI22_X1 U11059 ( .A1(n9951), .A2(n9946), .B1(n9945), .B2(n6296), .ZN(
        P2_U3466) );
  AOI22_X1 U11060 ( .A1(n9951), .A2(n9947), .B1(n5949), .B2(n6296), .ZN(
        P2_U3467) );
  AOI22_X1 U11061 ( .A1(n9951), .A2(n9948), .B1(n6302), .B2(n6296), .ZN(
        P2_U3468) );
  AOI22_X1 U11062 ( .A1(n9951), .A2(n9949), .B1(n5974), .B2(n6296), .ZN(
        P2_U3469) );
  AOI22_X1 U11063 ( .A1(n9951), .A2(n9950), .B1(n6300), .B2(n6296), .ZN(
        P2_U3470) );
  NOR2_X1 U11064 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  XOR2_X1 U11065 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9954), .Z(ADD_1068_U5) );
  XOR2_X1 U11066 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11067 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9956), .A(n9955), .ZN(
        n9957) );
  XOR2_X1 U11068 ( .A(n9957), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55) );
  XNOR2_X1 U11069 ( .A(n9959), .B(n9958), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11070 ( .A(n9961), .B(n9960), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11071 ( .A(n9963), .B(n9962), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11072 ( .A(n9965), .B(n9964), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11073 ( .A(n9967), .B(n9966), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11074 ( .A(n9969), .B(n9968), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11075 ( .A(n9971), .B(n9970), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11076 ( .A(n9973), .B(n9972), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11077 ( .A(n9975), .B(n9974), .ZN(ADD_1068_U50) );
  NOR4_X1 U11078 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        SI_7_), .A4(P2_REG1_REG_23__SCAN_IN), .ZN(n9979) );
  NOR4_X1 U11079 ( .A1(P2_REG0_REG_30__SCAN_IN), .A2(P2_REG1_REG_27__SCAN_IN), 
        .A3(P2_REG1_REG_26__SCAN_IN), .A4(P2_REG1_REG_24__SCAN_IN), .ZN(n9978)
         );
  NOR4_X1 U11080 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P1_DATAO_REG_18__SCAN_IN), 
        .A3(SI_3_), .A4(P2_REG2_REG_4__SCAN_IN), .ZN(n9977) );
  NOR4_X1 U11081 ( .A1(SI_8_), .A2(P2_REG0_REG_10__SCAN_IN), .A3(
        P2_REG0_REG_9__SCAN_IN), .A4(P2_REG0_REG_3__SCAN_IN), .ZN(n9976) );
  NAND4_X1 U11082 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n10020) );
  NOR2_X1 U11083 ( .A1(SI_12_), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U11084 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9980) );
  AND4_X1 U11085 ( .A1(n10185), .A2(n9981), .A3(P1_ADDR_REG_4__SCAN_IN), .A4(
        n9980), .ZN(n9984) );
  NOR4_X1 U11086 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P2_DATAO_REG_23__SCAN_IN), .A3(P1_DATAO_REG_22__SCAN_IN), .A4(P2_ADDR_REG_10__SCAN_IN), .ZN(n9983) );
  NOR4_X1 U11087 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_REG1_REG_30__SCAN_IN), 
        .A3(P1_DATAO_REG_21__SCAN_IN), .A4(P1_REG3_REG_10__SCAN_IN), .ZN(n9982) );
  NAND4_X1 U11088 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n10019) );
  NOR4_X1 U11089 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P1_DATAO_REG_28__SCAN_IN), .A3(P2_REG2_REG_10__SCAN_IN), .A4(P2_U3151), .ZN(n9996) );
  NOR4_X1 U11090 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG1_REG_17__SCAN_IN), 
        .A3(P2_REG1_REG_2__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n9995)
         );
  NAND4_X1 U11091 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .A3(P2_IR_REG_28__SCAN_IN), .A4(P2_REG3_REG_9__SCAN_IN), .ZN(n9993) );
  INV_X1 U11092 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9986) );
  INV_X1 U11093 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10148) );
  NAND4_X1 U11094 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(P2_REG0_REG_31__SCAN_IN), .A3(n9986), .A4(n10148), .ZN(n9992) );
  NOR4_X1 U11095 ( .A1(SI_0_), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        P1_IR_REG_2__SCAN_IN), .A4(P1_REG0_REG_7__SCAN_IN), .ZN(n9990) );
  NOR4_X1 U11096 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(P2_REG1_REG_18__SCAN_IN), 
        .A3(P1_REG0_REG_27__SCAN_IN), .A4(P1_REG0_REG_21__SCAN_IN), .ZN(n9989)
         );
  NOR4_X1 U11097 ( .A1(P2_RD_REG_SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), .A3(
        P1_ADDR_REG_17__SCAN_IN), .A4(P1_ADDR_REG_16__SCAN_IN), .ZN(n9988) );
  NOR4_X1 U11098 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG2_REG_11__SCAN_IN), 
        .A3(P1_REG2_REG_9__SCAN_IN), .A4(P1_REG2_REG_8__SCAN_IN), .ZN(n9987)
         );
  NAND4_X1 U11099 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n9991)
         );
  NOR3_X1 U11100 ( .A1(n9993), .A2(n9992), .A3(n9991), .ZN(n9994) );
  NAND3_X1 U11101 ( .A1(n9996), .A2(n9995), .A3(n9994), .ZN(n10018) );
  NAND4_X1 U11102 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(SI_21_), .A3(
        P2_DATAO_REG_15__SCAN_IN), .A4(P2_REG1_REG_10__SCAN_IN), .ZN(n10000)
         );
  NAND4_X1 U11103 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(SI_6_), .A3(
        P2_DATAO_REG_4__SCAN_IN), .A4(P2_REG0_REG_7__SCAN_IN), .ZN(n9999) );
  NAND4_X1 U11104 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9998) );
  NAND4_X1 U11105 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(P1_REG0_REG_29__SCAN_IN), .ZN(n9997)
         );
  NOR4_X1 U11106 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(n10016) );
  NAND4_X1 U11107 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(P1_D_REG_0__SCAN_IN), 
        .A3(P1_D_REG_1__SCAN_IN), .A4(P2_ADDR_REG_13__SCAN_IN), .ZN(n10004) );
  NAND4_X1 U11108 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .A3(P2_REG0_REG_29__SCAN_IN), .A4(P2_DATAO_REG_1__SCAN_IN), .ZN(n10003) );
  NAND4_X1 U11109 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        SI_10_), .A4(P1_DATAO_REG_7__SCAN_IN), .ZN(n10002) );
  NAND4_X1 U11110 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_REG0_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_20__SCAN_IN), .A4(P2_ADDR_REG_17__SCAN_IN), .ZN(n10001) );
  NOR4_X1 U11111 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10015) );
  NAND4_X1 U11112 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(P2_REG2_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_15__SCAN_IN), .A4(P1_REG3_REG_24__SCAN_IN), .ZN(n10008) );
  NAND4_X1 U11113 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(P1_REG0_REG_16__SCAN_IN), .A4(P1_REG2_REG_0__SCAN_IN), .ZN(n10007)
         );
  NAND4_X1 U11114 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_26__SCAN_IN), .A4(P1_ADDR_REG_10__SCAN_IN), .ZN(n10006) );
  NAND4_X1 U11115 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P2_REG2_REG_24__SCAN_IN), 
        .A3(P2_REG2_REG_17__SCAN_IN), .A4(P1_DATAO_REG_31__SCAN_IN), .ZN(
        n10005) );
  NOR4_X1 U11116 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10014) );
  NAND4_X1 U11117 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_REG3_REG_13__SCAN_IN), .A4(P1_REG3_REG_7__SCAN_IN), .ZN(n10012) );
  NAND4_X1 U11118 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .A3(P1_IR_REG_11__SCAN_IN), .A4(P1_IR_REG_27__SCAN_IN), .ZN(n10011) );
  NAND4_X1 U11119 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG2_REG_5__SCAN_IN), .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n10010)
         );
  NAND4_X1 U11120 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(P1_REG0_REG_3__SCAN_IN), .A4(P1_REG0_REG_1__SCAN_IN), .ZN(n10009)
         );
  NOR4_X1 U11121 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10013) );
  NAND4_X1 U11122 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10017) );
  NOR4_X1 U11123 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10279) );
  AOI22_X1 U11124 ( .A1(n10023), .A2(keyinput64), .B1(n10022), .B2(keyinput107), .ZN(n10021) );
  OAI221_X1 U11125 ( .B1(n10023), .B2(keyinput64), .C1(n10022), .C2(
        keyinput107), .A(n10021), .ZN(n10032) );
  XNOR2_X1 U11126 ( .A(keyinput70), .B(n8176), .ZN(n10031) );
  XNOR2_X1 U11127 ( .A(keyinput37), .B(n10024), .ZN(n10030) );
  XNOR2_X1 U11128 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput25), .ZN(n10028) );
  XNOR2_X1 U11129 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput19), .ZN(n10027) );
  XNOR2_X1 U11130 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput35), .ZN(n10026) );
  XNOR2_X1 U11131 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput22), .ZN(n10025)
         );
  NAND4_X1 U11132 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10029) );
  NOR4_X1 U11133 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        n10079) );
  AOI22_X1 U11134 ( .A1(n10035), .A2(keyinput52), .B1(keyinput84), .B2(n10034), 
        .ZN(n10033) );
  OAI221_X1 U11135 ( .B1(n10035), .B2(keyinput52), .C1(n10034), .C2(keyinput84), .A(n10033), .ZN(n10047) );
  AOI22_X1 U11136 ( .A1(n10037), .A2(keyinput15), .B1(n9891), .B2(keyinput20), 
        .ZN(n10036) );
  OAI221_X1 U11137 ( .B1(n10037), .B2(keyinput15), .C1(n9891), .C2(keyinput20), 
        .A(n10036), .ZN(n10046) );
  AOI22_X1 U11138 ( .A1(n10040), .A2(keyinput68), .B1(keyinput96), .B2(n10039), 
        .ZN(n10038) );
  OAI221_X1 U11139 ( .B1(n10040), .B2(keyinput68), .C1(n10039), .C2(keyinput96), .A(n10038), .ZN(n10045) );
  XOR2_X1 U11140 ( .A(n10041), .B(keyinput14), .Z(n10043) );
  XNOR2_X1 U11141 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput7), .ZN(n10042) );
  NAND2_X1 U11142 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  NOR4_X1 U11143 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n10078) );
  AOI22_X1 U11144 ( .A1(n5849), .A2(keyinput24), .B1(keyinput43), .B2(n10049), 
        .ZN(n10048) );
  OAI221_X1 U11145 ( .B1(n5849), .B2(keyinput24), .C1(n10049), .C2(keyinput43), 
        .A(n10048), .ZN(n10062) );
  AOI22_X1 U11146 ( .A1(n10052), .A2(keyinput112), .B1(n10051), .B2(keyinput89), .ZN(n10050) );
  OAI221_X1 U11147 ( .B1(n10052), .B2(keyinput112), .C1(n10051), .C2(
        keyinput89), .A(n10050), .ZN(n10061) );
  AOI22_X1 U11148 ( .A1(n10055), .A2(keyinput98), .B1(n10054), .B2(keyinput42), 
        .ZN(n10053) );
  OAI221_X1 U11149 ( .B1(n10055), .B2(keyinput98), .C1(n10054), .C2(keyinput42), .A(n10053), .ZN(n10060) );
  XOR2_X1 U11150 ( .A(n10056), .B(keyinput81), .Z(n10058) );
  XNOR2_X1 U11151 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput60), .ZN(n10057)
         );
  NAND2_X1 U11152 ( .A1(n10058), .A2(n10057), .ZN(n10059) );
  NOR4_X1 U11153 ( .A1(n10062), .A2(n10061), .A3(n10060), .A4(n10059), .ZN(
        n10077) );
  INV_X1 U11154 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U11155 ( .A1(n10065), .A2(keyinput100), .B1(keyinput71), .B2(n10064), .ZN(n10063) );
  OAI221_X1 U11156 ( .B1(n10065), .B2(keyinput100), .C1(n10064), .C2(
        keyinput71), .A(n10063), .ZN(n10069) );
  XNOR2_X1 U11157 ( .A(n10066), .B(keyinput118), .ZN(n10068) );
  XOR2_X1 U11158 ( .A(SI_0_), .B(keyinput27), .Z(n10067) );
  OR3_X1 U11159 ( .A1(n10069), .A2(n10068), .A3(n10067), .ZN(n10075) );
  INV_X1 U11160 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10071) );
  AOI22_X1 U11161 ( .A1(n10071), .A2(keyinput111), .B1(keyinput126), .B2(n5599), .ZN(n10070) );
  OAI221_X1 U11162 ( .B1(n10071), .B2(keyinput111), .C1(n5599), .C2(
        keyinput126), .A(n10070), .ZN(n10074) );
  AOI22_X1 U11163 ( .A1(n8290), .A2(keyinput57), .B1(P2_U3151), .B2(keyinput47), .ZN(n10072) );
  OAI221_X1 U11164 ( .B1(n8290), .B2(keyinput57), .C1(P2_U3151), .C2(
        keyinput47), .A(n10072), .ZN(n10073) );
  NOR3_X1 U11165 ( .A1(n10075), .A2(n10074), .A3(n10073), .ZN(n10076) );
  NAND4_X1 U11166 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10272) );
  AOI22_X1 U11167 ( .A1(n5779), .A2(keyinput45), .B1(keyinput58), .B2(n10081), 
        .ZN(n10080) );
  OAI221_X1 U11168 ( .B1(n5779), .B2(keyinput45), .C1(n10081), .C2(keyinput58), 
        .A(n10080), .ZN(n10091) );
  INV_X1 U11169 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U11170 ( .A1(n10084), .A2(keyinput104), .B1(n10083), .B2(keyinput44), .ZN(n10082) );
  OAI221_X1 U11171 ( .B1(n10084), .B2(keyinput104), .C1(n10083), .C2(
        keyinput44), .A(n10082), .ZN(n10090) );
  XNOR2_X1 U11172 ( .A(SI_8_), .B(keyinput80), .ZN(n10088) );
  XNOR2_X1 U11173 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput83), .ZN(n10087) );
  XNOR2_X1 U11174 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput66), .ZN(n10086) );
  XNOR2_X1 U11175 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput115), .ZN(n10085) );
  NAND4_X1 U11176 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10089) );
  NOR3_X1 U11177 ( .A1(n10091), .A2(n10090), .A3(n10089), .ZN(n10141) );
  XNOR2_X1 U11178 ( .A(n10092), .B(keyinput62), .ZN(n10097) );
  XNOR2_X1 U11179 ( .A(n10093), .B(keyinput85), .ZN(n10096) );
  XNOR2_X1 U11180 ( .A(n10094), .B(keyinput18), .ZN(n10095) );
  NOR3_X1 U11181 ( .A1(n10097), .A2(n10096), .A3(n10095), .ZN(n10100) );
  XNOR2_X1 U11182 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput6), .ZN(n10099) );
  XNOR2_X1 U11183 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput106), .ZN(n10098) );
  NAND3_X1 U11184 ( .A1(n10100), .A2(n10099), .A3(n10098), .ZN(n10107) );
  AOI22_X1 U11185 ( .A1(n10103), .A2(keyinput102), .B1(n10102), .B2(keyinput99), .ZN(n10101) );
  OAI221_X1 U11186 ( .B1(n10103), .B2(keyinput102), .C1(n10102), .C2(
        keyinput99), .A(n10101), .ZN(n10106) );
  XNOR2_X1 U11187 ( .A(n10104), .B(keyinput3), .ZN(n10105) );
  NOR3_X1 U11188 ( .A1(n10107), .A2(n10106), .A3(n10105), .ZN(n10140) );
  INV_X1 U11189 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U11190 ( .A1(n10110), .A2(keyinput101), .B1(keyinput65), .B2(n10109), .ZN(n10108) );
  OAI221_X1 U11191 ( .B1(n10110), .B2(keyinput101), .C1(n10109), .C2(
        keyinput65), .A(n10108), .ZN(n10122) );
  INV_X1 U11192 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11193 ( .A1(n10112), .A2(keyinput127), .B1(keyinput1), .B2(n5933), 
        .ZN(n10111) );
  OAI221_X1 U11194 ( .B1(n10112), .B2(keyinput127), .C1(n5933), .C2(keyinput1), 
        .A(n10111), .ZN(n10121) );
  AOI22_X1 U11195 ( .A1(n10115), .A2(keyinput92), .B1(n10114), .B2(keyinput88), 
        .ZN(n10113) );
  OAI221_X1 U11196 ( .B1(n10115), .B2(keyinput92), .C1(n10114), .C2(keyinput88), .A(n10113), .ZN(n10120) );
  INV_X1 U11197 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10116) );
  XOR2_X1 U11198 ( .A(n10116), .B(keyinput79), .Z(n10118) );
  XNOR2_X1 U11199 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput12), .ZN(n10117) );
  NAND2_X1 U11200 ( .A1(n10118), .A2(n10117), .ZN(n10119) );
  NOR4_X1 U11201 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10139) );
  AOI22_X1 U11202 ( .A1(n10125), .A2(keyinput36), .B1(keyinput63), .B2(n10124), 
        .ZN(n10123) );
  OAI221_X1 U11203 ( .B1(n10125), .B2(keyinput36), .C1(n10124), .C2(keyinput63), .A(n10123), .ZN(n10137) );
  AOI22_X1 U11204 ( .A1(n10128), .A2(keyinput59), .B1(keyinput13), .B2(n10127), 
        .ZN(n10126) );
  OAI221_X1 U11205 ( .B1(n10128), .B2(keyinput59), .C1(n10127), .C2(keyinput13), .A(n10126), .ZN(n10136) );
  AOI22_X1 U11206 ( .A1(n10131), .A2(keyinput75), .B1(n10130), .B2(keyinput93), 
        .ZN(n10129) );
  OAI221_X1 U11207 ( .B1(n10131), .B2(keyinput75), .C1(n10130), .C2(keyinput93), .A(n10129), .ZN(n10135) );
  XNOR2_X1 U11208 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput4), .ZN(n10133) );
  XNOR2_X1 U11209 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput23), .ZN(n10132)
         );
  NAND2_X1 U11210 ( .A1(n10133), .A2(n10132), .ZN(n10134) );
  NOR4_X1 U11211 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  NAND4_X1 U11212 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10271) );
  AOI22_X1 U11213 ( .A1(n10143), .A2(keyinput8), .B1(keyinput0), .B2(n5974), 
        .ZN(n10142) );
  OAI221_X1 U11214 ( .B1(n10143), .B2(keyinput8), .C1(n5974), .C2(keyinput0), 
        .A(n10142), .ZN(n10155) );
  AOI22_X1 U11215 ( .A1(n10146), .A2(keyinput110), .B1(keyinput29), .B2(n10145), .ZN(n10144) );
  OAI221_X1 U11216 ( .B1(n10146), .B2(keyinput110), .C1(n10145), .C2(
        keyinput29), .A(n10144), .ZN(n10154) );
  AOI22_X1 U11217 ( .A1(n5971), .A2(keyinput33), .B1(keyinput16), .B2(n10148), 
        .ZN(n10147) );
  OAI221_X1 U11218 ( .B1(n5971), .B2(keyinput33), .C1(n10148), .C2(keyinput16), 
        .A(n10147), .ZN(n10153) );
  INV_X1 U11219 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10149) );
  XOR2_X1 U11220 ( .A(n10149), .B(keyinput97), .Z(n10151) );
  XNOR2_X1 U11221 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput53), .ZN(n10150) );
  NAND2_X1 U11222 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  NOR4_X1 U11223 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10203) );
  AOI22_X1 U11224 ( .A1(n10158), .A2(keyinput77), .B1(n10157), .B2(keyinput17), 
        .ZN(n10156) );
  OAI221_X1 U11225 ( .B1(n10158), .B2(keyinput77), .C1(n10157), .C2(keyinput17), .A(n10156), .ZN(n10169) );
  AOI22_X1 U11226 ( .A1(n6164), .A2(keyinput116), .B1(n10160), .B2(keyinput55), 
        .ZN(n10159) );
  OAI221_X1 U11227 ( .B1(n6164), .B2(keyinput116), .C1(n10160), .C2(keyinput55), .A(n10159), .ZN(n10168) );
  INV_X1 U11228 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U11229 ( .A1(n10163), .A2(keyinput125), .B1(keyinput38), .B2(n10162), .ZN(n10161) );
  OAI221_X1 U11230 ( .B1(n10163), .B2(keyinput125), .C1(n10162), .C2(
        keyinput38), .A(n10161), .ZN(n10167) );
  XNOR2_X1 U11231 ( .A(P1_REG2_REG_23__SCAN_IN), .B(keyinput50), .ZN(n10165)
         );
  XNOR2_X1 U11232 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput61), .ZN(n10164) );
  NAND2_X1 U11233 ( .A1(n10165), .A2(n10164), .ZN(n10166) );
  NOR4_X1 U11234 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10202) );
  AOI22_X1 U11235 ( .A1(n10172), .A2(keyinput87), .B1(keyinput109), .B2(n10171), .ZN(n10170) );
  OAI221_X1 U11236 ( .B1(n10172), .B2(keyinput87), .C1(n10171), .C2(
        keyinput109), .A(n10170), .ZN(n10183) );
  INV_X1 U11237 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U11238 ( .A1(n10175), .A2(keyinput5), .B1(n10174), .B2(keyinput69), 
        .ZN(n10173) );
  OAI221_X1 U11239 ( .B1(n10175), .B2(keyinput5), .C1(n10174), .C2(keyinput69), 
        .A(n10173), .ZN(n10182) );
  XOR2_X1 U11240 ( .A(n10176), .B(keyinput30), .Z(n10180) );
  XNOR2_X1 U11241 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput113), .ZN(n10179) );
  XNOR2_X1 U11242 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput82), .ZN(n10178)
         );
  XNOR2_X1 U11243 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(keyinput10), .ZN(n10177)
         );
  NAND4_X1 U11244 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10181) );
  NOR3_X1 U11245 ( .A1(n10183), .A2(n10182), .A3(n10181), .ZN(n10201) );
  AOI22_X1 U11246 ( .A1(n10186), .A2(keyinput40), .B1(keyinput31), .B2(n10185), 
        .ZN(n10184) );
  OAI221_X1 U11247 ( .B1(n10186), .B2(keyinput40), .C1(n10185), .C2(keyinput31), .A(n10184), .ZN(n10199) );
  AOI22_X1 U11248 ( .A1(n10189), .A2(keyinput123), .B1(n10188), .B2(keyinput28), .ZN(n10187) );
  OAI221_X1 U11249 ( .B1(n10189), .B2(keyinput123), .C1(n10188), .C2(
        keyinput28), .A(n10187), .ZN(n10198) );
  INV_X1 U11250 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U11251 ( .A1(n10192), .A2(keyinput51), .B1(keyinput54), .B2(n10191), 
        .ZN(n10190) );
  OAI221_X1 U11252 ( .B1(n10192), .B2(keyinput51), .C1(n10191), .C2(keyinput54), .A(n10190), .ZN(n10197) );
  AOI22_X1 U11253 ( .A1(n10195), .A2(keyinput120), .B1(n10194), .B2(keyinput90), .ZN(n10193) );
  OAI221_X1 U11254 ( .B1(n10195), .B2(keyinput120), .C1(n10194), .C2(
        keyinput90), .A(n10193), .ZN(n10196) );
  NOR4_X1 U11255 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  NAND4_X1 U11256 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10270) );
  AOI22_X1 U11257 ( .A1(n10206), .A2(keyinput105), .B1(keyinput91), .B2(n10205), .ZN(n10204) );
  OAI221_X1 U11258 ( .B1(n10206), .B2(keyinput105), .C1(n10205), .C2(
        keyinput91), .A(n10204), .ZN(n10219) );
  AOI22_X1 U11259 ( .A1(n10209), .A2(keyinput48), .B1(n10208), .B2(keyinput78), 
        .ZN(n10207) );
  OAI221_X1 U11260 ( .B1(n10209), .B2(keyinput48), .C1(n10208), .C2(keyinput78), .A(n10207), .ZN(n10218) );
  INV_X1 U11261 ( .A(SI_7_), .ZN(n10212) );
  AOI22_X1 U11262 ( .A1(n10212), .A2(keyinput119), .B1(keyinput122), .B2(
        n10211), .ZN(n10210) );
  OAI221_X1 U11263 ( .B1(n10212), .B2(keyinput119), .C1(n10211), .C2(
        keyinput122), .A(n10210), .ZN(n10217) );
  XOR2_X1 U11264 ( .A(n10213), .B(keyinput121), .Z(n10215) );
  XNOR2_X1 U11265 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput46), .ZN(n10214) );
  NAND2_X1 U11266 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  NOR4_X1 U11267 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10268) );
  AOI22_X1 U11268 ( .A1(n10222), .A2(keyinput9), .B1(keyinput108), .B2(n10221), 
        .ZN(n10220) );
  OAI221_X1 U11269 ( .B1(n10222), .B2(keyinput9), .C1(n10221), .C2(keyinput108), .A(n10220), .ZN(n10235) );
  AOI22_X1 U11270 ( .A1(n10225), .A2(keyinput34), .B1(n10224), .B2(keyinput103), .ZN(n10223) );
  OAI221_X1 U11271 ( .B1(n10225), .B2(keyinput34), .C1(n10224), .C2(
        keyinput103), .A(n10223), .ZN(n10234) );
  AOI22_X1 U11272 ( .A1(n10228), .A2(keyinput117), .B1(keyinput32), .B2(n10227), .ZN(n10226) );
  OAI221_X1 U11273 ( .B1(n10228), .B2(keyinput117), .C1(n10227), .C2(
        keyinput32), .A(n10226), .ZN(n10233) );
  AOI22_X1 U11274 ( .A1(n10231), .A2(keyinput67), .B1(keyinput39), .B2(n10230), 
        .ZN(n10229) );
  OAI221_X1 U11275 ( .B1(n10231), .B2(keyinput67), .C1(n10230), .C2(keyinput39), .A(n10229), .ZN(n10232) );
  NOR4_X1 U11276 ( .A1(n10235), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10267) );
  AOI22_X1 U11277 ( .A1(n10238), .A2(keyinput74), .B1(n10237), .B2(keyinput72), 
        .ZN(n10236) );
  OAI221_X1 U11278 ( .B1(n10238), .B2(keyinput74), .C1(n10237), .C2(keyinput72), .A(n10236), .ZN(n10249) );
  AOI22_X1 U11279 ( .A1(n10241), .A2(keyinput41), .B1(keyinput26), .B2(n10240), 
        .ZN(n10239) );
  OAI221_X1 U11280 ( .B1(n10241), .B2(keyinput41), .C1(n10240), .C2(keyinput26), .A(n10239), .ZN(n10248) );
  XNOR2_X1 U11281 ( .A(n10242), .B(keyinput76), .ZN(n10247) );
  XOR2_X1 U11282 ( .A(n6977), .B(keyinput114), .Z(n10245) );
  XNOR2_X1 U11283 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput94), .ZN(n10244) );
  XNOR2_X1 U11284 ( .A(SI_3_), .B(keyinput56), .ZN(n10243) );
  NAND3_X1 U11285 ( .A1(n10245), .A2(n10244), .A3(n10243), .ZN(n10246) );
  NOR4_X1 U11286 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10266) );
  AOI22_X1 U11287 ( .A1(n10252), .A2(keyinput73), .B1(n10251), .B2(keyinput86), 
        .ZN(n10250) );
  OAI221_X1 U11288 ( .B1(n10252), .B2(keyinput73), .C1(n10251), .C2(keyinput86), .A(n10250), .ZN(n10264) );
  INV_X1 U11289 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U11290 ( .A1(n10255), .A2(keyinput124), .B1(keyinput95), .B2(n10254), .ZN(n10253) );
  OAI221_X1 U11291 ( .B1(n10255), .B2(keyinput124), .C1(n10254), .C2(
        keyinput95), .A(n10253), .ZN(n10263) );
  AOI22_X1 U11292 ( .A1(n10258), .A2(keyinput11), .B1(n10257), .B2(keyinput2), 
        .ZN(n10256) );
  OAI221_X1 U11293 ( .B1(n10258), .B2(keyinput11), .C1(n10257), .C2(keyinput2), 
        .A(n10256), .ZN(n10262) );
  XNOR2_X1 U11294 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput49), .ZN(n10260) );
  XNOR2_X1 U11295 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput21), .ZN(n10259)
         );
  NAND2_X1 U11296 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  NOR4_X1 U11297 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10265) );
  NAND4_X1 U11298 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10269) );
  NOR4_X1 U11299 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10277) );
  AOI21_X1 U11300 ( .B1(n10275), .B2(n10274), .A(n10273), .ZN(n10276) );
  XOR2_X1 U11301 ( .A(n10277), .B(n10276), .Z(n10278) );
  XNOR2_X1 U11302 ( .A(n10279), .B(n10278), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11303 ( .A(n10281), .B(n10280), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11304 ( .A(n10283), .B(n10282), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11305 ( .A(n10285), .B(n10284), .ZN(ADD_1068_U49) );
  XOR2_X1 U11306 ( .A(n10287), .B(n10286), .Z(ADD_1068_U54) );
  XOR2_X1 U11307 ( .A(n10289), .B(n10288), .Z(ADD_1068_U53) );
  XNOR2_X1 U11308 ( .A(n10291), .B(n10290), .ZN(ADD_1068_U52) );
  XNOR2_X1 U6572 ( .A(n5078), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5739) );
  INV_X1 U4911 ( .A(n5869), .ZN(n7894) );
  NAND4_X1 U4922 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n8991)
         );
  CLKBUF_X1 U4914 ( .A(n5719), .Z(n4530) );
  CLKBUF_X1 U5248 ( .A(n5868), .Z(n6109) );
  CLKBUF_X1 U5867 ( .A(n8730), .Z(n8733) );
endmodule

