

module b15_C_gen_AntiSAT_k_256_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123;

  AOI211_X1 U3605 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5972), .A(n5529), .B(n5528), .ZN(n5530) );
  AOI21_X1 U3606 ( .B1(n4453), .B2(n5523), .A(n4457), .ZN(n4229) );
  INV_X2 U3607 ( .A(n4260), .ZN(n5719) );
  NAND2_X1 U3608 ( .A1(n3506), .A2(n3505), .ZN(n4089) );
  AND2_X1 U3609 ( .A1(n4133), .A2(n4177), .ZN(n4386) );
  INV_X2 U3610 ( .A(n4481), .ZN(n4374) );
  INV_X2 U3611 ( .A(n5537), .ZN(n4133) );
  CLKBUF_X2 U3612 ( .A(n3441), .Z(n4024) );
  CLKBUF_X2 U3613 ( .A(n3428), .Z(n3994) );
  CLKBUF_X2 U3614 ( .A(n3315), .Z(n3157) );
  NOR2_X2 U3615 ( .A1(n4384), .A2(n4361), .ZN(n5493) );
  NOR2_X1 U3616 ( .A1(n4387), .A2(n4270), .ZN(n4357) );
  CLKBUF_X1 U3617 ( .A(n3331), .Z(n4661) );
  OR2_X1 U3618 ( .A1(n3266), .A2(n3265), .ZN(n4264) );
  CLKBUF_X2 U3619 ( .A(n3328), .Z(n4270) );
  AND2_X1 U3620 ( .A1(n3225), .A2(n3224), .ZN(n3159) );
  NAND2_X1 U3621 ( .A1(n3275), .A2(n3173), .ZN(n4385) );
  AND4_X1 U3622 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3215)
         );
  AND2_X2 U3623 ( .A1(n4543), .A2(n3209), .ZN(n3388) );
  INV_X1 U3624 ( .A(n6310), .ZN(n6317) );
  OAI21_X1 U3625 ( .B1(n4101), .B2(n3364), .A(n3345), .ZN(n3326) );
  AND2_X1 U3626 ( .A1(n4420), .A2(n3456), .ZN(n3349) );
  NAND2_X1 U3627 ( .A1(n4264), .A2(n3332), .ZN(n4387) );
  NAND2_X1 U3628 ( .A1(n3225), .A2(n3224), .ZN(n3327) );
  AND4_X1 U3629 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3293)
         );
  NAND2_X1 U3630 ( .A1(n4133), .A2(n4481), .ZN(n4217) );
  NAND2_X1 U3631 ( .A1(n4226), .A2(n4225), .ZN(n5523) );
  NAND2_X1 U3632 ( .A1(n3195), .A2(n4131), .ZN(n4590) );
  INV_X1 U3633 ( .A(n4361), .ZN(n4688) );
  INV_X1 U3634 ( .A(n4264), .ZN(n4679) );
  INV_X1 U3635 ( .A(n4008), .ZN(n4106) );
  NAND2_X1 U3636 ( .A1(n6352), .A2(n4462), .ZN(n6717) );
  INV_X1 U3637 ( .A(n3316), .ZN(n3394) );
  NOR4_X2 U3638 ( .A1(n6693), .A2(n6698), .A3(n6696), .A4(n6001), .ZN(n5981)
         );
  NAND2_X2 U3639 ( .A1(n5743), .A2(n4343), .ZN(n5736) );
  NAND2_X2 U3640 ( .A1(n5742), .A2(n5744), .ZN(n5743) );
  OAI21_X2 U3641 ( .B1(n5642), .B2(n4434), .A(n4433), .ZN(n4435) );
  CLKBUF_X1 U3643 ( .A(n5514), .Z(n5560) );
  NAND2_X1 U3644 ( .A1(n3170), .A2(n3925), .ZN(n5426) );
  AND2_X1 U3645 ( .A1(n3925), .A2(n3924), .ZN(n5424) );
  OAI21_X1 U3646 ( .B1(n5736), .B2(n3181), .A(n3178), .ZN(n5707) );
  OR2_X1 U3647 ( .A1(n4243), .A2(n6026), .ZN(n6001) );
  INV_X2 U3648 ( .A(n6278), .ZN(n6264) );
  XNOR2_X1 U3649 ( .A(n3409), .B(n3408), .ZN(n4647) );
  NAND2_X1 U3651 ( .A1(n4102), .A2(n3330), .ZN(n4534) );
  AND2_X1 U3652 ( .A1(n4506), .A2(n4507), .ZN(n3195) );
  INV_X2 U3653 ( .A(n4688), .ZN(n5497) );
  AND4_X1 U3654 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  AND4_X1 U3655 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3294)
         );
  AND4_X1 U3656 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(n3214)
         );
  BUF_X2 U3657 ( .A(n3393), .Z(n3948) );
  CLKBUF_X2 U3658 ( .A(n3297), .Z(n4014) );
  CLKBUF_X2 U3659 ( .A(n3421), .Z(n4012) );
  BUF_X2 U3660 ( .A(n3388), .Z(n4540) );
  BUF_X2 U3661 ( .A(n3423), .Z(n4022) );
  NOR2_X4 U3662 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4544) );
  XNOR2_X1 U3663 ( .A(n5682), .B(n5665), .ZN(n5794) );
  NAND2_X1 U3664 ( .A1(n5664), .A2(n5687), .ZN(n5681) );
  AND2_X1 U3665 ( .A1(n5561), .A2(n5560), .ZN(n5976) );
  NAND3_X2 U3666 ( .A1(n4354), .A2(n3200), .A3(n4353), .ZN(n4431) );
  INV_X1 U3667 ( .A(n5569), .ZN(n3925) );
  NOR2_X1 U3668 ( .A1(n5572), .A2(n5573), .ZN(n4210) );
  AND2_X1 U3669 ( .A1(n3165), .A2(n3166), .ZN(n5389) );
  NAND2_X1 U3670 ( .A1(n3698), .A2(n3697), .ZN(n5316) );
  NAND2_X1 U3671 ( .A1(n4321), .A2(n4320), .ZN(n5228) );
  NOR2_X1 U3672 ( .A1(n5584), .A2(n5585), .ZN(n4199) );
  AND2_X1 U3673 ( .A1(n3186), .A2(n5760), .ZN(n3185) );
  OR2_X1 U3674 ( .A1(n3187), .A2(n5334), .ZN(n3186) );
  NOR2_X1 U3675 ( .A1(n5539), .A2(n5611), .ZN(n4187) );
  CLKBUF_X1 U3676 ( .A(n5539), .Z(n5551) );
  AND2_X1 U3677 ( .A1(n5143), .A2(n3196), .ZN(n3678) );
  XNOR2_X1 U3678 ( .A(n4338), .B(n4337), .ZN(n5159) );
  NOR2_X1 U3679 ( .A1(n4503), .A2(n4588), .ZN(n4586) );
  NOR2_X1 U3680 ( .A1(n5425), .A2(n5571), .ZN(n3170) );
  AOI21_X1 U3681 ( .B1(n4323), .B2(n3712), .A(n3598), .ZN(n4890) );
  NAND2_X1 U3682 ( .A1(n3495), .A2(n3494), .ZN(n4488) );
  CLKBUF_X1 U3683 ( .A(n4972), .Z(n5966) );
  XNOR2_X1 U3684 ( .A(n4314), .B(n3591), .ZN(n4323) );
  NAND2_X1 U3685 ( .A1(n3162), .A2(n3488), .ZN(n4489) );
  AND2_X1 U3686 ( .A1(n3464), .A2(n3702), .ZN(n3162) );
  NAND2_X1 U3687 ( .A1(n6717), .A2(n4238), .ZN(n6278) );
  NAND2_X1 U3688 ( .A1(n3519), .A2(n3518), .ZN(n4720) );
  NAND2_X2 U3689 ( .A1(n6351), .A2(n4436), .ZN(n6161) );
  NAND2_X1 U3690 ( .A1(n6351), .A2(n4094), .ZN(n6352) );
  INV_X2 U3691 ( .A(n4469), .ZN(n6351) );
  XNOR2_X1 U3692 ( .A(n3468), .B(n3467), .ZN(n4572) );
  OR2_X2 U3693 ( .A1(n5495), .A2(n6642), .ZN(n4469) );
  XNOR2_X1 U3694 ( .A(n3466), .B(n3465), .ZN(n3468) );
  NAND2_X1 U3695 ( .A1(n3477), .A2(n3460), .ZN(n3467) );
  OAI21_X2 U3696 ( .B1(n4647), .B2(STATE2_REG_0__SCAN_IN), .A(n3420), .ZN(
        n3466) );
  NAND2_X1 U3697 ( .A1(n4146), .A2(n4145), .ZN(n4893) );
  XNOR2_X1 U3698 ( .A(n3440), .B(n3439), .ZN(n3480) );
  NAND3_X1 U3699 ( .A1(n3356), .A2(n3355), .A3(n3354), .ZN(n3377) );
  NAND2_X1 U3700 ( .A1(n3358), .A2(n3357), .ZN(n3439) );
  OAI22_X1 U3701 ( .A1(n4080), .A2(n4066), .B1(n4075), .B2(n4074), .ZN(n4071)
         );
  AND2_X1 U3702 ( .A1(n3343), .A2(n3342), .ZN(n3359) );
  AND2_X1 U3703 ( .A1(n4389), .A2(n4064), .ZN(n4102) );
  AOI21_X1 U3704 ( .B1(n3340), .B2(n4661), .A(n4387), .ZN(n3344) );
  CLKBUF_X1 U3705 ( .A(n4232), .Z(n6354) );
  NOR2_X1 U3706 ( .A1(n4360), .A2(n4361), .ZN(n4389) );
  OR2_X1 U3707 ( .A1(n3366), .A2(n3365), .ZN(n4553) );
  AND2_X1 U3708 ( .A1(n3363), .A2(n4449), .ZN(n4103) );
  AND2_X1 U3709 ( .A1(n3456), .A2(n4270), .ZN(n4064) );
  NAND2_X1 U3710 ( .A1(n3327), .A2(n4449), .ZN(n4360) );
  CLKBUF_X1 U3711 ( .A(n3158), .Z(n4425) );
  CLKBUF_X1 U3712 ( .A(n3456), .Z(n4666) );
  AND2_X1 U3714 ( .A1(n3159), .A2(n3328), .ZN(n3360) );
  CLKBUF_X1 U3715 ( .A(n3341), .Z(n3361) );
  INV_X1 U3716 ( .A(n3341), .ZN(n3456) );
  NAND4_X1 U3717 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3341)
         );
  AND4_X1 U3718 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3322)
         );
  AND4_X1 U3719 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  AND4_X1 U3720 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3324)
         );
  AND4_X1 U3721 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3295)
         );
  AND4_X1 U3722 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3323)
         );
  AND4_X1 U3723 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3173)
         );
  AND4_X1 U3724 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3275)
         );
  AND4_X1 U3725 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3244)
         );
  AND4_X1 U3726 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3245)
         );
  AND4_X1 U3727 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n3225)
         );
  AND4_X1 U3728 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3224)
         );
  AND4_X1 U3729 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3246)
         );
  AND4_X1 U3730 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3243)
         );
  NAND2_X2 U3731 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6716), .ZN(n6701) );
  NAND2_X2 U3732 ( .A1(n6716), .A2(n6671), .ZN(n6691) );
  OR2_X1 U3733 ( .A1(n3394), .A2(n3238), .ZN(n3240) );
  BUF_X2 U3734 ( .A(n3303), .Z(n4020) );
  BUF_X2 U3735 ( .A(n3422), .Z(n4023) );
  BUF_X2 U3736 ( .A(n3446), .Z(n4015) );
  BUF_X2 U3737 ( .A(n3304), .Z(n3989) );
  BUF_X2 U3738 ( .A(n3309), .Z(n4011) );
  AND2_X2 U3739 ( .A1(n4654), .A2(n4608), .ZN(n6719) );
  BUF_X2 U3740 ( .A(n3310), .Z(n4013) );
  AND2_X1 U3741 ( .A1(n3203), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3208)
         );
  NOR2_X2 U3742 ( .A1(n6845), .A2(n5547), .ZN(n6054) );
  NAND2_X1 U3743 ( .A1(n3159), .A2(n3328), .ZN(n3158) );
  CLKBUF_X1 U3744 ( .A(n4638), .Z(n3160) );
  OAI21_X1 U3745 ( .B1(n5736), .B2(n3181), .A(n3178), .ZN(n3161) );
  NOR2_X2 U3746 ( .A1(n5796), .A2(n5795), .ZN(n5579) );
  NAND2_X1 U3747 ( .A1(n4163), .A2(n4162), .ZN(n5297) );
  INV_X2 U3748 ( .A(n4505), .ZN(n4131) );
  BUF_X4 U3749 ( .A(n4112), .Z(n5537) );
  AND2_X2 U3750 ( .A1(n4264), .A2(n4384), .ZN(n4112) );
  NAND2_X1 U3751 ( .A1(n4293), .A2(n4292), .ZN(n4642) );
  NAND2_X2 U3752 ( .A1(n4431), .A2(n4355), .ZN(n5649) );
  OAI21_X2 U3753 ( .B1(n5332), .B2(n3187), .A(n3185), .ZN(n5749) );
  NAND2_X2 U3754 ( .A1(n3549), .A2(n3522), .ZN(n4290) );
  INV_X1 U3755 ( .A(n5610), .ZN(n3163) );
  NOR2_X2 U3756 ( .A1(n5531), .A2(n3164), .ZN(n5601) );
  NAND2_X1 U3757 ( .A1(n3783), .A2(n3163), .ZN(n3164) );
  NAND2_X1 U3758 ( .A1(n3698), .A2(n3697), .ZN(n3165) );
  AND2_X1 U3759 ( .A1(n3167), .A2(n5318), .ZN(n3166) );
  INV_X1 U3760 ( .A(n5396), .ZN(n3167) );
  NAND2_X1 U3761 ( .A1(n3925), .A2(n3924), .ZN(n3168) );
  NOR2_X2 U3762 ( .A1(n3168), .A2(n3169), .ZN(n5437) );
  OR2_X1 U3763 ( .A1(n5438), .A2(n5425), .ZN(n3169) );
  XNOR2_X1 U3764 ( .A(n3520), .B(n3463), .ZN(n3171) );
  XNOR2_X1 U3765 ( .A(n3520), .B(n3463), .ZN(n4262) );
  INV_X4 U3766 ( .A(n4385), .ZN(n3332) );
  OR2_X1 U3767 ( .A1(n3379), .A2(n5478), .ZN(n3358) );
  NAND3_X1 U3768 ( .A1(n3520), .A2(n3496), .A3(n4720), .ZN(n3549) );
  NAND2_X2 U3769 ( .A1(n3477), .A2(n3476), .ZN(n5077) );
  AND2_X2 U3770 ( .A1(n5894), .A2(n4546), .ZN(n3309) );
  CLKBUF_X2 U3771 ( .A(n3302), .Z(n4021) );
  INV_X1 U3772 ( .A(n3549), .ZN(n3194) );
  NAND2_X1 U3773 ( .A1(n3194), .A2(n3192), .ZN(n3581) );
  AND2_X1 U3774 ( .A1(n3193), .A2(n3550), .ZN(n3192) );
  INV_X1 U3775 ( .A(n3563), .ZN(n3193) );
  AND2_X1 U3776 ( .A1(n3580), .A2(n3579), .ZN(n3587) );
  NAND2_X1 U3777 ( .A1(n5437), .A2(n5559), .ZN(n5514) );
  NAND2_X1 U3778 ( .A1(n6351), .A2(n4517), .ZN(n6355) );
  AOI22_X1 U3779 ( .A1(n4038), .A2(n4037), .B1(n5505), .B2(n4106), .ZN(n4416)
         );
  AND2_X1 U3780 ( .A1(n4403), .A2(n6604), .ZN(n5863) );
  AND2_X1 U3781 ( .A1(n4403), .A2(n4399), .ZN(n5865) );
  INV_X1 U3782 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6619) );
  AND2_X2 U3783 ( .A1(n4543), .A2(n4544), .ZN(n3428) );
  AND2_X1 U3784 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  OR2_X1 U3785 ( .A1(n3400), .A2(n3399), .ZN(n3403) );
  OR2_X1 U3786 ( .A1(n3361), .A2(n4654), .ZN(n3506) );
  AND2_X2 U3787 ( .A1(n3500), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3209)
         );
  AOI21_X1 U3788 ( .B1(n3349), .B2(n3478), .A(n3332), .ZN(n3350) );
  NOR2_X1 U3789 ( .A1(n6603), .A2(n4654), .ZN(n4033) );
  NOR2_X1 U3790 ( .A1(n3327), .A2(n5115), .ZN(n3712) );
  INV_X1 U3791 ( .A(n4345), .ZN(n3183) );
  INV_X1 U3792 ( .A(n4344), .ZN(n3180) );
  INV_X1 U3793 ( .A(n5729), .ZN(n3179) );
  INV_X1 U3794 ( .A(n4217), .ZN(n4200) );
  INV_X1 U3795 ( .A(n4339), .ZN(n3190) );
  INV_X1 U3796 ( .A(n3587), .ZN(n3588) );
  INV_X1 U3797 ( .A(n3581), .ZN(n3589) );
  INV_X1 U3798 ( .A(n4211), .ZN(n5536) );
  CLKBUF_X1 U3799 ( .A(n4132), .Z(n4211) );
  NAND2_X1 U3800 ( .A1(n5537), .A2(n4481), .ZN(n4123) );
  NAND2_X2 U3801 ( .A1(n4270), .A2(n4384), .ZN(n4308) );
  INV_X1 U3802 ( .A(n3506), .ZN(n4258) );
  OR2_X1 U3803 ( .A1(n3434), .A2(n3433), .ZN(n4334) );
  OR2_X1 U3804 ( .A1(n3379), .A2(n3380), .ZN(n3387) );
  OR2_X1 U3805 ( .A1(n5497), .A2(n4654), .ZN(n3505) );
  NAND3_X1 U3806 ( .A1(n3361), .A2(n5497), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4078) );
  NOR2_X1 U3807 ( .A1(n4078), .A2(n4308), .ZN(n4069) );
  NAND2_X1 U3808 ( .A1(n5115), .A2(n7092), .ZN(n4008) );
  NAND2_X1 U3809 ( .A1(n4105), .A2(n4104), .ZN(n4462) );
  INV_X1 U3810 ( .A(n3702), .ZN(n4039) );
  NOR2_X1 U3811 ( .A1(n3985), .A2(n5654), .ZN(n3986) );
  AND2_X1 U3812 ( .A1(n5143), .A2(n5142), .ZN(n5209) );
  NAND2_X1 U3813 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3523) );
  AND2_X1 U3814 ( .A1(n4404), .A2(n6489), .ZN(n5829) );
  NAND2_X1 U3815 ( .A1(n3188), .A2(n5759), .ZN(n3187) );
  INV_X1 U3816 ( .A(n5287), .ZN(n4157) );
  OAI21_X1 U3817 ( .B1(n4469), .B2(n4373), .A(n4372), .ZN(n4403) );
  AND2_X1 U3818 ( .A1(n5352), .A2(n5917), .ZN(n5359) );
  CLKBUF_X1 U3819 ( .A(n4529), .Z(n4530) );
  OR2_X1 U3820 ( .A1(n4533), .A2(n6720), .ZN(n6632) );
  AND2_X1 U3821 ( .A1(n6232), .A2(n5177), .ZN(n6250) );
  AND2_X1 U3822 ( .A1(n5176), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5177) );
  AND2_X1 U3823 ( .A1(n4448), .A2(n6645), .ZN(n6322) );
  OAI21_X1 U3824 ( .B1(n4514), .B2(n4422), .A(n6645), .ZN(n4424) );
  CLKBUF_X2 U3825 ( .A(n6433), .Z(n6423) );
  INV_X1 U3826 ( .A(n4416), .ZN(n4417) );
  INV_X1 U3827 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6606) );
  CLKBUF_X1 U3828 ( .A(n4572), .Z(n4573) );
  CLKBUF_X1 U3829 ( .A(n3171), .Z(n4571) );
  AND2_X1 U3830 ( .A1(n6628), .A2(n6627), .ZN(n6643) );
  INV_X1 U3831 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4043) );
  AND2_X1 U3832 ( .A1(n4055), .A2(n4056), .ZN(n4053) );
  AOI22_X1 U3833 ( .A1(n3302), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3205) );
  OR2_X1 U3834 ( .A1(n4060), .A2(n4062), .ZN(n4046) );
  OR2_X1 U3835 ( .A1(n3578), .A2(n3577), .ZN(n4325) );
  OR2_X1 U3836 ( .A1(n3560), .A2(n3559), .ZN(n4305) );
  OR2_X1 U3837 ( .A1(n3538), .A2(n3537), .ZN(n4302) );
  INV_X1 U3838 ( .A(n4123), .ZN(n4132) );
  OR2_X1 U3839 ( .A1(n3419), .A2(n3418), .ZN(n4269) );
  NAND2_X1 U3840 ( .A1(n3316), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3289)
         );
  AOI22_X1 U3841 ( .A1(n3309), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U3842 ( .A1(n3303), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3216) );
  OR2_X1 U3843 ( .A1(n3517), .A2(n3516), .ZN(n4288) );
  INV_X1 U3844 ( .A(n4078), .ZN(n4085) );
  INV_X1 U3845 ( .A(n5534), .ZN(n3783) );
  AND2_X1 U3846 ( .A1(n5146), .A2(n5144), .ZN(n5145) );
  NAND2_X1 U3847 ( .A1(n3581), .A2(n3565), .ZN(n4309) );
  AND2_X1 U3848 ( .A1(n5563), .A2(n5562), .ZN(n4224) );
  NAND2_X1 U3849 ( .A1(n5333), .A2(n5334), .ZN(n3188) );
  INV_X1 U3850 ( .A(n4334), .ZN(n3453) );
  OR2_X1 U3851 ( .A1(n3452), .A2(n3451), .ZN(n4278) );
  NAND2_X1 U3852 ( .A1(n3439), .A2(n3438), .ZN(n3407) );
  AND2_X1 U3853 ( .A1(n3159), .A2(n3341), .ZN(n3364) );
  AND2_X1 U3854 ( .A1(n4395), .A2(n4394), .ZN(n4536) );
  NAND2_X1 U3855 ( .A1(n3499), .A2(n3498), .ZN(n4511) );
  OAI21_X1 U3856 ( .B1(n6723), .B2(n4608), .A(n5902), .ZN(n4655) );
  INV_X1 U3857 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5114) );
  INV_X1 U3858 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4838) );
  AND2_X1 U3859 ( .A1(n4562), .A2(n4561), .ZN(n6615) );
  AND2_X1 U3860 ( .A1(n4536), .A2(n4396), .ZN(n5487) );
  AND2_X1 U3861 ( .A1(n4166), .A2(n4165), .ZN(n5296) );
  NOR2_X1 U3862 ( .A1(n4469), .A2(n4468), .ZN(n6330) );
  AND2_X1 U3863 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3962), .ZN(n3963)
         );
  NAND2_X1 U3864 ( .A1(n3963), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3985)
         );
  AND2_X1 U3865 ( .A1(n3919), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3920)
         );
  CLKBUF_X1 U3866 ( .A(n5569), .Z(n5570) );
  AND2_X1 U3867 ( .A1(n3887), .A2(n3886), .ZN(n5675) );
  NOR2_X1 U3868 ( .A1(n3882), .A2(n5691), .ZN(n3883) );
  AND2_X1 U3869 ( .A1(n3883), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3919)
         );
  CLKBUF_X1 U3870 ( .A(n5588), .Z(n5589) );
  AND2_X1 U3871 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3834), .ZN(n3835)
         );
  INV_X1 U3872 ( .A(n3833), .ZN(n3834) );
  NAND2_X1 U3873 ( .A1(n3835), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3882)
         );
  CLKBUF_X1 U3874 ( .A(n5592), .Z(n5593) );
  NOR2_X1 U3875 ( .A1(n3799), .A2(n5713), .ZN(n3800) );
  CLKBUF_X1 U3876 ( .A(n5601), .Z(n5602) );
  AND2_X1 U3877 ( .A1(n3761), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3762)
         );
  NAND2_X1 U3878 ( .A1(n3762), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3799)
         );
  NOR2_X1 U3879 ( .A1(n3733), .A2(n6186), .ZN(n3761) );
  CLKBUF_X1 U3880 ( .A(n5391), .Z(n5392) );
  NAND2_X1 U3881 ( .A1(n3717), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3733)
         );
  CLKBUF_X1 U3882 ( .A(n5389), .Z(n5390) );
  NOR2_X1 U3883 ( .A1(n3700), .A2(n3699), .ZN(n3717) );
  NAND2_X1 U3884 ( .A1(n3680), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3700)
         );
  INV_X1 U3885 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U3886 ( .A1(n3663), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3630)
         );
  NAND2_X1 U3887 ( .A1(n3614), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3646)
         );
  INV_X1 U3888 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5216) );
  NOR2_X1 U3889 ( .A1(n3593), .A2(n3592), .ZN(n3594) );
  NAND2_X1 U3890 ( .A1(n3594), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3599)
         );
  AOI21_X1 U3891 ( .B1(n4313), .B2(n3712), .A(n3584), .ZN(n4709) );
  CLKBUF_X1 U3892 ( .A(n4707), .Z(n4708) );
  NOR2_X1 U3893 ( .A1(n3545), .A2(n6273), .ZN(n3566) );
  INV_X1 U3894 ( .A(n3523), .ZN(n3524) );
  NAND2_X1 U3895 ( .A1(n3524), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3545)
         );
  OAI211_X1 U3896 ( .C1(n3544), .C2(n3380), .A(n3491), .B(n3490), .ZN(n4490)
         );
  NAND2_X1 U3897 ( .A1(n4285), .A2(n4284), .ZN(n6438) );
  CLKBUF_X1 U3898 ( .A(n5572), .Z(n5582) );
  CLKBUF_X1 U3899 ( .A(n5579), .Z(n5798) );
  AND2_X1 U3900 ( .A1(n4198), .A2(n4197), .ZN(n5585) );
  NOR2_X1 U3901 ( .A1(n6115), .A2(n4401), .ZN(n5806) );
  OAI21_X1 U3902 ( .B1(n5702), .B2(n5703), .A(n5663), .ZN(n5696) );
  AND2_X1 U3903 ( .A1(n4186), .A2(n4185), .ZN(n5611) );
  AND2_X1 U3904 ( .A1(n4183), .A2(n4182), .ZN(n5548) );
  INV_X1 U3905 ( .A(n3182), .ZN(n3181) );
  AOI21_X1 U3906 ( .B1(n3182), .B2(n3180), .A(n3179), .ZN(n3178) );
  NOR2_X1 U3907 ( .A1(n5728), .A2(n3183), .ZN(n3182) );
  AND2_X1 U3908 ( .A1(n4260), .A2(n5848), .ZN(n5728) );
  NAND2_X1 U3909 ( .A1(n5736), .A2(n4344), .ZN(n3184) );
  INV_X1 U3910 ( .A(n5290), .ZN(n4163) );
  AND2_X1 U3911 ( .A1(n4156), .A2(n4155), .ZN(n5287) );
  NAND2_X1 U3912 ( .A1(n3191), .A2(n3189), .ZN(n4341) );
  NOR2_X1 U3913 ( .A1(n3175), .A2(n3190), .ZN(n3189) );
  AND2_X1 U3914 ( .A1(n4153), .A2(n4152), .ZN(n5212) );
  CLKBUF_X1 U3915 ( .A(n5211), .Z(n5288) );
  NAND2_X1 U3916 ( .A1(n5158), .A2(n5159), .ZN(n3191) );
  AND3_X1 U3917 ( .A1(n4322), .A2(n4258), .A3(n4334), .ZN(n4259) );
  XNOR2_X1 U3918 ( .A(n4330), .B(n6480), .ZN(n5229) );
  INV_X1 U3919 ( .A(n4713), .ZN(n4145) );
  INV_X1 U3920 ( .A(n4712), .ZN(n4146) );
  NOR2_X2 U3921 ( .A1(n4590), .A2(n4591), .ZN(n4634) );
  XNOR2_X1 U3922 ( .A(n4299), .B(n4298), .ZN(n4643) );
  NAND2_X1 U3923 ( .A1(n4120), .A2(n4119), .ZN(n4507) );
  NOR2_X1 U3924 ( .A1(n4405), .A2(n6486), .ZN(n5839) );
  NAND2_X1 U3925 ( .A1(n3459), .A2(n3473), .ZN(n3477) );
  OR2_X1 U3926 ( .A1(n4290), .A2(n4571), .ZN(n5112) );
  INV_X1 U3927 ( .A(n3404), .ZN(n3405) );
  INV_X1 U3928 ( .A(n4764), .ZN(n5038) );
  AND2_X2 U3929 ( .A1(n3202), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5893)
         );
  AND2_X2 U3930 ( .A1(n3177), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5894)
         );
  INV_X1 U3931 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3177) );
  OR2_X1 U3932 ( .A1(n4425), .A2(n3742), .ZN(n6603) );
  AND2_X2 U3934 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4546) );
  AND2_X1 U3935 ( .A1(n4786), .A2(n5917), .ZN(n5080) );
  NOR2_X1 U3936 ( .A1(n5112), .A2(n4573), .ZN(n5013) );
  INV_X1 U3937 ( .A(n5077), .ZN(n5012) );
  INV_X2 U3938 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U3939 ( .A1(n5402), .A2(n4655), .ZN(n4689) );
  INV_X1 U3940 ( .A(n5112), .ZN(n5122) );
  NAND2_X1 U3941 ( .A1(n4654), .A2(n4655), .ZN(n4764) );
  AOI21_X1 U3942 ( .B1(n6606), .B2(STATE2_REG_3__SCAN_IN), .A(n4764), .ZN(
        n5244) );
  AND2_X1 U3943 ( .A1(n5472), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4093) );
  INV_X1 U3944 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4654) );
  NOR2_X1 U3945 ( .A1(n5472), .A2(n5115), .ZN(n4608) );
  OR2_X1 U3946 ( .A1(n6656), .A2(n3325), .ZN(n4233) );
  OR2_X1 U3947 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  AND2_X1 U3948 ( .A1(n6025), .A2(n4245), .ZN(n5992) );
  INV_X1 U3949 ( .A(n6236), .ZN(n6252) );
  AND2_X1 U3950 ( .A1(n6232), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6245) );
  CLKBUF_X1 U3951 ( .A(n4479), .Z(n5308) );
  AND2_X1 U3952 ( .A1(n6717), .A2(n4231), .ZN(n6297) );
  INV_X1 U3953 ( .A(n6295), .ZN(n6246) );
  INV_X1 U3954 ( .A(n6322), .ZN(n5613) );
  INV_X1 U3955 ( .A(n5464), .ZN(n5513) );
  INV_X1 U3956 ( .A(n6021), .ZN(n6067) );
  INV_X1 U3957 ( .A(n5481), .ZN(n6326) );
  AND2_X1 U3958 ( .A1(n5481), .A2(n4426), .ZN(n6323) );
  NAND2_X1 U3959 ( .A1(n5481), .A2(n4594), .ZN(n5398) );
  BUF_X1 U3960 ( .A(n6347), .Z(n6344) );
  OAI21_X1 U3961 ( .B1(n6354), .B2(n6828), .A(n6353), .ZN(n6433) );
  INV_X1 U3962 ( .A(n6355), .ZN(n6432) );
  XNOR2_X1 U3963 ( .A(n4110), .B(n4109), .ZN(n5176) );
  OR2_X1 U3964 ( .A1(n4108), .A2(n5465), .ZN(n4110) );
  INV_X1 U3965 ( .A(n4040), .ZN(n4041) );
  INV_X1 U3966 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5713) );
  AND2_X1 U3967 ( .A1(n5286), .A2(n5285), .ZN(n6227) );
  INV_X1 U3968 ( .A(n6100), .ZN(n6448) );
  INV_X1 U3969 ( .A(n6161), .ZN(n6450) );
  NOR3_X1 U3970 ( .A1(n5711), .A2(n5843), .A3(n5847), .ZN(n6124) );
  NAND2_X1 U3971 ( .A1(n5838), .A2(n6458), .ZN(n5847) );
  INV_X1 U3972 ( .A(n6148), .ZN(n6458) );
  BUF_X1 U3973 ( .A(n6259), .Z(n6120) );
  NAND2_X1 U3974 ( .A1(n6495), .A2(n4400), .ZN(n6489) );
  INV_X1 U3975 ( .A(n5839), .ZN(n6497) );
  INV_X1 U3976 ( .A(n5863), .ZN(n6495) );
  CLKBUF_X1 U3977 ( .A(n4647), .Z(n4648) );
  CLKBUF_X1 U3978 ( .A(n4551), .Z(n4552) );
  INV_X1 U3979 ( .A(n5917), .ZN(n6517) );
  INV_X1 U3980 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5472) );
  INV_X1 U3981 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5478) );
  NOR2_X1 U3982 ( .A1(n5471), .A2(n5495), .ZN(n6635) );
  INV_X1 U3983 ( .A(n6635), .ZN(n5902) );
  NOR2_X1 U3984 ( .A1(n5402), .A2(n6151), .ZN(n6149) );
  INV_X1 U3985 ( .A(n6579), .ZN(n4924) );
  AOI22_X1 U3986 ( .A1(n5359), .A2(n5356), .B1(n6510), .B2(n5353), .ZN(n5388)
         );
  NOR2_X1 U3987 ( .A1(n4689), .A2(n3332), .ZN(n6570) );
  NOR2_X1 U3988 ( .A1(n4689), .A2(n5480), .ZN(n6561) );
  NAND2_X1 U3989 ( .A1(n5122), .A2(n5121), .ZN(n6601) );
  INV_X1 U3990 ( .A(n6596), .ZN(n5141) );
  NOR2_X1 U3991 ( .A1(n7063), .A2(n4764), .ZN(n6514) );
  NOR2_X1 U3992 ( .A1(n4827), .A2(n4764), .ZN(n6530) );
  NOR2_X1 U3993 ( .A1(n7089), .A2(n4764), .ZN(n6588) );
  NOR2_X1 U3994 ( .A1(n7090), .A2(n4764), .ZN(n6580) );
  NOR2_X1 U3995 ( .A1(n6829), .A2(n4764), .ZN(n6597) );
  NOR2_X1 U3996 ( .A1(n6981), .A2(n4764), .ZN(n6559) );
  INV_X1 U3997 ( .A(n6514), .ZN(n5919) );
  INV_X1 U3998 ( .A(n6530), .ZN(n5926) );
  INV_X1 U3999 ( .A(n6580), .ZN(n5943) );
  INV_X1 U4000 ( .A(n6597), .ZN(n5948) );
  INV_X1 U4001 ( .A(n6552), .ZN(n5953) );
  INV_X1 U4002 ( .A(n6559), .ZN(n5961) );
  INV_X1 U4003 ( .A(n6561), .ZN(n5964) );
  AND2_X1 U4004 ( .A1(n4759), .A2(n4571), .ZN(n5072) );
  AND2_X1 U4005 ( .A1(n6634), .A2(n6633), .ZN(n6651) );
  AND2_X1 U4006 ( .A1(n4093), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6645) );
  INV_X1 U4007 ( .A(n6651), .ZN(n6708) );
  INV_X1 U4008 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U4009 ( .A1(n4234), .A2(STATE_REG_1__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U4010 ( .A1(n5464), .A2(n6318), .ZN(n4461) );
  OAI22_X1 U4011 ( .A1(n5508), .A2(n6310), .B1(n4458), .B2(n6322), .ZN(n4459)
         );
  OR2_X1 U4012 ( .A1(n4532), .A2(n4360), .ZN(n3172) );
  OAI21_X1 U4013 ( .B1(n5749), .B2(n5752), .A(n5750), .ZN(n5742) );
  NAND2_X2 U4014 ( .A1(n4679), .A2(n4361), .ZN(n4177) );
  INV_X1 U4015 ( .A(n3328), .ZN(n3331) );
  NAND2_X1 U4016 ( .A1(n3387), .A2(n3386), .ZN(n3498) );
  NAND2_X1 U4017 ( .A1(n4351), .A2(n4350), .ZN(n5658) );
  NAND2_X1 U4018 ( .A1(n5696), .A2(n5697), .ZN(n5695) );
  OR2_X1 U4019 ( .A1(n3354), .A2(n3338), .ZN(n3174) );
  NOR2_X1 U4020 ( .A1(n4260), .A2(n6471), .ZN(n3175) );
  NAND2_X1 U4021 ( .A1(n3347), .A2(n4531), .ZN(n3371) );
  NOR2_X2 U4022 ( .A1(n5514), .A2(n5516), .ZN(n5515) );
  OAI21_X1 U4023 ( .B1(n5332), .B2(n5333), .A(n5334), .ZN(n5758) );
  NAND2_X1 U4024 ( .A1(n3191), .A2(n4339), .ZN(n5320) );
  NAND2_X1 U4025 ( .A1(n3184), .A2(n4345), .ZN(n5727) );
  INV_X1 U4026 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3500) );
  AND2_X1 U4027 ( .A1(n4286), .A2(n6438), .ZN(n4596) );
  AND3_X1 U4028 ( .A1(n5808), .A2(n5822), .A3(n4402), .ZN(n3176) );
  NAND2_X1 U4029 ( .A1(n4638), .A2(n4637), .ZN(n4312) );
  XNOR2_X1 U4030 ( .A(n4310), .B(n4397), .ZN(n4637) );
  NAND2_X1 U4032 ( .A1(n3194), .A2(n3550), .ZN(n3564) );
  NAND2_X1 U4033 ( .A1(n4354), .A2(n4353), .ZN(n5432) );
  AND2_X1 U4034 ( .A1(n4420), .A2(n4449), .ZN(n3343) );
  NAND2_X1 U4035 ( .A1(n3455), .A2(n3475), .ZN(n3459) );
  AND2_X1 U4036 ( .A1(n4403), .A2(n4379), .ZN(n6502) );
  AND2_X1 U4037 ( .A1(n3677), .A2(n5145), .ZN(n3196) );
  INV_X1 U4038 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3380) );
  NOR2_X1 U4039 ( .A1(n4552), .A2(n4648), .ZN(n3197) );
  INV_X1 U4040 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6186) );
  AND2_X1 U4041 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3198) );
  AND2_X2 U4042 ( .A1(n3208), .A2(n5893), .ZN(n3422) );
  AND2_X2 U4043 ( .A1(n5893), .A2(n4546), .ZN(n3421) );
  AND3_X1 U4044 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3199) );
  XOR2_X1 U4045 ( .A(n4260), .B(n6106), .Z(n3200) );
  AND2_X1 U4046 ( .A1(n4429), .A2(n4428), .ZN(n3201) );
  NAND2_X1 U4047 ( .A1(n4480), .A2(n4130), .ZN(n4505) );
  INV_X2 U4048 ( .A(n6318), .ZN(n6311) );
  AND2_X1 U4049 ( .A1(n6322), .A2(n4449), .ZN(n6318) );
  NAND2_X1 U4050 ( .A1(n3464), .A2(n3702), .ZN(n3493) );
  AND2_X1 U4051 ( .A1(n4477), .A2(n4478), .ZN(n3492) );
  NAND2_X1 U4052 ( .A1(n5114), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4049) );
  OR2_X1 U4053 ( .A1(n4058), .A2(n4057), .ZN(n4059) );
  INV_X1 U4054 ( .A(n4059), .ZN(n4095) );
  NAND2_X1 U4055 ( .A1(n3462), .A2(n3461), .ZN(n3496) );
  AND2_X1 U4056 ( .A1(n3336), .A2(n3335), .ZN(n3355) );
  AOI22_X1 U4057 ( .A1(n3302), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3267) );
  INV_X1 U4058 ( .A(n5595), .ZN(n3838) );
  INV_X1 U4059 ( .A(n5545), .ZN(n3765) );
  INV_X1 U4060 ( .A(n4709), .ZN(n3585) );
  INV_X1 U4061 ( .A(n3403), .ZN(n4263) );
  AOI21_X1 U4062 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6619), .A(n4053), 
        .ZN(n4051) );
  INV_X1 U4063 ( .A(n5571), .ZN(n3924) );
  NAND2_X1 U4064 ( .A1(n5115), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3702) );
  INV_X1 U4065 ( .A(n3599), .ZN(n3614) );
  INV_X1 U4066 ( .A(n3712), .ZN(n3731) );
  INV_X1 U4067 ( .A(n5149), .ZN(n4162) );
  INV_X1 U4068 ( .A(n4283), .ZN(n4285) );
  XNOR2_X1 U4069 ( .A(n4511), .B(n4897), .ZN(n4529) );
  AND2_X1 U4070 ( .A1(n4169), .A2(n4168), .ZN(n6137) );
  AND2_X1 U4072 ( .A1(n3345), .A2(n4361), .ZN(n4232) );
  AOI21_X1 U4073 ( .B1(n3984), .B2(n3983), .A(n3982), .ZN(n5559) );
  INV_X1 U4074 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5186) );
  INV_X1 U4076 ( .A(n5851), .ZN(n4176) );
  OR2_X1 U4077 ( .A1(n5865), .A2(n5863), .ZN(n4405) );
  INV_X1 U4078 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3202) );
  INV_X1 U4079 ( .A(n4720), .ZN(n4602) );
  INV_X1 U4080 ( .A(n3473), .ZN(n3474) );
  AND2_X1 U4081 ( .A1(n4571), .A2(n4603), .ZN(n5034) );
  AND2_X1 U4082 ( .A1(n6150), .A2(n4527), .ZN(n4564) );
  AND2_X1 U4083 ( .A1(n5511), .A2(REIP_REG_31__SCAN_IN), .ZN(n4253) );
  NOR2_X1 U4084 ( .A1(n3646), .A2(n5216), .ZN(n3663) );
  INV_X1 U4085 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3592) );
  AND2_X1 U4086 ( .A1(n4172), .A2(n4171), .ZN(n5329) );
  INV_X1 U4087 ( .A(n4033), .ZN(n4005) );
  NAND2_X1 U4088 ( .A1(n3472), .A2(n3471), .ZN(n4477) );
  NAND2_X1 U4089 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4108)
         );
  NOR2_X1 U4090 ( .A1(n3630), .A2(n5186), .ZN(n3680) );
  NOR2_X1 U4091 ( .A1(n4890), .A2(n5152), .ZN(n5143) );
  INV_X1 U4092 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6273) );
  AND2_X1 U4093 ( .A1(n3359), .A2(n4366), .ZN(n4377) );
  NOR2_X1 U4094 ( .A1(n5445), .A2(n5444), .ZN(n5563) );
  AND2_X1 U4095 ( .A1(n4622), .A2(n4282), .ZN(n6440) );
  INV_X1 U4096 ( .A(n6499), .ZN(n5869) );
  AND3_X1 U4097 ( .A1(n4525), .A2(n4524), .A3(n4523), .ZN(n6611) );
  NAND2_X1 U4098 ( .A1(n4719), .A2(n4963), .ZN(n4935) );
  NAND2_X1 U4099 ( .A1(n4904), .A2(n4835), .ZN(n6568) );
  NAND2_X1 U4100 ( .A1(n3504), .A2(n3503), .ZN(n4897) );
  INV_X1 U4101 ( .A(n6553), .ZN(n5954) );
  INV_X1 U4102 ( .A(n6354), .ZN(n6720) );
  OR2_X1 U4103 ( .A1(n6717), .A2(n4107), .ZN(n6232) );
  NAND2_X1 U4104 ( .A1(n3566), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3593)
         );
  AND2_X1 U4105 ( .A1(n4140), .A2(n4139), .ZN(n4633) );
  INV_X1 U4106 ( .A(n4386), .ZN(n4487) );
  AND2_X1 U4107 ( .A1(n5481), .A2(n4427), .ZN(n6327) );
  NOR2_X1 U4108 ( .A1(n6719), .A2(n6330), .ZN(n6347) );
  NAND2_X1 U4109 ( .A1(n3920), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3961)
         );
  NAND2_X1 U4110 ( .A1(n3800), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3833)
         );
  INV_X1 U4111 ( .A(n6446), .ZN(n6095) );
  AND2_X1 U4112 ( .A1(n4377), .A2(n4064), .ZN(n4436) );
  NAND2_X1 U4113 ( .A1(n4413), .A2(n4412), .ZN(n4414) );
  NOR2_X1 U4114 ( .A1(n5804), .A2(n4410), .ZN(n6107) );
  OAI21_X1 U4115 ( .B1(n5719), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5695), 
        .ZN(n5689) );
  NOR2_X1 U4116 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5474) );
  OAI21_X1 U4117 ( .B1(n5912), .B2(n5913), .A(n5911), .ZN(n5960) );
  OAI21_X1 U4118 ( .B1(n4976), .B2(n4975), .A(n4974), .ZN(n5000) );
  OAI21_X1 U4119 ( .B1(n5084), .B2(n5083), .A(n5082), .ZN(n5108) );
  INV_X1 U4120 ( .A(n6516), .ZN(n6562) );
  AND2_X1 U4121 ( .A1(n4571), .A2(n4602), .ZN(n4904) );
  INV_X1 U4122 ( .A(n5033), .ZN(n4876) );
  NOR2_X1 U4123 ( .A1(n4689), .A2(n3159), .ZN(n6553) );
  AND2_X1 U4124 ( .A1(n5013), .A2(n5012), .ZN(n5386) );
  NOR2_X1 U4125 ( .A1(n6964), .A2(n4764), .ZN(n6571) );
  NOR2_X1 U4126 ( .A1(n6841), .A2(n4764), .ZN(n6552) );
  INV_X1 U4127 ( .A(n4653), .ZN(n6593) );
  INV_X1 U4128 ( .A(n5233), .ZN(n5272) );
  INV_X1 U4129 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6671) );
  INV_X1 U4130 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7092) );
  NOR2_X1 U4131 ( .A1(n4255), .A2(n4254), .ZN(n4256) );
  INV_X1 U4132 ( .A(n6297), .ZN(n6198) );
  INV_X1 U4133 ( .A(n6245), .ZN(n6292) );
  NAND2_X1 U4134 ( .A1(n6232), .A2(n4111), .ZN(n6236) );
  INV_X1 U4135 ( .A(n6250), .ZN(n6291) );
  INV_X1 U4136 ( .A(n4459), .ZN(n4460) );
  NAND2_X1 U4137 ( .A1(n6322), .A2(n5480), .ZN(n6310) );
  INV_X1 U4138 ( .A(n5976), .ZN(n5625) );
  INV_X1 U4139 ( .A(n6227), .ZN(n5300) );
  NAND2_X1 U4140 ( .A1(n4424), .A2(n6355), .ZN(n5481) );
  NAND2_X1 U4141 ( .A1(n6330), .A2(n5497), .ZN(n4585) );
  INV_X1 U4142 ( .A(n6330), .ZN(n6349) );
  NAND2_X1 U4143 ( .A1(n6161), .A2(n4439), .ZN(n6100) );
  NAND2_X1 U4144 ( .A1(n6100), .A2(n6447), .ZN(n6446) );
  OR2_X1 U4145 ( .A1(n6652), .A2(n6517), .ZN(n6454) );
  AOI21_X1 U4146 ( .B1(n5995), .B2(n6499), .A(n4414), .ZN(n4415) );
  NOR2_X1 U4147 ( .A1(n5864), .A2(n5829), .ZN(n6148) );
  INV_X1 U4148 ( .A(n6502), .ZN(n6134) );
  NOR2_X1 U4149 ( .A1(n4570), .A2(n5038), .ZN(n6507) );
  AND2_X1 U4150 ( .A1(n4723), .A2(n4722), .ZN(n4758) );
  NAND2_X1 U4151 ( .A1(n4932), .A2(n5012), .ZN(n5971) );
  AND2_X1 U4152 ( .A1(n4789), .A2(n4788), .ZN(n4826) );
  NAND2_X1 U4153 ( .A1(n4904), .A2(n5121), .ZN(n6584) );
  NOR2_X1 U4154 ( .A1(n4841), .A2(n4840), .ZN(n4879) );
  NAND2_X1 U4155 ( .A1(n5013), .A2(n5077), .ZN(n5033) );
  INV_X1 U4156 ( .A(n6588), .ZN(n5938) );
  INV_X1 U4157 ( .A(n6571), .ZN(n5933) );
  NOR2_X1 U4158 ( .A1(n4652), .A2(n4651), .ZN(n4696) );
  INV_X1 U4159 ( .A(n5036), .ZN(n5274) );
  INV_X1 U4160 ( .A(n4724), .ZN(n4931) );
  INV_X1 U4161 ( .A(n6645), .ZN(n6642) );
  INV_X1 U4162 ( .A(n6705), .ZN(n6654) );
  NAND2_X1 U4163 ( .A1(n4461), .A2(n4460), .ZN(U2829) );
  OAI21_X1 U4164 ( .B1(n5431), .B2(n6134), .A(n4415), .ZN(U2992) );
  AND2_X2 U4165 ( .A1(n3209), .A2(n5893), .ZN(n3423) );
  NOR2_X4 U4166 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4528) );
  AND2_X2 U4167 ( .A1(n4528), .A2(n4546), .ZN(n3315) );
  AOI22_X1 U4168 ( .A1(n3423), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3207) );
  INV_X1 U4169 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3203) );
  AND2_X2 U4170 ( .A1(n3208), .A2(n5894), .ZN(n3446) );
  AOI22_X1 U4171 ( .A1(n3446), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3206) );
  AND2_X2 U4172 ( .A1(n3209), .A2(n5894), .ZN(n3302) );
  AND2_X4 U4173 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4543) );
  AND2_X2 U4174 ( .A1(n4528), .A2(n4544), .ZN(n3310) );
  AOI22_X1 U4175 ( .A1(n3388), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3204) );
  AND2_X2 U4176 ( .A1(n3208), .A2(n4528), .ZN(n3303) );
  AOI22_X1 U4177 ( .A1(n3303), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3213) );
  AND2_X2 U4178 ( .A1(n5894), .A2(n4544), .ZN(n3297) );
  AOI22_X1 U4179 ( .A1(n3309), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3212) );
  AND2_X2 U4180 ( .A1(n3208), .A2(n4543), .ZN(n3393) );
  AND2_X2 U4181 ( .A1(n5893), .A2(n4544), .ZN(n3304) );
  AOI22_X1 U4182 ( .A1(n3393), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4184 ( .A1(n3441), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3210) );
  NAND2_X2 U4185 ( .A1(n3215), .A2(n3214), .ZN(n3328) );
  AOI22_X1 U4186 ( .A1(n3441), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4187 ( .A1(n3297), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4188 ( .A1(n3309), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4189 ( .A1(n3423), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4190 ( .A1(n3421), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4191 ( .A1(n3446), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4192 ( .A1(n3302), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3220) );
  NAND2_X2 U4193 ( .A1(n3331), .A2(n3327), .ZN(n4420) );
  NAND2_X1 U4194 ( .A1(n3423), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4195 ( .A1(n3446), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4196 ( .A1(n3297), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4197 ( .A1(n3304), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4198 ( .A1(n3422), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4199 ( .A1(n3309), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3232)
         );
  NAND2_X1 U4200 ( .A1(n3388), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4201 ( .A1(n3310), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4202 ( .A1(n3302), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U4203 ( .A1(n3303), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U4204 ( .A1(n3421), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3235)
         );
  NAND2_X1 U4205 ( .A1(n3428), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4206 ( .A1(n3441), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4207 ( .A1(n3393), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3241)
         );
  INV_X1 U4208 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4209 ( .A1(n3315), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3239)
         );
  AOI22_X1 U4210 ( .A1(n3446), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4211 ( .A1(n3309), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4212 ( .A1(n3423), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4213 ( .A1(n3422), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3247) );
  NAND4_X1 U4214 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n3256)
         );
  AOI22_X1 U4215 ( .A1(n3303), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4216 ( .A1(n3302), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4217 ( .A1(n3393), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4218 ( .A1(n3441), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3251) );
  NAND4_X1 U4219 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3255)
         );
  OR2_X2 U4220 ( .A1(n3256), .A2(n3255), .ZN(n4449) );
  NAND2_X2 U4221 ( .A1(n3349), .A2(n4449), .ZN(n3346) );
  INV_X1 U4222 ( .A(n3346), .ZN(n4358) );
  AOI22_X1 U4223 ( .A1(n3393), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4224 ( .A1(n3446), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4225 ( .A1(n3441), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3258) );
  NAND4_X1 U4226 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3266)
         );
  AOI22_X1 U4227 ( .A1(n3423), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4228 ( .A1(n3303), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4229 ( .A1(n3388), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4230 ( .A1(n3302), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3261) );
  NAND4_X1 U4231 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3265)
         );
  AOI22_X1 U4232 ( .A1(n3309), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4233 ( .A1(n3446), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4234 ( .A1(n3441), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4235 ( .A1(n3303), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4236 ( .A1(n3423), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4237 ( .A1(n3297), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4238 ( .A1(n3428), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4239 ( .A1(n3446), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4240 ( .A1(n3423), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4241 ( .A1(n3297), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4242 ( .A1(n3310), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4243 ( .A1(n3422), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4244 ( .A1(n3309), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3282)
         );
  NAND2_X1 U4245 ( .A1(n3388), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4246 ( .A1(n3304), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4247 ( .A1(n3302), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U4248 ( .A1(n3303), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4249 ( .A1(n3421), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4250 ( .A1(n3315), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3284)
         );
  NAND2_X1 U4251 ( .A1(n3441), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4252 ( .A1(n3393), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3290)
         );
  NAND2_X1 U4253 ( .A1(n3428), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3288) );
  NAND4_X4 U4254 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n4361)
         );
  AND2_X1 U4255 ( .A1(n4357), .A2(n4361), .ZN(n3296) );
  NAND2_X1 U4256 ( .A1(n4358), .A2(n3296), .ZN(n5499) );
  NAND2_X1 U4257 ( .A1(n3423), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4258 ( .A1(n3393), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3300)
         );
  NAND2_X1 U4259 ( .A1(n3446), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4260 ( .A1(n3297), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U4261 ( .A1(n3302), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4262 ( .A1(n3303), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3307) );
  NAND2_X1 U4263 ( .A1(n3441), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4264 ( .A1(n3304), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4265 ( .A1(n3422), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3314)
         );
  NAND2_X1 U4266 ( .A1(n3309), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3313)
         );
  NAND2_X1 U4267 ( .A1(n3388), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4268 ( .A1(n3310), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4269 ( .A1(n3421), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3320)
         );
  NAND2_X1 U4270 ( .A1(n3428), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4271 ( .A1(n3315), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3318)
         );
  NAND2_X1 U4272 ( .A1(n3316), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3317)
         );
  NAND4_X4 U4273 ( .A1(n3324), .A2(n3323), .A3(n3322), .A4(n3321), .ZN(n4384)
         );
  INV_X2 U4274 ( .A(n4384), .ZN(n3345) );
  NOR2_X1 U4275 ( .A1(n6671), .A2(n6662), .ZN(n6656) );
  NOR2_X1 U4276 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n3325) );
  NAND2_X1 U4277 ( .A1(n3345), .A2(n4233), .ZN(n3340) );
  INV_X1 U4278 ( .A(n3340), .ZN(n3333) );
  NAND2_X1 U4279 ( .A1(n4420), .A2(n3332), .ZN(n4101) );
  INV_X1 U4280 ( .A(n3326), .ZN(n3329) );
  NAND2_X1 U4281 ( .A1(n3158), .A2(n4264), .ZN(n3363) );
  NAND2_X1 U4282 ( .A1(n3329), .A2(n4103), .ZN(n3351) );
  INV_X1 U4283 ( .A(n3351), .ZN(n3330) );
  NAND4_X1 U4284 ( .A1(n4661), .A2(n4679), .A3(n3332), .A4(n5493), .ZN(n4532)
         );
  OAI211_X1 U4285 ( .C1(n5499), .C2(n3333), .A(n4534), .B(n3172), .ZN(n3334)
         );
  NAND2_X1 U4286 ( .A1(n3334), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4287 ( .A1(n5474), .A2(n4654), .ZN(n4438) );
  INV_X1 U4288 ( .A(n4438), .ZN(n3385) );
  XNOR2_X1 U4289 ( .A(n6606), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6510)
         );
  NAND2_X1 U4290 ( .A1(n3385), .A2(n6510), .ZN(n3336) );
  INV_X1 U4291 ( .A(n4093), .ZN(n3384) );
  NAND2_X1 U4292 ( .A1(n3384), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3335) );
  INV_X1 U4293 ( .A(n3355), .ZN(n3337) );
  NOR2_X1 U4294 ( .A1(n3337), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3338)
         );
  AND2_X1 U4295 ( .A1(n3158), .A2(n4361), .ZN(n3339) );
  NAND2_X1 U4296 ( .A1(n3346), .A2(n3339), .ZN(n4364) );
  NAND2_X1 U4297 ( .A1(n3360), .A2(n3456), .ZN(n3342) );
  NAND3_X1 U4298 ( .A1(n4364), .A2(n3344), .A3(n3359), .ZN(n3348) );
  NAND2_X1 U4299 ( .A1(n3346), .A2(n4232), .ZN(n3347) );
  NAND2_X1 U4300 ( .A1(n4064), .A2(n4112), .ZN(n4531) );
  NOR2_X1 U4301 ( .A1(n3348), .A2(n3371), .ZN(n3352) );
  NAND2_X1 U4302 ( .A1(n3159), .A2(n4449), .ZN(n3478) );
  OAI21_X1 U4303 ( .B1(n3351), .B2(n3350), .A(n4688), .ZN(n3375) );
  NAND2_X1 U4304 ( .A1(n3352), .A2(n3375), .ZN(n3353) );
  NAND2_X1 U4305 ( .A1(n3353), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3379) );
  AND2_X2 U4307 ( .A1(n3174), .A2(n3377), .ZN(n3409) );
  MUX2_X1 U4308 ( .A(n4093), .B(n4438), .S(n6606), .Z(n3357) );
  AOI21_X1 U4309 ( .B1(n4425), .B2(n3361), .A(n4679), .ZN(n3362) );
  NAND2_X1 U4310 ( .A1(n3359), .A2(n3362), .ZN(n3370) );
  NAND2_X1 U4311 ( .A1(n3363), .A2(n4232), .ZN(n3368) );
  NAND3_X1 U4312 ( .A1(n3332), .A2(n4679), .A3(n4449), .ZN(n3366) );
  INV_X1 U4313 ( .A(n3364), .ZN(n3365) );
  NAND2_X1 U4314 ( .A1(n5474), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6644) );
  AOI21_X1 U4315 ( .B1(n4385), .B2(n5497), .A(n6644), .ZN(n3367) );
  NAND3_X1 U4316 ( .A1(n3368), .A2(n4553), .A3(n3367), .ZN(n3369) );
  AOI21_X1 U4317 ( .B1(n3370), .B2(n4384), .A(n3369), .ZN(n3373) );
  INV_X1 U4318 ( .A(n3371), .ZN(n3372) );
  AND2_X1 U4319 ( .A1(n3373), .A2(n3372), .ZN(n3376) );
  NOR2_X1 U4320 ( .A1(n4308), .A2(n3361), .ZN(n3374) );
  OR2_X1 U4321 ( .A1(n3375), .A2(n3374), .ZN(n4395) );
  NAND2_X1 U4322 ( .A1(n3376), .A2(n4395), .ZN(n3438) );
  NAND2_X1 U4323 ( .A1(n3409), .A2(n3407), .ZN(n3378) );
  NAND2_X1 U4324 ( .A1(n3378), .A2(n3377), .ZN(n3497) );
  AND2_X1 U4325 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4326 ( .A1(n3381), .A2(n5114), .ZN(n5113) );
  INV_X1 U4327 ( .A(n3381), .ZN(n3382) );
  NAND2_X1 U4328 ( .A1(n3382), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4329 ( .A1(n5113), .A2(n3383), .ZN(n4656) );
  AOI22_X1 U4330 ( .A1(n3385), .A2(n4656), .B1(n3384), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3386) );
  XNOR2_X1 U4331 ( .A(n3497), .B(n3498), .ZN(n4551) );
  NAND2_X1 U4332 ( .A1(n4551), .A2(n4654), .ZN(n3402) );
  AOI22_X1 U4333 ( .A1(n4015), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4334 ( .A1(n4011), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4335 ( .A1(n4022), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4336 ( .A1(n4023), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3389) );
  NAND4_X1 U4337 ( .A1(n3392), .A2(n3391), .A3(n3390), .A4(n3389), .ZN(n3400)
         );
  AOI22_X1 U4338 ( .A1(n4020), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4339 ( .A1(n4021), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4340 ( .A1(n3948), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3396) );
  INV_X2 U4341 ( .A(n3394), .ZN(n4539) );
  AOI22_X1 U4342 ( .A1(n4024), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3395) );
  NAND4_X1 U4343 ( .A1(n3398), .A2(n3397), .A3(n3396), .A4(n3395), .ZN(n3399)
         );
  NAND2_X1 U4344 ( .A1(n4258), .A2(n3403), .ZN(n3401) );
  INV_X1 U4345 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4747) );
  OAI22_X1 U4346 ( .A1(n4078), .A2(n4747), .B1(n4263), .B2(n3505), .ZN(n3404)
         );
  XNOR2_X2 U4347 ( .A(n3406), .B(n3405), .ZN(n3520) );
  INV_X1 U4348 ( .A(n3407), .ZN(n3408) );
  AOI22_X1 U4349 ( .A1(n4021), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4350 ( .A1(n4011), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4351 ( .A1(n4020), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4352 ( .A1(n4014), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3410) );
  NAND4_X1 U4353 ( .A1(n3413), .A2(n3412), .A3(n3411), .A4(n3410), .ZN(n3419)
         );
  AOI22_X1 U4354 ( .A1(n4015), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4355 ( .A1(n3948), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4356 ( .A1(n3994), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4357 ( .A1(n4024), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3414) );
  NAND4_X1 U4358 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3418)
         );
  NAND2_X1 U4359 ( .A1(n4258), .A2(n4269), .ZN(n3420) );
  INV_X1 U4360 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U4361 ( .A1(n3302), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4362 ( .A1(n4023), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4363 ( .A1(n4022), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4364 ( .A1(n3441), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4365 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3434)
         );
  AOI22_X1 U4366 ( .A1(n4015), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4367 ( .A1(n4020), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4368 ( .A1(n4011), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4369 ( .A1(n3948), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4370 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3433)
         );
  NAND2_X1 U4371 ( .A1(n4258), .A2(n3453), .ZN(n3437) );
  INV_X1 U4372 ( .A(n3505), .ZN(n3435) );
  NAND2_X1 U4373 ( .A1(n3435), .A2(n4269), .ZN(n3436) );
  OAI211_X1 U4374 ( .C1(n4078), .C2(n4728), .A(n3437), .B(n3436), .ZN(n3465)
         );
  INV_X1 U4375 ( .A(n3438), .ZN(n3440) );
  NAND2_X1 U4376 ( .A1(n3480), .A2(n4654), .ZN(n3455) );
  AOI22_X1 U4377 ( .A1(n3302), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4378 ( .A1(n4011), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4379 ( .A1(n3948), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4380 ( .A1(n3297), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4381 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3452)
         );
  AOI22_X1 U4382 ( .A1(n4015), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4383 ( .A1(n4020), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4384 ( .A1(n3994), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4385 ( .A1(n4022), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4386 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3451)
         );
  XNOR2_X1 U4387 ( .A(n3453), .B(n4278), .ZN(n3454) );
  NAND2_X1 U4388 ( .A1(n3454), .A2(n4258), .ZN(n3475) );
  INV_X1 U4389 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4739) );
  AOI21_X1 U4390 ( .B1(n4666), .B2(n4334), .A(n4654), .ZN(n3458) );
  NAND2_X1 U4391 ( .A1(n4688), .A2(n4278), .ZN(n3457) );
  OAI211_X1 U4392 ( .C1(n4078), .C2(n4739), .A(n3458), .B(n3457), .ZN(n3473)
         );
  NAND2_X1 U4393 ( .A1(n4258), .A2(n4334), .ZN(n3460) );
  OAI21_X1 U4394 ( .B1(n3466), .B2(n3465), .A(n3467), .ZN(n3462) );
  NAND2_X1 U4395 ( .A1(n3466), .A2(n3465), .ZN(n3461) );
  INV_X1 U4396 ( .A(n3496), .ZN(n3463) );
  NAND2_X1 U4397 ( .A1(n4262), .A2(n3712), .ZN(n3464) );
  NAND2_X1 U4398 ( .A1(n4572), .A2(n3712), .ZN(n3472) );
  INV_X1 U4399 ( .A(n4360), .ZN(n4426) );
  AND2_X1 U4400 ( .A1(n4426), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4401 ( .A1(n3481), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4402 ( .A1(n3489), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5115), .ZN(n3469) );
  AND2_X1 U4403 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  NAND2_X1 U4404 ( .A1(n3475), .A2(n3474), .ZN(n3476) );
  INV_X1 U4405 ( .A(n3478), .ZN(n3479) );
  AOI21_X1 U4406 ( .B1(n5077), .B2(n3479), .A(n5115), .ZN(n4485) );
  NAND2_X1 U4407 ( .A1(n6609), .A2(n3712), .ZN(n3486) );
  INV_X1 U4408 ( .A(n3481), .ZN(n3544) );
  NAND2_X1 U4409 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5115), .ZN(n3483)
         );
  NAND2_X1 U4410 ( .A1(n3489), .A2(EAX_REG_0__SCAN_IN), .ZN(n3482) );
  OAI211_X1 U4411 ( .C1(n3544), .C2(n5478), .A(n3483), .B(n3482), .ZN(n3484)
         );
  INV_X1 U4412 ( .A(n3484), .ZN(n3485) );
  NAND2_X1 U4413 ( .A1(n3486), .A2(n3485), .ZN(n4484) );
  NAND2_X1 U4414 ( .A1(n4485), .A2(n4484), .ZN(n4483) );
  OR2_X1 U4415 ( .A1(n4484), .A2(n4008), .ZN(n3487) );
  NAND2_X1 U4416 ( .A1(n4483), .A2(n3487), .ZN(n4478) );
  INV_X1 U4417 ( .A(n3492), .ZN(n3488) );
  OAI21_X1 U4418 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3523), .ZN(n6445) );
  AOI22_X1 U4419 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4106), 
        .B2(n6445), .ZN(n3491) );
  NAND2_X1 U4420 ( .A1(n4036), .A2(EAX_REG_2__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U4421 ( .A1(n4489), .A2(n4490), .ZN(n3495) );
  NAND2_X1 U4422 ( .A1(n3492), .A2(n3493), .ZN(n3494) );
  INV_X1 U4423 ( .A(n3497), .ZN(n3499) );
  OR2_X1 U4424 ( .A1(n3379), .A2(n3500), .ZN(n3504) );
  NOR3_X1 U4425 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5114), .A3(n4838), 
        .ZN(n6508) );
  NAND2_X1 U4426 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6508), .ZN(n4920) );
  NAND2_X1 U4427 ( .A1(n6619), .A2(n4920), .ZN(n3501) );
  NOR3_X1 U4428 ( .A1(n6619), .A2(n5114), .A3(n4838), .ZN(n5040) );
  NAND2_X1 U4429 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5040), .ZN(n4926) );
  NAND2_X1 U4430 ( .A1(n3501), .A2(n4926), .ZN(n4715) );
  OAI22_X1 U4431 ( .A1(n4438), .A2(n4715), .B1(n4093), .B2(n6619), .ZN(n3502)
         );
  INV_X1 U4432 ( .A(n3502), .ZN(n3503) );
  NAND2_X1 U4433 ( .A1(n4529), .A2(n4654), .ZN(n3519) );
  AOI22_X1 U4434 ( .A1(n4015), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4435 ( .A1(n4011), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4436 ( .A1(n4022), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4437 ( .A1(n4023), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4438 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3517)
         );
  AOI22_X1 U4439 ( .A1(n4020), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4440 ( .A1(n4021), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4441 ( .A1(n3948), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3513) );
  INV_X1 U4442 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4443 ( .A1(n4024), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4444 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3516)
         );
  AOI22_X1 U4445 ( .A1(n4085), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4089), 
        .B2(n4288), .ZN(n3518) );
  NAND2_X1 U4446 ( .A1(n3520), .A2(n3496), .ZN(n3521) );
  NAND2_X1 U4447 ( .A1(n3521), .A2(n4602), .ZN(n3522) );
  OAI21_X1 U4448 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3524), .A(n3545), 
        .ZN(n6290) );
  AOI22_X1 U4449 ( .A1(n4106), .A2(n6290), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4450 ( .A1(n4036), .A2(EAX_REG_3__SCAN_IN), .ZN(n3525) );
  OAI211_X1 U4451 ( .C1(n3544), .C2(n3500), .A(n3526), .B(n3525), .ZN(n3527)
         );
  INV_X1 U4452 ( .A(n3527), .ZN(n3528) );
  OAI21_X1 U4453 ( .B1(n4290), .B2(n3731), .A(n3528), .ZN(n4502) );
  NAND2_X1 U4454 ( .A1(n4488), .A2(n4502), .ZN(n4503) );
  AOI22_X1 U4455 ( .A1(n4021), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4456 ( .A1(n4011), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4457 ( .A1(n4015), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4458 ( .A1(n3948), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4459 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3538)
         );
  AOI22_X1 U4460 ( .A1(n4014), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4461 ( .A1(n4020), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4462 ( .A1(n4540), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4463 ( .A1(n3994), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3533) );
  NAND4_X1 U4464 ( .A1(n3536), .A2(n3535), .A3(n3534), .A4(n3533), .ZN(n3537)
         );
  NAND2_X1 U4465 ( .A1(n4089), .A2(n4302), .ZN(n3540) );
  INV_X1 U4466 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4757) );
  OR2_X1 U4467 ( .A1(n4078), .A2(n4757), .ZN(n3539) );
  NAND2_X1 U4468 ( .A1(n3540), .A2(n3539), .ZN(n3550) );
  XNOR2_X1 U4469 ( .A(n3549), .B(n3550), .ZN(n4294) );
  INV_X1 U4470 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3543) );
  OAI21_X1 U4471 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n7092), .A(n5115), 
        .ZN(n3542) );
  NAND2_X1 U4472 ( .A1(n4036), .A2(EAX_REG_4__SCAN_IN), .ZN(n3541) );
  OAI211_X1 U4473 ( .C1(n3544), .C2(n3543), .A(n3542), .B(n3541), .ZN(n3547)
         );
  AOI21_X1 U4474 ( .B1(n3545), .B2(n6273), .A(n3566), .ZN(n6270) );
  NAND2_X1 U4475 ( .A1(n6270), .A2(n4106), .ZN(n3546) );
  AND2_X1 U4476 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  AOI21_X1 U4477 ( .B1(n4294), .B2(n3712), .A(n3548), .ZN(n4588) );
  NAND2_X1 U4478 ( .A1(n4085), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4479 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4015), .B1(n4014), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4480 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n4540), .B1(n4011), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4481 ( .A1(n4022), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4482 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n4023), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4483 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3560)
         );
  AOI22_X1 U4484 ( .A1(n4020), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4485 ( .A1(n4021), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4486 ( .A1(n3948), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4487 ( .A1(n4024), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3555) );
  NAND4_X1 U4488 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3559)
         );
  NAND2_X1 U4489 ( .A1(n4089), .A2(n4305), .ZN(n3561) );
  NAND2_X1 U4490 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  AOI22_X1 U4491 ( .A1(n3489), .A2(EAX_REG_5__SCAN_IN), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3568) );
  OAI21_X1 U4492 ( .B1(n3566), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3593), 
        .ZN(n6269) );
  NAND2_X1 U4493 ( .A1(n6269), .A2(n4106), .ZN(n3567) );
  OAI211_X1 U4494 ( .C1(n4309), .C2(n3731), .A(n3568), .B(n3567), .ZN(n4631)
         );
  NAND2_X1 U4495 ( .A1(n4586), .A2(n4631), .ZN(n4630) );
  INV_X1 U4496 ( .A(n4630), .ZN(n3586) );
  NAND2_X1 U4497 ( .A1(n4085), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4498 ( .A1(n4021), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4499 ( .A1(n4011), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4500 ( .A1(n4015), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4501 ( .A1(n4022), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3569) );
  NAND4_X1 U4502 ( .A1(n3572), .A2(n3571), .A3(n3570), .A4(n3569), .ZN(n3578)
         );
  AOI22_X1 U4503 ( .A1(n3948), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4504 ( .A1(n4012), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4505 ( .A1(n4540), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4506 ( .A1(n4024), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4507 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3577)
         );
  NAND2_X1 U4508 ( .A1(n4089), .A2(n4325), .ZN(n3579) );
  NAND2_X1 U4509 ( .A1(n3581), .A2(n3587), .ZN(n4313) );
  NAND2_X1 U4510 ( .A1(n4036), .A2(EAX_REG_6__SCAN_IN), .ZN(n3583) );
  OAI21_X1 U4511 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n7092), .A(n5115), 
        .ZN(n3582) );
  XOR2_X1 U4512 ( .A(n3592), .B(n3593), .Z(n6251) );
  AOI22_X1 U4513 ( .A1(n3583), .A2(n3582), .B1(n4106), .B2(n6251), .ZN(n3584)
         );
  NAND2_X1 U4514 ( .A1(n3586), .A2(n3585), .ZN(n4707) );
  INV_X1 U4515 ( .A(n4707), .ZN(n3679) );
  NAND2_X1 U4516 ( .A1(n3589), .A2(n3588), .ZN(n4314) );
  INV_X1 U4517 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U4518 ( .A1(n4089), .A2(n4334), .ZN(n3590) );
  OAI21_X1 U4519 ( .B1(n4732), .B2(n4078), .A(n3590), .ZN(n3591) );
  OAI21_X1 U4520 ( .B1(n3594), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3599), 
        .ZN(n6235) );
  NAND2_X1 U4521 ( .A1(n6235), .A2(n4106), .ZN(n3597) );
  NAND2_X1 U4522 ( .A1(n4036), .A2(EAX_REG_7__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4523 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3595)
         );
  NAND3_X1 U4524 ( .A1(n3597), .A2(n3596), .A3(n3595), .ZN(n3598) );
  XOR2_X1 U4525 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3614), .Z(n5178) );
  INV_X1 U4526 ( .A(n5178), .ZN(n5222) );
  AOI22_X1 U4527 ( .A1(n4024), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4528 ( .A1(n4011), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4529 ( .A1(n4015), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4530 ( .A1(n3994), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3600) );
  NAND4_X1 U4531 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3609)
         );
  AOI22_X1 U4532 ( .A1(n4022), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4533 ( .A1(n4020), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4534 ( .A1(n4540), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4535 ( .A1(n4021), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3604) );
  NAND4_X1 U4536 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3608)
         );
  NOR2_X1 U4537 ( .A1(n3609), .A2(n3608), .ZN(n3612) );
  NAND2_X1 U4538 ( .A1(n3489), .A2(EAX_REG_8__SCAN_IN), .ZN(n3611) );
  NAND2_X1 U4539 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3610)
         );
  OAI211_X1 U4540 ( .C1(n3731), .C2(n3612), .A(n3611), .B(n3610), .ZN(n3613)
         );
  AOI21_X1 U4541 ( .B1(n5222), .B2(n4106), .A(n3613), .ZN(n5152) );
  XOR2_X1 U4542 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3680), .Z(n6216) );
  INV_X1 U4543 ( .A(n6216), .ZN(n3629) );
  AOI22_X1 U4544 ( .A1(n4020), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4545 ( .A1(n4015), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4546 ( .A1(n4022), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4547 ( .A1(n3948), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4548 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3624)
         );
  AOI22_X1 U4549 ( .A1(n4011), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4550 ( .A1(n4024), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4551 ( .A1(n4014), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4552 ( .A1(n4021), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4553 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3623)
         );
  NOR2_X1 U4554 ( .A1(n3624), .A2(n3623), .ZN(n3627) );
  NAND2_X1 U4555 ( .A1(n3489), .A2(EAX_REG_12__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4556 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3625)
         );
  OAI211_X1 U4557 ( .C1(n3731), .C2(n3627), .A(n3626), .B(n3625), .ZN(n3628)
         );
  AOI21_X1 U4558 ( .B1(n3629), .B2(n4106), .A(n3628), .ZN(n5295) );
  INV_X1 U4559 ( .A(n5295), .ZN(n3677) );
  XNOR2_X1 U4560 ( .A(n3630), .B(n5186), .ZN(n5762) );
  AOI22_X1 U4561 ( .A1(n3948), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4562 ( .A1(n4015), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4563 ( .A1(n4024), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4564 ( .A1(n4540), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3631) );
  NAND4_X1 U4565 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3640)
         );
  AOI22_X1 U4566 ( .A1(n4011), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4567 ( .A1(n4020), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4568 ( .A1(n4021), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4569 ( .A1(n3989), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3635) );
  NAND4_X1 U4570 ( .A1(n3638), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3639)
         );
  NOR2_X1 U4571 ( .A1(n3640), .A2(n3639), .ZN(n3643) );
  NAND2_X1 U4572 ( .A1(n4036), .A2(EAX_REG_11__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4573 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3641)
         );
  OAI211_X1 U4574 ( .C1(n3731), .C2(n3643), .A(n3642), .B(n3641), .ZN(n3644)
         );
  AOI21_X1 U4575 ( .B1(n5762), .B2(n4106), .A(n3644), .ZN(n3645) );
  INV_X1 U4576 ( .A(n3645), .ZN(n5146) );
  XNOR2_X1 U4577 ( .A(n3646), .B(n5216), .ZN(n5323) );
  NAND2_X1 U4578 ( .A1(n5323), .A2(n4106), .ZN(n3662) );
  AOI22_X1 U4579 ( .A1(n4024), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4580 ( .A1(n4014), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4581 ( .A1(n4021), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4582 ( .A1(n4015), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4583 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3656)
         );
  AOI22_X1 U4584 ( .A1(n4011), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4585 ( .A1(n4020), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4586 ( .A1(n3948), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4587 ( .A1(n3157), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4588 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3655)
         );
  NOR2_X1 U4589 ( .A1(n3656), .A2(n3655), .ZN(n3659) );
  NAND2_X1 U4590 ( .A1(n4036), .A2(EAX_REG_9__SCAN_IN), .ZN(n3658) );
  NAND2_X1 U4591 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3657)
         );
  OAI211_X1 U4592 ( .C1(n3731), .C2(n3659), .A(n3658), .B(n3657), .ZN(n3660)
         );
  INV_X1 U4593 ( .A(n3660), .ZN(n3661) );
  NAND2_X1 U4594 ( .A1(n3662), .A2(n3661), .ZN(n5208) );
  XOR2_X1 U4595 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3663), .Z(n6226) );
  AOI22_X1 U4596 ( .A1(n4021), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4597 ( .A1(n4014), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4598 ( .A1(n4011), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4599 ( .A1(n3948), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3664) );
  NAND4_X1 U4600 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3673)
         );
  AOI22_X1 U4601 ( .A1(n4020), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4602 ( .A1(n4015), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4603 ( .A1(n4540), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4604 ( .A1(n3994), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4605 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3672)
         );
  OR2_X1 U4606 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  AOI22_X1 U4607 ( .A1(n3712), .A2(n3674), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4608 ( .A1(n4036), .A2(EAX_REG_10__SCAN_IN), .ZN(n3675) );
  OAI211_X1 U4609 ( .C1(n6226), .C2(n4008), .A(n3676), .B(n3675), .ZN(n5283)
         );
  AND2_X1 U4610 ( .A1(n5208), .A2(n5283), .ZN(n5144) );
  NAND2_X1 U4611 ( .A1(n3679), .A2(n3678), .ZN(n3695) );
  XNOR2_X1 U4612 ( .A(n3700), .B(n3699), .ZN(n6206) );
  NAND2_X1 U4613 ( .A1(n6206), .A2(n4106), .ZN(n3683) );
  NOR2_X1 U4614 ( .A1(n3702), .A2(n3699), .ZN(n3681) );
  AOI21_X1 U4615 ( .B1(n4036), .B2(EAX_REG_13__SCAN_IN), .A(n3681), .ZN(n3682)
         );
  NAND2_X1 U4616 ( .A1(n3683), .A2(n3682), .ZN(n3696) );
  XNOR2_X2 U4617 ( .A(n3695), .B(n3696), .ZN(n5312) );
  AOI22_X1 U4618 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n4015), .B1(n4014), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4619 ( .A1(n4011), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4620 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n4022), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4621 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4023), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4622 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4623 ( .A1(n4020), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4624 ( .A1(n4021), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4625 ( .A1(n3948), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4626 ( .A1(n4024), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4627 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  OR2_X1 U4628 ( .A1(n3693), .A2(n3692), .ZN(n3694) );
  AND2_X1 U4629 ( .A1(n3712), .A2(n3694), .ZN(n5313) );
  NAND2_X1 U4630 ( .A1(n5312), .A2(n5313), .ZN(n3698) );
  INV_X1 U4631 ( .A(n3695), .ZN(n5293) );
  NAND2_X1 U4632 ( .A1(n5293), .A2(n3696), .ZN(n3697) );
  INV_X1 U4633 ( .A(n3717), .ZN(n3701) );
  XNOR2_X1 U4634 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3701), .ZN(n6201)
         );
  INV_X1 U4635 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5738) );
  OAI22_X1 U4636 ( .A1(n6201), .A2(n4008), .B1(n3702), .B2(n5738), .ZN(n3703)
         );
  AOI21_X1 U4637 ( .B1(n4036), .B2(EAX_REG_14__SCAN_IN), .A(n3703), .ZN(n3716)
         );
  AOI22_X1 U4638 ( .A1(n4024), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4639 ( .A1(n4022), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4640 ( .A1(n4540), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4641 ( .A1(n4021), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4642 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3714)
         );
  AOI22_X1 U4643 ( .A1(n4015), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4644 ( .A1(n4011), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4645 ( .A1(n4020), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4646 ( .A1(n3994), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4647 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3713)
         );
  OAI21_X1 U4648 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3715) );
  NAND2_X1 U4649 ( .A1(n3716), .A2(n3715), .ZN(n5318) );
  NAND2_X1 U4650 ( .A1(n5316), .A2(n5318), .ZN(n5317) );
  XOR2_X1 U4651 ( .A(n6186), .B(n3733), .Z(n5734) );
  INV_X1 U4652 ( .A(n5734), .ZN(n6189) );
  AOI22_X1 U4653 ( .A1(n4011), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4654 ( .A1(n4020), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4655 ( .A1(n4024), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4656 ( .A1(n4014), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3718) );
  NAND4_X1 U4657 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3727)
         );
  AOI22_X1 U4658 ( .A1(n3948), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4659 ( .A1(n4015), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4660 ( .A1(n4023), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4661 ( .A1(n4021), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3722) );
  NAND4_X1 U4662 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3726)
         );
  NOR2_X1 U4663 ( .A1(n3727), .A2(n3726), .ZN(n3730) );
  NAND2_X1 U4664 ( .A1(n3489), .A2(EAX_REG_15__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U4665 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3728)
         );
  OAI211_X1 U4666 ( .C1(n3731), .C2(n3730), .A(n3729), .B(n3728), .ZN(n3732)
         );
  AOI21_X1 U4667 ( .B1(n6189), .B2(n4106), .A(n3732), .ZN(n5396) );
  INV_X1 U4668 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5723) );
  XNOR2_X1 U4669 ( .A(n3761), .B(n5723), .ZN(n6179) );
  AOI22_X1 U4670 ( .A1(n3489), .A2(EAX_REG_16__SCAN_IN), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4671 ( .A1(n4011), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4672 ( .A1(n4015), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4673 ( .A1(n4024), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4674 ( .A1(n4022), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4675 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3744)
         );
  AOI22_X1 U4676 ( .A1(n3948), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4677 ( .A1(n4020), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4678 ( .A1(n4023), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4679 ( .A1(n4021), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4680 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3743)
         );
  NAND2_X1 U4681 ( .A1(n4449), .A2(n3361), .ZN(n3742) );
  OAI21_X1 U4682 ( .B1(n3744), .B2(n3743), .A(n4033), .ZN(n3745) );
  OAI211_X1 U4683 ( .C1(n6179), .C2(n4008), .A(n3746), .B(n3745), .ZN(n5393)
         );
  NAND2_X1 U4684 ( .A1(n5389), .A2(n5393), .ZN(n5391) );
  INV_X1 U4685 ( .A(n5391), .ZN(n3766) );
  AOI22_X1 U4686 ( .A1(n4015), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4687 ( .A1(n4011), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4688 ( .A1(n4021), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4689 ( .A1(n4022), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4690 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3756)
         );
  AOI22_X1 U4691 ( .A1(n3948), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4692 ( .A1(n4014), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4693 ( .A1(n4020), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4694 ( .A1(n4024), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4695 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3755)
         );
  NOR2_X1 U4696 ( .A1(n3756), .A2(n3755), .ZN(n3760) );
  NAND2_X1 U4697 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3757)
         );
  NAND2_X1 U4698 ( .A1(n4008), .A2(n3757), .ZN(n3758) );
  AOI21_X1 U4699 ( .B1(n4036), .B2(EAX_REG_17__SCAN_IN), .A(n3758), .ZN(n3759)
         );
  OAI21_X1 U4700 ( .B1(n4005), .B2(n3760), .A(n3759), .ZN(n3764) );
  OAI21_X1 U4701 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3762), .A(n3799), 
        .ZN(n6094) );
  OR2_X1 U4702 ( .A1(n4008), .A2(n6094), .ZN(n3763) );
  NAND2_X1 U4703 ( .A1(n3764), .A2(n3763), .ZN(n5545) );
  NAND2_X1 U4704 ( .A1(n3766), .A2(n3765), .ZN(n5531) );
  INV_X1 U4705 ( .A(n5531), .ZN(n3784) );
  AOI22_X1 U4706 ( .A1(n4022), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4707 ( .A1(n4021), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4708 ( .A1(n4024), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4709 ( .A1(n4014), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4710 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3778)
         );
  NAND2_X1 U4711 ( .A1(n4011), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4712 ( .A1(n4020), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3771)
         );
  AND3_X1 U4713 ( .A1(n3772), .A2(n3771), .A3(n4008), .ZN(n3776) );
  AOI22_X1 U4714 ( .A1(n4023), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4715 ( .A1(n3948), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4716 ( .A1(n4015), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4717 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3777)
         );
  NAND2_X1 U4718 ( .A1(n4005), .A2(n4008), .ZN(n3850) );
  OAI21_X1 U4719 ( .B1(n3778), .B2(n3777), .A(n3850), .ZN(n3780) );
  AOI22_X1 U4720 ( .A1(n3489), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5115), .ZN(n3779) );
  NAND2_X1 U4721 ( .A1(n3780), .A2(n3779), .ZN(n3782) );
  XNOR2_X1 U4722 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3799), .ZN(n5715)
         );
  NAND2_X1 U4723 ( .A1(n5715), .A2(n4106), .ZN(n3781) );
  NAND2_X1 U4724 ( .A1(n3782), .A2(n3781), .ZN(n5534) );
  NAND2_X1 U4725 ( .A1(n3784), .A2(n3783), .ZN(n5532) );
  AOI22_X1 U4726 ( .A1(n4024), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4727 ( .A1(n4015), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4728 ( .A1(n4021), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4729 ( .A1(n4540), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4730 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4731 ( .A1(n4020), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4732 ( .A1(n4011), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4733 ( .A1(n3948), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4734 ( .A1(n3994), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4735 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  NOR2_X1 U4736 ( .A1(n3794), .A2(n3793), .ZN(n3798) );
  NAND2_X1 U4737 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3795)
         );
  NAND2_X1 U4738 ( .A1(n4008), .A2(n3795), .ZN(n3796) );
  AOI21_X1 U4739 ( .B1(n4036), .B2(EAX_REG_19__SCAN_IN), .A(n3796), .ZN(n3797)
         );
  OAI21_X1 U4740 ( .B1(n4005), .B2(n3798), .A(n3797), .ZN(n3802) );
  OAI21_X1 U4741 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3800), .A(n3833), 
        .ZN(n6090) );
  OR2_X1 U4742 ( .A1(n4008), .A2(n6090), .ZN(n3801) );
  NAND2_X1 U4743 ( .A1(n3802), .A2(n3801), .ZN(n5610) );
  NAND2_X1 U4744 ( .A1(n4011), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4745 ( .A1(n4020), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3803)
         );
  AND3_X1 U4746 ( .A1(n3804), .A2(n3803), .A3(n4008), .ZN(n3808) );
  AOI22_X1 U4747 ( .A1(n4540), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4748 ( .A1(n3948), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4749 ( .A1(n4013), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4750 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3814)
         );
  AOI22_X1 U4751 ( .A1(n4022), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4752 ( .A1(n4024), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4753 ( .A1(n4021), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4754 ( .A1(n4015), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4755 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  OR2_X1 U4756 ( .A1(n3814), .A2(n3813), .ZN(n3815) );
  NAND2_X1 U4757 ( .A1(n3850), .A2(n3815), .ZN(n3818) );
  AOI22_X1 U4758 ( .A1(n3489), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5115), .ZN(n3817) );
  XNOR2_X1 U4759 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3833), .ZN(n6045)
         );
  AND2_X1 U4760 ( .A1(n6045), .A2(n4106), .ZN(n3816) );
  AOI21_X1 U4761 ( .B1(n3818), .B2(n3817), .A(n3816), .ZN(n5603) );
  NAND2_X1 U4762 ( .A1(n5601), .A2(n5603), .ZN(n5592) );
  INV_X1 U4763 ( .A(n5592), .ZN(n3839) );
  AOI22_X1 U4764 ( .A1(n4020), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4765 ( .A1(n4011), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4766 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4015), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4767 ( .A1(n4021), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4768 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3828)
         );
  AOI22_X1 U4769 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n3948), .B1(n4024), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4770 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n4014), .B1(n4022), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4771 ( .A1(n3994), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4772 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4023), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4773 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  NOR2_X1 U4774 ( .A1(n3828), .A2(n3827), .ZN(n3832) );
  NAND2_X1 U4775 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3829)
         );
  NAND2_X1 U4776 ( .A1(n4008), .A2(n3829), .ZN(n3830) );
  AOI21_X1 U4777 ( .B1(n4036), .B2(EAX_REG_21__SCAN_IN), .A(n3830), .ZN(n3831)
         );
  OAI21_X1 U4778 ( .B1(n4005), .B2(n3832), .A(n3831), .ZN(n3837) );
  OAI21_X1 U4779 ( .B1(n3835), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3882), 
        .ZN(n6036) );
  OR2_X1 U4780 ( .A1(n6036), .A2(n4008), .ZN(n3836) );
  NAND2_X1 U4781 ( .A1(n3837), .A2(n3836), .ZN(n5595) );
  NAND2_X1 U4782 ( .A1(n3839), .A2(n3838), .ZN(n5587) );
  AOI22_X1 U4783 ( .A1(n3948), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4784 ( .A1(n4024), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4785 ( .A1(n3994), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4786 ( .A1(n4012), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3840) );
  NAND4_X1 U4787 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n3852)
         );
  AOI22_X1 U4788 ( .A1(n4021), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4789 ( .A1(n4022), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4790 ( .A1(n4014), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3847) );
  NAND2_X1 U4791 ( .A1(n4011), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3845) );
  NAND2_X1 U4792 ( .A1(n4020), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3844)
         );
  AND3_X1 U4793 ( .A1(n3845), .A2(n3844), .A3(n4008), .ZN(n3846) );
  NAND4_X1 U4794 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3851)
         );
  OAI21_X1 U4795 ( .B1(n3852), .B2(n3851), .A(n3850), .ZN(n3855) );
  INV_X1 U4796 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5691) );
  NOR2_X1 U4797 ( .A1(n5691), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3853) );
  AOI21_X1 U4798 ( .B1(n4036), .B2(EAX_REG_22__SCAN_IN), .A(n3853), .ZN(n3854)
         );
  NAND2_X1 U4799 ( .A1(n3855), .A2(n3854), .ZN(n3857) );
  XNOR2_X1 U4800 ( .A(n3882), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6027)
         );
  NAND2_X1 U4801 ( .A1(n6027), .A2(n4106), .ZN(n3856) );
  NAND2_X1 U4802 ( .A1(n3857), .A2(n3856), .ZN(n5590) );
  NOR2_X2 U4803 ( .A1(n5587), .A2(n5590), .ZN(n5588) );
  AOI22_X1 U4804 ( .A1(n4021), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4805 ( .A1(n4015), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4806 ( .A1(n3157), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4807 ( .A1(n4540), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4808 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3867)
         );
  AOI22_X1 U4809 ( .A1(n4024), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4810 ( .A1(n4011), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4811 ( .A1(n4014), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4812 ( .A1(n4012), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4813 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3866)
         );
  NOR2_X1 U4814 ( .A1(n3867), .A2(n3866), .ZN(n3888) );
  AOI22_X1 U4815 ( .A1(n4020), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4816 ( .A1(n4540), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4817 ( .A1(n4023), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4818 ( .A1(n4024), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4819 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3877)
         );
  AOI22_X1 U4820 ( .A1(n3948), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4821 ( .A1(n4011), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4822 ( .A1(n4021), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4823 ( .A1(n4015), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4824 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3876)
         );
  NOR2_X1 U4825 ( .A1(n3877), .A2(n3876), .ZN(n3889) );
  XNOR2_X1 U4826 ( .A(n3888), .B(n3889), .ZN(n3881) );
  NAND2_X1 U4827 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3878)
         );
  NAND2_X1 U4828 ( .A1(n4008), .A2(n3878), .ZN(n3879) );
  AOI21_X1 U4829 ( .B1(n4036), .B2(EAX_REG_23__SCAN_IN), .A(n3879), .ZN(n3880)
         );
  OAI21_X1 U4830 ( .B1(n4005), .B2(n3881), .A(n3880), .ZN(n3887) );
  NOR2_X1 U4831 ( .A1(n3883), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3884)
         );
  OR2_X1 U4832 ( .A1(n3919), .A2(n3884), .ZN(n6018) );
  INV_X1 U4833 ( .A(n6018), .ZN(n3885) );
  NAND2_X1 U4834 ( .A1(n3885), .A2(n4106), .ZN(n3886) );
  AND2_X2 U4835 ( .A1(n5588), .A2(n5675), .ZN(n5577) );
  OR2_X1 U4836 ( .A1(n3889), .A2(n3888), .ZN(n3914) );
  AOI22_X1 U4837 ( .A1(n4020), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4838 ( .A1(n4023), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4839 ( .A1(n3948), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4840 ( .A1(n4021), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4841 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3899)
         );
  AOI22_X1 U4842 ( .A1(n4015), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4843 ( .A1(n4024), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4844 ( .A1(n4011), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4845 ( .A1(n4540), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4846 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  NOR2_X1 U4847 ( .A1(n3899), .A2(n3898), .ZN(n3913) );
  XNOR2_X1 U4848 ( .A(n3914), .B(n3913), .ZN(n3902) );
  AOI22_X1 U4849 ( .A1(n3489), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4039), .ZN(n3901) );
  XNOR2_X1 U4850 ( .A(n3919), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6007)
         );
  NAND2_X1 U4851 ( .A1(n6007), .A2(n4106), .ZN(n3900) );
  OAI211_X1 U4852 ( .C1(n3902), .C2(n4005), .A(n3901), .B(n3900), .ZN(n5578)
         );
  NAND2_X1 U4853 ( .A1(n5577), .A2(n5578), .ZN(n5569) );
  AOI22_X1 U4854 ( .A1(n4021), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4855 ( .A1(n4011), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4856 ( .A1(n4015), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4857 ( .A1(n4020), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4858 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3912)
         );
  AOI22_X1 U4859 ( .A1(n4014), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4860 ( .A1(n3948), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4861 ( .A1(n4023), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4862 ( .A1(n4012), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4863 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3911)
         );
  NOR2_X1 U4864 ( .A1(n3912), .A2(n3911), .ZN(n3927) );
  OR2_X1 U4865 ( .A1(n3914), .A2(n3913), .ZN(n3926) );
  XNOR2_X1 U4866 ( .A(n3927), .B(n3926), .ZN(n3918) );
  NAND2_X1 U4867 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3915)
         );
  NAND2_X1 U4868 ( .A1(n4008), .A2(n3915), .ZN(n3916) );
  AOI21_X1 U4869 ( .B1(n4036), .B2(EAX_REG_25__SCAN_IN), .A(n3916), .ZN(n3917)
         );
  OAI21_X1 U4870 ( .B1(n3918), .B2(n4005), .A(n3917), .ZN(n3923) );
  OR2_X1 U4871 ( .A1(n3920), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3921)
         );
  NAND2_X1 U4872 ( .A1(n3921), .A2(n3961), .ZN(n6084) );
  INV_X1 U4873 ( .A(n6084), .ZN(n6000) );
  NAND2_X1 U4874 ( .A1(n6000), .A2(n4106), .ZN(n3922) );
  NAND2_X1 U4875 ( .A1(n3923), .A2(n3922), .ZN(n5571) );
  NOR2_X1 U4876 ( .A1(n3927), .A2(n3926), .ZN(n3956) );
  AOI22_X1 U4877 ( .A1(n4015), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4878 ( .A1(n4011), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4879 ( .A1(n4022), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4880 ( .A1(n4023), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4881 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U4882 ( .A1(n4020), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4883 ( .A1(n4021), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4884 ( .A1(n3948), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4885 ( .A1(n4024), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4886 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  OR2_X1 U4887 ( .A1(n3937), .A2(n3936), .ZN(n3955) );
  XNOR2_X1 U4888 ( .A(n3956), .B(n3955), .ZN(n3941) );
  NAND2_X1 U4889 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3938)
         );
  NAND2_X1 U4890 ( .A1(n4008), .A2(n3938), .ZN(n3939) );
  AOI21_X1 U4891 ( .B1(n4036), .B2(EAX_REG_26__SCAN_IN), .A(n3939), .ZN(n3940)
         );
  OAI21_X1 U4892 ( .B1(n3941), .B2(n4005), .A(n3940), .ZN(n3943) );
  XNOR2_X1 U4893 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n3961), .ZN(n5990)
         );
  NAND2_X1 U4894 ( .A1(n5990), .A2(n4106), .ZN(n3942) );
  NAND2_X1 U4895 ( .A1(n3943), .A2(n3942), .ZN(n5425) );
  AOI22_X1 U4896 ( .A1(n4014), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4897 ( .A1(n4011), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4898 ( .A1(n4020), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4899 ( .A1(n4023), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4900 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3954)
         );
  AOI22_X1 U4901 ( .A1(n4021), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4902 ( .A1(n4015), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4903 ( .A1(n4012), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4904 ( .A1(n3948), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U4905 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3953)
         );
  NOR2_X1 U4906 ( .A1(n3954), .A2(n3953), .ZN(n3967) );
  NAND2_X1 U4907 ( .A1(n3956), .A2(n3955), .ZN(n3966) );
  XNOR2_X1 U4908 ( .A(n3967), .B(n3966), .ZN(n3960) );
  NAND2_X1 U4909 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3957)
         );
  NAND2_X1 U4910 ( .A1(n4008), .A2(n3957), .ZN(n3958) );
  AOI21_X1 U4911 ( .B1(n4036), .B2(EAX_REG_27__SCAN_IN), .A(n3958), .ZN(n3959)
         );
  OAI21_X1 U4912 ( .B1(n3960), .B2(n4005), .A(n3959), .ZN(n3965) );
  INV_X1 U4913 ( .A(n3961), .ZN(n3962) );
  OAI21_X1 U4914 ( .B1(n3963), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n3985), 
        .ZN(n5982) );
  OR2_X1 U4915 ( .A1(n5982), .A2(n4008), .ZN(n3964) );
  NAND2_X1 U4916 ( .A1(n3965), .A2(n3964), .ZN(n5438) );
  NOR2_X1 U4917 ( .A1(n3967), .A2(n3966), .ZN(n4002) );
  AOI22_X1 U4918 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4015), .B1(n4014), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4919 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n4540), .B1(n4011), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4920 ( .A1(n4022), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4921 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n4023), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3968) );
  NAND4_X1 U4922 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(n3977)
         );
  AOI22_X1 U4923 ( .A1(n4020), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4924 ( .A1(n4021), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4925 ( .A1(n3948), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4926 ( .A1(n4024), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4927 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976)
         );
  OR2_X1 U4928 ( .A1(n3977), .A2(n3976), .ZN(n4001) );
  INV_X1 U4929 ( .A(n4001), .ZN(n3978) );
  XNOR2_X1 U4930 ( .A(n4002), .B(n3978), .ZN(n3979) );
  NAND2_X1 U4931 ( .A1(n3979), .A2(n4033), .ZN(n3984) );
  NAND2_X1 U4932 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3980)
         );
  NAND2_X1 U4933 ( .A1(n4008), .A2(n3980), .ZN(n3981) );
  AOI21_X1 U4934 ( .B1(n4036), .B2(EAX_REG_28__SCAN_IN), .A(n3981), .ZN(n3983)
         );
  XNOR2_X1 U4935 ( .A(n3985), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5973)
         );
  AND2_X1 U4936 ( .A1(n5973), .A2(n4106), .ZN(n3982) );
  INV_X1 U4937 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5654) );
  INV_X1 U4938 ( .A(n3986), .ZN(n3987) );
  INV_X1 U4939 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U4940 ( .A1(n3987), .A2(n5524), .ZN(n3988) );
  NAND2_X1 U4941 ( .A1(n4108), .A2(n3988), .ZN(n5645) );
  AOI22_X1 U4942 ( .A1(n4014), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4023), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4943 ( .A1(n4015), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4944 ( .A1(n4540), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4945 ( .A1(n4024), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U4946 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n4000)
         );
  AOI22_X1 U4947 ( .A1(n4011), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4948 ( .A1(n4020), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4949 ( .A1(n4021), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4950 ( .A1(n3948), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4951 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  NOR2_X1 U4952 ( .A1(n4000), .A2(n3999), .ZN(n4010) );
  NAND2_X1 U4953 ( .A1(n4002), .A2(n4001), .ZN(n4009) );
  XNOR2_X1 U4954 ( .A(n4010), .B(n4009), .ZN(n4006) );
  AOI21_X1 U4955 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5115), .A(n4106), 
        .ZN(n4004) );
  NAND2_X1 U4956 ( .A1(n3489), .A2(EAX_REG_29__SCAN_IN), .ZN(n4003) );
  OAI211_X1 U4957 ( .C1(n4006), .C2(n4005), .A(n4004), .B(n4003), .ZN(n4007)
         );
  OAI21_X1 U4958 ( .B1(n4008), .B2(n5645), .A(n4007), .ZN(n5516) );
  NOR2_X1 U4959 ( .A1(n4010), .A2(n4009), .ZN(n4032) );
  AOI22_X1 U4960 ( .A1(n4011), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4961 ( .A1(n4012), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4962 ( .A1(n4014), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4963 ( .A1(n4015), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4964 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4030)
         );
  AOI22_X1 U4965 ( .A1(n4021), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4966 ( .A1(n3948), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4967 ( .A1(n4023), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4968 ( .A1(n4024), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U4969 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4029)
         );
  NOR2_X1 U4970 ( .A1(n4030), .A2(n4029), .ZN(n4031) );
  XNOR2_X1 U4971 ( .A(n4032), .B(n4031), .ZN(n4034) );
  NAND2_X1 U4972 ( .A1(n4034), .A2(n4033), .ZN(n4038) );
  INV_X1 U4973 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5465) );
  AOI21_X1 U4974 ( .B1(n5465), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4035) );
  AOI21_X1 U4975 ( .B1(n4036), .B2(EAX_REG_30__SCAN_IN), .A(n4035), .ZN(n4037)
         );
  XNOR2_X1 U4976 ( .A(n4108), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5505)
         );
  NAND2_X1 U4977 ( .A1(n5515), .A2(n4416), .ZN(n4042) );
  AOI22_X1 U4978 ( .A1(n4036), .A2(EAX_REG_31__SCAN_IN), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4040) );
  XNOR2_X2 U4979 ( .A(n4042), .B(n4041), .ZN(n5483) );
  INV_X1 U4980 ( .A(n5483), .ZN(n4257) );
  NAND2_X1 U4981 ( .A1(n4838), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U4982 ( .A1(n4043), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4044) );
  NAND2_X1 U4983 ( .A1(n4045), .A2(n4044), .ZN(n4060) );
  NAND2_X1 U4984 ( .A1(n6606), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U4985 ( .A1(n4046), .A2(n4045), .ZN(n4077) );
  NAND2_X1 U4986 ( .A1(n3380), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4047) );
  NAND2_X1 U4987 ( .A1(n4049), .A2(n4047), .ZN(n4076) );
  INV_X1 U4988 ( .A(n4076), .ZN(n4048) );
  NAND2_X1 U4989 ( .A1(n4077), .A2(n4048), .ZN(n4050) );
  NAND2_X1 U4990 ( .A1(n4050), .A2(n4049), .ZN(n4055) );
  XNOR2_X1 U4991 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4056) );
  OAI222_X1 U4992 ( .A1(n3543), .A2(n4051), .B1(n3543), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n4051), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4100) );
  NAND2_X1 U4993 ( .A1(n4100), .A2(n4069), .ZN(n4092) );
  NAND2_X1 U4994 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4051), .ZN(n4052) );
  NOR2_X1 U4995 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4052), .ZN(n4058)
         );
  INV_X1 U4996 ( .A(n4053), .ZN(n4054) );
  OAI21_X1 U4997 ( .B1(n4056), .B2(n4055), .A(n4054), .ZN(n4057) );
  AOI22_X1 U4998 ( .A1(n4069), .A2(n4059), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4654), .ZN(n4087) );
  XOR2_X1 U4999 ( .A(n4060), .B(n4062), .Z(n4096) );
  INV_X1 U5000 ( .A(n4096), .ZN(n4061) );
  NOR2_X1 U5001 ( .A1(n4654), .A2(n4061), .ZN(n4075) );
  INV_X1 U5002 ( .A(n4089), .ZN(n4068) );
  OAI21_X1 U5003 ( .B1(n3345), .B2(n4068), .A(n4270), .ZN(n4074) );
  INV_X1 U5004 ( .A(n4062), .ZN(n4063) );
  AOI21_X1 U5005 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n5478), .A(n4063), 
        .ZN(n4065) );
  INV_X1 U5006 ( .A(n4065), .ZN(n4067) );
  AOI21_X1 U5007 ( .B1(n4661), .B2(n4361), .A(n4384), .ZN(n4080) );
  INV_X1 U5008 ( .A(n4064), .ZN(n4376) );
  AOI21_X1 U5009 ( .B1(n4065), .B2(n4376), .A(n4688), .ZN(n4066) );
  NOR3_X1 U5010 ( .A1(n4068), .A2(n4067), .A3(n4071), .ZN(n4073) );
  INV_X1 U5011 ( .A(n4069), .ZN(n4070) );
  AOI21_X1 U5012 ( .B1(n4096), .B2(n4071), .A(n4070), .ZN(n4072) );
  AOI211_X1 U5013 ( .C1(n4075), .C2(n4074), .A(n4073), .B(n4072), .ZN(n4083)
         );
  XNOR2_X1 U5014 ( .A(n4077), .B(n4076), .ZN(n4098) );
  NOR2_X1 U5015 ( .A1(n4078), .A2(n4098), .ZN(n4079) );
  AOI211_X1 U5016 ( .C1(n4089), .C2(n4098), .A(n4079), .B(n4080), .ZN(n4082)
         );
  NAND3_X1 U5017 ( .A1(n4080), .A2(n4089), .A3(n4098), .ZN(n4081) );
  OAI21_X1 U5018 ( .B1(n4083), .B2(n4082), .A(n4081), .ZN(n4084) );
  OAI21_X1 U5019 ( .B1(n4085), .B2(n4095), .A(n4084), .ZN(n4086) );
  NAND2_X1 U5020 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  AOI21_X1 U5021 ( .B1(n4089), .B2(n4100), .A(n4088), .ZN(n4090) );
  INV_X1 U5022 ( .A(n4090), .ZN(n4091) );
  INV_X1 U5023 ( .A(n5499), .ZN(n4094) );
  AND2_X1 U5024 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  AND2_X1 U5025 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  OR2_X1 U5026 ( .A1(n4100), .A2(n4099), .ZN(n5501) );
  INV_X1 U5027 ( .A(n5501), .ZN(n4105) );
  NAND3_X1 U5028 ( .A1(n4103), .A2(n4102), .A3(n4101), .ZN(n5500) );
  NOR2_X1 U5029 ( .A1(n5500), .A2(n6642), .ZN(n4104) );
  NOR2_X1 U5030 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6723) );
  NAND3_X1 U5031 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), 
        .A3(n6723), .ZN(n6640) );
  OR2_X1 U5032 ( .A1(n4438), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6259) );
  AND2_X1 U5033 ( .A1(n4654), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U5034 ( .A1(n4106), .A2(n4437), .ZN(n6649) );
  NAND3_X1 U5035 ( .A1(n6640), .A2(n6120), .A3(n6649), .ZN(n4107) );
  INV_X1 U5036 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4109) );
  NOR2_X1 U5037 ( .A1(n5176), .A2(n5472), .ZN(n4111) );
  AND2_X2 U5038 ( .A1(n4361), .A2(n4384), .ZN(n4481) );
  AND2_X1 U5039 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4113)
         );
  AOI21_X1 U5040 ( .B1(n4487), .B2(EBX_REG_30__SCAN_IN), .A(n4113), .ZN(n4453)
         );
  MUX2_X1 U5041 ( .A(n4217), .B(n4133), .S(EBX_REG_3__SCAN_IN), .Z(n4116) );
  INV_X1 U5042 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U5043 ( .A1(n4386), .A2(n4114), .ZN(n4115) );
  AND2_X1 U5044 ( .A1(n4116), .A2(n4115), .ZN(n4506) );
  INV_X1 U5045 ( .A(n4177), .ZN(n4117) );
  MUX2_X1 U5046 ( .A(n4123), .B(n4177), .S(EBX_REG_2__SCAN_IN), .Z(n4120) );
  NAND2_X1 U5047 ( .A1(n4117), .A2(n4374), .ZN(n4205) );
  NAND2_X1 U5048 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4118)
         );
  AND2_X1 U5049 ( .A1(n4205), .A2(n4118), .ZN(n4119) );
  INV_X1 U5050 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U5051 ( .A1(n4177), .A2(n4281), .ZN(n4122) );
  INV_X1 U5052 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4124) );
  NAND2_X1 U5053 ( .A1(n4481), .A2(n4124), .ZN(n4121) );
  NAND3_X1 U5054 ( .A1(n4122), .A2(n4133), .A3(n4121), .ZN(n4126) );
  NAND2_X1 U5055 ( .A1(n4132), .A2(n4124), .ZN(n4125) );
  NAND2_X1 U5056 ( .A1(n4126), .A2(n4125), .ZN(n4128) );
  NAND2_X1 U5057 ( .A1(n4177), .A2(EBX_REG_0__SCAN_IN), .ZN(n4127) );
  OAI21_X1 U5058 ( .B1(n5537), .B2(EBX_REG_0__SCAN_IN), .A(n4127), .ZN(n4486)
         );
  XNOR2_X1 U5059 ( .A(n4128), .B(n4486), .ZN(n4479) );
  NAND2_X1 U5060 ( .A1(n4479), .A2(n4481), .ZN(n4480) );
  INV_X1 U5061 ( .A(n4128), .ZN(n4129) );
  NAND2_X1 U5062 ( .A1(n4129), .A2(n4486), .ZN(n4130) );
  INV_X1 U5063 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4134) );
  NAND2_X1 U5064 ( .A1(n4211), .A2(n4134), .ZN(n4138) );
  INV_X1 U5065 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U5066 ( .A1(n4177), .A2(n4298), .ZN(n4136) );
  NAND2_X1 U5067 ( .A1(n4481), .A2(n4134), .ZN(n4135) );
  NAND3_X1 U5068 ( .A1(n4136), .A2(n4133), .A3(n4135), .ZN(n4137) );
  AND2_X1 U5069 ( .A1(n4138), .A2(n4137), .ZN(n4591) );
  MUX2_X1 U5070 ( .A(n4217), .B(n4133), .S(EBX_REG_5__SCAN_IN), .Z(n4140) );
  INV_X1 U5071 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U5072 ( .A1(n4397), .A2(n4386), .ZN(n4139) );
  NAND2_X1 U5073 ( .A1(n4634), .A2(n4633), .ZN(n4712) );
  INV_X1 U5074 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U5075 ( .A1(n4211), .A2(n6247), .ZN(n4144) );
  INV_X1 U5076 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U5077 ( .A1(n4177), .A2(n4318), .ZN(n4142) );
  NAND2_X1 U5078 ( .A1(n4481), .A2(n6247), .ZN(n4141) );
  NAND3_X1 U5079 ( .A1(n4142), .A2(n4133), .A3(n4141), .ZN(n4143) );
  AND2_X1 U5080 ( .A1(n4144), .A2(n4143), .ZN(n4713) );
  INV_X1 U5081 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U5082 ( .A1(n6480), .A2(n4386), .ZN(n4148) );
  MUX2_X1 U5083 ( .A(n4217), .B(n4133), .S(EBX_REG_7__SCAN_IN), .Z(n4147) );
  NAND2_X1 U5084 ( .A1(n4148), .A2(n4147), .ZN(n4894) );
  NOR2_X2 U5085 ( .A1(n4893), .A2(n4894), .ZN(n4892) );
  INV_X1 U5086 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4337) );
  NAND2_X1 U5087 ( .A1(n4177), .A2(n4337), .ZN(n4150) );
  INV_X1 U5088 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U5089 ( .A1(n4481), .A2(n5174), .ZN(n4149) );
  NAND3_X1 U5090 ( .A1(n4150), .A2(n4133), .A3(n4149), .ZN(n4151) );
  OAI21_X1 U5091 ( .B1(n5536), .B2(EBX_REG_8__SCAN_IN), .A(n4151), .ZN(n5153)
         );
  AND2_X2 U5092 ( .A1(n4892), .A2(n5153), .ZN(n5213) );
  MUX2_X1 U5093 ( .A(n4217), .B(n4133), .S(EBX_REG_9__SCAN_IN), .Z(n4153) );
  INV_X1 U5094 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U5095 ( .A1(n6471), .A2(n4386), .ZN(n4152) );
  NAND2_X1 U5096 ( .A1(n5213), .A2(n5212), .ZN(n5211) );
  INV_X1 U5097 ( .A(n5211), .ZN(n4158) );
  MUX2_X1 U5098 ( .A(n5536), .B(n4177), .S(EBX_REG_10__SCAN_IN), .Z(n4156) );
  NAND2_X1 U5099 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4154) );
  AND2_X1 U5100 ( .A1(n4205), .A2(n4154), .ZN(n4155) );
  NAND2_X1 U5101 ( .A1(n4158), .A2(n4157), .ZN(n5290) );
  INV_X1 U5102 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U5103 ( .A1(n4200), .A2(n5187), .ZN(n4161) );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U5105 ( .A1(n4481), .A2(n5187), .ZN(n4159) );
  OAI211_X1 U5106 ( .C1(n5537), .C2(n6462), .A(n4159), .B(n4177), .ZN(n4160)
         );
  NAND2_X1 U5107 ( .A1(n4161), .A2(n4160), .ZN(n5149) );
  MUX2_X1 U5108 ( .A(n5536), .B(n4177), .S(EBX_REG_12__SCAN_IN), .Z(n4166) );
  NAND2_X1 U5109 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4164) );
  AND2_X1 U5110 ( .A1(n4205), .A2(n4164), .ZN(n4165) );
  NOR2_X2 U5111 ( .A1(n5297), .A2(n5296), .ZN(n6138) );
  INV_X1 U5112 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U5113 ( .A1(n4200), .A2(n6321), .ZN(n4169) );
  INV_X1 U5114 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U5115 ( .A1(n4481), .A2(n6321), .ZN(n4167) );
  OAI211_X1 U5116 ( .C1(n5537), .C2(n6142), .A(n4167), .B(n4177), .ZN(n4168)
         );
  NAND2_X1 U5117 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  MUX2_X1 U5118 ( .A(n5536), .B(n4177), .S(EBX_REG_14__SCAN_IN), .Z(n4172) );
  NAND2_X1 U5119 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4170) );
  AND2_X1 U5120 ( .A1(n4205), .A2(n4170), .ZN(n4171) );
  NOR2_X2 U5121 ( .A1(n6139), .A2(n5329), .ZN(n5328) );
  INV_X1 U5122 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U5123 ( .A1(n4200), .A2(n6315), .ZN(n4175) );
  INV_X1 U5124 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U5125 ( .A1(n4481), .A2(n6315), .ZN(n4173) );
  OAI211_X1 U5126 ( .C1(n5537), .C2(n5848), .A(n4173), .B(n4177), .ZN(n4174)
         );
  NAND2_X1 U5127 ( .A1(n4175), .A2(n4174), .ZN(n5851) );
  AND2_X2 U5128 ( .A1(n5328), .A2(n4176), .ZN(n5854) );
  MUX2_X1 U5129 ( .A(n5536), .B(n4177), .S(EBX_REG_16__SCAN_IN), .Z(n4180) );
  NAND2_X1 U5130 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4178) );
  AND2_X1 U5131 ( .A1(n4205), .A2(n4178), .ZN(n4179) );
  NAND2_X1 U5132 ( .A1(n4180), .A2(n4179), .ZN(n5399) );
  AND2_X2 U5133 ( .A1(n5854), .A2(n5399), .ZN(n5549) );
  INV_X1 U5134 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U5135 ( .A1(n4200), .A2(n5619), .ZN(n4183) );
  INV_X1 U5136 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U5137 ( .A1(n4481), .A2(n5619), .ZN(n4181) );
  OAI211_X1 U5138 ( .C1(n5537), .C2(n5711), .A(n4181), .B(n4177), .ZN(n4182)
         );
  NAND2_X1 U5139 ( .A1(n5549), .A2(n5548), .ZN(n5539) );
  MUX2_X1 U5140 ( .A(n5536), .B(n4177), .S(EBX_REG_19__SCAN_IN), .Z(n4186) );
  NAND2_X1 U5141 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4184) );
  AND2_X1 U5142 ( .A1(n4205), .A2(n4184), .ZN(n4185) );
  INV_X1 U5143 ( .A(n4187), .ZN(n5605) );
  INV_X1 U5144 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5662) );
  NOR2_X1 U5145 ( .A1(n4374), .A2(EBX_REG_20__SCAN_IN), .ZN(n4188) );
  AOI21_X1 U5146 ( .B1(n4386), .B2(n5662), .A(n4188), .ZN(n5607) );
  OR2_X1 U5147 ( .A1(n4487), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4190)
         );
  INV_X1 U5148 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U5149 ( .A1(n4481), .A2(n5617), .ZN(n4189) );
  NAND2_X1 U5150 ( .A1(n4190), .A2(n4189), .ZN(n5606) );
  NAND2_X1 U5151 ( .A1(n5537), .A2(EBX_REG_20__SCAN_IN), .ZN(n4192) );
  NAND2_X1 U5152 ( .A1(n5606), .A2(n4133), .ZN(n4191) );
  OAI211_X1 U5153 ( .C1(n5607), .C2(n5606), .A(n4192), .B(n4191), .ZN(n4193)
         );
  NOR2_X2 U5154 ( .A1(n5605), .A2(n4193), .ZN(n5597) );
  MUX2_X1 U5155 ( .A(n4200), .B(n5537), .S(EBX_REG_21__SCAN_IN), .Z(n4195) );
  NOR2_X1 U5156 ( .A1(n4487), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4194)
         );
  NOR2_X1 U5157 ( .A1(n4195), .A2(n4194), .ZN(n5596) );
  NAND2_X1 U5158 ( .A1(n5597), .A2(n5596), .ZN(n5584) );
  MUX2_X1 U5159 ( .A(n5536), .B(n4177), .S(EBX_REG_22__SCAN_IN), .Z(n4198) );
  NAND2_X1 U5160 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4196) );
  AND2_X1 U5161 ( .A1(n4205), .A2(n4196), .ZN(n4197) );
  INV_X1 U5162 ( .A(n4199), .ZN(n5796) );
  INV_X1 U5163 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U5164 ( .A1(n4200), .A2(n6065), .ZN(n4203) );
  NAND2_X1 U5165 ( .A1(n4481), .A2(n6065), .ZN(n4201) );
  OAI211_X1 U5166 ( .C1(n5537), .C2(n5665), .A(n4201), .B(n4177), .ZN(n4202)
         );
  NAND2_X1 U5167 ( .A1(n4203), .A2(n4202), .ZN(n5795) );
  MUX2_X1 U5168 ( .A(n5536), .B(n4177), .S(EBX_REG_24__SCAN_IN), .Z(n4207) );
  NAND2_X1 U5169 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4204) );
  AND2_X1 U5170 ( .A1(n4205), .A2(n4204), .ZN(n4206) );
  NAND2_X1 U5171 ( .A1(n4207), .A2(n4206), .ZN(n5580) );
  NAND2_X1 U5172 ( .A1(n5579), .A2(n5580), .ZN(n5572) );
  MUX2_X1 U5173 ( .A(n4217), .B(n4133), .S(EBX_REG_25__SCAN_IN), .Z(n4209) );
  INV_X1 U5174 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U5175 ( .A1(n4386), .A2(n6106), .ZN(n4208) );
  NAND2_X1 U5176 ( .A1(n4209), .A2(n4208), .ZN(n5573) );
  INV_X1 U5177 ( .A(n4210), .ZN(n5575) );
  INV_X1 U5178 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U5179 ( .A1(n4211), .A2(n5998), .ZN(n4216) );
  INV_X1 U5180 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U5181 ( .A1(n4177), .A2(n4212), .ZN(n4214) );
  NAND2_X1 U5182 ( .A1(n4481), .A2(n5998), .ZN(n4213) );
  NAND3_X1 U5183 ( .A1(n4214), .A2(n4133), .A3(n4213), .ZN(n4215) );
  AND2_X1 U5184 ( .A1(n4216), .A2(n4215), .ZN(n4381) );
  OR2_X2 U5185 ( .A1(n5575), .A2(n4381), .ZN(n5445) );
  MUX2_X1 U5186 ( .A(n4217), .B(n4133), .S(EBX_REG_27__SCAN_IN), .Z(n4218) );
  OAI21_X1 U5187 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4487), .A(n4218), 
        .ZN(n5444) );
  INV_X1 U5188 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U5189 ( .A1(n4177), .A2(n5652), .ZN(n4221) );
  INV_X1 U5190 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4219) );
  NAND2_X1 U5191 ( .A1(n4481), .A2(n4219), .ZN(n4220) );
  NAND3_X1 U5192 ( .A1(n4221), .A2(n4133), .A3(n4220), .ZN(n4222) );
  OAI21_X1 U5193 ( .B1(n5536), .B2(EBX_REG_28__SCAN_IN), .A(n4222), .ZN(n5562)
         );
  INV_X1 U5194 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5772) );
  NOR2_X1 U5195 ( .A1(n4374), .A2(EBX_REG_29__SCAN_IN), .ZN(n4223) );
  AOI21_X1 U5196 ( .B1(n4386), .B2(n5772), .A(n4223), .ZN(n5517) );
  NAND2_X1 U5197 ( .A1(n4224), .A2(n5517), .ZN(n4454) );
  OR2_X1 U5198 ( .A1(n4454), .A2(n5537), .ZN(n4226) );
  NOR2_X1 U5199 ( .A1(n5536), .A2(EBX_REG_29__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U5200 ( .A1(n5565), .A2(n5518), .ZN(n4225) );
  INV_X1 U5201 ( .A(n4454), .ZN(n4452) );
  NOR2_X1 U5202 ( .A1(n4452), .A2(n5537), .ZN(n4457) );
  OAI22_X1 U5203 ( .A1(n4487), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4374), .ZN(n4227) );
  INV_X1 U5204 ( .A(n4227), .ZN(n4228) );
  XNOR2_X2 U5205 ( .A(n4229), .B(n4228), .ZN(n5453) );
  NOR2_X1 U5206 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5168) );
  INV_X1 U5207 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5452) );
  OR2_X1 U5208 ( .A1(n5168), .A2(n5452), .ZN(n4230) );
  NOR2_X1 U5209 ( .A1(n4374), .A2(n4230), .ZN(n4231) );
  INV_X1 U5210 ( .A(n4233), .ZN(n4235) );
  INV_X1 U5211 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U5212 ( .A1(n4235), .A2(n4234), .ZN(n6660) );
  NOR3_X1 U5213 ( .A1(n6660), .A2(READY_N), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n5167) );
  NOR3_X1 U5214 ( .A1(n6720), .A2(n5167), .A3(n5452), .ZN(n4236) );
  AOI22_X1 U5215 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n6245), .B1(n6717), 
        .B2(n4236), .ZN(n4237) );
  OAI21_X1 U5216 ( .B1(n5453), .B2(n6198), .A(n4237), .ZN(n4255) );
  INV_X1 U5217 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6693) );
  INV_X1 U5218 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6698) );
  INV_X1 U5219 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6696) );
  NAND3_X1 U5220 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4243) );
  INV_X1 U5221 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6845) );
  INV_X1 U5222 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U5223 ( .A1(n3345), .A2(n6660), .ZN(n4359) );
  AND3_X1 U5224 ( .A1(n4359), .A2(n5168), .A3(n4361), .ZN(n4238) );
  INV_X1 U5225 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6685) );
  INV_X1 U5226 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6684) );
  INV_X1 U5227 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6681) );
  INV_X1 U5228 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6678) );
  INV_X1 U5229 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6674) );
  NAND3_X1 U5230 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6277) );
  NOR2_X1 U5231 ( .A1(n6674), .A2(n6277), .ZN(n6263) );
  NAND2_X1 U5232 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6263), .ZN(n6234) );
  NOR2_X1 U5233 ( .A1(n6678), .A2(n6234), .ZN(n6239) );
  NAND2_X1 U5234 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6239), .ZN(n5181) );
  NOR2_X1 U5235 ( .A1(n6681), .A2(n5181), .ZN(n5210) );
  NAND3_X1 U5236 ( .A1(n5210), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n6208) );
  NOR2_X1 U5237 ( .A1(n6684), .A2(n6208), .ZN(n5185) );
  NAND2_X1 U5238 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5185), .ZN(n6204) );
  NOR2_X1 U5239 ( .A1(n6685), .A2(n6204), .ZN(n4239) );
  NAND2_X1 U5240 ( .A1(n6264), .A2(n4239), .ZN(n6195) );
  NOR2_X2 U5241 ( .A1(n6686), .A2(n6195), .ZN(n6185) );
  NAND3_X1 U5242 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        n6185), .ZN(n5547) );
  NAND4_X1 U5243 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .A4(n6054), .ZN(n6026) );
  AND2_X1 U5244 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4246) );
  NAND2_X1 U5245 ( .A1(n5981), .A2(n4246), .ZN(n5527) );
  AND2_X1 U5246 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4250) );
  NAND2_X1 U5247 ( .A1(n6278), .A2(n6232), .ZN(n6271) );
  NAND3_X1 U5248 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4239), .A3(n6232), .ZN(
        n6175) );
  NAND2_X1 U5249 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6180) );
  OR2_X1 U5250 ( .A1(n6175), .A2(n6180), .ZN(n4240) );
  OAI21_X1 U5251 ( .B1(n4240), .B2(n6845), .A(n6271), .ZN(n6055) );
  NAND3_X1 U5252 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U5253 ( .A1(n6264), .A2(n4241), .ZN(n4242) );
  NAND2_X1 U5254 ( .A1(n6055), .A2(n4242), .ZN(n6046) );
  AOI21_X1 U5255 ( .B1(n6271), .B2(n4243), .A(n6046), .ZN(n6025) );
  NAND3_X1 U5256 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U5257 ( .A1(n6271), .A2(n4244), .ZN(n4245) );
  INV_X1 U5258 ( .A(n4246), .ZN(n4247) );
  NAND2_X1 U5259 ( .A1(n6264), .A2(n4247), .ZN(n4248) );
  NAND2_X1 U5260 ( .A1(n5992), .A2(n4248), .ZN(n5972) );
  INV_X1 U5261 ( .A(n5972), .ZN(n4249) );
  OAI21_X1 U5262 ( .B1(n5527), .B2(n4250), .A(n4249), .ZN(n5511) );
  INV_X1 U5263 ( .A(n4250), .ZN(n4251) );
  NOR3_X1 U5264 ( .A1(n5527), .A2(REIP_REG_31__SCAN_IN), .A3(n4251), .ZN(n4252) );
  OAI21_X1 U5265 ( .B1(n4257), .B2(n6236), .A(n4256), .ZN(U2796) );
  INV_X1 U5266 ( .A(n4308), .ZN(n4322) );
  NAND2_X4 U5267 ( .A1(n4314), .A2(n4259), .ZN(n4260) );
  NOR2_X1 U5268 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5433)
         );
  INV_X1 U5269 ( .A(n5433), .ZN(n4261) );
  NAND2_X1 U5270 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U5271 ( .A1(n4261), .A2(n4430), .ZN(n4356) );
  NAND2_X1 U5272 ( .A1(n3171), .A2(n4322), .ZN(n4267) );
  NAND2_X1 U5273 ( .A1(n4278), .A2(n4269), .ZN(n4268) );
  NAND2_X1 U5274 ( .A1(n4268), .A2(n4263), .ZN(n4287) );
  OAI21_X1 U5275 ( .B1(n4263), .B2(n4268), .A(n4287), .ZN(n4265) );
  AND2_X1 U5276 ( .A1(n4688), .A2(n4264), .ZN(n4276) );
  AOI21_X1 U5277 ( .B1(n4265), .B2(n6354), .A(n4276), .ZN(n4266) );
  NAND2_X1 U5278 ( .A1(n4267), .A2(n4266), .ZN(n4283) );
  NAND2_X1 U5279 ( .A1(n4283), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6437)
         );
  NAND2_X1 U5280 ( .A1(n4572), .A2(n4322), .ZN(n4275) );
  OAI21_X1 U5281 ( .B1(n4269), .B2(n4278), .A(n4268), .ZN(n4272) );
  INV_X1 U5282 ( .A(n4387), .ZN(n4271) );
  OAI211_X1 U5283 ( .C1(n4272), .C2(n6720), .A(n4271), .B(n4270), .ZN(n4273)
         );
  INV_X1 U5284 ( .A(n4273), .ZN(n4274) );
  NAND2_X1 U5285 ( .A1(n4275), .A2(n4274), .ZN(n4623) );
  INV_X1 U5286 ( .A(n4276), .ZN(n4277) );
  OAI21_X1 U5287 ( .B1(n6720), .B2(n4278), .A(n4277), .ZN(n4279) );
  INV_X1 U5288 ( .A(n4279), .ZN(n4280) );
  OAI21_X1 U5289 ( .B1(n5077), .B2(n4308), .A(n4280), .ZN(n4493) );
  NAND2_X1 U5290 ( .A1(n4493), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4495)
         );
  XNOR2_X1 U5291 ( .A(n4495), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4624)
         );
  NAND2_X1 U5292 ( .A1(n4623), .A2(n4624), .ZN(n4622) );
  OR2_X1 U5293 ( .A1(n4495), .A2(n4281), .ZN(n4282) );
  NAND2_X1 U5294 ( .A1(n6437), .A2(n6440), .ZN(n4286) );
  INV_X1 U5295 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U5296 ( .A1(n4287), .A2(n4288), .ZN(n4304) );
  OAI211_X1 U5297 ( .C1(n4288), .C2(n4287), .A(n4304), .B(n6354), .ZN(n4289)
         );
  OAI21_X2 U5298 ( .B1(n4290), .B2(n4308), .A(n4289), .ZN(n4291) );
  XNOR2_X1 U5299 ( .A(n4291), .B(n4114), .ZN(n4597) );
  NAND2_X1 U5300 ( .A1(n4596), .A2(n4597), .ZN(n4293) );
  NAND2_X1 U5301 ( .A1(n4291), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4292)
         );
  NAND2_X1 U5302 ( .A1(n4294), .A2(n4322), .ZN(n4297) );
  XNOR2_X1 U5303 ( .A(n4304), .B(n4302), .ZN(n4295) );
  NAND2_X1 U5304 ( .A1(n4295), .A2(n6354), .ZN(n4296) );
  NAND2_X1 U5305 ( .A1(n4297), .A2(n4296), .ZN(n4299) );
  NAND2_X1 U5306 ( .A1(n4642), .A2(n4643), .ZN(n4301) );
  NAND2_X1 U5307 ( .A1(n4299), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4300)
         );
  NAND2_X1 U5308 ( .A1(n4301), .A2(n4300), .ZN(n4638) );
  INV_X1 U5309 ( .A(n4302), .ZN(n4303) );
  NOR2_X1 U5310 ( .A1(n4304), .A2(n4303), .ZN(n4306) );
  NAND2_X1 U5311 ( .A1(n4306), .A2(n4305), .ZN(n4324) );
  OAI211_X1 U5312 ( .C1(n4306), .C2(n4305), .A(n4324), .B(n6354), .ZN(n4307)
         );
  OAI21_X1 U5313 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(n4310) );
  NAND2_X1 U5314 ( .A1(n4310), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4311)
         );
  NAND2_X1 U5315 ( .A1(n4312), .A2(n4311), .ZN(n4829) );
  NAND3_X1 U5316 ( .A1(n4314), .A2(n4322), .A3(n4313), .ZN(n4317) );
  XNOR2_X1 U5317 ( .A(n4324), .B(n4325), .ZN(n4315) );
  NAND2_X1 U5318 ( .A1(n4315), .A2(n6354), .ZN(n4316) );
  NAND2_X1 U5319 ( .A1(n4317), .A2(n4316), .ZN(n4319) );
  XNOR2_X1 U5320 ( .A(n4319), .B(n4318), .ZN(n4830) );
  NAND2_X1 U5321 ( .A1(n4829), .A2(n4830), .ZN(n4321) );
  NAND2_X1 U5322 ( .A1(n4319), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4320)
         );
  NAND2_X1 U5323 ( .A1(n4323), .A2(n4322), .ZN(n4329) );
  INV_X1 U5324 ( .A(n4324), .ZN(n4326) );
  NAND2_X1 U5325 ( .A1(n4326), .A2(n4325), .ZN(n4333) );
  XNOR2_X1 U5326 ( .A(n4333), .B(n4334), .ZN(n4327) );
  NAND2_X1 U5327 ( .A1(n4327), .A2(n6354), .ZN(n4328) );
  NAND2_X1 U5328 ( .A1(n4329), .A2(n4328), .ZN(n4330) );
  NAND2_X1 U5329 ( .A1(n5228), .A2(n5229), .ZN(n4332) );
  NAND2_X1 U5330 ( .A1(n4330), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4331)
         );
  NAND2_X1 U5331 ( .A1(n4332), .A2(n4331), .ZN(n5158) );
  INV_X1 U5332 ( .A(n4333), .ZN(n4335) );
  NAND3_X1 U5333 ( .A1(n4335), .A2(n6354), .A3(n4334), .ZN(n4336) );
  NAND2_X1 U5334 ( .A1(n4260), .A2(n4336), .ZN(n4338) );
  NAND2_X1 U5335 ( .A1(n4338), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4339)
         );
  NAND2_X1 U5336 ( .A1(n4260), .A2(n6471), .ZN(n4340) );
  NAND2_X1 U5337 ( .A1(n4341), .A2(n4340), .ZN(n5332) );
  INV_X1 U5338 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5347) );
  AND2_X1 U5339 ( .A1(n4260), .A2(n5347), .ZN(n5333) );
  NAND2_X1 U5340 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U5341 ( .A1(n4260), .A2(n6462), .ZN(n5759) );
  NAND2_X1 U5342 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5760) );
  INV_X1 U5343 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4342) );
  NOR2_X1 U5344 ( .A1(n4260), .A2(n4342), .ZN(n5752) );
  NAND2_X1 U5345 ( .A1(n4260), .A2(n4342), .ZN(n5750) );
  XNOR2_X1 U5346 ( .A(n4260), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5744)
         );
  NAND2_X1 U5347 ( .A1(n4260), .A2(n6142), .ZN(n4343) );
  NAND2_X1 U5348 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4344) );
  INV_X1 U5349 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U5350 ( .A1(n4260), .A2(n5866), .ZN(n4345) );
  NAND2_X1 U5351 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5729) );
  INV_X1 U5352 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5353 ( .A1(n4260), .A2(n5708), .ZN(n4346) );
  NAND2_X1 U5354 ( .A1(n5707), .A2(n4346), .ZN(n5677) );
  INV_X1 U5355 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6123) );
  AND3_X1 U5356 ( .A1(n5708), .A2(n6123), .A3(n5711), .ZN(n4347) );
  NAND2_X1 U5357 ( .A1(n5677), .A2(n4347), .ZN(n4348) );
  NAND2_X1 U5358 ( .A1(n4348), .A2(n5719), .ZN(n4351) );
  INV_X1 U5359 ( .A(n5677), .ZN(n4349) );
  NAND2_X1 U5360 ( .A1(n4349), .A2(n3198), .ZN(n4350) );
  NOR2_X1 U5361 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5821) );
  NOR2_X1 U5362 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5807) );
  INV_X1 U5363 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5788) );
  NAND4_X1 U5364 ( .A1(n5821), .A2(n5807), .A3(n5665), .A4(n5788), .ZN(n4352)
         );
  OAI21_X1 U5365 ( .B1(n5658), .B2(n4352), .A(n5719), .ZN(n4354) );
  AND2_X1 U5366 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5808) );
  AND2_X1 U5367 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5822) );
  AND2_X1 U5368 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U5369 ( .A1(n5658), .A2(n3176), .ZN(n4353) );
  NAND2_X1 U5370 ( .A1(n4260), .A2(n6106), .ZN(n4355) );
  XOR2_X1 U5371 ( .A(n4356), .B(n5649), .Z(n5431) );
  NAND2_X1 U5372 ( .A1(n4358), .A2(n4357), .ZN(n4533) );
  NAND2_X1 U5373 ( .A1(n4359), .A2(n6828), .ZN(n4362) );
  OAI211_X1 U5374 ( .C1(n4533), .C2(n4362), .A(n4361), .B(n4360), .ZN(n4363)
         );
  NAND2_X1 U5375 ( .A1(n4363), .A2(n3332), .ZN(n4373) );
  NOR2_X1 U5376 ( .A1(n6603), .A2(n3345), .ZN(n4396) );
  NAND2_X1 U5377 ( .A1(n5495), .A2(n4396), .ZN(n4370) );
  NAND2_X1 U5378 ( .A1(n3360), .A2(n6354), .ZN(n4365) );
  NAND2_X1 U5379 ( .A1(n4364), .A2(n4365), .ZN(n4392) );
  INV_X1 U5380 ( .A(n4392), .ZN(n4367) );
  AOI21_X1 U5381 ( .B1(n6603), .B2(n4688), .A(n4387), .ZN(n4366) );
  NAND2_X1 U5382 ( .A1(n4367), .A2(n4377), .ZN(n4368) );
  NAND2_X1 U5383 ( .A1(n4368), .A2(n5500), .ZN(n4520) );
  NAND2_X1 U5384 ( .A1(n4384), .A2(n6660), .ZN(n5498) );
  NOR2_X1 U5385 ( .A1(READY_N), .A2(n5501), .ZN(n4418) );
  NAND3_X1 U5386 ( .A1(n5498), .A2(n4418), .A3(n4385), .ZN(n4369) );
  NAND3_X1 U5387 ( .A1(n4370), .A2(n4520), .A3(n4369), .ZN(n4371) );
  NAND2_X1 U5388 ( .A1(n4371), .A2(n6645), .ZN(n4372) );
  NAND2_X1 U5389 ( .A1(n4377), .A2(n5493), .ZN(n5488) );
  OR2_X1 U5390 ( .A1(n4533), .A2(n4374), .ZN(n4423) );
  OAI211_X1 U5391 ( .C1(n4666), .C2(n3172), .A(n5488), .B(n4423), .ZN(n4375)
         );
  INV_X1 U5392 ( .A(n4375), .ZN(n4378) );
  INV_X1 U5393 ( .A(n4436), .ZN(n6621) );
  NAND3_X1 U5394 ( .A1(n4378), .A2(n6621), .A3(n4534), .ZN(n4379) );
  INV_X1 U5395 ( .A(n5445), .ZN(n4380) );
  AOI21_X1 U5396 ( .B1(n4381), .B2(n5575), .A(n4380), .ZN(n5995) );
  NAND2_X1 U5397 ( .A1(n4426), .A2(n4666), .ZN(n4382) );
  OAI21_X1 U5398 ( .B1(n4532), .B2(n4382), .A(n6632), .ZN(n4383) );
  AND2_X2 U5399 ( .A1(n4403), .A2(n4383), .ZN(n6499) );
  NAND2_X1 U5400 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5843) );
  NOR2_X1 U5401 ( .A1(n6462), .A2(n4342), .ZN(n6136) );
  NAND2_X1 U5402 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6136), .ZN(n5862) );
  NOR2_X1 U5403 ( .A1(n5866), .A2(n5862), .ZN(n5838) );
  NAND2_X1 U5404 ( .A1(n4688), .A2(n4384), .ZN(n5198) );
  OR2_X1 U5405 ( .A1(n5198), .A2(n4385), .ZN(n4519) );
  NAND2_X1 U5406 ( .A1(n4386), .A2(n4519), .ZN(n4388) );
  NAND2_X1 U5407 ( .A1(n4388), .A2(n4387), .ZN(n4391) );
  OR2_X1 U5408 ( .A1(n4389), .A2(n3332), .ZN(n4390) );
  OAI211_X1 U5409 ( .C1(n3359), .C2(n4133), .A(n4391), .B(n4390), .ZN(n4393)
         );
  NOR2_X1 U5410 ( .A1(n4393), .A2(n4392), .ZN(n4394) );
  NAND2_X1 U5411 ( .A1(n4403), .A2(n5487), .ZN(n5835) );
  NAND2_X1 U5412 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5882) );
  NOR2_X1 U5413 ( .A1(n4397), .A2(n5882), .ZN(n4883) );
  NAND2_X1 U5414 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4883), .ZN(n5160)
         );
  NOR2_X1 U5415 ( .A1(n6480), .A2(n4337), .ZN(n5162) );
  INV_X1 U5416 ( .A(n5162), .ZN(n5342) );
  NAND2_X1 U5417 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5343) );
  NOR3_X1 U5418 ( .A1(n5160), .A2(n5342), .A3(n5343), .ZN(n4398) );
  NAND2_X1 U5419 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U5420 ( .A1(n4284), .A2(n6483), .ZN(n6482) );
  NAND2_X1 U5421 ( .A1(n4398), .A2(n6482), .ZN(n5833) );
  NOR2_X1 U5422 ( .A1(n5835), .A2(n5833), .ZN(n5864) );
  NOR2_X1 U5423 ( .A1(n4284), .A2(n4281), .ZN(n4614) );
  AND2_X1 U5424 ( .A1(n4614), .A2(n4398), .ZN(n4404) );
  OR2_X1 U5425 ( .A1(n5500), .A2(n3345), .ZN(n5895) );
  INV_X1 U5426 ( .A(n5895), .ZN(n6604) );
  OAI211_X1 U5427 ( .C1(n4531), .C2(n5497), .A(n4536), .B(n4553), .ZN(n4399)
         );
  NAND2_X1 U5428 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4400)
         );
  NAND2_X1 U5429 ( .A1(n6124), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6115) );
  INV_X1 U5430 ( .A(n5822), .ZN(n4401) );
  NAND2_X1 U5431 ( .A1(n5806), .A2(n5808), .ZN(n5804) );
  INV_X1 U5432 ( .A(n4402), .ZN(n4410) );
  NAND2_X1 U5433 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5410) );
  OAI211_X1 U5434 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6107), .B(n5410), .ZN(n4413) );
  INV_X2 U5435 ( .A(n6259), .ZN(n6503) );
  NAND3_X1 U5436 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5838), .ZN(n5825) );
  INV_X1 U5437 ( .A(n4405), .ZN(n4615) );
  INV_X1 U5438 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6494) );
  NOR2_X1 U5439 ( .A1(n4403), .A2(n6503), .ZN(n4497) );
  AOI21_X1 U5440 ( .B1(n5865), .B2(n6494), .A(n4497), .ZN(n4613) );
  OAI21_X1 U5441 ( .B1(n4615), .B2(n4404), .A(n4613), .ZN(n5837) );
  AOI21_X1 U5442 ( .B1(n4405), .B2(n5825), .A(n5837), .ZN(n5827) );
  INV_X1 U5443 ( .A(n5835), .ZN(n6486) );
  NOR2_X1 U5444 ( .A1(n5825), .A2(n5833), .ZN(n4406) );
  NAND2_X1 U5445 ( .A1(n4406), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U5446 ( .A1(n5822), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5678) );
  NOR2_X1 U5447 ( .A1(n5826), .A2(n5678), .ZN(n4407) );
  OR2_X1 U5448 ( .A1(n5839), .A2(n4407), .ZN(n4408) );
  NAND2_X1 U5449 ( .A1(n5827), .A2(n4408), .ZN(n5816) );
  NOR2_X1 U5450 ( .A1(n5839), .A2(n5808), .ZN(n4409) );
  NOR2_X1 U5451 ( .A1(n5816), .A2(n4409), .ZN(n5799) );
  OAI21_X1 U5452 ( .B1(n6489), .B2(n6486), .A(n4410), .ZN(n4411) );
  NAND2_X1 U5453 ( .A1(n5799), .A2(n4411), .ZN(n6105) );
  AOI22_X1 U5454 ( .A1(n6503), .A2(REIP_REG_26__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6105), .ZN(n4412) );
  XNOR2_X1 U5455 ( .A(n5515), .B(n4417), .ZN(n5464) );
  INV_X1 U5456 ( .A(n4418), .ZN(n4419) );
  OAI22_X1 U5457 ( .A1(n5495), .A2(n5488), .B1(n4534), .B2(n4419), .ZN(n4514)
         );
  INV_X1 U5458 ( .A(n4449), .ZN(n5480) );
  NAND4_X1 U5459 ( .A1(n3332), .A2(n5480), .A3(n4679), .A4(n4666), .ZN(n4421)
         );
  NOR2_X1 U5460 ( .A1(n4421), .A2(n4420), .ZN(n4446) );
  AND2_X1 U5461 ( .A1(n5493), .A2(n4446), .ZN(n4422) );
  NOR2_X1 U5462 ( .A1(n4423), .A2(READY_N), .ZN(n4517) );
  NAND2_X1 U5463 ( .A1(n4425), .A2(n4449), .ZN(n4593) );
  NAND2_X2 U5464 ( .A1(n5481), .A2(n4593), .ZN(n6066) );
  AOI22_X1 U5465 ( .A1(n6323), .A2(DATAI_30_), .B1(n6326), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4429) );
  AND2_X1 U5466 ( .A1(n4661), .A2(n4449), .ZN(n4427) );
  NAND2_X1 U5467 ( .A1(n6327), .A2(DATAI_14_), .ZN(n4428) );
  OAI21_X1 U5468 ( .B1(n5513), .B2(n6066), .A(n3201), .ZN(U2861) );
  NOR2_X2 U5469 ( .A1(n5649), .A2(n4430), .ZN(n5435) );
  AND2_X1 U5470 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U5471 ( .A1(n5435), .A2(n5417), .ZN(n5642) );
  NAND2_X1 U5472 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4434) );
  INV_X1 U5473 ( .A(n4431), .ZN(n6079) );
  NOR2_X1 U5474 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4432) );
  AND2_X1 U5475 ( .A1(n5433), .A2(n4432), .ZN(n5454) );
  INV_X1 U5476 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5457) );
  NAND4_X1 U5477 ( .A1(n6079), .A2(n5454), .A3(n5457), .A4(n5772), .ZN(n4433)
         );
  XNOR2_X1 U5478 ( .A(n4435), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5422)
         );
  NAND2_X1 U5479 ( .A1(n4437), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6652) );
  NOR2_X2 U5480 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5917) );
  INV_X2 U5481 ( .A(n6454), .ZN(n6441) );
  NAND2_X1 U5482 ( .A1(n5483), .A2(n6441), .ZN(n4445) );
  NAND2_X1 U5483 ( .A1(n6517), .A2(n4438), .ZN(n6718) );
  NAND2_X1 U5484 ( .A1(n6718), .A2(n4654), .ZN(n4439) );
  NAND2_X1 U5485 ( .A1(n4654), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4441) );
  NAND2_X1 U5486 ( .A1(n7092), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4440) );
  NAND2_X1 U5487 ( .A1(n4441), .A2(n4440), .ZN(n6447) );
  INV_X1 U5488 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7057) );
  NOR2_X1 U5489 ( .A1(n6120), .A2(n7057), .ZN(n5415) );
  AOI21_X1 U5490 ( .B1(n6448), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5415), 
        .ZN(n4442) );
  OAI21_X1 U5491 ( .B1(n6446), .B2(n5176), .A(n4442), .ZN(n4443) );
  INV_X1 U5492 ( .A(n4443), .ZN(n4444) );
  OAI211_X1 U5493 ( .C1(n5422), .C2(n6161), .A(n4445), .B(n4444), .ZN(U2955)
         );
  NAND2_X1 U5494 ( .A1(n5487), .A2(n5495), .ZN(n4525) );
  NAND2_X1 U5495 ( .A1(n4446), .A2(n4481), .ZN(n4447) );
  NAND2_X1 U5496 ( .A1(n4525), .A2(n4447), .ZN(n4448) );
  INV_X1 U5497 ( .A(n5565), .ZN(n4451) );
  INV_X1 U5498 ( .A(n4453), .ZN(n4450) );
  OAI21_X1 U5499 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4456) );
  OAI211_X1 U5500 ( .C1(n5565), .C2(n4133), .A(n4454), .B(n4453), .ZN(n4455)
         );
  OAI21_X1 U5501 ( .B1(n4457), .B2(n4456), .A(n4455), .ZN(n5508) );
  INV_X1 U5502 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4458) );
  INV_X1 U5503 ( .A(n4462), .ZN(n6155) );
  INV_X1 U5504 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6884) );
  NOR2_X1 U5505 ( .A1(n6517), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4464) );
  INV_X1 U5506 ( .A(n4464), .ZN(n4463) );
  OAI211_X1 U5507 ( .C1(n6155), .C2(n6884), .A(n6352), .B(n4463), .ZN(U2788)
         );
  NOR2_X1 U5508 ( .A1(n4464), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4466) );
  NAND3_X1 U5509 ( .A1(n6717), .A2(n6720), .A3(n5198), .ZN(n4465) );
  OAI21_X1 U5510 ( .B1(n6717), .B2(n4466), .A(n4465), .ZN(U3474) );
  INV_X1 U5511 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U5512 ( .A1(n5895), .A2(n6632), .ZN(n4467) );
  INV_X1 U5513 ( .A(n6660), .ZN(n4515) );
  NAND2_X1 U5514 ( .A1(n4467), .A2(n4515), .ZN(n4468) );
  AOI22_X1 U5515 ( .A1(n6719), .A2(UWORD_REG_9__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5516 ( .B1(n6375), .B2(n4585), .A(n4470), .ZN(U2898) );
  INV_X1 U5517 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6377) );
  AOI22_X1 U5518 ( .A1(n6719), .A2(UWORD_REG_10__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4471) );
  OAI21_X1 U5519 ( .B1(n6377), .B2(n4585), .A(n4471), .ZN(U2897) );
  INV_X1 U5520 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6373) );
  AOI22_X1 U5521 ( .A1(n6719), .A2(UWORD_REG_8__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5522 ( .B1(n6373), .B2(n4585), .A(n4472), .ZN(U2899) );
  INV_X1 U5523 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6381) );
  AOI22_X1 U5524 ( .A1(n6719), .A2(UWORD_REG_12__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4473) );
  OAI21_X1 U5525 ( .B1(n6381), .B2(n4585), .A(n4473), .ZN(U2895) );
  INV_X1 U5526 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6383) );
  AOI22_X1 U5527 ( .A1(n6719), .A2(UWORD_REG_13__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5528 ( .B1(n6383), .B2(n4585), .A(n4474), .ZN(U2894) );
  INV_X1 U5529 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6379) );
  AOI22_X1 U5530 ( .A1(n6719), .A2(UWORD_REG_11__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4475) );
  OAI21_X1 U5531 ( .B1(n6379), .B2(n4585), .A(n4475), .ZN(U2896) );
  INV_X1 U5532 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6385) );
  AOI22_X1 U5533 ( .A1(n6719), .A2(UWORD_REG_14__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4476) );
  OAI21_X1 U5534 ( .B1(n6385), .B2(n4585), .A(n4476), .ZN(U2893) );
  OAI21_X1 U5535 ( .B1(n4478), .B2(n4477), .A(n3488), .ZN(n5311) );
  OAI21_X1 U5536 ( .B1(n5308), .B2(n4481), .A(n4480), .ZN(n6500) );
  AOI22_X1 U5537 ( .A1(n6317), .A2(n6500), .B1(EBX_REG_1__SCAN_IN), .B2(n5613), 
        .ZN(n4482) );
  OAI21_X1 U5538 ( .B1(n5311), .B2(n6311), .A(n4482), .ZN(U2858) );
  OAI21_X1 U5539 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(n6455) );
  INV_X1 U5540 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5279) );
  OAI21_X1 U5541 ( .B1(n4487), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4486), 
        .ZN(n5278) );
  OAI222_X1 U5542 ( .A1(n6455), .A2(n6311), .B1(n5279), .B2(n6322), .C1(n5278), 
        .C2(n6310), .ZN(U2859) );
  NOR2_X1 U5543 ( .A1(n4489), .A2(n4490), .ZN(n4491) );
  NOR2_X1 U5544 ( .A1(n4488), .A2(n4491), .ZN(n6442) );
  INV_X1 U5545 ( .A(n6442), .ZN(n5206) );
  XNOR2_X1 U5546 ( .A(n4505), .B(n4507), .ZN(n6484) );
  AOI22_X1 U5547 ( .A1(n6317), .A2(n6484), .B1(EBX_REG_2__SCAN_IN), .B2(n5613), 
        .ZN(n4492) );
  OAI21_X1 U5548 ( .B1(n5206), .B2(n6311), .A(n4492), .ZN(U2857) );
  OR2_X1 U5549 ( .A1(n4493), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4494)
         );
  AND2_X1 U5550 ( .A1(n4495), .A2(n4494), .ZN(n6451) );
  INV_X1 U5551 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4496) );
  OR2_X1 U5552 ( .A1(n6120), .A2(n4496), .ZN(n6452) );
  OAI21_X1 U5553 ( .B1(n5869), .B2(n5278), .A(n6452), .ZN(n4500) );
  NOR2_X1 U5554 ( .A1(n6486), .A2(n5865), .ZN(n5860) );
  INV_X1 U5555 ( .A(n5860), .ZN(n4498) );
  AOI21_X1 U5556 ( .B1(n6494), .B2(n4498), .A(n4497), .ZN(n6505) );
  AOI22_X1 U5557 ( .A1(n6505), .A2(n6495), .B1(n5860), .B2(n6494), .ZN(n4499)
         );
  AOI211_X1 U5558 ( .C1(n6502), .C2(n6451), .A(n4500), .B(n4499), .ZN(n4501)
         );
  INV_X1 U5559 ( .A(n4501), .ZN(U3018) );
  OR2_X1 U5560 ( .A1(n4488), .A2(n4502), .ZN(n4504) );
  AND2_X1 U5561 ( .A1(n4504), .A2(n4503), .ZN(n6304) );
  INV_X1 U5562 ( .A(n6304), .ZN(n4595) );
  AOI21_X1 U5563 ( .B1(n4131), .B2(n4507), .A(n4506), .ZN(n4509) );
  INV_X1 U5564 ( .A(n4590), .ZN(n4508) );
  NOR2_X1 U5565 ( .A1(n4509), .A2(n4508), .ZN(n6296) );
  AOI22_X1 U5566 ( .A1(n6317), .A2(n6296), .B1(EBX_REG_3__SCAN_IN), .B2(n5613), 
        .ZN(n4510) );
  OAI21_X1 U5567 ( .B1(n4595), .B2(n6311), .A(n4510), .ZN(U2856) );
  INV_X1 U5568 ( .A(n4897), .ZN(n4787) );
  NOR2_X1 U5569 ( .A1(n4511), .A2(n4787), .ZN(n4512) );
  XNOR2_X1 U5570 ( .A(n4512), .B(n3543), .ZN(n6276) );
  NOR2_X1 U5571 ( .A1(n4534), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5572 ( .A1(n6276), .A2(n4513), .ZN(n6150) );
  INV_X1 U5573 ( .A(n4514), .ZN(n4524) );
  INV_X1 U5574 ( .A(n5495), .ZN(n5486) );
  INV_X1 U5575 ( .A(READY_N), .ZN(n6828) );
  NAND2_X1 U5576 ( .A1(n4515), .A2(n6828), .ZN(n4516) );
  AOI21_X1 U5577 ( .B1(n5895), .B2(n4533), .A(n4516), .ZN(n4518) );
  OR2_X1 U5578 ( .A1(n4518), .A2(n4517), .ZN(n4522) );
  NAND2_X1 U5579 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  AOI21_X1 U5580 ( .B1(n5486), .B2(n4522), .A(n4521), .ZN(n4523) );
  MUX2_X1 U5581 ( .A(n6611), .B(n6858), .S(STATE2_REG_1__SCAN_IN), .Z(n4526)
         );
  NAND2_X1 U5582 ( .A1(n4526), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4527) );
  INV_X1 U5583 ( .A(n4564), .ZN(n4569) );
  INV_X1 U5584 ( .A(n4528), .ZN(n4568) );
  INV_X1 U5585 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6858) );
  NAND2_X1 U5586 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6858), .ZN(n4567) );
  INV_X1 U5587 ( .A(n4546), .ZN(n4566) );
  AND4_X1 U5588 ( .A1(n4534), .A2(n4533), .A3(n4532), .A4(n4531), .ZN(n4535)
         );
  NAND2_X1 U5589 ( .A1(n4536), .A2(n4535), .ZN(n6608) );
  NAND2_X1 U5590 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4538) );
  INV_X1 U5591 ( .A(n4538), .ZN(n4537) );
  MUX2_X1 U5592 ( .A(n4538), .B(n4537), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4541) );
  OAI21_X1 U5593 ( .B1(n4540), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3394), 
        .ZN(n5903) );
  OAI22_X1 U5594 ( .A1(n5895), .A2(n4541), .B1(n4553), .B2(n5903), .ZN(n4549)
         );
  INV_X1 U5595 ( .A(n5487), .ZN(n4542) );
  NAND2_X1 U5596 ( .A1(n4542), .A2(n5488), .ZN(n4557) );
  INV_X1 U5597 ( .A(n4557), .ZN(n4547) );
  MUX2_X1 U5598 ( .A(n4544), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4543), 
        .Z(n4545) );
  NOR3_X1 U5599 ( .A1(n4547), .A2(n4546), .A3(n4545), .ZN(n4548) );
  AOI211_X1 U5600 ( .C1(n4530), .C2(n6608), .A(n4549), .B(n4548), .ZN(n5905)
         );
  NAND2_X1 U5601 ( .A1(n6611), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4550) );
  OAI21_X1 U5602 ( .B1(n6611), .B2(n5905), .A(n4550), .ZN(n6618) );
  NAND2_X1 U5603 ( .A1(n4552), .A2(n6608), .ZN(n4559) );
  XNOR2_X1 U5604 ( .A(n4543), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4556)
         );
  XNOR2_X1 U5605 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4554) );
  OAI22_X1 U5606 ( .A1(n5895), .A2(n4554), .B1(n4553), .B2(n4556), .ZN(n4555)
         );
  AOI21_X1 U5607 ( .B1(n4557), .B2(n4556), .A(n4555), .ZN(n4558) );
  NAND2_X1 U5608 ( .A1(n4559), .A2(n4558), .ZN(n5407) );
  INV_X1 U5609 ( .A(n6611), .ZN(n4560) );
  NAND2_X1 U5610 ( .A1(n5407), .A2(n4560), .ZN(n4562) );
  NAND2_X1 U5611 ( .A1(n6611), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4561) );
  INV_X1 U5612 ( .A(n6615), .ZN(n4563) );
  NAND3_X1 U5613 ( .A1(n6618), .A2(n5472), .A3(n4563), .ZN(n4565) );
  OAI211_X1 U5614 ( .C1(n4567), .C2(n4566), .A(n4565), .B(n4564), .ZN(n6626)
         );
  OAI21_X1 U5615 ( .B1(n4569), .B2(n4568), .A(n6626), .ZN(n4609) );
  NAND2_X1 U5616 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4608), .ZN(n6706) );
  AOI21_X1 U5617 ( .B1(n4609), .B2(n6858), .A(n6706), .ZN(n4570) );
  NAND2_X1 U5618 ( .A1(n4573), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U5619 ( .A(n4571), .B(n5889), .ZN(n4574) );
  NAND2_X1 U5620 ( .A1(n5471), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5621 ( .A1(n4574), .A2(n5917), .B1(n4604), .B2(n4552), .ZN(n4576)
         );
  NAND2_X1 U5622 ( .A1(n6507), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5623 ( .B1(n6507), .B2(n4576), .A(n4575), .ZN(U3463) );
  INV_X1 U5624 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6371) );
  AOI22_X1 U5625 ( .A1(n6719), .A2(UWORD_REG_7__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5626 ( .B1(n6371), .B2(n4585), .A(n4577), .ZN(U2900) );
  INV_X1 U5627 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6369) );
  AOI22_X1 U5628 ( .A1(n6719), .A2(UWORD_REG_6__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U5629 ( .B1(n6369), .B2(n4585), .A(n4578), .ZN(U2901) );
  INV_X1 U5630 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6361) );
  AOI22_X1 U5631 ( .A1(n6719), .A2(UWORD_REG_2__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U5632 ( .B1(n6361), .B2(n4585), .A(n4579), .ZN(U2905) );
  INV_X1 U5633 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6367) );
  AOI22_X1 U5634 ( .A1(n6719), .A2(UWORD_REG_5__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4580) );
  OAI21_X1 U5635 ( .B1(n6367), .B2(n4585), .A(n4580), .ZN(U2902) );
  INV_X1 U5636 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6365) );
  AOI22_X1 U5637 ( .A1(n6719), .A2(UWORD_REG_4__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4581) );
  OAI21_X1 U5638 ( .B1(n6365), .B2(n4585), .A(n4581), .ZN(U2903) );
  INV_X1 U5639 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6363) );
  AOI22_X1 U5640 ( .A1(n6719), .A2(UWORD_REG_3__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4582) );
  OAI21_X1 U5641 ( .B1(n6363), .B2(n4585), .A(n4582), .ZN(U2904) );
  INV_X1 U5642 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6357) );
  AOI22_X1 U5643 ( .A1(n6719), .A2(UWORD_REG_0__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4583) );
  OAI21_X1 U5644 ( .B1(n6357), .B2(n4585), .A(n4583), .ZN(U2907) );
  INV_X1 U5645 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6359) );
  AOI22_X1 U5646 ( .A1(n6719), .A2(UWORD_REG_1__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4584) );
  OAI21_X1 U5647 ( .B1(n6359), .B2(n4585), .A(n4584), .ZN(U2906) );
  CLKBUF_X1 U5648 ( .A(n4586), .Z(n4587) );
  AND2_X1 U5649 ( .A1(n4503), .A2(n4588), .ZN(n4589) );
  OR2_X1 U5650 ( .A1(n4587), .A2(n4589), .ZN(n6275) );
  AOI21_X1 U5651 ( .B1(n4591), .B2(n4590), .A(n4634), .ZN(n6280) );
  AOI22_X1 U5652 ( .A1(n6317), .A2(n6280), .B1(EBX_REG_4__SCAN_IN), .B2(n5613), 
        .ZN(n4592) );
  OAI21_X1 U5653 ( .B1(n6275), .B2(n6311), .A(n4592), .ZN(U2855) );
  INV_X1 U5654 ( .A(n4593), .ZN(n4594) );
  INV_X1 U5655 ( .A(DATAI_2_), .ZN(n6964) );
  INV_X1 U5656 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6394) );
  OAI222_X1 U5657 ( .A1(n5206), .A2(n6066), .B1(n5398), .B2(n6964), .C1(n5481), 
        .C2(n6394), .ZN(U2889) );
  INV_X1 U5658 ( .A(DATAI_0_), .ZN(n7063) );
  INV_X1 U5659 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6388) );
  OAI222_X1 U5660 ( .A1(n6455), .A2(n6066), .B1(n5398), .B2(n7063), .C1(n5481), 
        .C2(n6388), .ZN(U2891) );
  INV_X1 U5661 ( .A(DATAI_3_), .ZN(n7089) );
  INV_X1 U5662 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6397) );
  OAI222_X1 U5663 ( .A1(n4595), .A2(n6066), .B1(n5398), .B2(n7089), .C1(n5481), 
        .C2(n6397), .ZN(U2888) );
  XNOR2_X1 U5664 ( .A(n4597), .B(n4596), .ZN(n4621) );
  NOR2_X1 U5665 ( .A1(n6446), .A2(n6290), .ZN(n4600) );
  INV_X1 U5666 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6293) );
  INV_X1 U5667 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6673) );
  NOR2_X1 U5668 ( .A1(n6120), .A2(n6673), .ZN(n4618) );
  INV_X1 U5669 ( .A(n4618), .ZN(n4598) );
  OAI21_X1 U5670 ( .B1(n6100), .B2(n6293), .A(n4598), .ZN(n4599) );
  AOI211_X1 U5671 ( .C1(n6304), .C2(n6441), .A(n4600), .B(n4599), .ZN(n4601)
         );
  OAI21_X1 U5672 ( .B1(n4621), .B2(n6161), .A(n4601), .ZN(U2983) );
  INV_X1 U5673 ( .A(n6507), .ZN(n4612) );
  NOR2_X1 U5674 ( .A1(n4573), .A2(n4602), .ZN(n4603) );
  NAND2_X1 U5675 ( .A1(n5034), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5239) );
  AND2_X1 U5676 ( .A1(n5239), .A2(n5112), .ZN(n4964) );
  INV_X1 U5677 ( .A(n5889), .ZN(n4962) );
  NAND2_X1 U5678 ( .A1(n4904), .A2(n4962), .ZN(n4896) );
  AOI21_X1 U5679 ( .B1(n4964), .B2(n4896), .A(n6517), .ZN(n4606) );
  NAND2_X1 U5680 ( .A1(n5917), .A2(n7092), .ZN(n5907) );
  INV_X1 U5681 ( .A(n4530), .ZN(n6301) );
  INV_X1 U5682 ( .A(n4604), .ZN(n5891) );
  OAI22_X1 U5683 ( .A1(n4290), .A2(n5907), .B1(n6301), .B2(n5891), .ZN(n4605)
         );
  OAI21_X1 U5684 ( .B1(n4606), .B2(n4605), .A(n4612), .ZN(n4607) );
  OAI21_X1 U5685 ( .B1(n4612), .B2(n6619), .A(n4607), .ZN(U3462) );
  AND2_X1 U5686 ( .A1(n4609), .A2(n4608), .ZN(n6637) );
  INV_X1 U5687 ( .A(n6609), .ZN(n5277) );
  OAI22_X1 U5688 ( .A1(n5077), .A2(n6517), .B1(n5277), .B2(n5891), .ZN(n4610)
         );
  OAI21_X1 U5689 ( .B1(n6637), .B2(n4610), .A(n4612), .ZN(n4611) );
  OAI21_X1 U5690 ( .B1(n4612), .B2(n6606), .A(n4611), .ZN(U3465) );
  NAND2_X1 U5691 ( .A1(n4614), .A2(n6489), .ZN(n4698) );
  INV_X1 U5692 ( .A(n6482), .ZN(n4701) );
  AOI21_X1 U5693 ( .B1(n5835), .B2(n4698), .A(n4701), .ZN(n5883) );
  INV_X1 U5694 ( .A(n5883), .ZN(n4617) );
  NOR2_X1 U5695 ( .A1(n5835), .A2(n6482), .ZN(n5884) );
  OAI21_X1 U5696 ( .B1(n4615), .B2(n4614), .A(n4613), .ZN(n6488) );
  NOR2_X1 U5697 ( .A1(n5884), .A2(n6488), .ZN(n4616) );
  MUX2_X1 U5698 ( .A(n4617), .B(n4616), .S(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .Z(n4620) );
  AOI21_X1 U5699 ( .B1(n6499), .B2(n6296), .A(n4618), .ZN(n4619) );
  OAI211_X1 U5700 ( .C1(n4621), .C2(n6134), .A(n4620), .B(n4619), .ZN(U3015)
         );
  OAI21_X1 U5701 ( .B1(n4624), .B2(n4623), .A(n4622), .ZN(n6498) );
  AOI22_X1 U5702 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6503), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4627) );
  INV_X1 U5703 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U5704 ( .A1(n6095), .A2(n4625), .ZN(n4626) );
  OAI211_X1 U5705 ( .C1(n5311), .C2(n6454), .A(n4627), .B(n4626), .ZN(n4628)
         );
  INV_X1 U5706 ( .A(n4628), .ZN(n4629) );
  OAI21_X1 U5707 ( .B1(n6161), .B2(n6498), .A(n4629), .ZN(U2985) );
  OR2_X1 U5708 ( .A1(n4587), .A2(n4631), .ZN(n4632) );
  AND2_X1 U5709 ( .A1(n4630), .A2(n4632), .ZN(n6262) );
  INV_X1 U5710 ( .A(n6262), .ZN(n4636) );
  INV_X1 U5711 ( .A(DATAI_5_), .ZN(n6829) );
  INV_X1 U5712 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6403) );
  OAI222_X1 U5713 ( .A1(n4636), .A2(n6066), .B1(n5398), .B2(n6829), .C1(n5481), 
        .C2(n6403), .ZN(U2886) );
  INV_X1 U5714 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4635) );
  OAI21_X1 U5715 ( .B1(n4634), .B2(n4633), .A(n4712), .ZN(n4697) );
  OAI222_X1 U5716 ( .A1(n4636), .A2(n6311), .B1(n4635), .B2(n6322), .C1(n6310), 
        .C2(n4697), .ZN(U2854) );
  XNOR2_X1 U5717 ( .A(n4637), .B(n3160), .ZN(n4706) );
  INV_X1 U5718 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U5719 ( .A1(n6120), .A2(n6676), .ZN(n4700) );
  AOI21_X1 U5720 ( .B1(n6448), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4700), 
        .ZN(n4639) );
  OAI21_X1 U5721 ( .B1(n6269), .B2(n6446), .A(n4639), .ZN(n4640) );
  AOI21_X1 U5722 ( .B1(n6262), .B2(n6441), .A(n4640), .ZN(n4641) );
  OAI21_X1 U5723 ( .B1(n6161), .B2(n4706), .A(n4641), .ZN(U2981) );
  XOR2_X1 U5724 ( .A(n4643), .B(n4642), .Z(n5881) );
  NAND2_X1 U5725 ( .A1(n5881), .A2(n6450), .ZN(n4646) );
  OAI22_X1 U5726 ( .A1(n6100), .A2(n6273), .B1(n6120), .B2(n6674), .ZN(n4644)
         );
  AOI21_X1 U5727 ( .B1(n6095), .B2(n6270), .A(n4644), .ZN(n4645) );
  OAI211_X1 U5728 ( .C1(n6454), .C2(n6275), .A(n4646), .B(n4645), .ZN(U2982)
         );
  INV_X1 U5729 ( .A(n4552), .ZN(n4649) );
  INV_X1 U5730 ( .A(n4648), .ZN(n5897) );
  NOR2_X1 U5731 ( .A1(n4649), .A2(n5897), .ZN(n5236) );
  AND2_X1 U5732 ( .A1(n4573), .A2(n5012), .ZN(n4835) );
  NAND2_X1 U5733 ( .A1(n5122), .A2(n4835), .ZN(n4653) );
  NAND2_X1 U5734 ( .A1(n5034), .A2(n5077), .ZN(n5233) );
  AOI21_X1 U5735 ( .B1(n4653), .B2(n5233), .A(n7092), .ZN(n4650) );
  AOI211_X1 U5736 ( .C1(n5236), .C2(n4897), .A(n6517), .B(n4650), .ZN(n4652)
         );
  NAND2_X1 U5737 ( .A1(n4838), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5237) );
  NOR2_X1 U5738 ( .A1(n6619), .A2(n5237), .ZN(n5241) );
  AND2_X1 U5739 ( .A1(n6606), .A2(n5241), .ZN(n4691) );
  NOR2_X1 U5740 ( .A1(n4656), .A2(n5115), .ZN(n5039) );
  INV_X1 U5741 ( .A(n5039), .ZN(n5915) );
  OR2_X1 U5742 ( .A1(n6510), .A2(n4715), .ZN(n4842) );
  AOI21_X1 U5743 ( .B1(n4842), .B2(STATE2_REG_2__SCAN_IN), .A(n4764), .ZN(
        n4839) );
  OAI211_X1 U5744 ( .C1(n5471), .C2(n4691), .A(n5915), .B(n4839), .ZN(n4651)
         );
  INV_X1 U5745 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U5746 ( .A1(n6441), .A2(DATAI_25_), .ZN(n5932) );
  INV_X1 U5747 ( .A(n5932), .ZN(n6532) );
  NAND2_X1 U5748 ( .A1(n6441), .A2(DATAI_17_), .ZN(n6535) );
  NAND2_X1 U5749 ( .A1(n4654), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6707) );
  INV_X1 U5750 ( .A(n6707), .ZN(n5402) );
  NOR2_X1 U5751 ( .A1(n4689), .A2(n3345), .ZN(n6531) );
  INV_X1 U5752 ( .A(DATAI_1_), .ZN(n4827) );
  NAND2_X1 U5753 ( .A1(n5236), .A2(n5917), .ZN(n4791) );
  AND2_X1 U5754 ( .A1(n4656), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6511) );
  INV_X1 U5755 ( .A(n6511), .ZN(n5045) );
  OAI22_X1 U5756 ( .A1(n4791), .A2(n6301), .B1(n5045), .B2(n4842), .ZN(n4690)
         );
  AOI22_X1 U5757 ( .A1(n6531), .A2(n4691), .B1(n6530), .B2(n4690), .ZN(n4657)
         );
  OAI21_X1 U5758 ( .B1(n6535), .B2(n5233), .A(n4657), .ZN(n4658) );
  AOI21_X1 U5759 ( .B1(n6532), .B2(n6593), .A(n4658), .ZN(n4659) );
  OAI21_X1 U5760 ( .B1(n4696), .B2(n4660), .A(n4659), .ZN(U3117) );
  INV_X1 U5761 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5762 ( .A1(n6441), .A2(DATAI_29_), .ZN(n6602) );
  INV_X1 U5763 ( .A(n6602), .ZN(n6548) );
  NAND2_X1 U5764 ( .A1(n6441), .A2(DATAI_21_), .ZN(n6551) );
  NOR2_X1 U5765 ( .A1(n4689), .A2(n4661), .ZN(n6595) );
  AOI22_X1 U5766 ( .A1(n6595), .A2(n4691), .B1(n6597), .B2(n4690), .ZN(n4662)
         );
  OAI21_X1 U5767 ( .B1(n6551), .B2(n5233), .A(n4662), .ZN(n4663) );
  AOI21_X1 U5768 ( .B1(n6548), .B2(n6593), .A(n4663), .ZN(n4664) );
  OAI21_X1 U5769 ( .B1(n4696), .B2(n4665), .A(n4664), .ZN(U3121) );
  INV_X1 U5770 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4670) );
  NAND2_X1 U5771 ( .A1(n6441), .A2(DATAI_28_), .ZN(n6585) );
  INV_X1 U5772 ( .A(n6585), .ZN(n6544) );
  NAND2_X1 U5773 ( .A1(n6441), .A2(DATAI_20_), .ZN(n6547) );
  NOR2_X1 U5774 ( .A1(n4689), .A2(n4666), .ZN(n6578) );
  INV_X1 U5775 ( .A(DATAI_4_), .ZN(n7090) );
  AOI22_X1 U5776 ( .A1(n6578), .A2(n4691), .B1(n6580), .B2(n4690), .ZN(n4667)
         );
  OAI21_X1 U5777 ( .B1(n6547), .B2(n5233), .A(n4667), .ZN(n4668) );
  AOI21_X1 U5778 ( .B1(n6544), .B2(n6593), .A(n4668), .ZN(n4669) );
  OAI21_X1 U5779 ( .B1(n4696), .B2(n4670), .A(n4669), .ZN(U3120) );
  INV_X1 U5780 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U5781 ( .A1(n6441), .A2(DATAI_26_), .ZN(n6574) );
  INV_X1 U5782 ( .A(n6574), .ZN(n6536) );
  NAND2_X1 U5783 ( .A1(n6441), .A2(DATAI_18_), .ZN(n6539) );
  AOI22_X1 U5784 ( .A1(n6570), .A2(n4691), .B1(n6571), .B2(n4690), .ZN(n4671)
         );
  OAI21_X1 U5785 ( .B1(n6539), .B2(n5233), .A(n4671), .ZN(n4672) );
  AOI21_X1 U5786 ( .B1(n6536), .B2(n6593), .A(n4672), .ZN(n4673) );
  OAI21_X1 U5787 ( .B1(n4696), .B2(n4674), .A(n4673), .ZN(U3118) );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U5789 ( .A1(n6441), .A2(DATAI_31_), .ZN(n5970) );
  INV_X1 U5790 ( .A(n5970), .ZN(n6563) );
  NAND2_X1 U5791 ( .A1(n6441), .A2(DATAI_23_), .ZN(n6567) );
  INV_X1 U5792 ( .A(DATAI_7_), .ZN(n6981) );
  AOI22_X1 U5793 ( .A1(n6561), .A2(n4691), .B1(n6559), .B2(n4690), .ZN(n4675)
         );
  OAI21_X1 U5794 ( .B1(n6567), .B2(n5233), .A(n4675), .ZN(n4676) );
  AOI21_X1 U5795 ( .B1(n6563), .B2(n6593), .A(n4676), .ZN(n4677) );
  OAI21_X1 U5796 ( .B1(n4696), .B2(n4678), .A(n4677), .ZN(U3123) );
  INV_X1 U5797 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5798 ( .A1(n6441), .A2(DATAI_27_), .ZN(n6591) );
  INV_X1 U5799 ( .A(n6591), .ZN(n6540) );
  NAND2_X1 U5800 ( .A1(n6441), .A2(DATAI_19_), .ZN(n6543) );
  NOR2_X1 U5801 ( .A1(n4689), .A2(n4679), .ZN(n6587) );
  AOI22_X1 U5802 ( .A1(n6587), .A2(n4691), .B1(n6588), .B2(n4690), .ZN(n4680)
         );
  OAI21_X1 U5803 ( .B1(n6543), .B2(n5233), .A(n4680), .ZN(n4681) );
  AOI21_X1 U5804 ( .B1(n6540), .B2(n6593), .A(n4681), .ZN(n4682) );
  OAI21_X1 U5805 ( .B1(n4696), .B2(n4683), .A(n4682), .ZN(U3119) );
  INV_X1 U5806 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4687) );
  NAND2_X1 U5807 ( .A1(n6441), .A2(DATAI_30_), .ZN(n5959) );
  INV_X1 U5808 ( .A(n5959), .ZN(n6554) );
  NAND2_X1 U5809 ( .A1(n6441), .A2(DATAI_22_), .ZN(n6557) );
  INV_X1 U5810 ( .A(DATAI_6_), .ZN(n6841) );
  AOI22_X1 U5811 ( .A1(n6553), .A2(n4691), .B1(n6552), .B2(n4690), .ZN(n4684)
         );
  OAI21_X1 U5812 ( .B1(n6557), .B2(n5233), .A(n4684), .ZN(n4685) );
  AOI21_X1 U5813 ( .B1(n6554), .B2(n6593), .A(n4685), .ZN(n4686) );
  OAI21_X1 U5814 ( .B1(n4696), .B2(n4687), .A(n4686), .ZN(U3122) );
  INV_X1 U5815 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5816 ( .A1(n6441), .A2(DATAI_24_), .ZN(n5925) );
  INV_X1 U5817 ( .A(n5925), .ZN(n6526) );
  NAND2_X1 U5818 ( .A1(n6441), .A2(DATAI_16_), .ZN(n6529) );
  NOR2_X1 U5819 ( .A1(n4689), .A2(n4688), .ZN(n6515) );
  AOI22_X1 U5820 ( .A1(n6515), .A2(n4691), .B1(n6514), .B2(n4690), .ZN(n4692)
         );
  OAI21_X1 U5821 ( .B1(n6529), .B2(n5233), .A(n4692), .ZN(n4693) );
  AOI21_X1 U5822 ( .B1(n6526), .B2(n6593), .A(n4693), .ZN(n4694) );
  OAI21_X1 U5823 ( .B1(n4696), .B2(n4695), .A(n4694), .ZN(U3116) );
  INV_X1 U5824 ( .A(n4697), .ZN(n6257) );
  NOR3_X1 U5825 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5882), .A3(n4698), 
        .ZN(n4699) );
  AOI211_X1 U5826 ( .C1(n6499), .C2(n6257), .A(n4700), .B(n4699), .ZN(n4705)
         );
  NOR3_X1 U5827 ( .A1(n4701), .A2(n5882), .A3(n5835), .ZN(n4703) );
  INV_X1 U5828 ( .A(n6488), .ZN(n4702) );
  OAI221_X1 U5829 ( .B1(n5839), .B2(n4883), .C1(n5839), .C2(n6482), .A(n4702), 
        .ZN(n4887) );
  OAI21_X1 U5830 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4703), .A(n4887), 
        .ZN(n4704) );
  OAI211_X1 U5831 ( .C1(n6134), .C2(n4706), .A(n4705), .B(n4704), .ZN(U3013)
         );
  NAND2_X1 U5832 ( .A1(n4630), .A2(n4709), .ZN(n4710) );
  AND2_X1 U5833 ( .A1(n4708), .A2(n4710), .ZN(n6253) );
  INV_X1 U5834 ( .A(n6253), .ZN(n4828) );
  INV_X1 U5835 ( .A(n4893), .ZN(n4711) );
  AOI21_X1 U5836 ( .B1(n4713), .B2(n4712), .A(n4711), .ZN(n6244) );
  AOI22_X1 U5837 ( .A1(n6244), .A2(n6317), .B1(EBX_REG_6__SCAN_IN), .B2(n5613), 
        .ZN(n4714) );
  OAI21_X1 U5838 ( .B1(n4828), .B2(n6311), .A(n4714), .ZN(U2853) );
  NAND3_X1 U5839 ( .A1(n6619), .A2(n5114), .A3(n4838), .ZN(n4939) );
  NOR2_X1 U5840 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4939), .ZN(n4753)
         );
  INV_X1 U5841 ( .A(n4753), .ZN(n4718) );
  INV_X1 U5842 ( .A(n4715), .ZN(n4716) );
  OR2_X1 U5843 ( .A1(n6510), .A2(n4716), .ZN(n4790) );
  INV_X1 U5844 ( .A(n4790), .ZN(n4717) );
  OAI21_X1 U5845 ( .B1(n4717), .B2(n5115), .A(n5038), .ZN(n4783) );
  AOI211_X1 U5846 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4718), .A(n6511), .B(
        n4783), .ZN(n4723) );
  INV_X1 U5847 ( .A(n4573), .ZN(n4785) );
  AND2_X1 U5848 ( .A1(n4290), .A2(n4785), .ZN(n4719) );
  INV_X1 U5849 ( .A(n4571), .ZN(n4963) );
  NOR2_X2 U5850 ( .A1(n4935), .A2(n5012), .ZN(n4958) );
  NAND3_X1 U5851 ( .A1(n4571), .A2(n4720), .A3(n4573), .ZN(n4761) );
  NOR2_X1 U5852 ( .A1(n4761), .A2(n5077), .ZN(n4724) );
  OAI21_X1 U5853 ( .B1(n4958), .B2(n4724), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4721) );
  NOR2_X1 U5854 ( .A1(n4552), .A2(n5897), .ZN(n5005) );
  NAND2_X1 U5855 ( .A1(n6301), .A2(n5005), .ZN(n4933) );
  NAND3_X1 U5856 ( .A1(n4721), .A2(n5917), .A3(n4933), .ZN(n4722) );
  INV_X1 U5857 ( .A(n6535), .ZN(n5929) );
  OAI22_X1 U5858 ( .A1(n4933), .A2(n6517), .B1(n5915), .B2(n4790), .ZN(n4752)
         );
  AOI22_X1 U5859 ( .A1(n6531), .A2(n4753), .B1(n6530), .B2(n4752), .ZN(n4725)
         );
  OAI21_X1 U5860 ( .B1(n5932), .B2(n4931), .A(n4725), .ZN(n4726) );
  AOI21_X1 U5861 ( .B1(n5929), .B2(n4958), .A(n4726), .ZN(n4727) );
  OAI21_X1 U5862 ( .B1(n4758), .B2(n4728), .A(n4727), .ZN(U3021) );
  INV_X1 U5863 ( .A(n6567), .ZN(n5967) );
  AOI22_X1 U5864 ( .A1(n6561), .A2(n4753), .B1(n6559), .B2(n4752), .ZN(n4729)
         );
  OAI21_X1 U5865 ( .B1(n5970), .B2(n4931), .A(n4729), .ZN(n4730) );
  AOI21_X1 U5866 ( .B1(n5967), .B2(n4958), .A(n4730), .ZN(n4731) );
  OAI21_X1 U5867 ( .B1(n4758), .B2(n4732), .A(n4731), .ZN(U3027) );
  INV_X1 U5868 ( .A(n6543), .ZN(n6586) );
  AOI22_X1 U5869 ( .A1(n6587), .A2(n4753), .B1(n6588), .B2(n4752), .ZN(n4733)
         );
  OAI21_X1 U5870 ( .B1(n6591), .B2(n4931), .A(n4733), .ZN(n4734) );
  AOI21_X1 U5871 ( .B1(n6586), .B2(n4958), .A(n4734), .ZN(n4735) );
  OAI21_X1 U5872 ( .B1(n4758), .B2(n3511), .A(n4735), .ZN(U3023) );
  INV_X1 U5873 ( .A(n6529), .ZN(n5922) );
  AOI22_X1 U5874 ( .A1(n6515), .A2(n4753), .B1(n6514), .B2(n4752), .ZN(n4736)
         );
  OAI21_X1 U5875 ( .B1(n5925), .B2(n4931), .A(n4736), .ZN(n4737) );
  AOI21_X1 U5876 ( .B1(n5922), .B2(n4958), .A(n4737), .ZN(n4738) );
  OAI21_X1 U5877 ( .B1(n4758), .B2(n4739), .A(n4738), .ZN(U3020) );
  INV_X1 U5878 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4743) );
  INV_X1 U5879 ( .A(n6557), .ZN(n5956) );
  AOI22_X1 U5880 ( .A1(n6553), .A2(n4753), .B1(n6552), .B2(n4752), .ZN(n4740)
         );
  OAI21_X1 U5881 ( .B1(n5959), .B2(n4931), .A(n4740), .ZN(n4741) );
  AOI21_X1 U5882 ( .B1(n5956), .B2(n4958), .A(n4741), .ZN(n4742) );
  OAI21_X1 U5883 ( .B1(n4758), .B2(n4743), .A(n4742), .ZN(U3026) );
  INV_X1 U5884 ( .A(n6539), .ZN(n6569) );
  AOI22_X1 U5885 ( .A1(n6570), .A2(n4753), .B1(n6571), .B2(n4752), .ZN(n4744)
         );
  OAI21_X1 U5886 ( .B1(n6574), .B2(n4931), .A(n4744), .ZN(n4745) );
  AOI21_X1 U5887 ( .B1(n6569), .B2(n4958), .A(n4745), .ZN(n4746) );
  OAI21_X1 U5888 ( .B1(n4758), .B2(n4747), .A(n4746), .ZN(U3022) );
  INV_X1 U5889 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4751) );
  INV_X1 U5890 ( .A(n6551), .ZN(n6592) );
  AOI22_X1 U5891 ( .A1(n6595), .A2(n4753), .B1(n6597), .B2(n4752), .ZN(n4748)
         );
  OAI21_X1 U5892 ( .B1(n6602), .B2(n4931), .A(n4748), .ZN(n4749) );
  AOI21_X1 U5893 ( .B1(n6592), .B2(n4958), .A(n4749), .ZN(n4750) );
  OAI21_X1 U5894 ( .B1(n4758), .B2(n4751), .A(n4750), .ZN(U3025) );
  INV_X1 U5895 ( .A(n6547), .ZN(n6576) );
  AOI22_X1 U5896 ( .A1(n6578), .A2(n4753), .B1(n6580), .B2(n4752), .ZN(n4754)
         );
  OAI21_X1 U5897 ( .B1(n6585), .B2(n4931), .A(n4754), .ZN(n4755) );
  AOI21_X1 U5898 ( .B1(n6576), .B2(n4958), .A(n4755), .ZN(n4756) );
  OAI21_X1 U5899 ( .B1(n4758), .B2(n4757), .A(n4756), .ZN(U3024) );
  NAND2_X1 U5900 ( .A1(n4573), .A2(n5077), .ZN(n4970) );
  NOR2_X1 U5901 ( .A1(n4970), .A2(n4602), .ZN(n4759) );
  INV_X1 U5902 ( .A(n6587), .ZN(n5939) );
  NAND2_X1 U5903 ( .A1(n4530), .A2(n6609), .ZN(n5004) );
  NAND2_X1 U5904 ( .A1(n4552), .A2(n5897), .ZN(n5044) );
  OAI21_X1 U5905 ( .B1(n5004), .B2(n5044), .A(n4926), .ZN(n4762) );
  AOI22_X1 U5906 ( .A1(n4762), .A2(n5917), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5040), .ZN(n4925) );
  OAI22_X1 U5907 ( .A1(n5939), .A2(n4926), .B1(n4925), .B2(n5938), .ZN(n4760)
         );
  AOI21_X1 U5908 ( .B1(n6540), .B2(n5072), .A(n4760), .ZN(n4767) );
  INV_X1 U5909 ( .A(n5907), .ZN(n6520) );
  AOI21_X1 U5910 ( .B1(n4761), .B2(n6441), .A(n6520), .ZN(n4763) );
  OR2_X1 U5911 ( .A1(n4763), .A2(n4762), .ZN(n4765) );
  OAI211_X1 U5912 ( .C1(n5040), .C2(n5917), .A(n4765), .B(n5244), .ZN(n4928)
         );
  NAND2_X1 U5913 ( .A1(n4928), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4766)
         );
  OAI211_X1 U5914 ( .C1(n4931), .C2(n6543), .A(n4767), .B(n4766), .ZN(U3143)
         );
  OAI22_X1 U5915 ( .A1(n5964), .A2(n4926), .B1(n4925), .B2(n5961), .ZN(n4768)
         );
  AOI21_X1 U5916 ( .B1(n6563), .B2(n5072), .A(n4768), .ZN(n4770) );
  NAND2_X1 U5917 ( .A1(n4928), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4769)
         );
  OAI211_X1 U5918 ( .C1(n4931), .C2(n6567), .A(n4770), .B(n4769), .ZN(U3147)
         );
  OAI22_X1 U5919 ( .A1(n5954), .A2(n4926), .B1(n4925), .B2(n5953), .ZN(n4771)
         );
  AOI21_X1 U5920 ( .B1(n6554), .B2(n5072), .A(n4771), .ZN(n4773) );
  NAND2_X1 U5921 ( .A1(n4928), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4772)
         );
  OAI211_X1 U5922 ( .C1(n4931), .C2(n6557), .A(n4773), .B(n4772), .ZN(U3146)
         );
  INV_X1 U5923 ( .A(n6570), .ZN(n5934) );
  OAI22_X1 U5924 ( .A1(n5934), .A2(n4926), .B1(n4925), .B2(n5933), .ZN(n4774)
         );
  AOI21_X1 U5925 ( .B1(n6536), .B2(n5072), .A(n4774), .ZN(n4776) );
  NAND2_X1 U5926 ( .A1(n4928), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4775)
         );
  OAI211_X1 U5927 ( .C1(n4931), .C2(n6539), .A(n4776), .B(n4775), .ZN(U3142)
         );
  INV_X1 U5928 ( .A(n6515), .ZN(n5920) );
  OAI22_X1 U5929 ( .A1(n5920), .A2(n4926), .B1(n4925), .B2(n5919), .ZN(n4777)
         );
  AOI21_X1 U5930 ( .B1(n6526), .B2(n5072), .A(n4777), .ZN(n4779) );
  NAND2_X1 U5931 ( .A1(n4928), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4778)
         );
  OAI211_X1 U5932 ( .C1(n4931), .C2(n6529), .A(n4779), .B(n4778), .ZN(U3140)
         );
  INV_X1 U5933 ( .A(n6595), .ZN(n5949) );
  OAI22_X1 U5934 ( .A1(n5949), .A2(n4926), .B1(n4925), .B2(n5948), .ZN(n4780)
         );
  AOI21_X1 U5935 ( .B1(n6548), .B2(n5072), .A(n4780), .ZN(n4782) );
  NAND2_X1 U5936 ( .A1(n4928), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4781)
         );
  OAI211_X1 U5937 ( .C1(n4931), .C2(n6551), .A(n4782), .B(n4781), .ZN(U3145)
         );
  OR2_X1 U5938 ( .A1(n5237), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5081)
         );
  NOR2_X1 U5939 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5081), .ZN(n4821)
         );
  INV_X1 U5940 ( .A(n4821), .ZN(n4784) );
  AOI211_X1 U5941 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4784), .A(n5039), .B(
        n4783), .ZN(n4789) );
  NAND3_X1 U5942 ( .A1(n4963), .A2(n4835), .A3(n4290), .ZN(n4997) );
  NAND2_X1 U5943 ( .A1(n4904), .A2(n4785), .ZN(n5078) );
  OR2_X1 U5944 ( .A1(n5078), .A2(n7092), .ZN(n4786) );
  NAND2_X1 U5945 ( .A1(n5236), .A2(n4787), .ZN(n5075) );
  OAI211_X1 U5946 ( .C1(n6520), .C2(n4997), .A(n5080), .B(n5075), .ZN(n4788)
         );
  INV_X1 U5947 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4795) );
  NOR2_X2 U5948 ( .A1(n5078), .A2(n5012), .ZN(n5107) );
  OAI22_X1 U5949 ( .A1(n4791), .A2(n4530), .B1(n4790), .B2(n5045), .ZN(n4820)
         );
  AOI22_X1 U5950 ( .A1(n6531), .A2(n4821), .B1(n6530), .B2(n4820), .ZN(n4792)
         );
  OAI21_X1 U5951 ( .B1(n5932), .B2(n4997), .A(n4792), .ZN(n4793) );
  AOI21_X1 U5952 ( .B1(n5929), .B2(n5107), .A(n4793), .ZN(n4794) );
  OAI21_X1 U5953 ( .B1(n4826), .B2(n4795), .A(n4794), .ZN(U3053) );
  INV_X1 U5954 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5955 ( .A1(n6578), .A2(n4821), .B1(n6580), .B2(n4820), .ZN(n4796)
         );
  OAI21_X1 U5956 ( .B1(n6585), .B2(n4997), .A(n4796), .ZN(n4797) );
  AOI21_X1 U5957 ( .B1(n6576), .B2(n5107), .A(n4797), .ZN(n4798) );
  OAI21_X1 U5958 ( .B1(n4826), .B2(n4799), .A(n4798), .ZN(U3056) );
  INV_X1 U5959 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U5960 ( .A1(n6515), .A2(n4821), .B1(n6514), .B2(n4820), .ZN(n4800)
         );
  OAI21_X1 U5961 ( .B1(n5925), .B2(n4997), .A(n4800), .ZN(n4801) );
  AOI21_X1 U5962 ( .B1(n5922), .B2(n5107), .A(n4801), .ZN(n4802) );
  OAI21_X1 U5963 ( .B1(n4826), .B2(n4803), .A(n4802), .ZN(U3052) );
  INV_X1 U5964 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4807) );
  AOI22_X1 U5965 ( .A1(n6553), .A2(n4821), .B1(n6552), .B2(n4820), .ZN(n4804)
         );
  OAI21_X1 U5966 ( .B1(n5959), .B2(n4997), .A(n4804), .ZN(n4805) );
  AOI21_X1 U5967 ( .B1(n5956), .B2(n5107), .A(n4805), .ZN(n4806) );
  OAI21_X1 U5968 ( .B1(n4826), .B2(n4807), .A(n4806), .ZN(U3058) );
  INV_X1 U5969 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4811) );
  AOI22_X1 U5970 ( .A1(n6595), .A2(n4821), .B1(n6597), .B2(n4820), .ZN(n4808)
         );
  OAI21_X1 U5971 ( .B1(n6602), .B2(n4997), .A(n4808), .ZN(n4809) );
  AOI21_X1 U5972 ( .B1(n6592), .B2(n5107), .A(n4809), .ZN(n4810) );
  OAI21_X1 U5973 ( .B1(n4826), .B2(n4811), .A(n4810), .ZN(U3057) );
  INV_X1 U5974 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U5975 ( .A1(n6561), .A2(n4821), .B1(n6559), .B2(n4820), .ZN(n4812)
         );
  OAI21_X1 U5976 ( .B1(n5970), .B2(n4997), .A(n4812), .ZN(n4813) );
  AOI21_X1 U5977 ( .B1(n5967), .B2(n5107), .A(n4813), .ZN(n4814) );
  OAI21_X1 U5978 ( .B1(n4826), .B2(n4815), .A(n4814), .ZN(U3059) );
  INV_X1 U5979 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U5980 ( .A1(n6587), .A2(n4821), .B1(n6588), .B2(n4820), .ZN(n4816)
         );
  OAI21_X1 U5981 ( .B1(n6591), .B2(n4997), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5982 ( .B1(n6586), .B2(n5107), .A(n4817), .ZN(n4818) );
  OAI21_X1 U5983 ( .B1(n4826), .B2(n4819), .A(n4818), .ZN(U3055) );
  INV_X1 U5984 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5985 ( .A1(n6570), .A2(n4821), .B1(n6571), .B2(n4820), .ZN(n4822)
         );
  OAI21_X1 U5986 ( .B1(n6574), .B2(n4997), .A(n4822), .ZN(n4823) );
  AOI21_X1 U5987 ( .B1(n6569), .B2(n5107), .A(n4823), .ZN(n4824) );
  OAI21_X1 U5988 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(U3054) );
  INV_X1 U5989 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6391) );
  OAI222_X1 U5990 ( .A1(n5311), .A2(n6066), .B1(n5398), .B2(n4827), .C1(n5481), 
        .C2(n6391), .ZN(U2890) );
  INV_X1 U5991 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6406) );
  OAI222_X1 U5992 ( .A1(n4828), .A2(n6066), .B1(n5398), .B2(n6841), .C1(n5481), 
        .C2(n6406), .ZN(U2885) );
  INV_X1 U5993 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6400) );
  OAI222_X1 U5994 ( .A1(n6275), .A2(n6066), .B1(n5398), .B2(n7090), .C1(n5481), 
        .C2(n6400), .ZN(U2887) );
  XNOR2_X1 U5995 ( .A(n4830), .B(n4829), .ZN(n4889) );
  INV_X1 U5996 ( .A(n6251), .ZN(n4832) );
  AOI22_X1 U5997 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6503), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4831) );
  OAI21_X1 U5998 ( .B1(n4832), .B2(n6446), .A(n4831), .ZN(n4833) );
  AOI21_X1 U5999 ( .B1(n6253), .B2(n6441), .A(n4833), .ZN(n4834) );
  OAI21_X1 U6000 ( .B1(n4889), .B2(n6161), .A(n4834), .ZN(U2980) );
  NAND3_X1 U6001 ( .A1(n5033), .A2(n5917), .A3(n6568), .ZN(n4837) );
  NAND2_X1 U6002 ( .A1(n5005), .A2(n4530), .ZN(n4843) );
  INV_X1 U6003 ( .A(n4843), .ZN(n4836) );
  AOI21_X1 U6004 ( .B1(n4837), .B2(n5907), .A(n4836), .ZN(n4841) );
  NAND3_X1 U6005 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5114), .A3(n4838), .ZN(n5009) );
  NOR2_X1 U6006 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5009), .ZN(n4873)
         );
  OAI211_X1 U6007 ( .C1(n5471), .C2(n4873), .A(n5045), .B(n4839), .ZN(n4840)
         );
  INV_X1 U6008 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4847) );
  OAI22_X1 U6009 ( .A1(n4843), .A2(n6517), .B1(n5915), .B2(n4842), .ZN(n4872)
         );
  AOI22_X1 U6010 ( .A1(n6515), .A2(n4873), .B1(n6514), .B2(n4872), .ZN(n4844)
         );
  OAI21_X1 U6011 ( .B1(n5925), .B2(n6568), .A(n4844), .ZN(n4845) );
  AOI21_X1 U6012 ( .B1(n4876), .B2(n5922), .A(n4845), .ZN(n4846) );
  OAI21_X1 U6013 ( .B1(n4879), .B2(n4847), .A(n4846), .ZN(U3084) );
  INV_X1 U6014 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4851) );
  AOI22_X1 U6015 ( .A1(n6561), .A2(n4873), .B1(n6559), .B2(n4872), .ZN(n4848)
         );
  OAI21_X1 U6016 ( .B1(n5970), .B2(n6568), .A(n4848), .ZN(n4849) );
  AOI21_X1 U6017 ( .B1(n4876), .B2(n5967), .A(n4849), .ZN(n4850) );
  OAI21_X1 U6018 ( .B1(n4879), .B2(n4851), .A(n4850), .ZN(U3091) );
  INV_X1 U6019 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4855) );
  AOI22_X1 U6020 ( .A1(n6531), .A2(n4873), .B1(n6530), .B2(n4872), .ZN(n4852)
         );
  OAI21_X1 U6021 ( .B1(n5932), .B2(n6568), .A(n4852), .ZN(n4853) );
  AOI21_X1 U6022 ( .B1(n4876), .B2(n5929), .A(n4853), .ZN(n4854) );
  OAI21_X1 U6023 ( .B1(n4879), .B2(n4855), .A(n4854), .ZN(U3085) );
  INV_X1 U6024 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4859) );
  AOI22_X1 U6025 ( .A1(n6595), .A2(n4873), .B1(n6597), .B2(n4872), .ZN(n4856)
         );
  OAI21_X1 U6026 ( .B1(n6602), .B2(n6568), .A(n4856), .ZN(n4857) );
  AOI21_X1 U6027 ( .B1(n4876), .B2(n6592), .A(n4857), .ZN(n4858) );
  OAI21_X1 U6028 ( .B1(n4879), .B2(n4859), .A(n4858), .ZN(U3089) );
  INV_X1 U6029 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U6030 ( .A1(n6578), .A2(n4873), .B1(n6580), .B2(n4872), .ZN(n4860)
         );
  OAI21_X1 U6031 ( .B1(n6585), .B2(n6568), .A(n4860), .ZN(n4861) );
  AOI21_X1 U6032 ( .B1(n4876), .B2(n6576), .A(n4861), .ZN(n4862) );
  OAI21_X1 U6033 ( .B1(n4879), .B2(n4863), .A(n4862), .ZN(U3088) );
  INV_X1 U6034 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4867) );
  AOI22_X1 U6035 ( .A1(n6553), .A2(n4873), .B1(n6552), .B2(n4872), .ZN(n4864)
         );
  OAI21_X1 U6036 ( .B1(n5959), .B2(n6568), .A(n4864), .ZN(n4865) );
  AOI21_X1 U6037 ( .B1(n4876), .B2(n5956), .A(n4865), .ZN(n4866) );
  OAI21_X1 U6038 ( .B1(n4879), .B2(n4867), .A(n4866), .ZN(U3090) );
  INV_X1 U6039 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U6040 ( .A1(n6570), .A2(n4873), .B1(n6571), .B2(n4872), .ZN(n4868)
         );
  OAI21_X1 U6041 ( .B1(n6574), .B2(n6568), .A(n4868), .ZN(n4869) );
  AOI21_X1 U6042 ( .B1(n4876), .B2(n6569), .A(n4869), .ZN(n4870) );
  OAI21_X1 U6043 ( .B1(n4879), .B2(n4871), .A(n4870), .ZN(U3086) );
  INV_X1 U6044 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4878) );
  AOI22_X1 U6045 ( .A1(n6587), .A2(n4873), .B1(n6588), .B2(n4872), .ZN(n4874)
         );
  OAI21_X1 U6046 ( .B1(n6591), .B2(n6568), .A(n4874), .ZN(n4875) );
  AOI21_X1 U6047 ( .B1(n4876), .B2(n6586), .A(n4875), .ZN(n4877) );
  OAI21_X1 U6048 ( .B1(n4879), .B2(n4878), .A(n4877), .ZN(U3087) );
  INV_X1 U6049 ( .A(n6531), .ZN(n5927) );
  OAI22_X1 U6050 ( .A1(n5927), .A2(n4926), .B1(n4925), .B2(n5926), .ZN(n4880)
         );
  AOI21_X1 U6051 ( .B1(n6532), .B2(n5072), .A(n4880), .ZN(n4882) );
  NAND2_X1 U6052 ( .A1(n4928), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4881)
         );
  OAI211_X1 U6053 ( .C1(n4931), .C2(n6535), .A(n4882), .B(n4881), .ZN(U3141)
         );
  NAND3_X1 U6054 ( .A1(n4883), .A2(n5883), .A3(n4318), .ZN(n4885) );
  NAND2_X1 U6055 ( .A1(n6244), .A2(n6499), .ZN(n4884) );
  OAI211_X1 U6056 ( .C1(n6678), .C2(n6120), .A(n4885), .B(n4884), .ZN(n4886)
         );
  AOI21_X1 U6057 ( .B1(n4887), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4886), 
        .ZN(n4888) );
  OAI21_X1 U6058 ( .B1(n6134), .B2(n4889), .A(n4888), .ZN(U3012) );
  INV_X1 U6059 ( .A(n4708), .ZN(n5142) );
  INV_X1 U6060 ( .A(n4890), .ZN(n4891) );
  OR2_X1 U6061 ( .A1(n4708), .A2(n4890), .ZN(n5151) );
  OAI21_X1 U6062 ( .B1(n5142), .B2(n4891), .A(n5151), .ZN(n6237) );
  CLKBUF_X1 U6063 ( .A(n4892), .Z(n5154) );
  AOI21_X1 U6064 ( .B1(n4894), .B2(n4893), .A(n5154), .ZN(n6474) );
  AOI22_X1 U6065 ( .A1(n6474), .A2(n6317), .B1(EBX_REG_7__SCAN_IN), .B2(n5613), 
        .ZN(n4895) );
  OAI21_X1 U6066 ( .B1(n6237), .B2(n6311), .A(n4895), .ZN(U2852) );
  NAND2_X1 U6067 ( .A1(n4896), .A2(n5917), .ZN(n4900) );
  OR2_X1 U6068 ( .A1(n5044), .A2(n4897), .ZN(n6519) );
  INV_X1 U6069 ( .A(n6519), .ZN(n4898) );
  INV_X1 U6070 ( .A(n4920), .ZN(n6577) );
  AOI21_X1 U6071 ( .B1(n4898), .B2(n6609), .A(n6577), .ZN(n4901) );
  INV_X1 U6072 ( .A(n6508), .ZN(n4899) );
  OAI22_X1 U6073 ( .A1(n4900), .A2(n4901), .B1(n5115), .B2(n4899), .ZN(n6579)
         );
  INV_X1 U6074 ( .A(n4900), .ZN(n4902) );
  NAND2_X1 U6075 ( .A1(n4902), .A2(n4901), .ZN(n4903) );
  OAI211_X1 U6076 ( .C1(n6508), .C2(n5917), .A(n4903), .B(n5244), .ZN(n6581)
         );
  INV_X1 U6077 ( .A(n4970), .ZN(n5121) );
  NOR2_X1 U6078 ( .A1(n6584), .A2(n6591), .ZN(n4906) );
  OAI22_X1 U6079 ( .A1(n5939), .A2(n4920), .B1(n6543), .B2(n6568), .ZN(n4905)
         );
  AOI211_X1 U6080 ( .C1(INSTQUEUE_REG_7__3__SCAN_IN), .C2(n6581), .A(n4906), 
        .B(n4905), .ZN(n4907) );
  OAI21_X1 U6081 ( .B1(n4924), .B2(n5938), .A(n4907), .ZN(U3079) );
  NOR2_X1 U6082 ( .A1(n6584), .A2(n5932), .ZN(n4909) );
  OAI22_X1 U6083 ( .A1(n5927), .A2(n4920), .B1(n6535), .B2(n6568), .ZN(n4908)
         );
  AOI211_X1 U6084 ( .C1(INSTQUEUE_REG_7__1__SCAN_IN), .C2(n6581), .A(n4909), 
        .B(n4908), .ZN(n4910) );
  OAI21_X1 U6085 ( .B1(n4924), .B2(n5926), .A(n4910), .ZN(U3077) );
  NOR2_X1 U6086 ( .A1(n6584), .A2(n6602), .ZN(n4912) );
  OAI22_X1 U6087 ( .A1(n5949), .A2(n4920), .B1(n6551), .B2(n6568), .ZN(n4911)
         );
  AOI211_X1 U6088 ( .C1(INSTQUEUE_REG_7__5__SCAN_IN), .C2(n6581), .A(n4912), 
        .B(n4911), .ZN(n4913) );
  OAI21_X1 U6089 ( .B1(n4924), .B2(n5948), .A(n4913), .ZN(U3081) );
  NOR2_X1 U6090 ( .A1(n6584), .A2(n5970), .ZN(n4915) );
  OAI22_X1 U6091 ( .A1(n5964), .A2(n4920), .B1(n6567), .B2(n6568), .ZN(n4914)
         );
  AOI211_X1 U6092 ( .C1(INSTQUEUE_REG_7__7__SCAN_IN), .C2(n6581), .A(n4915), 
        .B(n4914), .ZN(n4916) );
  OAI21_X1 U6093 ( .B1(n4924), .B2(n5961), .A(n4916), .ZN(U3083) );
  NOR2_X1 U6094 ( .A1(n6584), .A2(n5959), .ZN(n4918) );
  OAI22_X1 U6095 ( .A1(n5954), .A2(n4920), .B1(n6557), .B2(n6568), .ZN(n4917)
         );
  AOI211_X1 U6096 ( .C1(INSTQUEUE_REG_7__6__SCAN_IN), .C2(n6581), .A(n4918), 
        .B(n4917), .ZN(n4919) );
  OAI21_X1 U6097 ( .B1(n4924), .B2(n5953), .A(n4919), .ZN(U3082) );
  NOR2_X1 U6098 ( .A1(n6584), .A2(n5925), .ZN(n4922) );
  OAI22_X1 U6099 ( .A1(n5920), .A2(n4920), .B1(n6529), .B2(n6568), .ZN(n4921)
         );
  AOI211_X1 U6100 ( .C1(INSTQUEUE_REG_7__0__SCAN_IN), .C2(n6581), .A(n4922), 
        .B(n4921), .ZN(n4923) );
  OAI21_X1 U6101 ( .B1(n4924), .B2(n5919), .A(n4923), .ZN(U3076) );
  INV_X1 U6102 ( .A(n6578), .ZN(n5944) );
  OAI22_X1 U6103 ( .A1(n5944), .A2(n4926), .B1(n4925), .B2(n5943), .ZN(n4927)
         );
  AOI21_X1 U6104 ( .B1(n6544), .B2(n5072), .A(n4927), .ZN(n4930) );
  NAND2_X1 U6105 ( .A1(n4928), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4929)
         );
  OAI211_X1 U6106 ( .C1(n4931), .C2(n6547), .A(n4930), .B(n4929), .ZN(U3144)
         );
  INV_X1 U6107 ( .A(n4935), .ZN(n4932) );
  INV_X1 U6108 ( .A(n4933), .ZN(n4934) );
  NOR2_X1 U6109 ( .A1(n6606), .A2(n4939), .ZN(n4959) );
  AOI21_X1 U6110 ( .B1(n4934), .B2(n6609), .A(n4959), .ZN(n4941) );
  OR2_X1 U6111 ( .A1(n4935), .A2(n7092), .ZN(n4936) );
  NAND2_X1 U6112 ( .A1(n4936), .A2(n5917), .ZN(n4940) );
  INV_X1 U6113 ( .A(n4940), .ZN(n4937) );
  AOI22_X1 U6114 ( .A1(n4941), .A2(n4937), .B1(n6517), .B2(n4939), .ZN(n4938)
         );
  NAND2_X1 U6115 ( .A1(n5244), .A2(n4938), .ZN(n4957) );
  OAI22_X1 U6116 ( .A1(n4941), .A2(n4940), .B1(n5115), .B2(n4939), .ZN(n4956)
         );
  AOI22_X1 U6117 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4957), .B1(n6552), 
        .B2(n4956), .ZN(n4943) );
  AOI22_X1 U6118 ( .A1(n6553), .A2(n4959), .B1(n4958), .B2(n6554), .ZN(n4942)
         );
  OAI211_X1 U6119 ( .C1(n6557), .C2(n5971), .A(n4943), .B(n4942), .ZN(U3034)
         );
  AOI22_X1 U6120 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4957), .B1(n6571), 
        .B2(n4956), .ZN(n4945) );
  AOI22_X1 U6121 ( .A1(n6570), .A2(n4959), .B1(n4958), .B2(n6536), .ZN(n4944)
         );
  OAI211_X1 U6122 ( .C1(n6539), .C2(n5971), .A(n4945), .B(n4944), .ZN(U3030)
         );
  AOI22_X1 U6123 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4957), .B1(n6588), 
        .B2(n4956), .ZN(n4947) );
  AOI22_X1 U6124 ( .A1(n6587), .A2(n4959), .B1(n4958), .B2(n6540), .ZN(n4946)
         );
  OAI211_X1 U6125 ( .C1(n6543), .C2(n5971), .A(n4947), .B(n4946), .ZN(U3031)
         );
  AOI22_X1 U6126 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4957), .B1(n6597), 
        .B2(n4956), .ZN(n4949) );
  AOI22_X1 U6127 ( .A1(n6595), .A2(n4959), .B1(n4958), .B2(n6548), .ZN(n4948)
         );
  OAI211_X1 U6128 ( .C1(n6551), .C2(n5971), .A(n4949), .B(n4948), .ZN(U3033)
         );
  AOI22_X1 U6129 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4957), .B1(n6559), 
        .B2(n4956), .ZN(n4951) );
  AOI22_X1 U6130 ( .A1(n6561), .A2(n4959), .B1(n4958), .B2(n6563), .ZN(n4950)
         );
  OAI211_X1 U6131 ( .C1(n6567), .C2(n5971), .A(n4951), .B(n4950), .ZN(U3035)
         );
  AOI22_X1 U6132 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4957), .B1(n6514), 
        .B2(n4956), .ZN(n4953) );
  AOI22_X1 U6133 ( .A1(n6515), .A2(n4959), .B1(n4958), .B2(n6526), .ZN(n4952)
         );
  OAI211_X1 U6134 ( .C1(n6529), .C2(n5971), .A(n4953), .B(n4952), .ZN(U3028)
         );
  AOI22_X1 U6135 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4957), .B1(n6580), 
        .B2(n4956), .ZN(n4955) );
  AOI22_X1 U6136 ( .A1(n6578), .A2(n4959), .B1(n4958), .B2(n6544), .ZN(n4954)
         );
  OAI211_X1 U6137 ( .C1(n6547), .C2(n5971), .A(n4955), .B(n4954), .ZN(U3032)
         );
  AOI22_X1 U6138 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4957), .B1(n6530), 
        .B2(n4956), .ZN(n4961) );
  AOI22_X1 U6139 ( .A1(n6531), .A2(n4959), .B1(n4958), .B2(n6532), .ZN(n4960)
         );
  OAI211_X1 U6140 ( .C1(n6535), .C2(n5971), .A(n4961), .B(n4960), .ZN(U3029)
         );
  NAND3_X1 U6141 ( .A1(n4964), .A2(n4963), .A3(n4962), .ZN(n4965) );
  NAND2_X1 U6142 ( .A1(n4965), .A2(n5917), .ZN(n4976) );
  INV_X1 U6143 ( .A(n4976), .ZN(n4969) );
  NAND2_X1 U6144 ( .A1(n6301), .A2(n3197), .ZN(n5914) );
  OR2_X1 U6145 ( .A1(n5914), .A2(n5277), .ZN(n4967) );
  INV_X1 U6146 ( .A(n5113), .ZN(n4966) );
  NAND2_X1 U6147 ( .A1(n4966), .A2(n6619), .ZN(n4998) );
  NAND2_X1 U6148 ( .A1(n4967), .A2(n4998), .ZN(n4975) );
  NAND3_X1 U6149 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6619), .A3(n5114), .ZN(n5910) );
  INV_X1 U6150 ( .A(n5910), .ZN(n4968) );
  AOI22_X1 U6151 ( .A1(n4969), .A2(n4975), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4968), .ZN(n5003) );
  INV_X1 U6152 ( .A(n4290), .ZN(n4971) );
  NOR3_X1 U6153 ( .A1(n4971), .A2(n4571), .A3(n4970), .ZN(n4972) );
  OAI22_X1 U6154 ( .A1(n5934), .A2(n4998), .B1(n6539), .B2(n4997), .ZN(n4973)
         );
  AOI21_X1 U6155 ( .B1(n6536), .B2(n5966), .A(n4973), .ZN(n4978) );
  INV_X1 U6156 ( .A(n5244), .ZN(n5117) );
  AOI21_X1 U6157 ( .B1(n6517), .B2(n5910), .A(n5117), .ZN(n4974) );
  NAND2_X1 U6158 ( .A1(n5000), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4977) );
  OAI211_X1 U6159 ( .C1(n5003), .C2(n5933), .A(n4978), .B(n4977), .ZN(U3046)
         );
  OAI22_X1 U6160 ( .A1(n5954), .A2(n4998), .B1(n6557), .B2(n4997), .ZN(n4979)
         );
  AOI21_X1 U6161 ( .B1(n6554), .B2(n5966), .A(n4979), .ZN(n4981) );
  NAND2_X1 U6162 ( .A1(n5000), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4980) );
  OAI211_X1 U6163 ( .C1(n5003), .C2(n5953), .A(n4981), .B(n4980), .ZN(U3050)
         );
  OAI22_X1 U6164 ( .A1(n5920), .A2(n4998), .B1(n6529), .B2(n4997), .ZN(n4982)
         );
  AOI21_X1 U6165 ( .B1(n6526), .B2(n5966), .A(n4982), .ZN(n4984) );
  NAND2_X1 U6166 ( .A1(n5000), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4983) );
  OAI211_X1 U6167 ( .C1(n5003), .C2(n5919), .A(n4984), .B(n4983), .ZN(U3044)
         );
  OAI22_X1 U6168 ( .A1(n5964), .A2(n4998), .B1(n6567), .B2(n4997), .ZN(n4985)
         );
  AOI21_X1 U6169 ( .B1(n6563), .B2(n5966), .A(n4985), .ZN(n4987) );
  NAND2_X1 U6170 ( .A1(n5000), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4986) );
  OAI211_X1 U6171 ( .C1(n5003), .C2(n5961), .A(n4987), .B(n4986), .ZN(U3051)
         );
  OAI22_X1 U6172 ( .A1(n5944), .A2(n4998), .B1(n6547), .B2(n4997), .ZN(n4988)
         );
  AOI21_X1 U6173 ( .B1(n6544), .B2(n5966), .A(n4988), .ZN(n4990) );
  NAND2_X1 U6174 ( .A1(n5000), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4989) );
  OAI211_X1 U6175 ( .C1(n5003), .C2(n5943), .A(n4990), .B(n4989), .ZN(U3048)
         );
  OAI22_X1 U6176 ( .A1(n5927), .A2(n4998), .B1(n6535), .B2(n4997), .ZN(n4991)
         );
  AOI21_X1 U6177 ( .B1(n6532), .B2(n5966), .A(n4991), .ZN(n4993) );
  NAND2_X1 U6178 ( .A1(n5000), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4992) );
  OAI211_X1 U6179 ( .C1(n5003), .C2(n5926), .A(n4993), .B(n4992), .ZN(U3045)
         );
  OAI22_X1 U6180 ( .A1(n5949), .A2(n4998), .B1(n6551), .B2(n4997), .ZN(n4994)
         );
  AOI21_X1 U6181 ( .B1(n6548), .B2(n5966), .A(n4994), .ZN(n4996) );
  NAND2_X1 U6182 ( .A1(n5000), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4995) );
  OAI211_X1 U6183 ( .C1(n5003), .C2(n5948), .A(n4996), .B(n4995), .ZN(U3049)
         );
  OAI22_X1 U6184 ( .A1(n5939), .A2(n4998), .B1(n6543), .B2(n4997), .ZN(n4999)
         );
  AOI21_X1 U6185 ( .B1(n6540), .B2(n5966), .A(n4999), .ZN(n5002) );
  NAND2_X1 U6186 ( .A1(n5000), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5001) );
  OAI211_X1 U6187 ( .C1(n5003), .C2(n5938), .A(n5002), .B(n5001), .ZN(U3047)
         );
  INV_X1 U6188 ( .A(n5004), .ZN(n5235) );
  NOR2_X1 U6189 ( .A1(n6606), .A2(n5009), .ZN(n5030) );
  AOI21_X1 U6190 ( .B1(n5235), .B2(n5005), .A(n5030), .ZN(n5011) );
  NOR2_X1 U6191 ( .A1(n4573), .A2(n7092), .ZN(n5006) );
  AOI21_X1 U6192 ( .B1(n5122), .B2(n5006), .A(n6517), .ZN(n5008) );
  AOI22_X1 U6193 ( .A1(n5011), .A2(n5008), .B1(n6517), .B2(n5009), .ZN(n5007)
         );
  NAND2_X1 U6194 ( .A1(n5244), .A2(n5007), .ZN(n5029) );
  INV_X1 U6195 ( .A(n5008), .ZN(n5010) );
  OAI22_X1 U6196 ( .A1(n5011), .A2(n5010), .B1(n5115), .B2(n5009), .ZN(n5028)
         );
  AOI22_X1 U6197 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5029), .B1(n6514), 
        .B2(n5028), .ZN(n5015) );
  AOI22_X1 U6198 ( .A1(n5922), .A2(n5386), .B1(n6515), .B2(n5030), .ZN(n5014)
         );
  OAI211_X1 U6199 ( .C1(n5033), .C2(n5925), .A(n5015), .B(n5014), .ZN(U3092)
         );
  AOI22_X1 U6200 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5029), .B1(n6588), 
        .B2(n5028), .ZN(n5017) );
  AOI22_X1 U6201 ( .A1(n5386), .A2(n6586), .B1(n6587), .B2(n5030), .ZN(n5016)
         );
  OAI211_X1 U6202 ( .C1(n5033), .C2(n6591), .A(n5017), .B(n5016), .ZN(U3095)
         );
  AOI22_X1 U6203 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5029), .B1(n6580), 
        .B2(n5028), .ZN(n5019) );
  AOI22_X1 U6204 ( .A1(n5386), .A2(n6576), .B1(n6578), .B2(n5030), .ZN(n5018)
         );
  OAI211_X1 U6205 ( .C1(n5033), .C2(n6585), .A(n5019), .B(n5018), .ZN(U3096)
         );
  AOI22_X1 U6206 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5029), .B1(n6597), 
        .B2(n5028), .ZN(n5021) );
  AOI22_X1 U6207 ( .A1(n5386), .A2(n6592), .B1(n6595), .B2(n5030), .ZN(n5020)
         );
  OAI211_X1 U6208 ( .C1(n5033), .C2(n6602), .A(n5021), .B(n5020), .ZN(U3097)
         );
  AOI22_X1 U6209 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5029), .B1(n6552), 
        .B2(n5028), .ZN(n5023) );
  AOI22_X1 U6210 ( .A1(n5386), .A2(n5956), .B1(n6553), .B2(n5030), .ZN(n5022)
         );
  OAI211_X1 U6211 ( .C1(n5033), .C2(n5959), .A(n5023), .B(n5022), .ZN(U3098)
         );
  AOI22_X1 U6212 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5029), .B1(n6559), 
        .B2(n5028), .ZN(n5025) );
  AOI22_X1 U6213 ( .A1(n5386), .A2(n5967), .B1(n6561), .B2(n5030), .ZN(n5024)
         );
  OAI211_X1 U6214 ( .C1(n5033), .C2(n5970), .A(n5025), .B(n5024), .ZN(U3099)
         );
  AOI22_X1 U6215 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5029), .B1(n6530), 
        .B2(n5028), .ZN(n5027) );
  AOI22_X1 U6216 ( .A1(n5386), .A2(n5929), .B1(n6531), .B2(n5030), .ZN(n5026)
         );
  OAI211_X1 U6217 ( .C1(n5033), .C2(n5932), .A(n5027), .B(n5026), .ZN(U3093)
         );
  AOI22_X1 U6218 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5029), .B1(n6571), 
        .B2(n5028), .ZN(n5032) );
  AOI22_X1 U6219 ( .A1(n5386), .A2(n6569), .B1(n6570), .B2(n5030), .ZN(n5031)
         );
  OAI211_X1 U6220 ( .C1(n5033), .C2(n6574), .A(n5032), .B(n5031), .ZN(U3094)
         );
  INV_X1 U6221 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6409) );
  OAI222_X1 U6222 ( .A1(n6237), .A2(n6066), .B1(n5398), .B2(n6981), .C1(n5481), 
        .C2(n6409), .ZN(U2884) );
  INV_X1 U6223 ( .A(n5034), .ZN(n5035) );
  NOR2_X1 U6224 ( .A1(n5035), .A2(n5077), .ZN(n5036) );
  NOR3_X1 U6225 ( .A1(n5036), .A2(n5072), .A3(n6517), .ZN(n5037) );
  OAI22_X1 U6226 ( .A1(n5037), .A2(n6520), .B1(n6301), .B2(n5044), .ZN(n5043)
         );
  OAI21_X1 U6227 ( .B1(n6510), .B2(n5115), .A(n5038), .ZN(n5355) );
  NOR2_X1 U6228 ( .A1(n5039), .A2(n5355), .ZN(n6524) );
  INV_X1 U6229 ( .A(n5040), .ZN(n5041) );
  OR2_X1 U6230 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5041), .ZN(n5070)
         );
  NOR2_X1 U6231 ( .A1(n5115), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5357)
         );
  AOI21_X1 U6232 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5070), .A(n5357), .ZN(
        n5042) );
  NAND3_X1 U6233 ( .A1(n5043), .A2(n6524), .A3(n5042), .ZN(n5068) );
  NAND2_X1 U6234 ( .A1(n5068), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5049)
         );
  NOR2_X1 U6235 ( .A1(n5044), .A2(n6517), .ZN(n6509) );
  NOR2_X1 U6236 ( .A1(n5045), .A2(n6619), .ZN(n5046) );
  AOI22_X1 U6237 ( .A1(n6509), .A2(n4530), .B1(n6510), .B2(n5046), .ZN(n5069)
         );
  OAI22_X1 U6238 ( .A1(n5954), .A2(n5070), .B1(n5069), .B2(n5953), .ZN(n5047)
         );
  AOI21_X1 U6239 ( .B1(n5956), .B2(n5072), .A(n5047), .ZN(n5048) );
  OAI211_X1 U6240 ( .C1(n5274), .C2(n5959), .A(n5049), .B(n5048), .ZN(U3138)
         );
  NAND2_X1 U6241 ( .A1(n5068), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5052)
         );
  OAI22_X1 U6242 ( .A1(n5939), .A2(n5070), .B1(n5069), .B2(n5938), .ZN(n5050)
         );
  AOI21_X1 U6243 ( .B1(n6586), .B2(n5072), .A(n5050), .ZN(n5051) );
  OAI211_X1 U6244 ( .C1(n5274), .C2(n6591), .A(n5052), .B(n5051), .ZN(U3135)
         );
  NAND2_X1 U6245 ( .A1(n5068), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5055)
         );
  OAI22_X1 U6246 ( .A1(n5927), .A2(n5070), .B1(n5069), .B2(n5926), .ZN(n5053)
         );
  AOI21_X1 U6247 ( .B1(n5929), .B2(n5072), .A(n5053), .ZN(n5054) );
  OAI211_X1 U6248 ( .C1(n5274), .C2(n5932), .A(n5055), .B(n5054), .ZN(U3133)
         );
  NAND2_X1 U6249 ( .A1(n5068), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5058)
         );
  OAI22_X1 U6250 ( .A1(n5920), .A2(n5070), .B1(n5069), .B2(n5919), .ZN(n5056)
         );
  AOI21_X1 U6251 ( .B1(n5922), .B2(n5072), .A(n5056), .ZN(n5057) );
  OAI211_X1 U6252 ( .C1(n5274), .C2(n5925), .A(n5058), .B(n5057), .ZN(U3132)
         );
  NAND2_X1 U6253 ( .A1(n5068), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5061)
         );
  OAI22_X1 U6254 ( .A1(n5964), .A2(n5070), .B1(n5069), .B2(n5961), .ZN(n5059)
         );
  AOI21_X1 U6255 ( .B1(n5967), .B2(n5072), .A(n5059), .ZN(n5060) );
  OAI211_X1 U6256 ( .C1(n5274), .C2(n5970), .A(n5061), .B(n5060), .ZN(U3139)
         );
  NAND2_X1 U6257 ( .A1(n5068), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5064)
         );
  OAI22_X1 U6258 ( .A1(n5944), .A2(n5070), .B1(n5069), .B2(n5943), .ZN(n5062)
         );
  AOI21_X1 U6259 ( .B1(n6576), .B2(n5072), .A(n5062), .ZN(n5063) );
  OAI211_X1 U6260 ( .C1(n5274), .C2(n6585), .A(n5064), .B(n5063), .ZN(U3136)
         );
  NAND2_X1 U6261 ( .A1(n5068), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5067)
         );
  OAI22_X1 U6262 ( .A1(n5934), .A2(n5070), .B1(n5069), .B2(n5933), .ZN(n5065)
         );
  AOI21_X1 U6263 ( .B1(n6569), .B2(n5072), .A(n5065), .ZN(n5066) );
  OAI211_X1 U6264 ( .C1(n5274), .C2(n6574), .A(n5067), .B(n5066), .ZN(U3134)
         );
  NAND2_X1 U6265 ( .A1(n5068), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5074)
         );
  OAI22_X1 U6266 ( .A1(n5949), .A2(n5070), .B1(n5069), .B2(n5948), .ZN(n5071)
         );
  AOI21_X1 U6267 ( .B1(n6592), .B2(n5072), .A(n5071), .ZN(n5073) );
  OAI211_X1 U6268 ( .C1(n5274), .C2(n6602), .A(n5074), .B(n5073), .ZN(U3137)
         );
  OR2_X1 U6269 ( .A1(n6606), .A2(n5081), .ZN(n5105) );
  OAI21_X1 U6270 ( .B1(n5075), .B2(n5277), .A(n5105), .ZN(n5083) );
  INV_X1 U6271 ( .A(n5081), .ZN(n5076) );
  AOI22_X1 U6272 ( .A1(n5080), .A2(n5083), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5076), .ZN(n5111) );
  OR2_X1 U6273 ( .A1(n5078), .A2(n5077), .ZN(n6516) );
  OAI22_X1 U6274 ( .A1(n5954), .A2(n5105), .B1(n6557), .B2(n6516), .ZN(n5079)
         );
  AOI21_X1 U6275 ( .B1(n6554), .B2(n5107), .A(n5079), .ZN(n5086) );
  INV_X1 U6276 ( .A(n5080), .ZN(n5084) );
  AOI21_X1 U6277 ( .B1(n6517), .B2(n5081), .A(n5117), .ZN(n5082) );
  NAND2_X1 U6278 ( .A1(n5108), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5085) );
  OAI211_X1 U6279 ( .C1(n5111), .C2(n5953), .A(n5086), .B(n5085), .ZN(U3066)
         );
  OAI22_X1 U6280 ( .A1(n5964), .A2(n5105), .B1(n6567), .B2(n6516), .ZN(n5087)
         );
  AOI21_X1 U6281 ( .B1(n6563), .B2(n5107), .A(n5087), .ZN(n5089) );
  NAND2_X1 U6282 ( .A1(n5108), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5088) );
  OAI211_X1 U6283 ( .C1(n5111), .C2(n5961), .A(n5089), .B(n5088), .ZN(U3067)
         );
  OAI22_X1 U6284 ( .A1(n5934), .A2(n5105), .B1(n6539), .B2(n6516), .ZN(n5090)
         );
  AOI21_X1 U6285 ( .B1(n6536), .B2(n5107), .A(n5090), .ZN(n5092) );
  NAND2_X1 U6286 ( .A1(n5108), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5091) );
  OAI211_X1 U6287 ( .C1(n5111), .C2(n5933), .A(n5092), .B(n5091), .ZN(U3062)
         );
  OAI22_X1 U6288 ( .A1(n5939), .A2(n5105), .B1(n6543), .B2(n6516), .ZN(n5093)
         );
  AOI21_X1 U6289 ( .B1(n6540), .B2(n5107), .A(n5093), .ZN(n5095) );
  NAND2_X1 U6290 ( .A1(n5108), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5094) );
  OAI211_X1 U6291 ( .C1(n5111), .C2(n5938), .A(n5095), .B(n5094), .ZN(U3063)
         );
  OAI22_X1 U6292 ( .A1(n5920), .A2(n5105), .B1(n6529), .B2(n6516), .ZN(n5096)
         );
  AOI21_X1 U6293 ( .B1(n6526), .B2(n5107), .A(n5096), .ZN(n5098) );
  NAND2_X1 U6294 ( .A1(n5108), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5097) );
  OAI211_X1 U6295 ( .C1(n5111), .C2(n5919), .A(n5098), .B(n5097), .ZN(U3060)
         );
  OAI22_X1 U6296 ( .A1(n5944), .A2(n5105), .B1(n6547), .B2(n6516), .ZN(n5099)
         );
  AOI21_X1 U6297 ( .B1(n6544), .B2(n5107), .A(n5099), .ZN(n5101) );
  NAND2_X1 U6298 ( .A1(n5108), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5100) );
  OAI211_X1 U6299 ( .C1(n5111), .C2(n5943), .A(n5101), .B(n5100), .ZN(U3064)
         );
  OAI22_X1 U6300 ( .A1(n5927), .A2(n5105), .B1(n6535), .B2(n6516), .ZN(n5102)
         );
  AOI21_X1 U6301 ( .B1(n6532), .B2(n5107), .A(n5102), .ZN(n5104) );
  NAND2_X1 U6302 ( .A1(n5108), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5103) );
  OAI211_X1 U6303 ( .C1(n5111), .C2(n5926), .A(n5104), .B(n5103), .ZN(U3061)
         );
  OAI22_X1 U6304 ( .A1(n5949), .A2(n5105), .B1(n6551), .B2(n6516), .ZN(n5106)
         );
  AOI21_X1 U6305 ( .B1(n6548), .B2(n5107), .A(n5106), .ZN(n5110) );
  NAND2_X1 U6306 ( .A1(n5108), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5109) );
  OAI211_X1 U6307 ( .C1(n5111), .C2(n5948), .A(n5110), .B(n5109), .ZN(U3065)
         );
  OAI21_X1 U6308 ( .B1(n5112), .B2(n5889), .A(n5917), .ZN(n5120) );
  AND2_X1 U6309 ( .A1(n3197), .A2(n4530), .ZN(n5356) );
  NOR2_X1 U6310 ( .A1(n5113), .A2(n6619), .ZN(n6594) );
  AOI21_X1 U6311 ( .B1(n5356), .B2(n6609), .A(n6594), .ZN(n5116) );
  NAND3_X1 U6312 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5114), .ZN(n5354) );
  OAI22_X1 U6313 ( .A1(n5120), .A2(n5116), .B1(n5354), .B2(n5115), .ZN(n6596)
         );
  INV_X1 U6314 ( .A(n5116), .ZN(n5119) );
  AOI21_X1 U6315 ( .B1(n6517), .B2(n5354), .A(n5117), .ZN(n5118) );
  OAI21_X1 U6316 ( .B1(n5120), .B2(n5119), .A(n5118), .ZN(n6598) );
  AOI22_X1 U6317 ( .A1(n6578), .A2(n6594), .B1(n6593), .B2(n6576), .ZN(n5123)
         );
  OAI21_X1 U6318 ( .B1(n6585), .B2(n6601), .A(n5123), .ZN(n5124) );
  AOI21_X1 U6319 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n6598), .A(n5124), 
        .ZN(n5125) );
  OAI21_X1 U6320 ( .B1(n5141), .B2(n5943), .A(n5125), .ZN(U3112) );
  AOI22_X1 U6321 ( .A1(n6531), .A2(n6594), .B1(n6593), .B2(n5929), .ZN(n5126)
         );
  OAI21_X1 U6322 ( .B1(n5932), .B2(n6601), .A(n5126), .ZN(n5127) );
  AOI21_X1 U6323 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(n6598), .A(n5127), 
        .ZN(n5128) );
  OAI21_X1 U6324 ( .B1(n5141), .B2(n5926), .A(n5128), .ZN(U3109) );
  AOI22_X1 U6325 ( .A1(n6570), .A2(n6594), .B1(n6593), .B2(n6569), .ZN(n5129)
         );
  OAI21_X1 U6326 ( .B1(n6574), .B2(n6601), .A(n5129), .ZN(n5130) );
  AOI21_X1 U6327 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(n6598), .A(n5130), 
        .ZN(n5131) );
  OAI21_X1 U6328 ( .B1(n5141), .B2(n5933), .A(n5131), .ZN(U3110) );
  AOI22_X1 U6329 ( .A1(n6553), .A2(n6594), .B1(n6593), .B2(n5956), .ZN(n5132)
         );
  OAI21_X1 U6330 ( .B1(n5959), .B2(n6601), .A(n5132), .ZN(n5133) );
  AOI21_X1 U6331 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n6598), .A(n5133), 
        .ZN(n5134) );
  OAI21_X1 U6332 ( .B1(n5141), .B2(n5953), .A(n5134), .ZN(U3114) );
  AOI22_X1 U6333 ( .A1(n6515), .A2(n6594), .B1(n6593), .B2(n5922), .ZN(n5135)
         );
  OAI21_X1 U6334 ( .B1(n5925), .B2(n6601), .A(n5135), .ZN(n5136) );
  AOI21_X1 U6335 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n6598), .A(n5136), 
        .ZN(n5137) );
  OAI21_X1 U6336 ( .B1(n5141), .B2(n5919), .A(n5137), .ZN(U3108) );
  AOI22_X1 U6337 ( .A1(n6561), .A2(n6594), .B1(n6593), .B2(n5967), .ZN(n5138)
         );
  OAI21_X1 U6338 ( .B1(n5970), .B2(n6601), .A(n5138), .ZN(n5139) );
  AOI21_X1 U6339 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6598), .A(n5139), 
        .ZN(n5140) );
  OAI21_X1 U6340 ( .B1(n5141), .B2(n5961), .A(n5140), .ZN(U3115) );
  NAND2_X1 U6341 ( .A1(n5209), .A2(n5144), .ZN(n5286) );
  INV_X1 U6342 ( .A(n5286), .ZN(n5147) );
  NAND2_X1 U6343 ( .A1(n5209), .A2(n5145), .ZN(n5294) );
  OAI21_X1 U6344 ( .B1(n5147), .B2(n5146), .A(n5294), .ZN(n5766) );
  INV_X1 U6345 ( .A(n5297), .ZN(n5148) );
  AOI21_X1 U6346 ( .B1(n5149), .B2(n5290), .A(n5148), .ZN(n6457) );
  AOI22_X1 U6347 ( .A1(n6457), .A2(n6317), .B1(EBX_REG_11__SCAN_IN), .B2(n5613), .ZN(n5150) );
  OAI21_X1 U6348 ( .B1(n5766), .B2(n6311), .A(n5150), .ZN(U2848) );
  AOI21_X1 U6349 ( .B1(n5152), .B2(n5151), .A(n5209), .ZN(n5224) );
  NOR2_X1 U6350 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  OR2_X1 U6351 ( .A1(n5213), .A2(n5155), .ZN(n5173) );
  OAI22_X1 U6352 ( .A1(n5173), .A2(n6310), .B1(n5174), .B2(n6322), .ZN(n5156)
         );
  AOI21_X1 U6353 ( .B1(n5224), .B2(n6318), .A(n5156), .ZN(n5157) );
  INV_X1 U6354 ( .A(n5157), .ZN(U2851) );
  XNOR2_X1 U6355 ( .A(n5158), .B(n5159), .ZN(n5226) );
  AOI211_X1 U6356 ( .C1(n6497), .C2(n5160), .A(n5884), .B(n6488), .ZN(n6481)
         );
  INV_X1 U6357 ( .A(n6481), .ZN(n5341) );
  OAI22_X1 U6358 ( .A1(n5173), .A2(n5869), .B1(n6681), .B2(n6120), .ZN(n5164)
         );
  INV_X1 U6359 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6360 ( .A1(n5161), .A2(n5883), .ZN(n6476) );
  AOI211_X1 U6361 ( .C1(n6480), .C2(n4337), .A(n5162), .B(n6476), .ZN(n5163)
         );
  AOI211_X1 U6362 ( .C1(n5341), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5164), 
        .B(n5163), .ZN(n5165) );
  OAI21_X1 U6363 ( .B1(n6134), .B2(n5226), .A(n5165), .ZN(U3010) );
  INV_X1 U6364 ( .A(n5224), .ZN(n5227) );
  INV_X1 U6365 ( .A(n5210), .ZN(n5166) );
  NAND2_X1 U6366 ( .A1(n6264), .A2(n5166), .ZN(n5182) );
  NAND2_X1 U6367 ( .A1(n5182), .A2(n6232), .ZN(n6225) );
  INV_X1 U6368 ( .A(n5167), .ZN(n6631) );
  NAND2_X1 U6369 ( .A1(n6354), .A2(n6631), .ZN(n5171) );
  NOR2_X1 U6370 ( .A1(n5168), .A2(EBX_REG_31__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6371 ( .A1(n5497), .A2(n5169), .ZN(n5170) );
  NAND2_X1 U6372 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  AND2_X2 U6373 ( .A1(n6717), .A2(n5172), .ZN(n6295) );
  OAI22_X1 U6374 ( .A1(n5174), .A2(n6246), .B1(n6198), .B2(n5173), .ZN(n5175)
         );
  AOI211_X1 U6375 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5175), 
        .B(n6503), .ZN(n5180) );
  NAND2_X1 U6376 ( .A1(n6250), .A2(n5178), .ZN(n5179) );
  OAI211_X1 U6377 ( .C1(n5182), .C2(n5181), .A(n5180), .B(n5179), .ZN(n5183)
         );
  AOI21_X1 U6378 ( .B1(REIP_REG_8__SCAN_IN), .B2(n6225), .A(n5183), .ZN(n5184)
         );
  OAI21_X1 U6379 ( .B1(n5227), .B2(n6236), .A(n5184), .ZN(U2819) );
  OR2_X1 U6380 ( .A1(n6278), .A2(n5185), .ZN(n5192) );
  NAND2_X1 U6381 ( .A1(n5192), .A2(n6232), .ZN(n6215) );
  NAND2_X1 U6382 ( .A1(n6215), .A2(REIP_REG_11__SCAN_IN), .ZN(n5191) );
  INV_X1 U6383 ( .A(n5762), .ZN(n5189) );
  OAI22_X1 U6384 ( .A1(n5187), .A2(n6246), .B1(n5186), .B2(n6292), .ZN(n5188)
         );
  AOI211_X1 U6385 ( .C1(n6250), .C2(n5189), .A(n5188), .B(n6503), .ZN(n5190)
         );
  OAI211_X1 U6386 ( .C1(n6208), .C2(n5192), .A(n5191), .B(n5190), .ZN(n5193)
         );
  AOI21_X1 U6387 ( .B1(n6457), .B2(n6297), .A(n5193), .ZN(n5194) );
  OAI21_X1 U6388 ( .B1(n5766), .B2(n6236), .A(n5194), .ZN(U2816) );
  NAND2_X1 U6389 ( .A1(n6717), .A2(n5493), .ZN(n5195) );
  NAND2_X1 U6390 ( .A1(n5195), .A2(n6236), .ZN(n6303) );
  INV_X1 U6391 ( .A(n6303), .ZN(n5310) );
  INV_X1 U6392 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6393 ( .A1(n6264), .A2(n5196), .ZN(n5302) );
  NAND2_X1 U6394 ( .A1(n5302), .A2(n6232), .ZN(n6289) );
  AOI22_X1 U6395 ( .A1(n6297), .A2(n6484), .B1(n6295), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5203) );
  INV_X1 U6396 ( .A(n6445), .ZN(n5197) );
  AOI22_X1 U6397 ( .A1(n6245), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6250), 
        .B2(n5197), .ZN(n5202) );
  INV_X1 U6398 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6288) );
  NAND3_X1 U6399 ( .A1(n6264), .A2(REIP_REG_1__SCAN_IN), .A3(n6288), .ZN(n5201) );
  INV_X1 U6400 ( .A(n5198), .ZN(n5199) );
  NAND2_X1 U6401 ( .A1(n6717), .A2(n5199), .ZN(n6300) );
  INV_X1 U6402 ( .A(n6300), .ZN(n5303) );
  NAND2_X1 U6403 ( .A1(n5303), .A2(n4552), .ZN(n5200) );
  NAND4_X1 U6404 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n5204)
         );
  AOI21_X1 U6405 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6289), .A(n5204), .ZN(n5205)
         );
  OAI21_X1 U6406 ( .B1(n5206), .B2(n5310), .A(n5205), .ZN(U2825) );
  AND2_X1 U6407 ( .A1(n5209), .A2(n5208), .ZN(n5284) );
  INV_X1 U6408 ( .A(n5284), .ZN(n5207) );
  OAI21_X1 U6409 ( .B1(n5209), .B2(n5208), .A(n5207), .ZN(n5327) );
  INV_X1 U6410 ( .A(n5323), .ZN(n5219) );
  NAND2_X1 U6411 ( .A1(n6264), .A2(n5210), .ZN(n6222) );
  OR2_X1 U6412 ( .A1(n5213), .A2(n5212), .ZN(n5214) );
  NAND2_X1 U6413 ( .A1(n5288), .A2(n5214), .ZN(n6464) );
  OAI22_X1 U6414 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6222), .B1(n6198), .B2(n6464), .ZN(n5218) );
  AOI22_X1 U6415 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6295), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6225), .ZN(n5215) );
  OAI211_X1 U6416 ( .C1(n6292), .C2(n5216), .A(n5215), .B(n6259), .ZN(n5217)
         );
  AOI211_X1 U6417 ( .C1(n6250), .C2(n5219), .A(n5218), .B(n5217), .ZN(n5220)
         );
  OAI21_X1 U6418 ( .B1(n6236), .B2(n5327), .A(n5220), .ZN(U2818) );
  AOI22_X1 U6419 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6503), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5221) );
  OAI21_X1 U6420 ( .B1(n6446), .B2(n5222), .A(n5221), .ZN(n5223) );
  AOI21_X1 U6421 ( .B1(n5224), .B2(n6441), .A(n5223), .ZN(n5225) );
  OAI21_X1 U6422 ( .B1(n6161), .B2(n5226), .A(n5225), .ZN(U2978) );
  INV_X1 U6423 ( .A(DATAI_8_), .ZN(n7067) );
  INV_X1 U6424 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6412) );
  OAI222_X1 U6425 ( .A1(n5227), .A2(n6066), .B1(n5398), .B2(n7067), .C1(n5481), 
        .C2(n6412), .ZN(U2883) );
  INV_X1 U6426 ( .A(DATAI_11_), .ZN(n6856) );
  INV_X1 U6427 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6421) );
  OAI222_X1 U6428 ( .A1(n5766), .A2(n6066), .B1(n5398), .B2(n6856), .C1(n5481), 
        .C2(n6421), .ZN(U2880) );
  XOR2_X1 U6429 ( .A(n5229), .B(n5228), .Z(n6478) );
  NAND2_X1 U6430 ( .A1(n6478), .A2(n6450), .ZN(n5232) );
  INV_X1 U6431 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6680) );
  NOR2_X1 U6432 ( .A1(n6120), .A2(n6680), .ZN(n6473) );
  NOR2_X1 U6433 ( .A1(n6446), .A2(n6235), .ZN(n5230) );
  AOI211_X1 U6434 ( .C1(n6448), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6473), 
        .B(n5230), .ZN(n5231) );
  OAI211_X1 U6435 ( .C1(n6454), .C2(n6237), .A(n5232), .B(n5231), .ZN(U2979)
         );
  AND2_X1 U6436 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5241), .ZN(n5234)
         );
  INV_X1 U6437 ( .A(n5234), .ZN(n5270) );
  AOI21_X1 U6438 ( .B1(n5236), .B2(n5235), .A(n5234), .ZN(n5240) );
  NAND2_X1 U6439 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5238) );
  OAI22_X1 U6440 ( .A1(n5240), .A2(n6517), .B1(n5238), .B2(n5237), .ZN(n5268)
         );
  NAND2_X1 U6441 ( .A1(n5240), .A2(n5239), .ZN(n5245) );
  INV_X1 U6442 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6443 ( .A1(n6517), .A2(n5242), .ZN(n5243) );
  OAI211_X1 U6444 ( .C1(n6517), .C2(n5245), .A(n5244), .B(n5243), .ZN(n5267)
         );
  AOI22_X1 U6445 ( .A1(n5268), .A2(n6559), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n5267), .ZN(n5246) );
  OAI21_X1 U6446 ( .B1(n5964), .B2(n5270), .A(n5246), .ZN(n5247) );
  AOI21_X1 U6447 ( .B1(n6563), .B2(n5272), .A(n5247), .ZN(n5248) );
  OAI21_X1 U6448 ( .B1(n6567), .B2(n5274), .A(n5248), .ZN(U3131) );
  AOI22_X1 U6449 ( .A1(n5268), .A2(n6588), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n5267), .ZN(n5249) );
  OAI21_X1 U6450 ( .B1(n5939), .B2(n5270), .A(n5249), .ZN(n5250) );
  AOI21_X1 U6451 ( .B1(n6540), .B2(n5272), .A(n5250), .ZN(n5251) );
  OAI21_X1 U6452 ( .B1(n6543), .B2(n5274), .A(n5251), .ZN(U3127) );
  AOI22_X1 U6453 ( .A1(n5268), .A2(n6552), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n5267), .ZN(n5252) );
  OAI21_X1 U6454 ( .B1(n5954), .B2(n5270), .A(n5252), .ZN(n5253) );
  AOI21_X1 U6455 ( .B1(n6554), .B2(n5272), .A(n5253), .ZN(n5254) );
  OAI21_X1 U6456 ( .B1(n6557), .B2(n5274), .A(n5254), .ZN(U3130) );
  AOI22_X1 U6457 ( .A1(n5268), .A2(n6571), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n5267), .ZN(n5255) );
  OAI21_X1 U6458 ( .B1(n5934), .B2(n5270), .A(n5255), .ZN(n5256) );
  AOI21_X1 U6459 ( .B1(n6536), .B2(n5272), .A(n5256), .ZN(n5257) );
  OAI21_X1 U6460 ( .B1(n6539), .B2(n5274), .A(n5257), .ZN(U3126) );
  AOI22_X1 U6461 ( .A1(n5268), .A2(n6514), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n5267), .ZN(n5258) );
  OAI21_X1 U6462 ( .B1(n5920), .B2(n5270), .A(n5258), .ZN(n5259) );
  AOI21_X1 U6463 ( .B1(n6526), .B2(n5272), .A(n5259), .ZN(n5260) );
  OAI21_X1 U6464 ( .B1(n6529), .B2(n5274), .A(n5260), .ZN(U3124) );
  AOI22_X1 U6465 ( .A1(n5268), .A2(n6580), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n5267), .ZN(n5261) );
  OAI21_X1 U6466 ( .B1(n5944), .B2(n5270), .A(n5261), .ZN(n5262) );
  AOI21_X1 U6467 ( .B1(n6544), .B2(n5272), .A(n5262), .ZN(n5263) );
  OAI21_X1 U6468 ( .B1(n6547), .B2(n5274), .A(n5263), .ZN(U3128) );
  AOI22_X1 U6469 ( .A1(n5268), .A2(n6530), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n5267), .ZN(n5264) );
  OAI21_X1 U6470 ( .B1(n5927), .B2(n5270), .A(n5264), .ZN(n5265) );
  AOI21_X1 U6471 ( .B1(n6532), .B2(n5272), .A(n5265), .ZN(n5266) );
  OAI21_X1 U6472 ( .B1(n6535), .B2(n5274), .A(n5266), .ZN(U3125) );
  AOI22_X1 U6473 ( .A1(n5268), .A2(n6597), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n5267), .ZN(n5269) );
  OAI21_X1 U6474 ( .B1(n5949), .B2(n5270), .A(n5269), .ZN(n5271) );
  AOI21_X1 U6475 ( .B1(n6548), .B2(n5272), .A(n5271), .ZN(n5273) );
  OAI21_X1 U6476 ( .B1(n6551), .B2(n5274), .A(n5273), .ZN(U3129) );
  INV_X1 U6477 ( .A(DATAI_9_), .ZN(n5275) );
  INV_X1 U6478 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6415) );
  OAI222_X1 U6479 ( .A1(n5327), .A2(n6066), .B1(n5398), .B2(n5275), .C1(n5481), 
        .C2(n6415), .ZN(U2882) );
  OAI21_X1 U6480 ( .B1(n6245), .B2(n6250), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5276) );
  OAI21_X1 U6481 ( .B1(n6300), .B2(n5277), .A(n5276), .ZN(n5281) );
  OAI22_X1 U6482 ( .A1(n5279), .A2(n6246), .B1(n6198), .B2(n5278), .ZN(n5280)
         );
  AOI211_X1 U6483 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6271), .A(n5281), .B(n5280), 
        .ZN(n5282) );
  OAI21_X1 U6484 ( .B1(n5310), .B2(n6455), .A(n5282), .ZN(U2827) );
  OR2_X1 U6485 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  NAND2_X1 U6486 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  AND2_X1 U6487 ( .A1(n5290), .A2(n5289), .ZN(n6224) );
  AOI22_X1 U6488 ( .A1(n6224), .A2(n6317), .B1(EBX_REG_10__SCAN_IN), .B2(n5613), .ZN(n5291) );
  OAI21_X1 U6489 ( .B1(n5300), .B2(n6311), .A(n5291), .ZN(U2849) );
  INV_X1 U6490 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5292) );
  OAI222_X1 U6491 ( .A1(n6464), .A2(n6310), .B1(n6322), .B2(n5292), .C1(n5327), 
        .C2(n6311), .ZN(U2850) );
  AOI21_X1 U6492 ( .B1(n5295), .B2(n5294), .A(n5293), .ZN(n6217) );
  INV_X1 U6493 ( .A(n6217), .ZN(n5301) );
  AND2_X1 U6494 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  NOR2_X1 U6495 ( .A1(n6138), .A2(n5298), .ZN(n6214) );
  AOI22_X1 U6496 ( .A1(n6214), .A2(n6317), .B1(EBX_REG_12__SCAN_IN), .B2(n5613), .ZN(n5299) );
  OAI21_X1 U6497 ( .B1(n5301), .B2(n6311), .A(n5299), .ZN(U2847) );
  INV_X1 U6498 ( .A(DATAI_10_), .ZN(n6885) );
  INV_X1 U6499 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6418) );
  OAI222_X1 U6500 ( .A1(n5300), .A2(n6066), .B1(n5398), .B2(n6885), .C1(n5481), 
        .C2(n6418), .ZN(U2881) );
  INV_X1 U6501 ( .A(DATAI_12_), .ZN(n7079) );
  INV_X1 U6502 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6425) );
  OAI222_X1 U6503 ( .A1(n5301), .A2(n6066), .B1(n5398), .B2(n7079), .C1(n5481), 
        .C2(n6425), .ZN(U2879) );
  INV_X1 U6504 ( .A(n5302), .ZN(n5307) );
  AOI22_X1 U6505 ( .A1(n5897), .A2(n5303), .B1(n6295), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5305) );
  INV_X1 U6506 ( .A(n6232), .ZN(n6272) );
  AOI22_X1 U6507 ( .A1(n6245), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6272), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5304) );
  OAI211_X1 U6508 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6291), .A(n5305), 
        .B(n5304), .ZN(n5306) );
  AOI211_X1 U6509 ( .C1(n6297), .C2(n5308), .A(n5307), .B(n5306), .ZN(n5309)
         );
  OAI21_X1 U6510 ( .B1(n5311), .B2(n5310), .A(n5309), .ZN(U2826) );
  INV_X1 U6511 ( .A(n5313), .ZN(n5314) );
  XNOR2_X1 U6512 ( .A(n5312), .B(n5314), .ZN(n6319) );
  INV_X1 U6513 ( .A(n6319), .ZN(n5315) );
  INV_X1 U6514 ( .A(DATAI_13_), .ZN(n6804) );
  INV_X1 U6515 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6428) );
  OAI222_X1 U6516 ( .A1(n6066), .A2(n5315), .B1(n5398), .B2(n6804), .C1(n5481), 
        .C2(n6428), .ZN(U2878) );
  OAI21_X1 U6517 ( .B1(n5316), .B2(n5318), .A(n5317), .ZN(n6199) );
  INV_X1 U6518 ( .A(DATAI_14_), .ZN(n5319) );
  INV_X1 U6519 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6431) );
  OAI222_X1 U6520 ( .A1(n6199), .A2(n6066), .B1(n5398), .B2(n5319), .C1(n5481), 
        .C2(n6431), .ZN(U2877) );
  XNOR2_X1 U6521 ( .A(n4260), .B(n6471), .ZN(n5321) );
  XNOR2_X1 U6522 ( .A(n5320), .B(n5321), .ZN(n6468) );
  NAND2_X1 U6523 ( .A1(n6468), .A2(n6450), .ZN(n5326) );
  INV_X1 U6524 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5322) );
  NOR2_X1 U6525 ( .A1(n6120), .A2(n5322), .ZN(n6465) );
  NOR2_X1 U6526 ( .A1(n6446), .A2(n5323), .ZN(n5324) );
  AOI211_X1 U6527 ( .C1(n6448), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6465), 
        .B(n5324), .ZN(n5325) );
  OAI211_X1 U6528 ( .C1(n6454), .C2(n5327), .A(n5326), .B(n5325), .ZN(U2977)
         );
  INV_X1 U6529 ( .A(n5328), .ZN(n5852) );
  NAND2_X1 U6530 ( .A1(n6139), .A2(n5329), .ZN(n5330) );
  NAND2_X1 U6531 ( .A1(n5852), .A2(n5330), .ZN(n6197) );
  INV_X1 U6532 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5331) );
  OAI222_X1 U6533 ( .A1(n6197), .A2(n6310), .B1(n6322), .B2(n5331), .C1(n6199), 
        .C2(n6311), .ZN(U2845) );
  INV_X1 U6534 ( .A(n5333), .ZN(n5335) );
  NAND2_X1 U6535 ( .A1(n5335), .A2(n5334), .ZN(n5336) );
  XNOR2_X1 U6536 ( .A(n5332), .B(n5336), .ZN(n5350) );
  INV_X1 U6537 ( .A(n6226), .ZN(n5338) );
  AOI22_X1 U6538 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6503), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5337) );
  OAI21_X1 U6539 ( .B1(n6446), .B2(n5338), .A(n5337), .ZN(n5339) );
  AOI21_X1 U6540 ( .B1(n6227), .B2(n6441), .A(n5339), .ZN(n5340) );
  OAI21_X1 U6541 ( .B1(n5350), .B2(n6161), .A(n5340), .ZN(U2976) );
  AOI21_X1 U6542 ( .B1(n6497), .B2(n5342), .A(n5341), .ZN(n6472) );
  NOR2_X1 U6543 ( .A1(n5342), .A2(n6476), .ZN(n6467) );
  OAI211_X1 U6544 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6467), .B(n5343), .ZN(n5346) );
  INV_X1 U6545 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U6546 ( .A1(n6120), .A2(n6682), .ZN(n5344) );
  AOI21_X1 U6547 ( .B1(n6224), .B2(n6499), .A(n5344), .ZN(n5345) );
  OAI211_X1 U6548 ( .C1(n6472), .C2(n5347), .A(n5346), .B(n5345), .ZN(n5348)
         );
  INV_X1 U6549 ( .A(n5348), .ZN(n5349) );
  OAI21_X1 U6550 ( .B1(n5350), .B2(n6134), .A(n5349), .ZN(U3008) );
  INV_X1 U6551 ( .A(n6601), .ZN(n5351) );
  OAI21_X1 U6552 ( .B1(n5386), .B2(n5351), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5352) );
  NOR2_X1 U6553 ( .A1(n5915), .A2(n6619), .ZN(n5353) );
  NOR2_X1 U6554 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5354), .ZN(n5383)
         );
  NOR2_X1 U6555 ( .A1(n6511), .A2(n5355), .ZN(n5911) );
  INV_X1 U6556 ( .A(n5356), .ZN(n5358) );
  AOI21_X1 U6557 ( .B1(n5359), .B2(n5358), .A(n5357), .ZN(n5360) );
  OAI211_X1 U6558 ( .C1(n5383), .C2(n5471), .A(n5911), .B(n5360), .ZN(n5382)
         );
  AOI22_X1 U6559 ( .A1(n6587), .A2(n5383), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5382), .ZN(n5361) );
  OAI21_X1 U6560 ( .B1(n6543), .B2(n6601), .A(n5361), .ZN(n5362) );
  AOI21_X1 U6561 ( .B1(n5386), .B2(n6540), .A(n5362), .ZN(n5363) );
  OAI21_X1 U6562 ( .B1(n5388), .B2(n5938), .A(n5363), .ZN(U3103) );
  AOI22_X1 U6563 ( .A1(n6570), .A2(n5383), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5382), .ZN(n5364) );
  OAI21_X1 U6564 ( .B1(n6539), .B2(n6601), .A(n5364), .ZN(n5365) );
  AOI21_X1 U6565 ( .B1(n5386), .B2(n6536), .A(n5365), .ZN(n5366) );
  OAI21_X1 U6566 ( .B1(n5388), .B2(n5933), .A(n5366), .ZN(U3102) );
  AOI22_X1 U6567 ( .A1(n6561), .A2(n5383), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5382), .ZN(n5367) );
  OAI21_X1 U6568 ( .B1(n6567), .B2(n6601), .A(n5367), .ZN(n5368) );
  AOI21_X1 U6569 ( .B1(n5386), .B2(n6563), .A(n5368), .ZN(n5369) );
  OAI21_X1 U6570 ( .B1(n5388), .B2(n5961), .A(n5369), .ZN(U3107) );
  AOI22_X1 U6571 ( .A1(n6553), .A2(n5383), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5382), .ZN(n5370) );
  OAI21_X1 U6572 ( .B1(n6557), .B2(n6601), .A(n5370), .ZN(n5371) );
  AOI21_X1 U6573 ( .B1(n5386), .B2(n6554), .A(n5371), .ZN(n5372) );
  OAI21_X1 U6574 ( .B1(n5388), .B2(n5953), .A(n5372), .ZN(U3106) );
  AOI22_X1 U6575 ( .A1(n6595), .A2(n5383), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5382), .ZN(n5373) );
  OAI21_X1 U6576 ( .B1(n6551), .B2(n6601), .A(n5373), .ZN(n5374) );
  AOI21_X1 U6577 ( .B1(n5386), .B2(n6548), .A(n5374), .ZN(n5375) );
  OAI21_X1 U6578 ( .B1(n5388), .B2(n5948), .A(n5375), .ZN(U3105) );
  AOI22_X1 U6579 ( .A1(n6531), .A2(n5383), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5382), .ZN(n5376) );
  OAI21_X1 U6580 ( .B1(n6535), .B2(n6601), .A(n5376), .ZN(n5377) );
  AOI21_X1 U6581 ( .B1(n5386), .B2(n6532), .A(n5377), .ZN(n5378) );
  OAI21_X1 U6582 ( .B1(n5388), .B2(n5926), .A(n5378), .ZN(U3101) );
  AOI22_X1 U6583 ( .A1(n6515), .A2(n5383), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5382), .ZN(n5379) );
  OAI21_X1 U6584 ( .B1(n6529), .B2(n6601), .A(n5379), .ZN(n5380) );
  AOI21_X1 U6585 ( .B1(n6526), .B2(n5386), .A(n5380), .ZN(n5381) );
  OAI21_X1 U6586 ( .B1(n5388), .B2(n5919), .A(n5381), .ZN(U3100) );
  AOI22_X1 U6587 ( .A1(n6578), .A2(n5383), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5382), .ZN(n5384) );
  OAI21_X1 U6588 ( .B1(n6547), .B2(n6601), .A(n5384), .ZN(n5385) );
  AOI21_X1 U6589 ( .B1(n5386), .B2(n6544), .A(n5385), .ZN(n5387) );
  OAI21_X1 U6590 ( .B1(n5388), .B2(n5943), .A(n5387), .ZN(U3104) );
  OAI21_X1 U6591 ( .B1(n5390), .B2(n5393), .A(n5392), .ZN(n6177) );
  AOI22_X1 U6592 ( .A1(n6323), .A2(DATAI_16_), .B1(n6326), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6593 ( .A1(n6327), .A2(DATAI_0_), .ZN(n5394) );
  OAI211_X1 U6594 ( .C1(n6177), .C2(n6066), .A(n5395), .B(n5394), .ZN(U2875)
         );
  AND2_X1 U6595 ( .A1(n5317), .A2(n5396), .ZN(n5397) );
  OR2_X1 U6596 ( .A1(n5397), .A2(n5390), .ZN(n6312) );
  INV_X1 U6597 ( .A(DATAI_15_), .ZN(n6975) );
  INV_X1 U6598 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6436) );
  OAI222_X1 U6599 ( .A1(n6312), .A2(n6066), .B1(n5398), .B2(n6975), .C1(n5481), 
        .C2(n6436), .ZN(U2876) );
  NOR2_X1 U6600 ( .A1(n5854), .A2(n5399), .ZN(n5400) );
  OR2_X1 U6601 ( .A1(n5549), .A2(n5400), .ZN(n6176) );
  INV_X1 U6602 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5401) );
  OAI222_X1 U6603 ( .A1(n6176), .A2(n6310), .B1(n6322), .B2(n5401), .C1(n6177), 
        .C2(n6311), .ZN(U2843) );
  INV_X1 U6604 ( .A(n4543), .ZN(n5404) );
  OAI22_X1 U6605 ( .A1(n6611), .A2(n6642), .B1(n6706), .B2(n6858), .ZN(n6151)
         );
  AOI21_X1 U6606 ( .B1(n6635), .B2(n5404), .A(n6149), .ZN(n5409) );
  INV_X1 U6607 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5419) );
  AOI22_X1 U6608 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5419), .B2(n4281), .ZN(n5899)
         );
  NAND2_X1 U6609 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5898) );
  INV_X1 U6610 ( .A(n5898), .ZN(n5403) );
  AND2_X1 U6611 ( .A1(n5899), .A2(n5403), .ZN(n5406) );
  NOR3_X1 U6612 ( .A1(n5404), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5902), 
        .ZN(n5405) );
  AOI211_X1 U6613 ( .C1(n5407), .C2(n5474), .A(n5406), .B(n5405), .ZN(n5408)
         );
  OAI22_X1 U6614 ( .A1(n5409), .A2(n3380), .B1(n6149), .B2(n5408), .ZN(U3459)
         );
  INV_X1 U6615 ( .A(n5453), .ZN(n5416) );
  OR2_X1 U6616 ( .A1(n6105), .A2(n6497), .ZN(n5412) );
  INV_X1 U6617 ( .A(n5412), .ZN(n5413) );
  OR2_X1 U6618 ( .A1(n6105), .A2(n5410), .ZN(n5411) );
  NAND2_X1 U6619 ( .A1(n5412), .A2(n5411), .ZN(n5782) );
  OAI21_X1 U6620 ( .B1(n5413), .B2(n5417), .A(n5782), .ZN(n5768) );
  AOI211_X1 U6621 ( .C1(n5772), .C2(n6497), .A(n5457), .B(n5768), .ZN(n5459)
         );
  NOR3_X1 U6622 ( .A1(n5459), .A2(n5413), .A3(n5419), .ZN(n5414) );
  AOI211_X2 U6623 ( .C1(n5416), .C2(n6499), .A(n5415), .B(n5414), .ZN(n5421)
         );
  NAND3_X1 U6624 ( .A1(n6107), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5777) );
  INV_X1 U6625 ( .A(n5417), .ZN(n5418) );
  NOR2_X1 U6626 ( .A1(n5777), .A2(n5418), .ZN(n5773) );
  NAND4_X1 U6627 ( .A1(n5773), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5419), .ZN(n5420) );
  OAI211_X1 U6628 ( .C1(n5422), .C2(n6134), .A(n5421), .B(n5420), .ZN(U2987)
         );
  INV_X1 U6629 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5423) );
  OAI22_X1 U6630 ( .A1(n6100), .A2(n5423), .B1(n6120), .B2(n6698), .ZN(n5429)
         );
  INV_X1 U6631 ( .A(n5425), .ZN(n5427) );
  OAI21_X1 U6632 ( .B1(n5424), .B2(n5427), .A(n5426), .ZN(n5993) );
  NOR2_X1 U6633 ( .A1(n5993), .A2(n6454), .ZN(n5428) );
  AOI211_X1 U6634 ( .C1(n6095), .C2(n5990), .A(n5429), .B(n5428), .ZN(n5430)
         );
  OAI21_X1 U6635 ( .B1(n5431), .B2(n6161), .A(n5430), .ZN(U2960) );
  NAND2_X1 U6636 ( .A1(n5433), .A2(n6106), .ZN(n5434) );
  NOR2_X1 U6637 ( .A1(n5432), .A2(n5434), .ZN(n5650) );
  NOR2_X1 U6638 ( .A1(n5435), .A2(n5650), .ZN(n5436) );
  XOR2_X1 U6639 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(n5436), .Z(n5451) );
  AND2_X1 U6640 ( .A1(n5426), .A2(n5438), .ZN(n5439) );
  NOR2_X1 U6641 ( .A1(n5437), .A2(n5439), .ZN(n5986) );
  NOR2_X1 U6642 ( .A1(n6446), .A2(n5982), .ZN(n5442) );
  INV_X1 U6643 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5440) );
  INV_X1 U6644 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6699) );
  OR2_X1 U6645 ( .A1(n6120), .A2(n6699), .ZN(n5447) );
  OAI21_X1 U6646 ( .B1(n6100), .B2(n5440), .A(n5447), .ZN(n5441) );
  AOI211_X1 U6647 ( .C1(n5986), .C2(n6441), .A(n5442), .B(n5441), .ZN(n5443)
         );
  OAI21_X1 U6648 ( .B1(n5451), .B2(n6161), .A(n5443), .ZN(U2959) );
  AND2_X1 U6649 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  NOR2_X1 U6650 ( .A1(n5563), .A2(n5446), .ZN(n5985) );
  INV_X1 U6651 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5776) );
  NOR2_X1 U6652 ( .A1(n5782), .A2(n5776), .ZN(n5449) );
  INV_X1 U6653 ( .A(n5447), .ZN(n5448) );
  AOI211_X1 U6654 ( .C1(n5985), .C2(n6499), .A(n5449), .B(n5448), .ZN(n5450)
         );
  OR2_X1 U6655 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5781)
         );
  OAI211_X1 U6656 ( .C1(n5451), .C2(n6134), .A(n5450), .B(n5781), .ZN(U2991)
         );
  OAI22_X1 U6657 ( .A1(n5453), .A2(n6310), .B1(n6322), .B2(n5452), .ZN(U2828)
         );
  NAND2_X1 U6658 ( .A1(n5642), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6659 ( .A1(n5649), .A2(n5454), .ZN(n5641) );
  NAND2_X1 U6660 ( .A1(n5641), .A2(n5772), .ZN(n5455) );
  NAND2_X1 U6661 ( .A1(n5456), .A2(n5455), .ZN(n5458) );
  XNOR2_X1 U6662 ( .A(n5458), .B(n5457), .ZN(n5470) );
  INV_X1 U6663 ( .A(n5508), .ZN(n5462) );
  INV_X1 U6664 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6814) );
  NOR2_X1 U6665 ( .A1(n6120), .A2(n6814), .ZN(n5467) );
  AOI21_X1 U6666 ( .B1(n5773), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5460) );
  NOR2_X1 U6667 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  AOI211_X1 U6668 ( .C1(n6499), .C2(n5462), .A(n5467), .B(n5461), .ZN(n5463)
         );
  OAI21_X1 U6669 ( .B1(n5470), .B2(n6134), .A(n5463), .ZN(U2988) );
  NAND2_X1 U6670 ( .A1(n5464), .A2(n6441), .ZN(n5469) );
  NOR2_X1 U6671 ( .A1(n6100), .A2(n5465), .ZN(n5466) );
  AOI211_X1 U6672 ( .C1(n5505), .C2(n6095), .A(n5467), .B(n5466), .ZN(n5468)
         );
  OAI211_X1 U6673 ( .C1(n5470), .C2(n6161), .A(n5469), .B(n5468), .ZN(U2956)
         );
  AOI21_X1 U6674 ( .B1(n6604), .B2(n5474), .A(n6149), .ZN(n5479) );
  INV_X1 U6675 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5471) );
  NAND3_X1 U6676 ( .A1(n6609), .A2(n5471), .A3(n6608), .ZN(n5473) );
  NAND2_X1 U6677 ( .A1(n5473), .A2(n5472), .ZN(n5476) );
  INV_X1 U6678 ( .A(n5474), .ZN(n5904) );
  OAI21_X1 U6679 ( .B1(n6603), .B2(n5904), .A(n5902), .ZN(n5475) );
  AOI22_X1 U6680 ( .A1(n5476), .A2(n5898), .B1(n5478), .B2(n5475), .ZN(n5477)
         );
  OAI22_X1 U6681 ( .A1(n5479), .A2(n5478), .B1(n6149), .B2(n5477), .ZN(U3461)
         );
  AND2_X1 U6682 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U6683 ( .A1(n5483), .A2(n5482), .ZN(n5485) );
  AOI22_X1 U6684 ( .A1(n6323), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6326), .ZN(n5484) );
  NAND2_X1 U6685 ( .A1(n5485), .A2(n5484), .ZN(U2860) );
  NAND2_X1 U6686 ( .A1(n5487), .A2(n5486), .ZN(n5492) );
  NAND3_X1 U6687 ( .A1(n6621), .A2(n5488), .A3(n5499), .ZN(n5490) );
  INV_X1 U6688 ( .A(n5500), .ZN(n5489) );
  AOI22_X1 U6689 ( .A1(n5490), .A2(n5495), .B1(n5489), .B2(n5501), .ZN(n5491)
         );
  AND2_X1 U6690 ( .A1(n5492), .A2(n5491), .ZN(n6622) );
  INV_X1 U6691 ( .A(n6622), .ZN(n5504) );
  INV_X1 U6692 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U6693 ( .A1(n5495), .A2(n5494), .ZN(n5503) );
  NAND2_X1 U6694 ( .A1(n6354), .A2(n6660), .ZN(n5496) );
  OAI211_X1 U6695 ( .C1(n5498), .C2(n5497), .A(n5496), .B(n6828), .ZN(n6721)
         );
  OAI21_X1 U6696 ( .B1(n5501), .B2(n5500), .A(n5499), .ZN(n5502) );
  NAND3_X1 U6697 ( .A1(n5503), .A2(n6721), .A3(n5502), .ZN(n6623) );
  AND2_X1 U6698 ( .A1(n6623), .A2(n6645), .ZN(n6162) );
  MUX2_X1 U6699 ( .A(MORE_REG_SCAN_IN), .B(n5504), .S(n6162), .Z(U3471) );
  INV_X1 U6700 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6702) );
  OAI21_X1 U6701 ( .B1(n5527), .B2(n6702), .A(n6814), .ZN(n5510) );
  AOI22_X1 U6702 ( .A1(n5505), .A2(n6250), .B1(n6245), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6703 ( .A1(n6295), .A2(EBX_REG_30__SCAN_IN), .ZN(n5506) );
  OAI211_X1 U6704 ( .C1(n5508), .C2(n6198), .A(n5507), .B(n5506), .ZN(n5509)
         );
  AOI21_X1 U6705 ( .B1(n5511), .B2(n5510), .A(n5509), .ZN(n5512) );
  OAI21_X1 U6706 ( .B1(n5513), .B2(n6236), .A(n5512), .ZN(U2797) );
  AOI21_X1 U6707 ( .B1(n5516), .B2(n5560), .A(n5515), .ZN(n5647) );
  INV_X1 U6708 ( .A(n5647), .ZN(n5622) );
  NAND2_X1 U6709 ( .A1(n5517), .A2(n4133), .ZN(n5520) );
  INV_X1 U6710 ( .A(n5518), .ZN(n5519) );
  NAND2_X1 U6711 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  NOR2_X1 U6712 ( .A1(n5565), .A2(n5521), .ZN(n5522) );
  NOR2_X1 U6713 ( .A1(n5523), .A2(n5522), .ZN(n5557) );
  INV_X1 U6714 ( .A(n5557), .ZN(n5770) );
  OAI22_X1 U6715 ( .A1(n5524), .A2(n6292), .B1(n6291), .B2(n5645), .ZN(n5525)
         );
  AOI21_X1 U6716 ( .B1(n6295), .B2(EBX_REG_29__SCAN_IN), .A(n5525), .ZN(n5526)
         );
  OAI21_X1 U6717 ( .B1(n5770), .B2(n6198), .A(n5526), .ZN(n5529) );
  NOR2_X1 U6718 ( .A1(n5527), .A2(REIP_REG_29__SCAN_IN), .ZN(n5528) );
  OAI21_X1 U6719 ( .B1(n5622), .B2(n6236), .A(n5530), .ZN(U2798) );
  INV_X1 U6720 ( .A(n5532), .ZN(n5533) );
  AOI21_X1 U6721 ( .B1(n5534), .B2(n5531), .A(n5533), .ZN(n5716) );
  INV_X1 U6722 ( .A(n5716), .ZN(n5640) );
  INV_X1 U6723 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U6724 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6295), .B1(n5715), .B2(n6250), .ZN(n5535) );
  OAI21_X1 U6725 ( .B1(n6055), .B2(n6882), .A(n5535), .ZN(n5543) );
  OAI22_X1 U6726 ( .A1(n5606), .A2(n5537), .B1(EBX_REG_18__SCAN_IN), .B2(n5536), .ZN(n5538) );
  INV_X1 U6727 ( .A(n5538), .ZN(n5540) );
  NOR2_X1 U6728 ( .A1(n5551), .A2(n5540), .ZN(n5612) );
  AOI21_X1 U6729 ( .B1(n5540), .B2(n5551), .A(n5612), .ZN(n6117) );
  INV_X1 U6730 ( .A(n6117), .ZN(n5616) );
  AOI21_X1 U6731 ( .B1(n6245), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6503), 
        .ZN(n5541) );
  OAI21_X1 U6732 ( .B1(n5616), .B2(n6198), .A(n5541), .ZN(n5542) );
  AOI211_X1 U6733 ( .C1(n6054), .C2(n6882), .A(n5543), .B(n5542), .ZN(n5544)
         );
  OAI21_X1 U6734 ( .B1(n5640), .B2(n6236), .A(n5544), .ZN(U2809) );
  NAND2_X1 U6735 ( .A1(n5392), .A2(n5545), .ZN(n5546) );
  AND2_X1 U6736 ( .A1(n5531), .A2(n5546), .ZN(n6325) );
  INV_X1 U6737 ( .A(n6325), .ZN(n5618) );
  AOI21_X1 U6738 ( .B1(n6845), .B2(n5547), .A(n6055), .ZN(n5555) );
  INV_X1 U6739 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6101) );
  OAI22_X1 U6740 ( .A1(n6101), .A2(n6292), .B1(n6094), .B2(n6291), .ZN(n5554)
         );
  OR2_X1 U6741 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U6742 ( .A1(n5551), .A2(n5550), .ZN(n6129) );
  AOI21_X1 U6743 ( .B1(n6295), .B2(EBX_REG_17__SCAN_IN), .A(n6503), .ZN(n5552)
         );
  OAI21_X1 U6744 ( .B1(n6129), .B2(n6198), .A(n5552), .ZN(n5553) );
  NOR3_X1 U6745 ( .A1(n5555), .A2(n5554), .A3(n5553), .ZN(n5556) );
  OAI21_X1 U6746 ( .B1(n5618), .B2(n6236), .A(n5556), .ZN(U2810) );
  AOI22_X1 U6747 ( .A1(n5557), .A2(n6317), .B1(EBX_REG_29__SCAN_IN), .B2(n5613), .ZN(n5558) );
  OAI21_X1 U6748 ( .B1(n5622), .B2(n6311), .A(n5558), .ZN(U2830) );
  OR2_X1 U6749 ( .A1(n5437), .A2(n5559), .ZN(n5561) );
  NOR2_X1 U6750 ( .A1(n5563), .A2(n5562), .ZN(n5564) );
  OR2_X1 U6751 ( .A1(n5565), .A2(n5564), .ZN(n5974) );
  INV_X1 U6752 ( .A(n5974), .ZN(n5780) );
  AOI22_X1 U6753 ( .A1(n5780), .A2(n6317), .B1(EBX_REG_28__SCAN_IN), .B2(n5613), .ZN(n5566) );
  OAI21_X1 U6754 ( .B1(n5625), .B2(n6311), .A(n5566), .ZN(U2831) );
  INV_X1 U6755 ( .A(n5986), .ZN(n5628) );
  AOI22_X1 U6756 ( .A1(n5985), .A2(n6317), .B1(EBX_REG_27__SCAN_IN), .B2(n5613), .ZN(n5567) );
  OAI21_X1 U6757 ( .B1(n5628), .B2(n6311), .A(n5567), .ZN(U2832) );
  AOI22_X1 U6758 ( .A1(n5995), .A2(n6317), .B1(EBX_REG_26__SCAN_IN), .B2(n5613), .ZN(n5568) );
  OAI21_X1 U6759 ( .B1(n5993), .B2(n6311), .A(n5568), .ZN(U2833) );
  AOI21_X1 U6760 ( .B1(n5571), .B2(n5570), .A(n5424), .ZN(n6081) );
  INV_X1 U6761 ( .A(n6081), .ZN(n5633) );
  NAND2_X1 U6762 ( .A1(n5582), .A2(n5573), .ZN(n5574) );
  AND2_X1 U6763 ( .A1(n5575), .A2(n5574), .ZN(n6102) );
  AOI22_X1 U6764 ( .A1(n6102), .A2(n6317), .B1(EBX_REG_25__SCAN_IN), .B2(n5613), .ZN(n5576) );
  OAI21_X1 U6765 ( .B1(n5633), .B2(n6311), .A(n5576), .ZN(U2834) );
  OAI21_X1 U6766 ( .B1(n5577), .B2(n5578), .A(n5570), .ZN(n5671) );
  INV_X1 U6767 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5583) );
  OR2_X1 U6768 ( .A1(n5798), .A2(n5580), .ZN(n5581) );
  NAND2_X1 U6769 ( .A1(n5582), .A2(n5581), .ZN(n6017) );
  OAI222_X1 U6770 ( .A1(n6311), .A2(n5671), .B1(n6322), .B2(n5583), .C1(n6017), 
        .C2(n6310), .ZN(U2835) );
  NAND2_X1 U6771 ( .A1(n5584), .A2(n5585), .ZN(n5586) );
  NAND2_X1 U6772 ( .A1(n5796), .A2(n5586), .ZN(n6035) );
  INV_X1 U6773 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5591) );
  AOI21_X1 U6774 ( .B1(n5590), .B2(n5587), .A(n5589), .ZN(n5693) );
  INV_X1 U6775 ( .A(n5693), .ZN(n6032) );
  OAI222_X1 U6776 ( .A1(n6035), .A2(n6310), .B1(n6322), .B2(n5591), .C1(n6032), 
        .C2(n6311), .ZN(U2837) );
  INV_X1 U6777 ( .A(n5587), .ZN(n5594) );
  AOI21_X1 U6778 ( .B1(n5595), .B2(n5593), .A(n5594), .ZN(n6070) );
  INV_X1 U6779 ( .A(n6070), .ZN(n5600) );
  INV_X1 U6780 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5599) );
  OR2_X1 U6781 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  NAND2_X1 U6782 ( .A1(n5584), .A2(n5598), .ZN(n6038) );
  OAI222_X1 U6783 ( .A1(n5600), .A2(n6311), .B1(n5599), .B2(n6322), .C1(n6310), 
        .C2(n6038), .ZN(U2838) );
  OR2_X1 U6784 ( .A1(n5602), .A2(n5603), .ZN(n5604) );
  NAND2_X1 U6785 ( .A1(n5593), .A2(n5604), .ZN(n6073) );
  MUX2_X1 U6786 ( .A(n5606), .B(n4133), .S(n5605), .Z(n5608) );
  XNOR2_X1 U6787 ( .A(n5608), .B(n5607), .ZN(n6050) );
  AOI22_X1 U6788 ( .A1(n6050), .A2(n6317), .B1(EBX_REG_20__SCAN_IN), .B2(n5613), .ZN(n5609) );
  OAI21_X1 U6789 ( .B1(n6073), .B2(n6311), .A(n5609), .ZN(U2839) );
  AOI21_X1 U6790 ( .B1(n5610), .B2(n5532), .A(n5602), .ZN(n6087) );
  INV_X1 U6791 ( .A(n6087), .ZN(n5615) );
  XNOR2_X1 U6792 ( .A(n5612), .B(n5611), .ZN(n6111) );
  AOI22_X1 U6793 ( .A1(n6111), .A2(n6317), .B1(EBX_REG_19__SCAN_IN), .B2(n5613), .ZN(n5614) );
  OAI21_X1 U6794 ( .B1(n5615), .B2(n6311), .A(n5614), .ZN(U2840) );
  OAI222_X1 U6795 ( .A1(n5640), .A2(n6311), .B1(n5617), .B2(n6322), .C1(n6310), 
        .C2(n5616), .ZN(U2841) );
  OAI222_X1 U6796 ( .A1(n6129), .A2(n6310), .B1(n5619), .B2(n6322), .C1(n5618), 
        .C2(n6311), .ZN(U2842) );
  AOI22_X1 U6797 ( .A1(n6323), .A2(DATAI_29_), .B1(n6326), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U6798 ( .A1(n6327), .A2(DATAI_13_), .ZN(n5620) );
  OAI211_X1 U6799 ( .C1(n5622), .C2(n6066), .A(n5621), .B(n5620), .ZN(U2862)
         );
  AOI22_X1 U6800 ( .A1(n6327), .A2(DATAI_12_), .B1(n6326), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U6801 ( .A1(n6323), .A2(DATAI_28_), .ZN(n5623) );
  OAI211_X1 U6802 ( .C1(n5625), .C2(n6066), .A(n5624), .B(n5623), .ZN(U2863)
         );
  AOI22_X1 U6803 ( .A1(n6327), .A2(DATAI_11_), .B1(n6326), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6804 ( .A1(n6323), .A2(DATAI_27_), .ZN(n5626) );
  OAI211_X1 U6805 ( .C1(n5628), .C2(n6066), .A(n5627), .B(n5626), .ZN(U2864)
         );
  AOI22_X1 U6806 ( .A1(n6327), .A2(DATAI_10_), .B1(n6326), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U6807 ( .A1(n6323), .A2(DATAI_26_), .ZN(n5629) );
  OAI211_X1 U6808 ( .C1(n5993), .C2(n6066), .A(n5630), .B(n5629), .ZN(U2865)
         );
  AOI22_X1 U6809 ( .A1(n6327), .A2(DATAI_9_), .B1(n6326), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U6810 ( .A1(n6323), .A2(DATAI_25_), .ZN(n5631) );
  OAI211_X1 U6811 ( .C1(n5633), .C2(n6066), .A(n5632), .B(n5631), .ZN(U2866)
         );
  AOI22_X1 U6812 ( .A1(n6327), .A2(DATAI_8_), .B1(n6326), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6813 ( .A1(n6323), .A2(DATAI_24_), .ZN(n5634) );
  OAI211_X1 U6814 ( .C1(n5671), .C2(n6066), .A(n5635), .B(n5634), .ZN(U2867)
         );
  AOI22_X1 U6815 ( .A1(n6327), .A2(DATAI_6_), .B1(n6326), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U6816 ( .A1(n6323), .A2(DATAI_22_), .ZN(n5636) );
  OAI211_X1 U6817 ( .C1(n6032), .C2(n6066), .A(n5637), .B(n5636), .ZN(U2869)
         );
  AOI22_X1 U6818 ( .A1(n6323), .A2(DATAI_18_), .B1(n6326), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6819 ( .A1(n6327), .A2(DATAI_2_), .ZN(n5638) );
  OAI211_X1 U6820 ( .C1(n5640), .C2(n6066), .A(n5639), .B(n5638), .ZN(U2873)
         );
  NAND2_X1 U6821 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  XNOR2_X1 U6822 ( .A(n5643), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5775)
         );
  NOR2_X1 U6823 ( .A1(n6120), .A2(n6702), .ZN(n5767) );
  AOI21_X1 U6824 ( .B1(n6448), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5767), 
        .ZN(n5644) );
  OAI21_X1 U6825 ( .B1(n5645), .B2(n6446), .A(n5644), .ZN(n5646) );
  AOI21_X1 U6826 ( .B1(n5647), .B2(n6441), .A(n5646), .ZN(n5648) );
  OAI21_X1 U6827 ( .B1(n5775), .B2(n6161), .A(n5648), .ZN(U2957) );
  NOR3_X1 U6828 ( .A1(n5649), .A2(n5719), .A3(n5776), .ZN(n5651) );
  OAI22_X1 U6829 ( .A1(n5651), .A2(n5650), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5776), .ZN(n5653) );
  XNOR2_X1 U6830 ( .A(n5653), .B(n5652), .ZN(n5787) );
  NAND2_X1 U6831 ( .A1(n5976), .A2(n6441), .ZN(n5657) );
  INV_X1 U6832 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6960) );
  NOR2_X1 U6833 ( .A1(n6120), .A2(n6960), .ZN(n5779) );
  NOR2_X1 U6834 ( .A1(n6100), .A2(n5654), .ZN(n5655) );
  AOI211_X1 U6835 ( .C1(n6095), .C2(n5973), .A(n5779), .B(n5655), .ZN(n5656)
         );
  OAI211_X1 U6836 ( .C1(n5787), .C2(n6161), .A(n5657), .B(n5656), .ZN(U2958)
         );
  INV_X1 U6837 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U6838 ( .A1(n4260), .A2(n6085), .ZN(n5659) );
  NAND2_X1 U6839 ( .A1(n5658), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U6840 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6841 ( .A1(n5661), .A2(n5660), .ZN(n5702) );
  XNOR2_X1 U6842 ( .A(n4260), .B(n5662), .ZN(n5703) );
  NAND2_X1 U6843 ( .A1(n4260), .A2(n5662), .ZN(n5663) );
  XNOR2_X1 U6844 ( .A(n4260), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5697)
         );
  INV_X1 U6845 ( .A(n5695), .ZN(n5664) );
  NOR2_X1 U6846 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5687)
         );
  INV_X1 U6847 ( .A(n5681), .ZN(n5666) );
  INV_X1 U6848 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6849 ( .A1(n5666), .A2(n5665), .ZN(n5669) );
  INV_X1 U6850 ( .A(n5689), .ZN(n5667) );
  NAND2_X1 U6851 ( .A1(n5667), .A2(n3199), .ZN(n5668) );
  NAND2_X1 U6852 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U6853 ( .A(n5670), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5793)
         );
  INV_X1 U6854 ( .A(n5671), .ZN(n6012) );
  NAND2_X1 U6855 ( .A1(n6503), .A2(REIP_REG_24__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6856 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5672)
         );
  OAI211_X1 U6857 ( .C1(n6446), .C2(n6007), .A(n5789), .B(n5672), .ZN(n5673)
         );
  AOI21_X1 U6858 ( .B1(n6012), .B2(n6441), .A(n5673), .ZN(n5674) );
  OAI21_X1 U6859 ( .B1(n5793), .B2(n6161), .A(n5674), .ZN(U2962) );
  NOR2_X1 U6860 ( .A1(n5589), .A2(n5675), .ZN(n5676) );
  OR2_X1 U6861 ( .A1(n5577), .A2(n5676), .ZN(n6021) );
  NOR3_X1 U6862 ( .A1(n5677), .A2(n5719), .A3(n5711), .ZN(n5710) );
  INV_X1 U6863 ( .A(n5678), .ZN(n5679) );
  NAND3_X1 U6864 ( .A1(n5710), .A2(n5808), .A3(n5679), .ZN(n5680) );
  NAND2_X1 U6865 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  NAND2_X1 U6866 ( .A1(n5794), .A2(n6450), .ZN(n5686) );
  INV_X1 U6867 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5683) );
  NOR2_X1 U6868 ( .A1(n6120), .A2(n5683), .ZN(n5801) );
  NOR2_X1 U6869 ( .A1(n6446), .A2(n6018), .ZN(n5684) );
  AOI211_X1 U6870 ( .C1(n6448), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5801), 
        .B(n5684), .ZN(n5685) );
  OAI211_X1 U6871 ( .C1(n6454), .C2(n6021), .A(n5686), .B(n5685), .ZN(U2963)
         );
  AOI21_X1 U6872 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4260), .A(n5687), 
        .ZN(n5688) );
  XNOR2_X1 U6873 ( .A(n5689), .B(n5688), .ZN(n5812) );
  NAND2_X1 U6874 ( .A1(n6095), .A2(n6027), .ZN(n5690) );
  NAND2_X1 U6875 ( .A1(n6503), .A2(REIP_REG_22__SCAN_IN), .ZN(n5805) );
  OAI211_X1 U6876 ( .C1(n6100), .C2(n5691), .A(n5690), .B(n5805), .ZN(n5692)
         );
  AOI21_X1 U6877 ( .B1(n5693), .B2(n6441), .A(n5692), .ZN(n5694) );
  OAI21_X1 U6878 ( .B1(n5812), .B2(n6161), .A(n5694), .ZN(U2964) );
  OAI21_X1 U6879 ( .B1(n5697), .B2(n5696), .A(n5695), .ZN(n5813) );
  INV_X1 U6880 ( .A(n5813), .ZN(n5701) );
  NAND2_X1 U6881 ( .A1(n6503), .A2(REIP_REG_21__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U6882 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5698)
         );
  OAI211_X1 U6883 ( .C1(n6446), .C2(n6036), .A(n5814), .B(n5698), .ZN(n5699)
         );
  AOI21_X1 U6884 ( .B1(n6070), .B2(n6441), .A(n5699), .ZN(n5700) );
  OAI21_X1 U6885 ( .B1(n5701), .B2(n6161), .A(n5700), .ZN(U2965) );
  XOR2_X1 U6886 ( .A(n5703), .B(n5702), .Z(n5832) );
  INV_X1 U6887 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U6888 ( .A1(n6503), .A2(REIP_REG_20__SCAN_IN), .ZN(n5820) );
  OAI21_X1 U6889 ( .B1(n6100), .B2(n6053), .A(n5820), .ZN(n5705) );
  NOR2_X1 U6890 ( .A1(n6073), .A2(n6454), .ZN(n5704) );
  AOI211_X1 U6891 ( .C1(n6095), .C2(n6045), .A(n5705), .B(n5704), .ZN(n5706)
         );
  OAI21_X1 U6892 ( .B1(n5832), .B2(n6161), .A(n5706), .ZN(U2966) );
  NAND2_X1 U6893 ( .A1(n5719), .A2(n5708), .ZN(n5709) );
  NOR2_X1 U6894 ( .A1(n3161), .A2(n5709), .ZN(n6092) );
  AOI21_X1 U6895 ( .B1(n6092), .B2(n5711), .A(n5710), .ZN(n5712) );
  XNOR2_X1 U6896 ( .A(n5712), .B(n6123), .ZN(n6116) );
  OAI22_X1 U6897 ( .A1(n6100), .A2(n5713), .B1(n6120), .B2(n6882), .ZN(n5714)
         );
  AOI21_X1 U6898 ( .B1(n6095), .B2(n5715), .A(n5714), .ZN(n5718) );
  NAND2_X1 U6899 ( .A1(n5716), .A2(n6441), .ZN(n5717) );
  OAI211_X1 U6900 ( .C1(n6116), .C2(n6161), .A(n5718), .B(n5717), .ZN(U2968)
         );
  NOR2_X1 U6901 ( .A1(n5719), .A2(n5708), .ZN(n5721) );
  MUX2_X1 U6902 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n5708), .S(n4260), 
        .Z(n5720) );
  MUX2_X1 U6903 ( .A(n5721), .B(n5720), .S(n3161), .Z(n5722) );
  NOR2_X1 U6904 ( .A1(n5722), .A2(n6092), .ZN(n5846) );
  NAND2_X1 U6905 ( .A1(n6503), .A2(REIP_REG_16__SCAN_IN), .ZN(n5840) );
  OAI21_X1 U6906 ( .B1(n6100), .B2(n5723), .A(n5840), .ZN(n5725) );
  NOR2_X1 U6907 ( .A1(n6177), .A2(n6454), .ZN(n5724) );
  AOI211_X1 U6908 ( .C1(n6095), .C2(n6179), .A(n5725), .B(n5724), .ZN(n5726)
         );
  OAI21_X1 U6909 ( .B1(n5846), .B2(n6161), .A(n5726), .ZN(U2970) );
  INV_X1 U6910 ( .A(n5728), .ZN(n5730) );
  NAND2_X1 U6911 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  XNOR2_X1 U6912 ( .A(n5727), .B(n5731), .ZN(n5859) );
  NAND2_X1 U6913 ( .A1(n6503), .A2(REIP_REG_15__SCAN_IN), .ZN(n5855) );
  OAI21_X1 U6914 ( .B1(n6100), .B2(n6186), .A(n5855), .ZN(n5733) );
  NOR2_X1 U6915 ( .A1(n6312), .A2(n6454), .ZN(n5732) );
  AOI211_X1 U6916 ( .C1(n6095), .C2(n5734), .A(n5733), .B(n5732), .ZN(n5735)
         );
  OAI21_X1 U6917 ( .B1(n6161), .B2(n5859), .A(n5735), .ZN(U2971) );
  XNOR2_X1 U6918 ( .A(n4260), .B(n5866), .ZN(n5737) );
  XNOR2_X1 U6919 ( .A(n5736), .B(n5737), .ZN(n5874) );
  NAND2_X1 U6920 ( .A1(n6503), .A2(REIP_REG_14__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U6921 ( .B1(n6100), .B2(n5738), .A(n5868), .ZN(n5740) );
  NOR2_X1 U6922 ( .A1(n6199), .A2(n6454), .ZN(n5739) );
  AOI211_X1 U6923 ( .C1(n6095), .C2(n6201), .A(n5740), .B(n5739), .ZN(n5741)
         );
  OAI21_X1 U6924 ( .B1(n6161), .B2(n5874), .A(n5741), .ZN(U2972) );
  OAI21_X1 U6925 ( .B1(n5742), .B2(n5744), .A(n5743), .ZN(n6145) );
  INV_X1 U6926 ( .A(n6145), .ZN(n5748) );
  AOI22_X1 U6927 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6503), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5745) );
  OAI21_X1 U6928 ( .B1(n6206), .B2(n6446), .A(n5745), .ZN(n5746) );
  AOI21_X1 U6929 ( .B1(n6319), .B2(n6441), .A(n5746), .ZN(n5747) );
  OAI21_X1 U6930 ( .B1(n5748), .B2(n6161), .A(n5747), .ZN(U2973) );
  INV_X1 U6931 ( .A(n5750), .ZN(n5751) );
  NOR2_X1 U6932 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  XNOR2_X1 U6933 ( .A(n5749), .B(n5753), .ZN(n5875) );
  INV_X1 U6934 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5754) );
  NOR2_X1 U6935 ( .A1(n6120), .A2(n5754), .ZN(n5876) );
  AND2_X1 U6936 ( .A1(n6448), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5755)
         );
  AOI211_X1 U6937 ( .C1(n6095), .C2(n6216), .A(n5876), .B(n5755), .ZN(n5757)
         );
  NAND2_X1 U6938 ( .A1(n6217), .A2(n6441), .ZN(n5756) );
  OAI211_X1 U6939 ( .C1(n5875), .C2(n6161), .A(n5757), .B(n5756), .ZN(U2974)
         );
  NAND2_X1 U6940 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  XNOR2_X1 U6941 ( .A(n5758), .B(n5761), .ZN(n6459) );
  NAND2_X1 U6942 ( .A1(n6459), .A2(n6450), .ZN(n5765) );
  NOR2_X1 U6943 ( .A1(n6120), .A2(n6684), .ZN(n6456) );
  NOR2_X1 U6944 ( .A1(n6446), .A2(n5762), .ZN(n5763) );
  AOI211_X1 U6945 ( .C1(n6448), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6456), 
        .B(n5763), .ZN(n5764) );
  OAI211_X1 U6946 ( .C1(n6454), .C2(n5766), .A(n5765), .B(n5764), .ZN(U2975)
         );
  AOI21_X1 U6947 ( .B1(n5768), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5767), 
        .ZN(n5769) );
  OAI21_X1 U6948 ( .B1(n5770), .B2(n5869), .A(n5769), .ZN(n5771) );
  AOI21_X1 U6949 ( .B1(n5773), .B2(n5772), .A(n5771), .ZN(n5774) );
  OAI21_X1 U6950 ( .B1(n5775), .B2(n6134), .A(n5774), .ZN(U2989) );
  NOR3_X1 U6951 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5776), 
        .ZN(n5778) );
  AOI211_X1 U6952 ( .C1(n6499), .C2(n5780), .A(n5779), .B(n5778), .ZN(n5786)
         );
  INV_X1 U6953 ( .A(n5781), .ZN(n5784) );
  INV_X1 U6954 ( .A(n5782), .ZN(n5783) );
  OAI21_X1 U6955 ( .B1(n5784), .B2(n5783), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n5785) );
  OAI211_X1 U6956 ( .C1(n5787), .C2(n6134), .A(n5786), .B(n5785), .ZN(U2990)
         );
  OAI21_X1 U6957 ( .B1(n5804), .B2(n5665), .A(n5788), .ZN(n5791) );
  OAI21_X1 U6958 ( .B1(n6017), .B2(n5869), .A(n5789), .ZN(n5790) );
  AOI21_X1 U6959 ( .B1(n5791), .B2(n6105), .A(n5790), .ZN(n5792) );
  OAI21_X1 U6960 ( .B1(n5793), .B2(n6134), .A(n5792), .ZN(U2994) );
  NAND2_X1 U6961 ( .A1(n5794), .A2(n6502), .ZN(n5803) );
  AND2_X1 U6962 ( .A1(n5796), .A2(n5795), .ZN(n5797) );
  NOR2_X1 U6963 ( .A1(n5798), .A2(n5797), .ZN(n6063) );
  NOR2_X1 U6964 ( .A1(n5799), .A2(n5665), .ZN(n5800) );
  AOI211_X1 U6965 ( .C1(n6063), .C2(n6499), .A(n5801), .B(n5800), .ZN(n5802)
         );
  OAI211_X1 U6966 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5804), .A(n5803), .B(n5802), .ZN(U2995) );
  OAI21_X1 U6967 ( .B1(n6035), .B2(n5869), .A(n5805), .ZN(n5810) );
  INV_X1 U6968 ( .A(n5806), .ZN(n5819) );
  NOR3_X1 U6969 ( .A1(n5819), .A2(n5808), .A3(n5807), .ZN(n5809) );
  AOI211_X1 U6970 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5816), .A(n5810), .B(n5809), .ZN(n5811) );
  OAI21_X1 U6971 ( .B1(n5812), .B2(n6134), .A(n5811), .ZN(U2996) );
  NAND2_X1 U6972 ( .A1(n5813), .A2(n6502), .ZN(n5818) );
  OAI21_X1 U6973 ( .B1(n6038), .B2(n5869), .A(n5814), .ZN(n5815) );
  AOI21_X1 U6974 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5816), .A(n5815), 
        .ZN(n5817) );
  OAI211_X1 U6975 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5819), .A(n5818), .B(n5817), .ZN(U2997) );
  INV_X1 U6976 ( .A(n5820), .ZN(n5824) );
  NOR3_X1 U6977 ( .A1(n5822), .A2(n5821), .A3(n6115), .ZN(n5823) );
  AOI211_X1 U6978 ( .C1(n6050), .C2(n6499), .A(n5824), .B(n5823), .ZN(n5831)
         );
  NOR2_X1 U6979 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5825), .ZN(n6128)
         );
  INV_X1 U6980 ( .A(n5826), .ZN(n5828) );
  OAI21_X1 U6981 ( .B1(n5828), .B2(n5835), .A(n5827), .ZN(n6131) );
  AOI21_X1 U6982 ( .B1(n5829), .B2(n6128), .A(n6131), .ZN(n6119) );
  OAI21_X1 U6983 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5839), .A(n6119), 
        .ZN(n6110) );
  NAND2_X1 U6984 ( .A1(n6110), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5830) );
  OAI211_X1 U6985 ( .C1(n5832), .C2(n6134), .A(n5831), .B(n5830), .ZN(U2998)
         );
  AOI21_X1 U6986 ( .B1(n5848), .B2(n5708), .A(n5847), .ZN(n5844) );
  INV_X1 U6987 ( .A(n5833), .ZN(n5834) );
  NOR2_X1 U6988 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NOR2_X1 U6989 ( .A1(n5837), .A2(n5836), .ZN(n6463) );
  OAI21_X1 U6990 ( .B1(n5839), .B2(n5838), .A(n6463), .ZN(n5850) );
  NAND2_X1 U6991 ( .A1(n5850), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U6992 ( .C1(n5869), .C2(n6176), .A(n5841), .B(n5840), .ZN(n5842)
         );
  AOI21_X1 U6993 ( .B1(n5844), .B2(n5843), .A(n5842), .ZN(n5845) );
  OAI21_X1 U6994 ( .B1(n5846), .B2(n6134), .A(n5845), .ZN(U3002) );
  INV_X1 U6995 ( .A(n5847), .ZN(n5849) );
  AOI22_X1 U6996 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5850), .B1(n5849), .B2(n5848), .ZN(n5858) );
  AND2_X1 U6997 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NOR2_X1 U6998 ( .A1(n5854), .A2(n5853), .ZN(n6308) );
  INV_X1 U6999 ( .A(n5855), .ZN(n5856) );
  AOI21_X1 U7000 ( .B1(n6308), .B2(n6499), .A(n5856), .ZN(n5857) );
  OAI211_X1 U7001 ( .C1(n5859), .C2(n6134), .A(n5858), .B(n5857), .ZN(U3003)
         );
  NOR3_X1 U7002 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6148), .A3(n5862), 
        .ZN(n5872) );
  OAI21_X1 U7003 ( .B1(n6136), .B2(n5860), .A(n6463), .ZN(n5861) );
  AOI21_X1 U7004 ( .B1(n5863), .B2(n5862), .A(n5861), .ZN(n6143) );
  OAI21_X1 U7005 ( .B1(n5865), .B2(n5864), .A(n6142), .ZN(n5867) );
  AOI21_X1 U7006 ( .B1(n6143), .B2(n5867), .A(n5866), .ZN(n5871) );
  OAI21_X1 U7007 ( .B1(n6197), .B2(n5869), .A(n5868), .ZN(n5870) );
  NOR3_X1 U7008 ( .A1(n5872), .A2(n5871), .A3(n5870), .ZN(n5873) );
  OAI21_X1 U7009 ( .B1(n5874), .B2(n6134), .A(n5873), .ZN(U3004) );
  NOR2_X1 U7010 ( .A1(n5875), .A2(n6134), .ZN(n5880) );
  AOI211_X1 U7011 ( .C1(n6462), .C2(n4342), .A(n6148), .B(n6136), .ZN(n5879)
         );
  AOI21_X1 U7012 ( .B1(n6214), .B2(n6499), .A(n5876), .ZN(n5877) );
  OAI21_X1 U7013 ( .B1(n6463), .B2(n4342), .A(n5877), .ZN(n5878) );
  OR3_X1 U7014 ( .A1(n5880), .A2(n5879), .A3(n5878), .ZN(U3006) );
  NAND2_X1 U7015 ( .A1(n5881), .A2(n6502), .ZN(n5888) );
  OAI211_X1 U7016 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5883), .B(n5882), .ZN(n5887) );
  AOI22_X1 U7017 ( .A1(n6280), .A2(n6499), .B1(n6503), .B2(REIP_REG_4__SCAN_IN), .ZN(n5886) );
  OAI21_X1 U7018 ( .B1(n6488), .B2(n5884), .A(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .ZN(n5885) );
  NAND4_X1 U7019 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(U3014)
         );
  OAI211_X1 U7020 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4573), .A(n5889), .B(
        n5917), .ZN(n5890) );
  OAI21_X1 U7021 ( .B1(n5891), .B2(n4648), .A(n5890), .ZN(n5892) );
  MUX2_X1 U7022 ( .A(n5892), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(n6507), 
        .Z(U3464) );
  NOR2_X1 U7023 ( .A1(n5894), .A2(n5893), .ZN(n5900) );
  OAI22_X1 U7024 ( .A1(n5895), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n5900), .B2(n6603), .ZN(n5896) );
  AOI21_X1 U7025 ( .B1(n5897), .B2(n6608), .A(n5896), .ZN(n6612) );
  OAI222_X1 U7026 ( .A1(n5902), .A2(n5900), .B1(n5904), .B2(n6612), .C1(n5899), 
        .C2(n5898), .ZN(n5901) );
  MUX2_X1 U7027 ( .A(n5901), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n6149), 
        .Z(U3460) );
  OAI22_X1 U7028 ( .A1(n5905), .A2(n5904), .B1(n5903), .B2(n5902), .ZN(n5906)
         );
  MUX2_X1 U7029 ( .A(n5906), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6149), 
        .Z(U3456) );
  INV_X1 U7030 ( .A(n5971), .ZN(n5908) );
  OAI21_X1 U7031 ( .B1(n5908), .B2(n5966), .A(n5907), .ZN(n5909) );
  AOI21_X1 U7032 ( .B1(n5909), .B2(n5914), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5912) );
  NOR2_X1 U7033 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5910), .ZN(n5913)
         );
  NAND2_X1 U7034 ( .A1(n5960), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5924) );
  INV_X1 U7035 ( .A(n5913), .ZN(n5963) );
  INV_X1 U7036 ( .A(n5914), .ZN(n5918) );
  NOR2_X1 U7037 ( .A1(n5915), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5916)
         );
  AOI22_X1 U7038 ( .A1(n5918), .A2(n5917), .B1(n6510), .B2(n5916), .ZN(n5962)
         );
  OAI22_X1 U7039 ( .A1(n5920), .A2(n5963), .B1(n5962), .B2(n5919), .ZN(n5921)
         );
  AOI21_X1 U7040 ( .B1(n5922), .B2(n5966), .A(n5921), .ZN(n5923) );
  OAI211_X1 U7041 ( .C1(n5971), .C2(n5925), .A(n5924), .B(n5923), .ZN(U3036)
         );
  NAND2_X1 U7042 ( .A1(n5960), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5931) );
  OAI22_X1 U7043 ( .A1(n5927), .A2(n5963), .B1(n5962), .B2(n5926), .ZN(n5928)
         );
  AOI21_X1 U7044 ( .B1(n5929), .B2(n5966), .A(n5928), .ZN(n5930) );
  OAI211_X1 U7045 ( .C1(n5971), .C2(n5932), .A(n5931), .B(n5930), .ZN(U3037)
         );
  NAND2_X1 U7046 ( .A1(n5960), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5937) );
  OAI22_X1 U7047 ( .A1(n5934), .A2(n5963), .B1(n5962), .B2(n5933), .ZN(n5935)
         );
  AOI21_X1 U7048 ( .B1(n6569), .B2(n5966), .A(n5935), .ZN(n5936) );
  OAI211_X1 U7049 ( .C1(n5971), .C2(n6574), .A(n5937), .B(n5936), .ZN(U3038)
         );
  NAND2_X1 U7050 ( .A1(n5960), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5942) );
  OAI22_X1 U7051 ( .A1(n5939), .A2(n5963), .B1(n5962), .B2(n5938), .ZN(n5940)
         );
  AOI21_X1 U7052 ( .B1(n6586), .B2(n5966), .A(n5940), .ZN(n5941) );
  OAI211_X1 U7053 ( .C1(n5971), .C2(n6591), .A(n5942), .B(n5941), .ZN(U3039)
         );
  NAND2_X1 U7054 ( .A1(n5960), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5947) );
  OAI22_X1 U7055 ( .A1(n5944), .A2(n5963), .B1(n5962), .B2(n5943), .ZN(n5945)
         );
  AOI21_X1 U7056 ( .B1(n6576), .B2(n5966), .A(n5945), .ZN(n5946) );
  OAI211_X1 U7057 ( .C1(n5971), .C2(n6585), .A(n5947), .B(n5946), .ZN(U3040)
         );
  NAND2_X1 U7058 ( .A1(n5960), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5952) );
  OAI22_X1 U7059 ( .A1(n5949), .A2(n5963), .B1(n5962), .B2(n5948), .ZN(n5950)
         );
  AOI21_X1 U7060 ( .B1(n6592), .B2(n5966), .A(n5950), .ZN(n5951) );
  OAI211_X1 U7061 ( .C1(n5971), .C2(n6602), .A(n5952), .B(n5951), .ZN(U3041)
         );
  NAND2_X1 U7062 ( .A1(n5960), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5958) );
  OAI22_X1 U7063 ( .A1(n5954), .A2(n5963), .B1(n5962), .B2(n5953), .ZN(n5955)
         );
  AOI21_X1 U7064 ( .B1(n5956), .B2(n5966), .A(n5955), .ZN(n5957) );
  OAI211_X1 U7065 ( .C1(n5971), .C2(n5959), .A(n5958), .B(n5957), .ZN(U3042)
         );
  NAND2_X1 U7066 ( .A1(n5960), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5969) );
  OAI22_X1 U7067 ( .A1(n5964), .A2(n5963), .B1(n5962), .B2(n5961), .ZN(n5965)
         );
  AOI21_X1 U7068 ( .B1(n5967), .B2(n5966), .A(n5965), .ZN(n5968) );
  OAI211_X1 U7069 ( .C1(n5971), .C2(n5970), .A(n5969), .B(n5968), .ZN(U3043)
         );
  AND2_X1 U7070 ( .A1(n6344), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7071 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6295), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6245), .ZN(n5980) );
  AOI22_X1 U7072 ( .A1(n5973), .A2(n6250), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5972), .ZN(n5979) );
  NOR2_X1 U7073 ( .A1(n5974), .A2(n6198), .ZN(n5975) );
  AOI21_X1 U7074 ( .B1(n5976), .B2(n6252), .A(n5975), .ZN(n5978) );
  NAND3_X1 U7075 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5981), .A3(n6960), .ZN(
        n5977) );
  NAND4_X1 U7076 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(U2799)
         );
  INV_X1 U7077 ( .A(n5981), .ZN(n5989) );
  NOR2_X1 U7078 ( .A1(n5982), .A2(n6291), .ZN(n5984) );
  OAI22_X1 U7079 ( .A1(n5992), .A2(n6699), .B1(n5440), .B2(n6292), .ZN(n5983)
         );
  AOI211_X1 U7080 ( .C1(n6295), .C2(EBX_REG_27__SCAN_IN), .A(n5984), .B(n5983), 
        .ZN(n5988) );
  AOI22_X1 U7081 ( .A1(n5986), .A2(n6252), .B1(n6297), .B2(n5985), .ZN(n5987)
         );
  OAI211_X1 U7082 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5989), .A(n5988), .B(n5987), .ZN(U2800) );
  AOI22_X1 U7083 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6245), .B1(n5990), 
        .B2(n6250), .ZN(n5997) );
  NOR2_X1 U7084 ( .A1(n6693), .A2(n6001), .ZN(n5999) );
  AOI21_X1 U7085 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5999), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5991) );
  OAI22_X1 U7086 ( .A1(n5993), .A2(n6236), .B1(n5992), .B2(n5991), .ZN(n5994)
         );
  AOI21_X1 U7087 ( .B1(n5995), .B2(n6297), .A(n5994), .ZN(n5996) );
  OAI211_X1 U7088 ( .C1(n5998), .C2(n6246), .A(n5997), .B(n5996), .ZN(U2801)
         );
  AOI22_X1 U7089 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6295), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6245), .ZN(n6006) );
  AOI22_X1 U7090 ( .A1(n6000), .A2(n6250), .B1(n5999), .B2(n6696), .ZN(n6005)
         );
  AOI22_X1 U7091 ( .A1(n6081), .A2(n6252), .B1(n6297), .B2(n6102), .ZN(n6004)
         );
  NOR2_X1 U7092 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6001), .ZN(n6014) );
  INV_X1 U7093 ( .A(n6025), .ZN(n6002) );
  OAI21_X1 U7094 ( .B1(n6014), .B2(n6002), .A(REIP_REG_25__SCAN_IN), .ZN(n6003) );
  NAND4_X1 U7095 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(U2802)
         );
  INV_X1 U7096 ( .A(n6007), .ZN(n6008) );
  AOI22_X1 U7097 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6245), .B1(n6250), 
        .B2(n6008), .ZN(n6010) );
  NAND2_X1 U7098 ( .A1(n6295), .A2(EBX_REG_24__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U7099 ( .C1(n6025), .C2(n6693), .A(n6010), .B(n6009), .ZN(n6011)
         );
  AOI21_X1 U7100 ( .B1(n6012), .B2(n6252), .A(n6011), .ZN(n6013) );
  INV_X1 U7101 ( .A(n6013), .ZN(n6015) );
  NOR2_X1 U7102 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  OAI21_X1 U7103 ( .B1(n6017), .B2(n6198), .A(n6016), .ZN(U2803) );
  INV_X1 U7104 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U7105 ( .A1(n6902), .A2(n6026), .ZN(n6030) );
  AOI21_X1 U7106 ( .B1(REIP_REG_22__SCAN_IN), .B2(n6030), .A(
        REIP_REG_23__SCAN_IN), .ZN(n6024) );
  INV_X1 U7107 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6019) );
  OAI22_X1 U7108 ( .A1(n6019), .A2(n6292), .B1(n6018), .B2(n6291), .ZN(n6020)
         );
  AOI21_X1 U7109 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6295), .A(n6020), .ZN(n6023)
         );
  AOI22_X1 U7110 ( .A1(n6067), .A2(n6252), .B1(n6297), .B2(n6063), .ZN(n6022)
         );
  OAI211_X1 U7111 ( .C1(n6025), .C2(n6024), .A(n6023), .B(n6022), .ZN(U2804)
         );
  NOR2_X1 U7112 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6026), .ZN(n6040) );
  INV_X1 U7113 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7093) );
  AOI22_X1 U7114 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6245), .B1(n6250), 
        .B2(n6027), .ZN(n6028) );
  OAI21_X1 U7115 ( .B1(n6246), .B2(n5591), .A(n6028), .ZN(n6029) );
  AOI21_X1 U7116 ( .B1(n6030), .B2(n7093), .A(n6029), .ZN(n6031) );
  OAI21_X1 U7117 ( .B1(n6032), .B2(n6236), .A(n6031), .ZN(n6033) );
  AOI221_X1 U7118 ( .B1(n6040), .B2(REIP_REG_22__SCAN_IN), .C1(n6046), .C2(
        REIP_REG_22__SCAN_IN), .A(n6033), .ZN(n6034) );
  OAI21_X1 U7119 ( .B1(n6035), .B2(n6198), .A(n6034), .ZN(U2805) );
  AOI22_X1 U7120 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6295), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6245), .ZN(n6044) );
  INV_X1 U7121 ( .A(n6036), .ZN(n6037) );
  AOI22_X1 U7122 ( .A1(n6037), .A2(n6250), .B1(REIP_REG_21__SCAN_IN), .B2(
        n6046), .ZN(n6043) );
  INV_X1 U7123 ( .A(n6038), .ZN(n6039) );
  AOI22_X1 U7124 ( .A1(n6070), .A2(n6252), .B1(n6297), .B2(n6039), .ZN(n6042)
         );
  INV_X1 U7125 ( .A(n6040), .ZN(n6041) );
  NAND4_X1 U7126 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(U2806)
         );
  AOI22_X1 U7127 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6295), .B1(n6045), .B2(n6250), .ZN(n6052) );
  INV_X1 U7128 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6692) );
  NOR2_X1 U7129 ( .A1(n6882), .A2(n6692), .ZN(n6062) );
  AOI21_X1 U7130 ( .B1(n6062), .B2(n6054), .A(REIP_REG_20__SCAN_IN), .ZN(n6048) );
  INV_X1 U7131 ( .A(n6046), .ZN(n6047) );
  OAI22_X1 U7132 ( .A1(n6073), .A2(n6236), .B1(n6048), .B2(n6047), .ZN(n6049)
         );
  AOI21_X1 U7133 ( .B1(n6297), .B2(n6050), .A(n6049), .ZN(n6051) );
  OAI211_X1 U7134 ( .C1(n6053), .C2(n6292), .A(n6052), .B(n6051), .ZN(U2807)
         );
  OAI21_X1 U7135 ( .B1(REIP_REG_18__SCAN_IN), .B2(REIP_REG_19__SCAN_IN), .A(
        n6054), .ZN(n6061) );
  INV_X1 U7136 ( .A(n6055), .ZN(n6056) );
  AOI22_X1 U7137 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6295), .B1(n6056), .B2(
        REIP_REG_19__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7138 ( .B1(n6090), .B2(n6291), .A(n6057), .ZN(n6058) );
  AOI211_X1 U7139 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6503), 
        .B(n6058), .ZN(n6060) );
  AOI22_X1 U7140 ( .A1(n6087), .A2(n6252), .B1(n6297), .B2(n6111), .ZN(n6059)
         );
  OAI211_X1 U7141 ( .C1(n6062), .C2(n6061), .A(n6060), .B(n6059), .ZN(U2808)
         );
  AOI22_X1 U7142 ( .A1(n6067), .A2(n6318), .B1(n6063), .B2(n6317), .ZN(n6064)
         );
  OAI21_X1 U7143 ( .B1(n6322), .B2(n6065), .A(n6064), .ZN(U2836) );
  INV_X1 U7144 ( .A(n6066), .ZN(n6324) );
  AOI22_X1 U7145 ( .A1(n6067), .A2(n6324), .B1(n6323), .B2(DATAI_23_), .ZN(
        n6069) );
  AOI22_X1 U7146 ( .A1(n6327), .A2(DATAI_7_), .B1(n6326), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7147 ( .A1(n6069), .A2(n6068), .ZN(U2868) );
  AOI22_X1 U7148 ( .A1(n6070), .A2(n6324), .B1(n6323), .B2(DATAI_21_), .ZN(
        n6072) );
  AOI22_X1 U7149 ( .A1(n6327), .A2(DATAI_5_), .B1(n6326), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7150 ( .A1(n6072), .A2(n6071), .ZN(U2870) );
  INV_X1 U7151 ( .A(n6073), .ZN(n6074) );
  AOI22_X1 U7152 ( .A1(n6074), .A2(n6324), .B1(n6323), .B2(DATAI_20_), .ZN(
        n6076) );
  AOI22_X1 U7153 ( .A1(n6327), .A2(DATAI_4_), .B1(n6326), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7154 ( .A1(n6076), .A2(n6075), .ZN(U2871) );
  AOI22_X1 U7155 ( .A1(n6087), .A2(n6324), .B1(n6323), .B2(DATAI_19_), .ZN(
        n6078) );
  AOI22_X1 U7156 ( .A1(n6327), .A2(DATAI_3_), .B1(n6326), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7157 ( .A1(n6078), .A2(n6077), .ZN(U2872) );
  AOI22_X1 U7158 ( .A1(n6503), .A2(REIP_REG_25__SCAN_IN), .B1(n6448), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6083) );
  INV_X1 U7159 ( .A(n5432), .ZN(n6080) );
  OAI21_X1 U7160 ( .B1(n6080), .B2(n3200), .A(n4431), .ZN(n6103) );
  AOI22_X1 U7161 ( .A1(n6081), .A2(n6441), .B1(n6450), .B2(n6103), .ZN(n6082)
         );
  OAI211_X1 U7162 ( .C1(n6446), .C2(n6084), .A(n6083), .B(n6082), .ZN(U2961)
         );
  AOI22_X1 U7163 ( .A1(n6503), .A2(REIP_REG_19__SCAN_IN), .B1(n6448), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6089) );
  XNOR2_X1 U7164 ( .A(n4260), .B(n6085), .ZN(n6086) );
  XNOR2_X1 U7165 ( .A(n5658), .B(n6086), .ZN(n6112) );
  AOI22_X1 U7166 ( .A1(n6450), .A2(n6112), .B1(n6087), .B2(n6441), .ZN(n6088)
         );
  OAI211_X1 U7167 ( .C1(n6446), .C2(n6090), .A(n6089), .B(n6088), .ZN(U2967)
         );
  AND3_X1 U7168 ( .A1(n3161), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n4260), 
        .ZN(n6091) );
  OR2_X1 U7169 ( .A1(n6092), .A2(n6091), .ZN(n6093) );
  XNOR2_X1 U7170 ( .A(n6093), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6135)
         );
  INV_X1 U7171 ( .A(n6135), .ZN(n6097) );
  INV_X1 U7172 ( .A(n6094), .ZN(n6096) );
  AOI222_X1 U7173 ( .A1(n6097), .A2(n6450), .B1(n6096), .B2(n6095), .C1(n6441), 
        .C2(n6325), .ZN(n6099) );
  NOR2_X1 U7174 ( .A1(n6120), .A2(n6845), .ZN(n6127) );
  INV_X1 U7175 ( .A(n6127), .ZN(n6098) );
  OAI211_X1 U7176 ( .C1(n6101), .C2(n6100), .A(n6099), .B(n6098), .ZN(U2969)
         );
  AOI22_X1 U7177 ( .A1(n6103), .A2(n6502), .B1(n6499), .B2(n6102), .ZN(n6109)
         );
  NOR2_X1 U7178 ( .A1(n6120), .A2(n6696), .ZN(n6104) );
  AOI221_X1 U7179 ( .B1(n6107), .B2(n6106), .C1(n6105), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6104), .ZN(n6108) );
  NAND2_X1 U7180 ( .A1(n6109), .A2(n6108), .ZN(U2993) );
  AOI22_X1 U7181 ( .A1(n6503), .A2(REIP_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n6110), .ZN(n6114) );
  AOI22_X1 U7182 ( .A1(n6112), .A2(n6502), .B1(n6499), .B2(n6111), .ZN(n6113)
         );
  OAI211_X1 U7183 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6115), .A(n6114), .B(n6113), .ZN(U2999) );
  INV_X1 U7184 ( .A(n6116), .ZN(n6118) );
  AOI22_X1 U7185 ( .A1(n6118), .A2(n6502), .B1(n6499), .B2(n6117), .ZN(n6126)
         );
  INV_X1 U7186 ( .A(n6119), .ZN(n6122) );
  NOR2_X1 U7187 ( .A1(n6120), .A2(n6882), .ZN(n6121) );
  AOI221_X1 U7188 ( .B1(n6124), .B2(n6123), .C1(n6122), .C2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6121), .ZN(n6125) );
  NAND2_X1 U7189 ( .A1(n6126), .A2(n6125), .ZN(U3000) );
  AOI21_X1 U7190 ( .B1(n6128), .B2(n6458), .A(n6127), .ZN(n6133) );
  INV_X1 U7191 ( .A(n6129), .ZN(n6130) );
  AOI22_X1 U7192 ( .A1(n6131), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n6499), .B2(n6130), .ZN(n6132) );
  OAI211_X1 U7193 ( .C1(n6135), .C2(n6134), .A(n6133), .B(n6132), .ZN(U3001)
         );
  NAND2_X1 U7194 ( .A1(n6136), .A2(n6142), .ZN(n6147) );
  OR2_X1 U7195 ( .A1(n6138), .A2(n6137), .ZN(n6140) );
  AND2_X1 U7196 ( .A1(n6140), .A2(n6139), .ZN(n6316) );
  AOI22_X1 U7197 ( .A1(n6316), .A2(n6499), .B1(n6503), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n6141) );
  OAI21_X1 U7198 ( .B1(n6143), .B2(n6142), .A(n6141), .ZN(n6144) );
  AOI21_X1 U7199 ( .B1(n6145), .B2(n6502), .A(n6144), .ZN(n6146) );
  OAI21_X1 U7200 ( .B1(n6148), .B2(n6147), .A(n6146), .ZN(U3005) );
  INV_X1 U7201 ( .A(n6149), .ZN(n6154) );
  INV_X1 U7202 ( .A(n6150), .ZN(n6152) );
  NAND3_X1 U7203 ( .A1(n6152), .A2(n5471), .A3(n6151), .ZN(n6153) );
  OAI21_X1 U7204 ( .B1(n6154), .B2(n3543), .A(n6153), .ZN(U3455) );
  AOI21_X1 U7205 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6671), .A(n4234), .ZN(n6159) );
  INV_X1 U7206 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6777) );
  INV_X2 U7207 ( .A(n7121), .ZN(n6716) );
  AOI21_X1 U7208 ( .B1(n6159), .B2(n6777), .A(n6716), .ZN(U2789) );
  INV_X1 U7209 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6825) );
  NOR2_X1 U7210 ( .A1(n6155), .A2(n6825), .ZN(n6156) );
  NAND2_X1 U7211 ( .A1(n6352), .A2(n6156), .ZN(n6157) );
  OAI21_X1 U7212 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6644), .A(n6157), .ZN(
        U2790) );
  NOR2_X1 U7213 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6160) );
  OAI21_X1 U7214 ( .B1(n6160), .B2(D_C_N_REG_SCAN_IN), .A(n7121), .ZN(n6158)
         );
  OAI21_X1 U7215 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7121), .A(n6158), .ZN(
        U2791) );
  NOR2_X2 U7216 ( .A1(n6716), .A2(n6159), .ZN(n6705) );
  OAI21_X1 U7217 ( .B1(BS16_N), .B2(n6160), .A(n6705), .ZN(n6704) );
  OAI21_X1 U7218 ( .B1(n6705), .B2(n7092), .A(n6704), .ZN(U2792) );
  OAI21_X1 U7219 ( .B1(n6162), .B2(n6858), .A(n6161), .ZN(U2793) );
  NOR4_X1 U7220 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6172)
         );
  AOI211_X1 U7221 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_7__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n6171) );
  NOR4_X1 U7222 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6163)
         );
  INV_X1 U7223 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6815) );
  INV_X1 U7224 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6843) );
  NAND3_X1 U7225 ( .A1(n6163), .A2(n6815), .A3(n6843), .ZN(n6169) );
  NOR4_X1 U7226 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6167) );
  NOR4_X1 U7227 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6166) );
  NOR4_X1 U7228 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6165) );
  NOR4_X1 U7229 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7230 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n6168)
         );
  NOR4_X1 U7231 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(n6169), .A4(n6168), .ZN(n6170) );
  NAND3_X1 U7232 ( .A1(n6172), .A2(n6171), .A3(n6170), .ZN(n6711) );
  INV_X1 U7233 ( .A(n6711), .ZN(n6713) );
  INV_X1 U7234 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7064) );
  OR4_X1 U7235 ( .A1(n6711), .A2(REIP_REG_0__SCAN_IN), .A3(
        DATAWIDTH_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6173)
         );
  OAI221_X1 U7236 ( .B1(n6713), .B2(n7064), .C1(n6711), .C2(n5196), .A(n6173), 
        .ZN(U2794) );
  NAND2_X1 U7237 ( .A1(n6713), .A2(n5196), .ZN(n6714) );
  NAND2_X1 U7238 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6711), .ZN(n6174) );
  OAI211_X1 U7239 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(n6714), .A(n6174), .B(
        n6173), .ZN(U2795) );
  AOI21_X1 U7240 ( .B1(n6245), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6503), 
        .ZN(n6184) );
  NAND2_X1 U7241 ( .A1(n6271), .A2(n6175), .ZN(n6194) );
  INV_X1 U7242 ( .A(n6194), .ZN(n6188) );
  AOI22_X1 U7243 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6295), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6188), .ZN(n6183) );
  OAI22_X1 U7244 ( .A1(n6177), .A2(n6236), .B1(n6198), .B2(n6176), .ZN(n6178)
         );
  AOI21_X1 U7245 ( .B1(n6179), .B2(n6250), .A(n6178), .ZN(n6182) );
  OAI211_X1 U7246 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n6185), .B(n6180), .ZN(n6181) );
  NAND4_X1 U7247 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(U2811)
         );
  INV_X1 U7248 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U7249 ( .A1(n6297), .A2(n6308), .B1(n6185), .B2(n6689), .ZN(n6193)
         );
  OAI22_X1 U7250 ( .A1(n6315), .A2(n6246), .B1(n6186), .B2(n6292), .ZN(n6187)
         );
  AOI211_X1 U7251 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6188), .A(n6503), .B(n6187), .ZN(n6192) );
  OAI22_X1 U7252 ( .A1(n6312), .A2(n6236), .B1(n6291), .B2(n6189), .ZN(n6190)
         );
  INV_X1 U7253 ( .A(n6190), .ZN(n6191) );
  NAND3_X1 U7254 ( .A1(n6193), .A2(n6192), .A3(n6191), .ZN(U2812) );
  AOI21_X1 U7255 ( .B1(n6686), .B2(n6195), .A(n6194), .ZN(n6196) );
  AOI211_X1 U7256 ( .C1(n6295), .C2(EBX_REG_14__SCAN_IN), .A(n6503), .B(n6196), 
        .ZN(n6203) );
  OAI22_X1 U7257 ( .A1(n6199), .A2(n6236), .B1(n6198), .B2(n6197), .ZN(n6200)
         );
  AOI21_X1 U7258 ( .B1(n6201), .B2(n6250), .A(n6200), .ZN(n6202) );
  OAI211_X1 U7259 ( .C1(n5738), .C2(n6292), .A(n6203), .B(n6202), .ZN(U2813)
         );
  AOI22_X1 U7260 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6295), .B1(n6297), .B2(n6316), .ZN(n6212) );
  NOR3_X1 U7261 ( .A1(n6278), .A2(REIP_REG_13__SCAN_IN), .A3(n6204), .ZN(n6205) );
  AOI211_X1 U7262 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6503), 
        .B(n6205), .ZN(n6211) );
  INV_X1 U7263 ( .A(n6206), .ZN(n6207) );
  AOI22_X1 U7264 ( .A1(n6319), .A2(n6252), .B1(n6250), .B2(n6207), .ZN(n6210)
         );
  NOR4_X1 U7265 ( .A1(n6278), .A2(n6684), .A3(REIP_REG_12__SCAN_IN), .A4(n6208), .ZN(n6213) );
  OAI21_X1 U7266 ( .B1(n6215), .B2(n6213), .A(REIP_REG_13__SCAN_IN), .ZN(n6209) );
  NAND4_X1 U7267 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(U2814)
         );
  AOI21_X1 U7268 ( .B1(n6214), .B2(n6297), .A(n6213), .ZN(n6221) );
  AOI22_X1 U7269 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6245), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6215), .ZN(n6220) );
  AOI21_X1 U7270 ( .B1(n6295), .B2(EBX_REG_12__SCAN_IN), .A(n6503), .ZN(n6219)
         );
  AOI22_X1 U7271 ( .A1(n6217), .A2(n6252), .B1(n6250), .B2(n6216), .ZN(n6218)
         );
  NAND4_X1 U7272 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(U2815)
         );
  AOI221_X1 U7273 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .C1(
        n6682), .C2(n5322), .A(n6222), .ZN(n6223) );
  AOI21_X1 U7274 ( .B1(n6224), .B2(n6297), .A(n6223), .ZN(n6231) );
  AOI22_X1 U7275 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6295), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6245), .ZN(n6230) );
  AOI21_X1 U7276 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6225), .A(n6503), .ZN(n6229) );
  AOI22_X1 U7277 ( .A1(n6227), .A2(n6252), .B1(n6250), .B2(n6226), .ZN(n6228)
         );
  NAND4_X1 U7278 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(U2817)
         );
  AOI21_X1 U7279 ( .B1(n6245), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6503), 
        .ZN(n6243) );
  AOI22_X1 U7280 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6295), .B1(n6297), .B2(n6474), 
        .ZN(n6242) );
  INV_X1 U7281 ( .A(n6234), .ZN(n6233) );
  OAI21_X1 U7282 ( .B1(n6278), .B2(n6233), .A(n6232), .ZN(n6265) );
  NOR3_X1 U7283 ( .A1(n6278), .A2(REIP_REG_6__SCAN_IN), .A3(n6234), .ZN(n6249)
         );
  OAI22_X1 U7284 ( .A1(n6237), .A2(n6236), .B1(n6235), .B2(n6291), .ZN(n6238)
         );
  AOI221_X1 U7285 ( .B1(n6265), .B2(REIP_REG_7__SCAN_IN), .C1(n6249), .C2(
        REIP_REG_7__SCAN_IN), .A(n6238), .ZN(n6241) );
  NAND3_X1 U7286 ( .A1(n6264), .A2(n6680), .A3(n6239), .ZN(n6240) );
  NAND4_X1 U7287 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(U2820)
         );
  AOI22_X1 U7288 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6245), .B1(n6297), 
        .B2(n6244), .ZN(n6256) );
  NOR2_X1 U7289 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  AOI211_X1 U7290 ( .C1(n6265), .C2(REIP_REG_6__SCAN_IN), .A(n6249), .B(n6248), 
        .ZN(n6255) );
  AOI22_X1 U7291 ( .A1(n6253), .A2(n6252), .B1(n6251), .B2(n6250), .ZN(n6254)
         );
  NAND4_X1 U7292 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6259), .ZN(U2821)
         );
  INV_X1 U7293 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6260) );
  AOI22_X1 U7294 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6295), .B1(n6297), .B2(n6257), 
        .ZN(n6258) );
  OAI211_X1 U7295 ( .C1(n6292), .C2(n6260), .A(n6259), .B(n6258), .ZN(n6261)
         );
  AOI21_X1 U7296 ( .B1(n6262), .B2(n6303), .A(n6261), .ZN(n6268) );
  AND2_X1 U7297 ( .A1(n6264), .A2(n6263), .ZN(n6266) );
  OAI21_X1 U7298 ( .B1(n6266), .B2(REIP_REG_5__SCAN_IN), .A(n6265), .ZN(n6267)
         );
  OAI211_X1 U7299 ( .C1(n6291), .C2(n6269), .A(n6268), .B(n6267), .ZN(U2822)
         );
  INV_X1 U7300 ( .A(n6270), .ZN(n6287) );
  OAI21_X1 U7301 ( .B1(n6272), .B2(n6277), .A(n6271), .ZN(n6307) );
  OAI22_X1 U7302 ( .A1(n6307), .A2(n6674), .B1(n6273), .B2(n6292), .ZN(n6274)
         );
  AOI211_X1 U7303 ( .C1(n6295), .C2(EBX_REG_4__SCAN_IN), .A(n6503), .B(n6274), 
        .ZN(n6286) );
  INV_X1 U7304 ( .A(n6275), .ZN(n6284) );
  INV_X1 U7305 ( .A(n6276), .ZN(n6282) );
  NOR3_X1 U7306 ( .A1(n6278), .A2(REIP_REG_4__SCAN_IN), .A3(n6277), .ZN(n6279)
         );
  AOI21_X1 U7307 ( .B1(n6280), .B2(n6297), .A(n6279), .ZN(n6281) );
  OAI21_X1 U7308 ( .B1(n6282), .B2(n6300), .A(n6281), .ZN(n6283) );
  AOI21_X1 U7309 ( .B1(n6284), .B2(n6303), .A(n6283), .ZN(n6285) );
  OAI211_X1 U7310 ( .C1(n6287), .C2(n6291), .A(n6286), .B(n6285), .ZN(U2823)
         );
  OR2_X1 U7311 ( .A1(n6289), .A2(n6288), .ZN(n6306) );
  OAI22_X1 U7312 ( .A1(n6293), .A2(n6292), .B1(n6291), .B2(n6290), .ZN(n6294)
         );
  AOI21_X1 U7313 ( .B1(n6295), .B2(EBX_REG_3__SCAN_IN), .A(n6294), .ZN(n6299)
         );
  NAND2_X1 U7314 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  OAI211_X1 U7315 ( .C1(n6301), .C2(n6300), .A(n6299), .B(n6298), .ZN(n6302)
         );
  AOI21_X1 U7316 ( .B1(n6304), .B2(n6303), .A(n6302), .ZN(n6305) );
  OAI221_X1 U7317 ( .B1(n6307), .B2(n6673), .C1(n6307), .C2(n6306), .A(n6305), 
        .ZN(U2824) );
  INV_X1 U7318 ( .A(n6308), .ZN(n6309) );
  OAI22_X1 U7319 ( .A1(n6312), .A2(n6311), .B1(n6310), .B2(n6309), .ZN(n6313)
         );
  INV_X1 U7320 ( .A(n6313), .ZN(n6314) );
  OAI21_X1 U7321 ( .B1(n6322), .B2(n6315), .A(n6314), .ZN(U2844) );
  AOI22_X1 U7322 ( .A1(n6319), .A2(n6318), .B1(n6317), .B2(n6316), .ZN(n6320)
         );
  OAI21_X1 U7323 ( .B1(n6322), .B2(n6321), .A(n6320), .ZN(U2846) );
  AOI22_X1 U7324 ( .A1(n6325), .A2(n6324), .B1(n6323), .B2(DATAI_17_), .ZN(
        n6329) );
  AOI22_X1 U7325 ( .A1(n6327), .A2(DATAI_1_), .B1(n6326), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7326 ( .A1(n6329), .A2(n6328), .ZN(U2874) );
  AOI22_X1 U7327 ( .A1(n6719), .A2(LWORD_REG_15__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6331) );
  OAI21_X1 U7328 ( .B1(n6436), .B2(n6349), .A(n6331), .ZN(U2908) );
  AOI22_X1 U7329 ( .A1(n6719), .A2(LWORD_REG_14__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6332) );
  OAI21_X1 U7330 ( .B1(n6431), .B2(n6349), .A(n6332), .ZN(U2909) );
  AOI22_X1 U7331 ( .A1(n6719), .A2(LWORD_REG_13__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6333) );
  OAI21_X1 U7332 ( .B1(n6428), .B2(n6349), .A(n6333), .ZN(U2910) );
  AOI22_X1 U7333 ( .A1(n6719), .A2(LWORD_REG_12__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6334) );
  OAI21_X1 U7334 ( .B1(n6425), .B2(n6349), .A(n6334), .ZN(U2911) );
  AOI22_X1 U7335 ( .A1(n6719), .A2(LWORD_REG_11__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6335) );
  OAI21_X1 U7336 ( .B1(n6421), .B2(n6349), .A(n6335), .ZN(U2912) );
  AOI22_X1 U7337 ( .A1(n6719), .A2(LWORD_REG_10__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6336) );
  OAI21_X1 U7338 ( .B1(n6418), .B2(n6349), .A(n6336), .ZN(U2913) );
  AOI22_X1 U7339 ( .A1(n6719), .A2(LWORD_REG_9__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7340 ( .B1(n6415), .B2(n6349), .A(n6337), .ZN(U2914) );
  AOI22_X1 U7341 ( .A1(n6719), .A2(LWORD_REG_8__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7342 ( .B1(n6412), .B2(n6349), .A(n6338), .ZN(U2915) );
  AOI22_X1 U7343 ( .A1(n6719), .A2(LWORD_REG_7__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U7344 ( .B1(n6409), .B2(n6349), .A(n6339), .ZN(U2916) );
  AOI22_X1 U7345 ( .A1(n6719), .A2(LWORD_REG_6__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U7346 ( .B1(n6406), .B2(n6349), .A(n6340), .ZN(U2917) );
  AOI22_X1 U7347 ( .A1(n6719), .A2(LWORD_REG_5__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7348 ( .B1(n6403), .B2(n6349), .A(n6341), .ZN(U2918) );
  AOI22_X1 U7349 ( .A1(n6719), .A2(LWORD_REG_4__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U7350 ( .B1(n6400), .B2(n6349), .A(n6342), .ZN(U2919) );
  AOI22_X1 U7351 ( .A1(n6719), .A2(LWORD_REG_3__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6343) );
  OAI21_X1 U7352 ( .B1(n6397), .B2(n6349), .A(n6343), .ZN(U2920) );
  AOI22_X1 U7353 ( .A1(n6719), .A2(LWORD_REG_2__SCAN_IN), .B1(n6344), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U7354 ( .B1(n6394), .B2(n6349), .A(n6345), .ZN(U2921) );
  AOI22_X1 U7355 ( .A1(n6719), .A2(LWORD_REG_1__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6346) );
  OAI21_X1 U7356 ( .B1(n6391), .B2(n6349), .A(n6346), .ZN(U2922) );
  AOI22_X1 U7357 ( .A1(n6719), .A2(LWORD_REG_0__SCAN_IN), .B1(n6347), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7358 ( .B1(n6388), .B2(n6349), .A(n6348), .ZN(U2923) );
  INV_X1 U7359 ( .A(n6632), .ZN(n6350) );
  NAND2_X2 U7360 ( .A1(n6351), .A2(n6350), .ZN(n6435) );
  INV_X1 U7361 ( .A(n6352), .ZN(n6353) );
  AND2_X1 U7362 ( .A1(n6432), .A2(DATAI_0_), .ZN(n6386) );
  AOI21_X1 U7363 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6433), .A(n6386), .ZN(n6356) );
  OAI21_X1 U7364 ( .B1(n6357), .B2(n6435), .A(n6356), .ZN(U2924) );
  AND2_X1 U7365 ( .A1(n6432), .A2(DATAI_1_), .ZN(n6389) );
  AOI21_X1 U7366 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6423), .A(n6389), .ZN(n6358) );
  OAI21_X1 U7367 ( .B1(n6359), .B2(n6435), .A(n6358), .ZN(U2925) );
  AND2_X1 U7368 ( .A1(n6432), .A2(DATAI_2_), .ZN(n6392) );
  AOI21_X1 U7369 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6433), .A(n6392), .ZN(n6360) );
  OAI21_X1 U7370 ( .B1(n6361), .B2(n6435), .A(n6360), .ZN(U2926) );
  AND2_X1 U7371 ( .A1(n6432), .A2(DATAI_3_), .ZN(n6395) );
  AOI21_X1 U7372 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6423), .A(n6395), .ZN(n6362) );
  OAI21_X1 U7373 ( .B1(n6363), .B2(n6435), .A(n6362), .ZN(U2927) );
  AND2_X1 U7374 ( .A1(n6432), .A2(DATAI_4_), .ZN(n6398) );
  AOI21_X1 U7375 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6423), .A(n6398), .ZN(n6364) );
  OAI21_X1 U7376 ( .B1(n6365), .B2(n6435), .A(n6364), .ZN(U2928) );
  AND2_X1 U7377 ( .A1(n6432), .A2(DATAI_5_), .ZN(n6401) );
  AOI21_X1 U7378 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6423), .A(n6401), .ZN(n6366) );
  OAI21_X1 U7379 ( .B1(n6367), .B2(n6435), .A(n6366), .ZN(U2929) );
  AND2_X1 U7380 ( .A1(n6432), .A2(DATAI_6_), .ZN(n6404) );
  AOI21_X1 U7381 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6423), .A(n6404), .ZN(n6368) );
  OAI21_X1 U7382 ( .B1(n6369), .B2(n6435), .A(n6368), .ZN(U2930) );
  AND2_X1 U7383 ( .A1(n6432), .A2(DATAI_7_), .ZN(n6407) );
  AOI21_X1 U7384 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6423), .A(n6407), .ZN(n6370) );
  OAI21_X1 U7385 ( .B1(n6371), .B2(n6435), .A(n6370), .ZN(U2931) );
  AND2_X1 U7386 ( .A1(n6432), .A2(DATAI_8_), .ZN(n6410) );
  AOI21_X1 U7387 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6423), .A(n6410), .ZN(n6372) );
  OAI21_X1 U7388 ( .B1(n6373), .B2(n6435), .A(n6372), .ZN(U2932) );
  AND2_X1 U7389 ( .A1(n6432), .A2(DATAI_9_), .ZN(n6413) );
  AOI21_X1 U7390 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6423), .A(n6413), .ZN(n6374) );
  OAI21_X1 U7391 ( .B1(n6375), .B2(n6435), .A(n6374), .ZN(U2933) );
  AND2_X1 U7392 ( .A1(n6432), .A2(DATAI_10_), .ZN(n6416) );
  AOI21_X1 U7393 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6423), .A(n6416), .ZN(
        n6376) );
  OAI21_X1 U7394 ( .B1(n6377), .B2(n6435), .A(n6376), .ZN(U2934) );
  AND2_X1 U7395 ( .A1(n6432), .A2(DATAI_11_), .ZN(n6419) );
  AOI21_X1 U7396 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6423), .A(n6419), .ZN(
        n6378) );
  OAI21_X1 U7397 ( .B1(n6379), .B2(n6435), .A(n6378), .ZN(U2935) );
  AND2_X1 U7398 ( .A1(n6432), .A2(DATAI_12_), .ZN(n6422) );
  AOI21_X1 U7399 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6423), .A(n6422), .ZN(
        n6380) );
  OAI21_X1 U7400 ( .B1(n6381), .B2(n6435), .A(n6380), .ZN(U2936) );
  AND2_X1 U7401 ( .A1(n6432), .A2(DATAI_13_), .ZN(n6426) );
  AOI21_X1 U7402 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6423), .A(n6426), .ZN(
        n6382) );
  OAI21_X1 U7403 ( .B1(n6383), .B2(n6435), .A(n6382), .ZN(U2937) );
  AND2_X1 U7404 ( .A1(n6432), .A2(DATAI_14_), .ZN(n6429) );
  AOI21_X1 U7405 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6423), .A(n6429), .ZN(
        n6384) );
  OAI21_X1 U7406 ( .B1(n6385), .B2(n6435), .A(n6384), .ZN(U2938) );
  AOI21_X1 U7407 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6423), .A(n6386), .ZN(n6387) );
  OAI21_X1 U7408 ( .B1(n6388), .B2(n6435), .A(n6387), .ZN(U2939) );
  AOI21_X1 U7409 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6423), .A(n6389), .ZN(n6390) );
  OAI21_X1 U7410 ( .B1(n6391), .B2(n6435), .A(n6390), .ZN(U2940) );
  AOI21_X1 U7411 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6423), .A(n6392), .ZN(n6393) );
  OAI21_X1 U7412 ( .B1(n6394), .B2(n6435), .A(n6393), .ZN(U2941) );
  AOI21_X1 U7413 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6423), .A(n6395), .ZN(n6396) );
  OAI21_X1 U7414 ( .B1(n6397), .B2(n6435), .A(n6396), .ZN(U2942) );
  AOI21_X1 U7415 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6423), .A(n6398), .ZN(n6399) );
  OAI21_X1 U7416 ( .B1(n6400), .B2(n6435), .A(n6399), .ZN(U2943) );
  AOI21_X1 U7417 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6423), .A(n6401), .ZN(n6402) );
  OAI21_X1 U7418 ( .B1(n6403), .B2(n6435), .A(n6402), .ZN(U2944) );
  AOI21_X1 U7419 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6423), .A(n6404), .ZN(n6405) );
  OAI21_X1 U7420 ( .B1(n6406), .B2(n6435), .A(n6405), .ZN(U2945) );
  AOI21_X1 U7421 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6423), .A(n6407), .ZN(n6408) );
  OAI21_X1 U7422 ( .B1(n6409), .B2(n6435), .A(n6408), .ZN(U2946) );
  AOI21_X1 U7423 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6423), .A(n6410), .ZN(n6411) );
  OAI21_X1 U7424 ( .B1(n6412), .B2(n6435), .A(n6411), .ZN(U2947) );
  AOI21_X1 U7425 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6423), .A(n6413), .ZN(n6414) );
  OAI21_X1 U7426 ( .B1(n6415), .B2(n6435), .A(n6414), .ZN(U2948) );
  AOI21_X1 U7427 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6423), .A(n6416), .ZN(
        n6417) );
  OAI21_X1 U7428 ( .B1(n6418), .B2(n6435), .A(n6417), .ZN(U2949) );
  AOI21_X1 U7429 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6423), .A(n6419), .ZN(
        n6420) );
  OAI21_X1 U7430 ( .B1(n6421), .B2(n6435), .A(n6420), .ZN(U2950) );
  AOI21_X1 U7431 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6423), .A(n6422), .ZN(
        n6424) );
  OAI21_X1 U7432 ( .B1(n6425), .B2(n6435), .A(n6424), .ZN(U2951) );
  AOI21_X1 U7433 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6433), .A(n6426), .ZN(
        n6427) );
  OAI21_X1 U7434 ( .B1(n6428), .B2(n6435), .A(n6427), .ZN(U2952) );
  AOI21_X1 U7435 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6433), .A(n6429), .ZN(
        n6430) );
  OAI21_X1 U7436 ( .B1(n6431), .B2(n6435), .A(n6430), .ZN(U2953) );
  AOI22_X1 U7437 ( .A1(n6433), .A2(LWORD_REG_15__SCAN_IN), .B1(n6432), .B2(
        DATAI_15_), .ZN(n6434) );
  OAI21_X1 U7438 ( .B1(n6436), .B2(n6435), .A(n6434), .ZN(U2954) );
  AOI22_X1 U7439 ( .A1(n6503), .A2(REIP_REG_2__SCAN_IN), .B1(n6448), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U7440 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  XOR2_X1 U7441 ( .A(n6440), .B(n6439), .Z(n6487) );
  AOI22_X1 U7442 ( .A1(n6487), .A2(n6450), .B1(n6442), .B2(n6441), .ZN(n6443)
         );
  OAI211_X1 U7443 ( .C1(n6446), .C2(n6445), .A(n6444), .B(n6443), .ZN(U2984)
         );
  OR2_X1 U7444 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  AOI22_X1 U7445 ( .A1(n6451), .A2(n6450), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6449), .ZN(n6453) );
  OAI211_X1 U7446 ( .C1(n6455), .C2(n6454), .A(n6453), .B(n6452), .ZN(U2986)
         );
  AOI21_X1 U7447 ( .B1(n6457), .B2(n6499), .A(n6456), .ZN(n6461) );
  AOI22_X1 U7448 ( .A1(n6502), .A2(n6459), .B1(n6462), .B2(n6458), .ZN(n6460)
         );
  OAI211_X1 U7449 ( .C1(n6463), .C2(n6462), .A(n6461), .B(n6460), .ZN(U3007)
         );
  INV_X1 U7450 ( .A(n6464), .ZN(n6466) );
  AOI21_X1 U7451 ( .B1(n6466), .B2(n6499), .A(n6465), .ZN(n6470) );
  AOI22_X1 U7452 ( .A1(n6468), .A2(n6502), .B1(n6467), .B2(n6471), .ZN(n6469)
         );
  OAI211_X1 U7453 ( .C1(n6472), .C2(n6471), .A(n6470), .B(n6469), .ZN(U3009)
         );
  AOI21_X1 U7454 ( .B1(n6474), .B2(n6499), .A(n6473), .ZN(n6475) );
  OAI21_X1 U7455 ( .B1(n6476), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6475), 
        .ZN(n6477) );
  AOI21_X1 U7456 ( .B1(n6478), .B2(n6502), .A(n6477), .ZN(n6479) );
  OAI21_X1 U7457 ( .B1(n6481), .B2(n6480), .A(n6479), .ZN(U3011) );
  OAI21_X1 U7458 ( .B1(n6483), .B2(n4284), .A(n6482), .ZN(n6485) );
  AOI22_X1 U7459 ( .A1(n6486), .A2(n6485), .B1(n6499), .B2(n6484), .ZN(n6493)
         );
  AOI22_X1 U7460 ( .A1(n6488), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6502), 
        .B2(n6487), .ZN(n6492) );
  NAND2_X1 U7461 ( .A1(n6503), .A2(REIP_REG_2__SCAN_IN), .ZN(n6491) );
  NAND3_X1 U7462 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6489), .A3(n4284), 
        .ZN(n6490) );
  NAND4_X1 U7463 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(U3016)
         );
  NAND2_X1 U7464 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  NAND2_X1 U7465 ( .A1(n6497), .A2(n6496), .ZN(n6506) );
  INV_X1 U7466 ( .A(n6498), .ZN(n6501) );
  AOI222_X1 U7467 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6503), .B1(n6502), .B2(
        n6501), .C1(n6500), .C2(n6499), .ZN(n6504) );
  OAI221_X1 U7468 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6506), .C1(n4281), .C2(n6505), .A(n6504), .ZN(U3017) );
  AND2_X1 U7469 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6507), .ZN(U3019)
         );
  NAND2_X1 U7470 ( .A1(n6606), .A2(n6508), .ZN(n6522) );
  INV_X1 U7471 ( .A(n6522), .ZN(n6560) );
  INV_X1 U7472 ( .A(n6509), .ZN(n6513) );
  NAND3_X1 U7473 ( .A1(n6511), .A2(n6510), .A3(n6619), .ZN(n6512) );
  OAI21_X1 U7474 ( .B1(n6513), .B2(n4530), .A(n6512), .ZN(n6558) );
  AOI22_X1 U7475 ( .A1(n6515), .A2(n6560), .B1(n6514), .B2(n6558), .ZN(n6528)
         );
  INV_X1 U7476 ( .A(n6584), .ZN(n6518) );
  NOR3_X1 U7477 ( .A1(n6562), .A2(n6518), .A3(n6517), .ZN(n6521) );
  OAI21_X1 U7478 ( .B1(n6521), .B2(n6520), .A(n6519), .ZN(n6525) );
  AOI21_X1 U7479 ( .B1(n6522), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6523) );
  NAND3_X1 U7480 ( .A1(n6525), .A2(n6524), .A3(n6523), .ZN(n6564) );
  AOI22_X1 U7481 ( .A1(n6564), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6526), 
        .B2(n6562), .ZN(n6527) );
  OAI211_X1 U7482 ( .C1(n6529), .C2(n6584), .A(n6528), .B(n6527), .ZN(U3068)
         );
  AOI22_X1 U7483 ( .A1(n6531), .A2(n6560), .B1(n6530), .B2(n6558), .ZN(n6534)
         );
  AOI22_X1 U7484 ( .A1(n6564), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6532), 
        .B2(n6562), .ZN(n6533) );
  OAI211_X1 U7485 ( .C1(n6535), .C2(n6584), .A(n6534), .B(n6533), .ZN(U3069)
         );
  AOI22_X1 U7486 ( .A1(n6570), .A2(n6560), .B1(n6571), .B2(n6558), .ZN(n6538)
         );
  AOI22_X1 U7487 ( .A1(n6564), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6536), 
        .B2(n6562), .ZN(n6537) );
  OAI211_X1 U7488 ( .C1(n6539), .C2(n6584), .A(n6538), .B(n6537), .ZN(U3070)
         );
  AOI22_X1 U7489 ( .A1(n6587), .A2(n6560), .B1(n6588), .B2(n6558), .ZN(n6542)
         );
  AOI22_X1 U7490 ( .A1(n6564), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6540), 
        .B2(n6562), .ZN(n6541) );
  OAI211_X1 U7491 ( .C1(n6543), .C2(n6584), .A(n6542), .B(n6541), .ZN(U3071)
         );
  AOI22_X1 U7492 ( .A1(n6578), .A2(n6560), .B1(n6580), .B2(n6558), .ZN(n6546)
         );
  AOI22_X1 U7493 ( .A1(n6564), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6544), 
        .B2(n6562), .ZN(n6545) );
  OAI211_X1 U7494 ( .C1(n6547), .C2(n6584), .A(n6546), .B(n6545), .ZN(U3072)
         );
  AOI22_X1 U7495 ( .A1(n6595), .A2(n6560), .B1(n6597), .B2(n6558), .ZN(n6550)
         );
  AOI22_X1 U7496 ( .A1(n6564), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6548), 
        .B2(n6562), .ZN(n6549) );
  OAI211_X1 U7497 ( .C1(n6551), .C2(n6584), .A(n6550), .B(n6549), .ZN(U3073)
         );
  AOI22_X1 U7498 ( .A1(n6553), .A2(n6560), .B1(n6552), .B2(n6558), .ZN(n6556)
         );
  AOI22_X1 U7499 ( .A1(n6564), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6554), 
        .B2(n6562), .ZN(n6555) );
  OAI211_X1 U7500 ( .C1(n6557), .C2(n6584), .A(n6556), .B(n6555), .ZN(U3074)
         );
  AOI22_X1 U7501 ( .A1(n6561), .A2(n6560), .B1(n6559), .B2(n6558), .ZN(n6566)
         );
  AOI22_X1 U7502 ( .A1(n6564), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6563), 
        .B2(n6562), .ZN(n6565) );
  OAI211_X1 U7503 ( .C1(n6567), .C2(n6584), .A(n6566), .B(n6565), .ZN(U3075)
         );
  INV_X1 U7504 ( .A(n6568), .ZN(n6575) );
  AOI22_X1 U7505 ( .A1(n6570), .A2(n6577), .B1(n6569), .B2(n6575), .ZN(n6573)
         );
  AOI22_X1 U7506 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6581), .B1(n6571), 
        .B2(n6579), .ZN(n6572) );
  OAI211_X1 U7507 ( .C1(n6574), .C2(n6584), .A(n6573), .B(n6572), .ZN(U3078)
         );
  AOI22_X1 U7508 ( .A1(n6578), .A2(n6577), .B1(n6576), .B2(n6575), .ZN(n6583)
         );
  AOI22_X1 U7509 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6581), .B1(n6580), 
        .B2(n6579), .ZN(n6582) );
  OAI211_X1 U7510 ( .C1(n6585), .C2(n6584), .A(n6583), .B(n6582), .ZN(U3080)
         );
  AOI22_X1 U7511 ( .A1(n6587), .A2(n6594), .B1(n6593), .B2(n6586), .ZN(n6590)
         );
  AOI22_X1 U7512 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6598), .B1(n6588), 
        .B2(n6596), .ZN(n6589) );
  OAI211_X1 U7513 ( .C1(n6591), .C2(n6601), .A(n6590), .B(n6589), .ZN(U3111)
         );
  AOI22_X1 U7514 ( .A1(n6595), .A2(n6594), .B1(n6593), .B2(n6592), .ZN(n6600)
         );
  AOI22_X1 U7515 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6598), .B1(n6597), 
        .B2(n6596), .ZN(n6599) );
  OAI211_X1 U7516 ( .C1(n6602), .C2(n6601), .A(n6600), .B(n6599), .ZN(U3113)
         );
  INV_X1 U7517 ( .A(n6603), .ZN(n6605) );
  MUX2_X1 U7518 ( .A(n6605), .B(n6604), .S(INSTQUEUERD_ADDR_REG_0__SCAN_IN), 
        .Z(n6607) );
  AOI211_X1 U7519 ( .C1(n6609), .C2(n6608), .A(n6607), .B(n6606), .ZN(n6610)
         );
  NAND2_X1 U7520 ( .A1(n6610), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6614) );
  OAI22_X1 U7521 ( .A1(n6612), .A2(n6611), .B1(n6610), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U7522 ( .A1(n6614), .A2(n6613), .ZN(n6616) );
  AOI222_X1 U7523 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6616), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6615), .C1(n6616), .C2(n6615), 
        .ZN(n6617) );
  AOI222_X1 U7524 ( .A1(n6619), .A2(n6618), .B1(n6619), .B2(n6617), .C1(n6618), 
        .C2(n6617), .ZN(n6620) );
  OR2_X1 U7525 ( .A1(n6620), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6628)
         );
  NOR2_X1 U7526 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6624) );
  OAI211_X1 U7527 ( .C1(n6624), .C2(n6623), .A(n6622), .B(n6621), .ZN(n6625)
         );
  NOR2_X1 U7528 ( .A1(n6626), .A2(n6625), .ZN(n6627) );
  NAND2_X1 U7529 ( .A1(n6643), .A2(n6645), .ZN(n6630) );
  NAND2_X1 U7530 ( .A1(READY_N), .A2(n6719), .ZN(n6629) );
  NAND2_X1 U7531 ( .A1(n6630), .A2(n6629), .ZN(n6634) );
  OR2_X1 U7532 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  AOI21_X1 U7533 ( .B1(n6635), .B2(n6723), .A(n6651), .ZN(n6636) );
  INV_X1 U7534 ( .A(n6636), .ZN(n6639) );
  OAI21_X1 U7535 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6828), .A(n6708), .ZN(
        n6647) );
  NOR2_X1 U7536 ( .A1(n6637), .A2(n6647), .ZN(n6638) );
  MUX2_X1 U7537 ( .A(n6639), .B(n6638), .S(STATE2_REG_0__SCAN_IN), .Z(n6641)
         );
  OAI211_X1 U7538 ( .C1(n6643), .C2(n6642), .A(n6641), .B(n6640), .ZN(U3148)
         );
  INV_X1 U7539 ( .A(n6644), .ZN(n6646) );
  AOI21_X1 U7540 ( .B1(n6646), .B2(n6828), .A(n6645), .ZN(n6650) );
  OAI211_X1 U7541 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6647), .ZN(n6648) );
  OAI211_X1 U7542 ( .C1(n6651), .C2(n6650), .A(n6649), .B(n6648), .ZN(U3149)
         );
  OAI221_X1 U7543 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6828), .A(n6706), .ZN(n6653) );
  OAI21_X1 U7544 ( .B1(n6723), .B2(n6653), .A(n6652), .ZN(U3150) );
  AND2_X1 U7545 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6654), .ZN(U3151) );
  AND2_X1 U7546 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6654), .ZN(U3152) );
  AND2_X1 U7547 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6654), .ZN(U3153) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6654), .ZN(U3154) );
  AND2_X1 U7549 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6654), .ZN(U3155) );
  AND2_X1 U7550 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6654), .ZN(U3156) );
  AND2_X1 U7551 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6654), .ZN(U3157) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6654), .ZN(U3158) );
  AND2_X1 U7553 ( .A1(n6654), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  INV_X1 U7554 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6826) );
  NOR2_X1 U7555 ( .A1(n6705), .A2(n6826), .ZN(U3160) );
  AND2_X1 U7556 ( .A1(n6654), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  NOR2_X1 U7557 ( .A1(n6705), .A2(n6843), .ZN(U3162) );
  INV_X1 U7558 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6972) );
  NOR2_X1 U7559 ( .A1(n6705), .A2(n6972), .ZN(U3163) );
  INV_X1 U7560 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6967) );
  NOR2_X1 U7561 ( .A1(n6705), .A2(n6967), .ZN(U3164) );
  AND2_X1 U7562 ( .A1(n6654), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  INV_X1 U7563 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U7564 ( .A1(n6705), .A2(n7047), .ZN(U3166) );
  INV_X1 U7565 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6978) );
  NOR2_X1 U7566 ( .A1(n6705), .A2(n6978), .ZN(U3167) );
  AND2_X1 U7567 ( .A1(n6654), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  INV_X1 U7568 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U7569 ( .A1(n6705), .A2(n6980), .ZN(U3169) );
  INV_X1 U7570 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7073) );
  NOR2_X1 U7571 ( .A1(n6705), .A2(n7073), .ZN(U3170) );
  AND2_X1 U7572 ( .A1(n6654), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  INV_X1 U7573 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U7574 ( .A1(n6705), .A2(n6894), .ZN(U3172) );
  INV_X1 U7575 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6819) );
  NOR2_X1 U7576 ( .A1(n6705), .A2(n6819), .ZN(U3173) );
  NOR2_X1 U7577 ( .A1(n6705), .A2(n6815), .ZN(U3174) );
  INV_X1 U7578 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6900) );
  NOR2_X1 U7579 ( .A1(n6705), .A2(n6900), .ZN(U3175) );
  INV_X1 U7580 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7051) );
  NOR2_X1 U7581 ( .A1(n6705), .A2(n7051), .ZN(U3176) );
  INV_X1 U7582 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U7583 ( .A1(n6705), .A2(n6875), .ZN(U3177) );
  INV_X1 U7584 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6799) );
  NOR2_X1 U7585 ( .A1(n6705), .A2(n6799), .ZN(U3178) );
  AND2_X1 U7586 ( .A1(n6654), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7587 ( .A1(n6654), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  AOI22_X1 U7588 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6670) );
  INV_X1 U7589 ( .A(HOLD), .ZN(n6988) );
  NOR2_X1 U7590 ( .A1(n6662), .A2(n6988), .ZN(n6658) );
  INV_X1 U7591 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7061) );
  OAI21_X1 U7592 ( .B1(n6658), .B2(n7061), .A(n7121), .ZN(n6655) );
  INV_X1 U7593 ( .A(n6656), .ZN(n6669) );
  OAI211_X1 U7594 ( .C1(NA_N), .C2(n6671), .A(n4234), .B(n6669), .ZN(n6665) );
  OAI211_X1 U7595 ( .C1(n6656), .C2(n6670), .A(n6655), .B(n6665), .ZN(U3181)
         );
  NOR2_X1 U7596 ( .A1(n4234), .A2(n7061), .ZN(n6661) );
  NAND2_X1 U7597 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6657) );
  OAI21_X1 U7598 ( .B1(n6661), .B2(n6658), .A(n6657), .ZN(n6659) );
  OAI211_X1 U7599 ( .C1(n6662), .C2(n6828), .A(n6660), .B(n6659), .ZN(U3182)
         );
  INV_X1 U7600 ( .A(NA_N), .ZN(n6996) );
  NAND4_X1 U7601 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .A3(n6661), .A4(
        n6996), .ZN(n6668) );
  NOR2_X1 U7602 ( .A1(NA_N), .A2(n6828), .ZN(n6663) );
  OAI21_X1 U7603 ( .B1(n6663), .B2(n6662), .A(n7061), .ZN(n6664) );
  AOI21_X1 U7604 ( .B1(n6671), .B2(n6664), .A(n6988), .ZN(n6666) );
  OAI21_X1 U7605 ( .B1(n4234), .B2(n6666), .A(n6665), .ZN(n6667) );
  OAI211_X1 U7606 ( .C1(n6670), .C2(n6669), .A(n6668), .B(n6667), .ZN(U3183)
         );
  INV_X1 U7607 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6966) );
  OAI222_X1 U7608 ( .A1(n6691), .A2(n6288), .B1(n6966), .B2(n6716), .C1(n5196), 
        .C2(n6701), .ZN(U3184) );
  INV_X1 U7609 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6672) );
  OAI222_X1 U7610 ( .A1(n6701), .A2(n6288), .B1(n6672), .B2(n6716), .C1(n6673), 
        .C2(n6691), .ZN(U3185) );
  INV_X1 U7611 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7041) );
  OAI222_X1 U7612 ( .A1(n6701), .A2(n6673), .B1(n7041), .B2(n6716), .C1(n6674), 
        .C2(n6691), .ZN(U3186) );
  INV_X1 U7613 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6862) );
  OAI222_X1 U7614 ( .A1(n6701), .A2(n6674), .B1(n6862), .B2(n6716), .C1(n6676), 
        .C2(n6691), .ZN(U3187) );
  INV_X1 U7615 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6675) );
  OAI222_X1 U7616 ( .A1(n6701), .A2(n6676), .B1(n6675), .B2(n6716), .C1(n6678), 
        .C2(n6691), .ZN(U3188) );
  INV_X1 U7617 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6677) );
  OAI222_X1 U7618 ( .A1(n6701), .A2(n6678), .B1(n6677), .B2(n6716), .C1(n6680), 
        .C2(n6691), .ZN(U3189) );
  INV_X1 U7619 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6679) );
  OAI222_X1 U7620 ( .A1(n6701), .A2(n6680), .B1(n6679), .B2(n6716), .C1(n6681), 
        .C2(n6691), .ZN(U3190) );
  INV_X1 U7621 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7058) );
  OAI222_X1 U7622 ( .A1(n6691), .A2(n5322), .B1(n7058), .B2(n6716), .C1(n6681), 
        .C2(n6701), .ZN(U3191) );
  INV_X1 U7623 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7082) );
  OAI222_X1 U7624 ( .A1(n6701), .A2(n5322), .B1(n7082), .B2(n6716), .C1(n6682), 
        .C2(n6691), .ZN(U3192) );
  INV_X1 U7625 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7050) );
  OAI222_X1 U7626 ( .A1(n6701), .A2(n6682), .B1(n7050), .B2(n6716), .C1(n6684), 
        .C2(n6691), .ZN(U3193) );
  INV_X1 U7627 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6683) );
  OAI222_X1 U7628 ( .A1(n6701), .A2(n6684), .B1(n6683), .B2(n6716), .C1(n5754), 
        .C2(n6691), .ZN(U3194) );
  INV_X1 U7629 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6868) );
  OAI222_X1 U7630 ( .A1(n6701), .A2(n5754), .B1(n6868), .B2(n6716), .C1(n6685), 
        .C2(n6691), .ZN(U3195) );
  INV_X1 U7631 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7083) );
  OAI222_X1 U7632 ( .A1(n6701), .A2(n6685), .B1(n7083), .B2(n6716), .C1(n6686), 
        .C2(n6691), .ZN(U3196) );
  INV_X1 U7633 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U7634 ( .A1(n6691), .A2(n6689), .B1(n6687), .B2(n6716), .C1(n6686), 
        .C2(n6701), .ZN(U3197) );
  INV_X1 U7635 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6688) );
  INV_X1 U7636 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6871) );
  OAI222_X1 U7637 ( .A1(n6701), .A2(n6689), .B1(n6688), .B2(n6716), .C1(n6871), 
        .C2(n6691), .ZN(U3198) );
  INV_X1 U7638 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6895) );
  OAI222_X1 U7639 ( .A1(n6701), .A2(n6871), .B1(n6895), .B2(n6716), .C1(n6845), 
        .C2(n6691), .ZN(U3199) );
  INV_X1 U7640 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6690) );
  OAI222_X1 U7641 ( .A1(n6691), .A2(n6882), .B1(n6690), .B2(n6716), .C1(n6845), 
        .C2(n6701), .ZN(U3200) );
  INV_X1 U7642 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7076) );
  OAI222_X1 U7643 ( .A1(n6691), .A2(n6692), .B1(n7076), .B2(n6716), .C1(n6882), 
        .C2(n6701), .ZN(U3201) );
  INV_X1 U7644 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6992) );
  INV_X1 U7645 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7048) );
  OAI222_X1 U7646 ( .A1(n6701), .A2(n6692), .B1(n6992), .B2(n6716), .C1(n7048), 
        .C2(n6691), .ZN(U3202) );
  INV_X1 U7647 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6801) );
  OAI222_X1 U7648 ( .A1(n6701), .A2(n7048), .B1(n6801), .B2(n6716), .C1(n6902), 
        .C2(n6691), .ZN(U3203) );
  INV_X1 U7649 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U7650 ( .A1(n6701), .A2(n6902), .B1(n6831), .B2(n6716), .C1(n7093), 
        .C2(n6691), .ZN(U3204) );
  INV_X1 U7651 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6888) );
  OAI222_X1 U7652 ( .A1(n6701), .A2(n7093), .B1(n6888), .B2(n6716), .C1(n5683), 
        .C2(n6691), .ZN(U3205) );
  INV_X1 U7653 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6897) );
  OAI222_X1 U7654 ( .A1(n6701), .A2(n5683), .B1(n6897), .B2(n6716), .C1(n6693), 
        .C2(n6691), .ZN(U3206) );
  INV_X1 U7655 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6694) );
  OAI222_X1 U7656 ( .A1(n6691), .A2(n6696), .B1(n6694), .B2(n6716), .C1(n6693), 
        .C2(n6701), .ZN(U3207) );
  INV_X1 U7657 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U7658 ( .A1(n6701), .A2(n6696), .B1(n6695), .B2(n6716), .C1(n6698), 
        .C2(n6691), .ZN(U3208) );
  INV_X1 U7659 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6697) );
  OAI222_X1 U7660 ( .A1(n6701), .A2(n6698), .B1(n6697), .B2(n6716), .C1(n6699), 
        .C2(n6691), .ZN(U3209) );
  INV_X1 U7661 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6961) );
  OAI222_X1 U7662 ( .A1(n6701), .A2(n6699), .B1(n6961), .B2(n6716), .C1(n6960), 
        .C2(n6691), .ZN(U3210) );
  INV_X1 U7663 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6700) );
  OAI222_X1 U7664 ( .A1(n6701), .A2(n6960), .B1(n6700), .B2(n6716), .C1(n6702), 
        .C2(n6691), .ZN(U3211) );
  INV_X1 U7665 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6807) );
  OAI222_X1 U7666 ( .A1(n6701), .A2(n6702), .B1(n6807), .B2(n6716), .C1(n6814), 
        .C2(n6691), .ZN(U3212) );
  INV_X1 U7667 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7044) );
  OAI222_X1 U7668 ( .A1(n6691), .A2(n7057), .B1(n7044), .B2(n6716), .C1(n6814), 
        .C2(n6701), .ZN(U3213) );
  INV_X1 U7669 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6839) );
  INV_X1 U7670 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7060) );
  AOI22_X1 U7671 ( .A1(n6716), .A2(n6839), .B1(n7060), .B2(n7121), .ZN(U3446)
         );
  INV_X1 U7672 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U7673 ( .A1(n6716), .A2(n7064), .B1(n6987), .B2(n7121), .ZN(U3447)
         );
  INV_X1 U7674 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6869) );
  INV_X1 U7675 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6899) );
  AOI22_X1 U7676 ( .A1(n6716), .A2(n6869), .B1(n6899), .B2(n7121), .ZN(U3448)
         );
  OAI21_X1 U7677 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6705), .A(n6704), .ZN(
        n6703) );
  INV_X1 U7678 ( .A(n6703), .ZN(U3451) );
  INV_X1 U7679 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7116) );
  OAI21_X1 U7680 ( .B1(n6705), .B2(n7116), .A(n6704), .ZN(U3452) );
  OAI211_X1 U7681 ( .C1(n5471), .C2(n6708), .A(n6707), .B(n6706), .ZN(U3453)
         );
  NAND2_X1 U7682 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6712) );
  AOI211_X1 U7683 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(n6714), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6709) );
  AOI21_X1 U7684 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6711), .A(n6709), .ZN(
        n6710) );
  OAI21_X1 U7685 ( .B1(n6712), .B2(n6711), .A(n6710), .ZN(U3468) );
  OAI22_X1 U7686 ( .A1(n6714), .A2(REIP_REG_0__SCAN_IN), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(n6713), .ZN(n6715) );
  INV_X1 U7687 ( .A(n6715), .ZN(U3469) );
  INV_X1 U7688 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7045) );
  AOI22_X1 U7689 ( .A1(n6716), .A2(READREQUEST_REG_SCAN_IN), .B1(n7045), .B2(
        n7121), .ZN(U3470) );
  AOI211_X1 U7690 ( .C1(n6719), .C2(n6828), .A(n6718), .B(n6717), .ZN(n6726)
         );
  OAI21_X1 U7691 ( .B1(n6720), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6722) );
  OAI21_X1 U7692 ( .B1(n6722), .B2(n6721), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6725) );
  NOR2_X1 U7693 ( .A1(n6726), .A2(n6723), .ZN(n6724) );
  AOI22_X1 U7694 ( .A1(n7061), .A2(n6726), .B1(n6725), .B2(n6724), .ZN(U3472)
         );
  INV_X1 U7695 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6977) );
  AOI22_X1 U7696 ( .A1(n6716), .A2(n6884), .B1(n6977), .B2(n7121), .ZN(U3473)
         );
  OAI22_X1 U7697 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_g54), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput_g77), .ZN(n6727) );
  AOI221_X1 U7698 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .C1(
        keyinput_g77), .C2(ADDRESS_REG_23__SCAN_IN), .A(n6727), .ZN(n6734) );
  OAI22_X1 U7699 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_g53), .B1(
        keyinput_g1), .B2(DATAI_30_), .ZN(n6728) );
  AOI221_X1 U7700 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_g53), .C1(
        DATAI_30_), .C2(keyinput_g1), .A(n6728), .ZN(n6733) );
  OAI22_X1 U7701 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_g101), .B1(
        keyinput_g28), .B2(DATAI_3_), .ZN(n6729) );
  AOI221_X1 U7702 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_g101), .C1(
        DATAI_3_), .C2(keyinput_g28), .A(n6729), .ZN(n6732) );
  OAI22_X1 U7703 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(keyinput_g118), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(keyinput_g73), .ZN(n6730) );
  AOI221_X1 U7704 ( .B1(DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput_g118), .C1(
        keyinput_g73), .C2(ADDRESS_REG_27__SCAN_IN), .A(n6730), .ZN(n6731) );
  NAND4_X1 U7705 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n6762)
         );
  OAI22_X1 U7706 ( .A1(ADDRESS_REG_5__SCAN_IN), .A2(keyinput_g95), .B1(
        keyinput_g87), .B2(ADDRESS_REG_13__SCAN_IN), .ZN(n6735) );
  AOI221_X1 U7707 ( .B1(ADDRESS_REG_5__SCAN_IN), .B2(keyinput_g95), .C1(
        ADDRESS_REG_13__SCAN_IN), .C2(keyinput_g87), .A(n6735), .ZN(n6742) );
  OAI22_X1 U7708 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput_g102), .B1(
        keyinput_g120), .B2(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6736) );
  AOI221_X1 U7709 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput_g102), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput_g120), .A(n6736), .ZN(n6741)
         );
  OAI22_X1 U7710 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput_g117), .B1(
        keyinput_g46), .B2(W_R_N_REG_SCAN_IN), .ZN(n6737) );
  AOI221_X1 U7711 ( .B1(DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_g117), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_g46), .A(n6737), .ZN(n6740) );
  OAI22_X1 U7712 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_g121), .ZN(n6738) );
  AOI221_X1 U7713 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(keyinput_g121), .C2(
        DATAWIDTH_REG_17__SCAN_IN), .A(n6738), .ZN(n6739) );
  NAND4_X1 U7714 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6761)
         );
  OAI22_X1 U7715 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(keyinput_g104), .B2(
        DATAWIDTH_REG_0__SCAN_IN), .ZN(n6743) );
  AOI221_X1 U7716 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput_g104), .A(n6743), .ZN(n6750)
         );
  OAI22_X1 U7717 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput_g94), .B1(
        keyinput_g34), .B2(BS16_N), .ZN(n6744) );
  AOI221_X1 U7718 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput_g94), .C1(BS16_N), .C2(keyinput_g34), .A(n6744), .ZN(n6749) );
  OAI22_X1 U7719 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g99), .B2(ADDRESS_REG_1__SCAN_IN), .ZN(n6745) );
  AOI221_X1 U7720 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .C1(
        ADDRESS_REG_1__SCAN_IN), .C2(keyinput_g99), .A(n6745), .ZN(n6748) );
  OAI22_X1 U7721 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_g63), .B1(
        keyinput_g107), .B2(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6746) );
  AOI221_X1 U7722 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .C1(
        DATAWIDTH_REG_3__SCAN_IN), .C2(keyinput_g107), .A(n6746), .ZN(n6747)
         );
  NAND4_X1 U7723 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6760)
         );
  OAI22_X1 U7724 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        keyinput_g88), .B2(ADDRESS_REG_12__SCAN_IN), .ZN(n6751) );
  AOI221_X1 U7725 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        ADDRESS_REG_12__SCAN_IN), .C2(keyinput_g88), .A(n6751), .ZN(n6758) );
  OAI22_X1 U7726 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(keyinput_g106), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput_g93), .ZN(n6752) );
  AOI221_X1 U7727 ( .B1(DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput_g106), .C1(
        keyinput_g93), .C2(ADDRESS_REG_7__SCAN_IN), .A(n6752), .ZN(n6757) );
  OAI22_X1 U7728 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput_g76), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(keyinput_g92), .ZN(n6753) );
  AOI221_X1 U7729 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput_g76), .C1(
        keyinput_g92), .C2(ADDRESS_REG_8__SCAN_IN), .A(n6753), .ZN(n6756) );
  OAI22_X1 U7730 ( .A1(n7073), .A2(keyinput_g116), .B1(n7051), .B2(
        keyinput_g110), .ZN(n6754) );
  AOI221_X1 U7731 ( .B1(n7073), .B2(keyinput_g116), .C1(keyinput_g110), .C2(
        n7051), .A(n6754), .ZN(n6755) );
  NAND4_X1 U7732 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6759)
         );
  NOR4_X1 U7733 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n7120)
         );
  OAI22_X1 U7734 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(HOLD), .B2(
        keyinput_g36), .ZN(n6763) );
  AOI221_X1 U7735 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(keyinput_g36), .C2(
        HOLD), .A(n6763), .ZN(n6770) );
  OAI22_X1 U7736 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput_g84), .B1(
        keyinput_g41), .B2(D_C_N_REG_SCAN_IN), .ZN(n6764) );
  AOI221_X1 U7737 ( .B1(ADDRESS_REG_16__SCAN_IN), .B2(keyinput_g84), .C1(
        D_C_N_REG_SCAN_IN), .C2(keyinput_g41), .A(n6764), .ZN(n6769) );
  OAI22_X1 U7738 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(keyinput_g86), .B1(
        keyinput_g96), .B2(ADDRESS_REG_4__SCAN_IN), .ZN(n6765) );
  AOI221_X1 U7739 ( .B1(ADDRESS_REG_14__SCAN_IN), .B2(keyinput_g86), .C1(
        ADDRESS_REG_4__SCAN_IN), .C2(keyinput_g96), .A(n6765), .ZN(n6768) );
  OAI22_X1 U7740 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(DATAI_8_), .B2(
        keyinput_g23), .ZN(n6766) );
  AOI221_X1 U7741 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(keyinput_g23), .C2(
        DATAI_8_), .A(n6766), .ZN(n6767) );
  NAND4_X1 U7742 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6914)
         );
  OAI22_X1 U7743 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .ZN(n6771) );
  AOI221_X1 U7744 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(keyinput_g48), .C2(
        BYTEENABLE_REG_1__SCAN_IN), .A(n6771), .ZN(n6797) );
  OAI22_X1 U7745 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(keyinput_g37), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n6772) );
  AOI221_X1 U7746 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(
        READREQUEST_REG_SCAN_IN), .C2(keyinput_g37), .A(n6772), .ZN(n6775) );
  OAI22_X1 U7747 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_g60), .B1(DATAI_19_), .B2(keyinput_g12), .ZN(n6773) );
  AOI221_X1 U7748 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g12), .C2(DATAI_19_), .A(n6773), .ZN(n6774) );
  OAI211_X1 U7749 ( .C1(n6777), .C2(keyinput_g38), .A(n6775), .B(n6774), .ZN(
        n6776) );
  AOI21_X1 U7750 ( .B1(n6777), .B2(keyinput_g38), .A(n6776), .ZN(n6796) );
  AOI22_X1 U7751 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_g75), .B1(
        DATAI_1_), .B2(keyinput_g30), .ZN(n6778) );
  OAI221_X1 U7752 ( .B1(ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .C1(
        DATAI_1_), .C2(keyinput_g30), .A(n6778), .ZN(n6785) );
  AOI22_X1 U7753 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_g55), .ZN(n6779) );
  OAI221_X1 U7754 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6779), .ZN(n6784) );
  AOI22_X1 U7755 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6780) );
  OAI221_X1 U7756 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6780), .ZN(n6783) );
  AOI22_X1 U7757 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(DATAI_21_), .B2(
        keyinput_g10), .ZN(n6781) );
  OAI221_X1 U7758 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(DATAI_21_), .C2(
        keyinput_g10), .A(n6781), .ZN(n6782) );
  NOR4_X1 U7759 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6795)
         );
  AOI22_X1 U7760 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput_g82), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6786) );
  OAI221_X1 U7761 ( .B1(ADDRESS_REG_18__SCAN_IN), .B2(keyinput_g82), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6786), .ZN(n6793) );
  AOI22_X1 U7762 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput_g127), .B1(
        BE_N_REG_3__SCAN_IN), .B2(keyinput_g67), .ZN(n6787) );
  OAI221_X1 U7763 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .C1(
        BE_N_REG_3__SCAN_IN), .C2(keyinput_g67), .A(n6787), .ZN(n6792) );
  AOI22_X1 U7764 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput_g115), .B1(
        DATAI_22_), .B2(keyinput_g9), .ZN(n6788) );
  OAI221_X1 U7765 ( .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput_g115), .C1(
        DATAI_22_), .C2(keyinput_g9), .A(n6788), .ZN(n6791) );
  AOI22_X1 U7766 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(keyinput_g90), .B1(
        DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_g125), .ZN(n6789) );
  OAI221_X1 U7767 ( .B1(ADDRESS_REG_10__SCAN_IN), .B2(keyinput_g90), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput_g125), .A(n6789), .ZN(n6790)
         );
  NOR4_X1 U7768 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6794)
         );
  NAND4_X1 U7769 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6913)
         );
  AOI22_X1 U7770 ( .A1(n4234), .A2(keyinput_g103), .B1(keyinput_g108), .B2(
        n6799), .ZN(n6798) );
  OAI221_X1 U7771 ( .B1(n4234), .B2(keyinput_g103), .C1(n6799), .C2(
        keyinput_g108), .A(n6798), .ZN(n6811) );
  AOI22_X1 U7772 ( .A1(n7050), .A2(keyinput_g91), .B1(n6801), .B2(keyinput_g81), .ZN(n6800) );
  OAI221_X1 U7773 ( .B1(n7050), .B2(keyinput_g91), .C1(n6801), .C2(
        keyinput_g81), .A(n6800), .ZN(n6810) );
  INV_X1 U7774 ( .A(DATAI_24_), .ZN(n6803) );
  AOI22_X1 U7775 ( .A1(n6804), .A2(keyinput_g18), .B1(keyinput_g7), .B2(n6803), 
        .ZN(n6802) );
  OAI221_X1 U7776 ( .B1(n6804), .B2(keyinput_g18), .C1(n6803), .C2(keyinput_g7), .A(n6802), .ZN(n6809) );
  INV_X1 U7777 ( .A(DATAI_26_), .ZN(n6806) );
  AOI22_X1 U7778 ( .A1(n6807), .A2(keyinput_g72), .B1(n6806), .B2(keyinput_g5), 
        .ZN(n6805) );
  OAI221_X1 U7779 ( .B1(n6807), .B2(keyinput_g72), .C1(n6806), .C2(keyinput_g5), .A(n6805), .ZN(n6808) );
  NOR4_X1 U7780 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6853)
         );
  AOI22_X1 U7781 ( .A1(n6981), .A2(keyinput_g24), .B1(keyinput_g40), .B2(n6977), .ZN(n6812) );
  OAI221_X1 U7782 ( .B1(n6981), .B2(keyinput_g24), .C1(n6977), .C2(
        keyinput_g40), .A(n6812), .ZN(n6823) );
  AOI22_X1 U7783 ( .A1(n6815), .A2(keyinput_g112), .B1(n6814), .B2(
        keyinput_g52), .ZN(n6813) );
  OAI221_X1 U7784 ( .B1(n6815), .B2(keyinput_g112), .C1(n6814), .C2(
        keyinput_g52), .A(n6813), .ZN(n6822) );
  INV_X1 U7785 ( .A(DATAI_27_), .ZN(n6817) );
  AOI22_X1 U7786 ( .A1(n7060), .A2(keyinput_g68), .B1(n6817), .B2(keyinput_g4), 
        .ZN(n6816) );
  OAI221_X1 U7787 ( .B1(n7060), .B2(keyinput_g68), .C1(n6817), .C2(keyinput_g4), .A(n6816), .ZN(n6821) );
  AOI22_X1 U7788 ( .A1(n7063), .A2(keyinput_g31), .B1(keyinput_g113), .B2(
        n6819), .ZN(n6818) );
  OAI221_X1 U7789 ( .B1(n7063), .B2(keyinput_g31), .C1(n6819), .C2(
        keyinput_g113), .A(n6818), .ZN(n6820) );
  NOR4_X1 U7790 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6852)
         );
  AOI22_X1 U7791 ( .A1(n6826), .A2(keyinput_g126), .B1(n6825), .B2(
        keyinput_g39), .ZN(n6824) );
  OAI221_X1 U7792 ( .B1(n6826), .B2(keyinput_g126), .C1(n6825), .C2(
        keyinput_g39), .A(n6824), .ZN(n6837) );
  AOI22_X1 U7793 ( .A1(n6829), .A2(keyinput_g26), .B1(n6828), .B2(keyinput_g35), .ZN(n6827) );
  OAI221_X1 U7794 ( .B1(n6829), .B2(keyinput_g26), .C1(n6828), .C2(
        keyinput_g35), .A(n6827), .ZN(n6836) );
  AOI22_X1 U7795 ( .A1(n6831), .A2(keyinput_g80), .B1(keyinput_g74), .B2(n6961), .ZN(n6830) );
  OAI221_X1 U7796 ( .B1(n6831), .B2(keyinput_g80), .C1(n6961), .C2(
        keyinput_g74), .A(n6830), .ZN(n6835) );
  INV_X1 U7797 ( .A(DATAI_29_), .ZN(n6833) );
  AOI22_X1 U7798 ( .A1(n6833), .A2(keyinput_g2), .B1(keyinput_g19), .B2(n7079), 
        .ZN(n6832) );
  OAI221_X1 U7799 ( .B1(n6833), .B2(keyinput_g2), .C1(n7079), .C2(keyinput_g19), .A(n6832), .ZN(n6834) );
  NOR4_X1 U7800 ( .A1(n6837), .A2(n6836), .A3(n6835), .A4(n6834), .ZN(n6851)
         );
  AOI22_X1 U7801 ( .A1(n6996), .A2(keyinput_g33), .B1(n6839), .B2(keyinput_g49), .ZN(n6838) );
  OAI221_X1 U7802 ( .B1(n6996), .B2(keyinput_g33), .C1(n6839), .C2(
        keyinput_g49), .A(n6838), .ZN(n6849) );
  AOI22_X1 U7803 ( .A1(n5683), .A2(keyinput_g59), .B1(keyinput_g25), .B2(n6841), .ZN(n6840) );
  OAI221_X1 U7804 ( .B1(n5683), .B2(keyinput_g59), .C1(n6841), .C2(
        keyinput_g25), .A(n6840), .ZN(n6848) );
  AOI22_X1 U7805 ( .A1(n6972), .A2(keyinput_g123), .B1(n6843), .B2(
        keyinput_g124), .ZN(n6842) );
  OAI221_X1 U7806 ( .B1(n6972), .B2(keyinput_g123), .C1(n6843), .C2(
        keyinput_g124), .A(n6842), .ZN(n6847) );
  AOI22_X1 U7807 ( .A1(n6967), .A2(keyinput_g122), .B1(n6845), .B2(
        keyinput_g65), .ZN(n6844) );
  OAI221_X1 U7808 ( .B1(n6967), .B2(keyinput_g122), .C1(n6845), .C2(
        keyinput_g65), .A(n6844), .ZN(n6846) );
  NOR4_X1 U7809 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6850)
         );
  NAND4_X1 U7810 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6912)
         );
  INV_X1 U7811 ( .A(DATAI_28_), .ZN(n6855) );
  AOI22_X1 U7812 ( .A1(n6856), .A2(keyinput_g20), .B1(n6855), .B2(keyinput_g3), 
        .ZN(n6854) );
  OAI221_X1 U7813 ( .B1(n6856), .B2(keyinput_g20), .C1(n6855), .C2(keyinput_g3), .A(n6854), .ZN(n6866) );
  AOI22_X1 U7814 ( .A1(n6987), .A2(keyinput_g69), .B1(n6858), .B2(keyinput_g45), .ZN(n6857) );
  OAI221_X1 U7815 ( .B1(n6987), .B2(keyinput_g69), .C1(n6858), .C2(
        keyinput_g45), .A(n6857), .ZN(n6865) );
  INV_X1 U7816 ( .A(MORE_REG_SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7817 ( .A1(n6860), .A2(keyinput_g44), .B1(keyinput_g98), .B2(n7041), .ZN(n6859) );
  OAI221_X1 U7818 ( .B1(n6860), .B2(keyinput_g44), .C1(n7041), .C2(
        keyinput_g98), .A(n6859), .ZN(n6864) );
  AOI22_X1 U7819 ( .A1(n6966), .A2(keyinput_g100), .B1(n6862), .B2(
        keyinput_g97), .ZN(n6861) );
  OAI221_X1 U7820 ( .B1(n6966), .B2(keyinput_g100), .C1(n6862), .C2(
        keyinput_g97), .A(n6861), .ZN(n6863) );
  NOR4_X1 U7821 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6910)
         );
  AOI22_X1 U7822 ( .A1(n6869), .A2(keyinput_g47), .B1(n6868), .B2(keyinput_g89), .ZN(n6867) );
  OAI221_X1 U7823 ( .B1(n6869), .B2(keyinput_g47), .C1(n6868), .C2(
        keyinput_g89), .A(n6867), .ZN(n6879) );
  AOI22_X1 U7824 ( .A1(n6871), .A2(keyinput_g66), .B1(keyinput_g71), .B2(n7044), .ZN(n6870) );
  OAI221_X1 U7825 ( .B1(n6871), .B2(keyinput_g66), .C1(n7044), .C2(
        keyinput_g71), .A(n6870), .ZN(n6878) );
  INV_X1 U7826 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U7827 ( .A1(n6873), .A2(keyinput_g50), .B1(keyinput_g83), .B2(n7076), .ZN(n6872) );
  OAI221_X1 U7828 ( .B1(n6873), .B2(keyinput_g50), .C1(n7076), .C2(
        keyinput_g83), .A(n6872), .ZN(n6877) );
  INV_X1 U7829 ( .A(DATAI_18_), .ZN(n7042) );
  AOI22_X1 U7830 ( .A1(n6875), .A2(keyinput_g109), .B1(n7042), .B2(
        keyinput_g13), .ZN(n6874) );
  OAI221_X1 U7831 ( .B1(n6875), .B2(keyinput_g109), .C1(n7042), .C2(
        keyinput_g13), .A(n6874), .ZN(n6876) );
  NOR4_X1 U7832 ( .A1(n6879), .A2(n6878), .A3(n6877), .A4(n6876), .ZN(n6909)
         );
  AOI22_X1 U7833 ( .A1(n7048), .A2(keyinput_g62), .B1(n7057), .B2(keyinput_g51), .ZN(n6880) );
  OAI221_X1 U7834 ( .B1(n7048), .B2(keyinput_g62), .C1(n7057), .C2(
        keyinput_g51), .A(n6880), .ZN(n6892) );
  AOI22_X1 U7835 ( .A1(n6882), .A2(keyinput_g64), .B1(keyinput_g27), .B2(n7090), .ZN(n6881) );
  OAI221_X1 U7836 ( .B1(n6882), .B2(keyinput_g64), .C1(n7090), .C2(
        keyinput_g27), .A(n6881), .ZN(n6891) );
  AOI22_X1 U7837 ( .A1(n6885), .A2(keyinput_g21), .B1(keyinput_g32), .B2(n6884), .ZN(n6883) );
  OAI221_X1 U7838 ( .B1(n6885), .B2(keyinput_g21), .C1(n6884), .C2(
        keyinput_g32), .A(n6883), .ZN(n6890) );
  INV_X1 U7839 ( .A(DATAI_25_), .ZN(n6887) );
  AOI22_X1 U7840 ( .A1(n6888), .A2(keyinput_g79), .B1(n6887), .B2(keyinput_g6), 
        .ZN(n6886) );
  OAI221_X1 U7841 ( .B1(n6888), .B2(keyinput_g79), .C1(n6887), .C2(keyinput_g6), .A(n6886), .ZN(n6889) );
  NOR4_X1 U7842 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6908)
         );
  AOI22_X1 U7843 ( .A1(n6895), .A2(keyinput_g85), .B1(keyinput_g114), .B2(
        n6894), .ZN(n6893) );
  OAI221_X1 U7844 ( .B1(n6895), .B2(keyinput_g85), .C1(n6894), .C2(
        keyinput_g114), .A(n6893), .ZN(n6906) );
  AOI22_X1 U7845 ( .A1(n6978), .A2(keyinput_g119), .B1(n6897), .B2(
        keyinput_g78), .ZN(n6896) );
  OAI221_X1 U7846 ( .B1(n6978), .B2(keyinput_g119), .C1(n6897), .C2(
        keyinput_g78), .A(n6896), .ZN(n6905) );
  AOI22_X1 U7847 ( .A1(n6900), .A2(keyinput_g111), .B1(keyinput_g70), .B2(
        n6899), .ZN(n6898) );
  OAI221_X1 U7848 ( .B1(n6900), .B2(keyinput_g111), .C1(n6899), .C2(
        keyinput_g70), .A(n6898), .ZN(n6904) );
  AOI22_X1 U7849 ( .A1(n7092), .A2(keyinput_g43), .B1(keyinput_g61), .B2(n6902), .ZN(n6901) );
  OAI221_X1 U7850 ( .B1(n7092), .B2(keyinput_g43), .C1(n6902), .C2(
        keyinput_g61), .A(n6901), .ZN(n6903) );
  NOR4_X1 U7851 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n6907)
         );
  NAND4_X1 U7852 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6911)
         );
  NOR4_X1 U7853 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n7119)
         );
  OAI22_X1 U7854 ( .A1(keyinput_f38), .A2(ADS_N_REG_SCAN_IN), .B1(
        keyinput_f114), .B2(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6915) );
  AOI221_X1 U7855 ( .B1(keyinput_f38), .B2(ADS_N_REG_SCAN_IN), .C1(
        DATAWIDTH_REG_10__SCAN_IN), .C2(keyinput_f114), .A(n6915), .ZN(n6922)
         );
  OAI22_X1 U7856 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_f56), .B1(DATAI_5_), 
        .B2(keyinput_f26), .ZN(n6916) );
  AOI221_X1 U7857 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_f56), .C1(
        keyinput_f26), .C2(DATAI_5_), .A(n6916), .ZN(n6921) );
  OAI22_X1 U7858 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(
        DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_f125), .ZN(n6917) );
  AOI221_X1 U7859 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(keyinput_f125), .C2(
        DATAWIDTH_REG_21__SCAN_IN), .A(n6917), .ZN(n6920) );
  OAI22_X1 U7860 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(keyinput_f3), .B2(
        DATAI_28_), .ZN(n6918) );
  AOI221_X1 U7861 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(DATAI_28_), .C2(
        keyinput_f3), .A(n6918), .ZN(n6919) );
  NAND4_X1 U7862 ( .A1(n6922), .A2(n6921), .A3(n6920), .A4(n6919), .ZN(n6950)
         );
  OAI22_X1 U7863 ( .A1(keyinput_f96), .A2(ADDRESS_REG_4__SCAN_IN), .B1(
        keyinput_f121), .B2(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6923) );
  AOI221_X1 U7864 ( .B1(keyinput_f96), .B2(ADDRESS_REG_4__SCAN_IN), .C1(
        DATAWIDTH_REG_17__SCAN_IN), .C2(keyinput_f121), .A(n6923), .ZN(n6930)
         );
  OAI22_X1 U7865 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(keyinput_f95), .ZN(n6924) );
  AOI221_X1 U7866 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        keyinput_f95), .C2(ADDRESS_REG_5__SCAN_IN), .A(n6924), .ZN(n6929) );
  OAI22_X1 U7867 ( .A1(keyinput_f126), .A2(DATAWIDTH_REG_22__SCAN_IN), .B1(
        keyinput_f87), .B2(ADDRESS_REG_13__SCAN_IN), .ZN(n6925) );
  AOI221_X1 U7868 ( .B1(keyinput_f126), .B2(DATAWIDTH_REG_22__SCAN_IN), .C1(
        ADDRESS_REG_13__SCAN_IN), .C2(keyinput_f87), .A(n6925), .ZN(n6928) );
  OAI22_X1 U7869 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_f65), .B1(
        keyinput_f17), .B2(DATAI_14_), .ZN(n6926) );
  AOI221_X1 U7870 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .C1(
        DATAI_14_), .C2(keyinput_f17), .A(n6926), .ZN(n6927) );
  NAND4_X1 U7871 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n6949)
         );
  OAI22_X1 U7872 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(BS16_N), .B2(
        keyinput_f34), .ZN(n6931) );
  AOI221_X1 U7873 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(keyinput_f34), .C2(
        BS16_N), .A(n6931), .ZN(n6938) );
  OAI22_X1 U7874 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f22), .B2(DATAI_9_), .ZN(n6932) );
  AOI221_X1 U7875 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_f101), .C1(
        DATAI_9_), .C2(keyinput_f22), .A(n6932), .ZN(n6937) );
  OAI22_X1 U7876 ( .A1(keyinput_f79), .A2(ADDRESS_REG_21__SCAN_IN), .B1(
        keyinput_f73), .B2(ADDRESS_REG_27__SCAN_IN), .ZN(n6933) );
  AOI221_X1 U7877 ( .B1(keyinput_f79), .B2(ADDRESS_REG_21__SCAN_IN), .C1(
        ADDRESS_REG_27__SCAN_IN), .C2(keyinput_f73), .A(n6933), .ZN(n6936) );
  OAI22_X1 U7878 ( .A1(keyinput_f81), .A2(ADDRESS_REG_19__SCAN_IN), .B1(
        keyinput_f84), .B2(ADDRESS_REG_16__SCAN_IN), .ZN(n6934) );
  AOI221_X1 U7879 ( .B1(keyinput_f81), .B2(ADDRESS_REG_19__SCAN_IN), .C1(
        ADDRESS_REG_16__SCAN_IN), .C2(keyinput_f84), .A(n6934), .ZN(n6935) );
  NAND4_X1 U7880 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n6948)
         );
  OAI22_X1 U7881 ( .A1(keyinput_f77), .A2(ADDRESS_REG_23__SCAN_IN), .B1(
        keyinput_f49), .B2(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6939) );
  AOI221_X1 U7882 ( .B1(keyinput_f77), .B2(ADDRESS_REG_23__SCAN_IN), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_f49), .A(n6939), .ZN(n6946)
         );
  OAI22_X1 U7883 ( .A1(keyinput_f90), .A2(ADDRESS_REG_10__SCAN_IN), .B1(
        keyinput_f112), .B2(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6940) );
  AOI221_X1 U7884 ( .B1(keyinput_f90), .B2(ADDRESS_REG_10__SCAN_IN), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput_f112), .A(n6940), .ZN(n6945)
         );
  OAI22_X1 U7885 ( .A1(keyinput_f76), .A2(ADDRESS_REG_24__SCAN_IN), .B1(
        keyinput_f124), .B2(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6941) );
  AOI221_X1 U7886 ( .B1(keyinput_f76), .B2(ADDRESS_REG_24__SCAN_IN), .C1(
        DATAWIDTH_REG_20__SCAN_IN), .C2(keyinput_f124), .A(n6941), .ZN(n6944)
         );
  OAI22_X1 U7887 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(keyinput_f99), .ZN(n6942) );
  AOI221_X1 U7888 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(keyinput_f99), .C2(
        ADDRESS_REG_1__SCAN_IN), .A(n6942), .ZN(n6943) );
  NAND4_X1 U7889 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(n6947)
         );
  NOR4_X1 U7890 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(n7112)
         );
  AOI22_X1 U7891 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f32), .B1(
        DATAI_11_), .B2(keyinput_f20), .ZN(n6951) );
  OAI221_X1 U7892 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        DATAI_11_), .C2(keyinput_f20), .A(n6951), .ZN(n6958) );
  AOI22_X1 U7893 ( .A1(keyinput_f67), .A2(BE_N_REG_3__SCAN_IN), .B1(DATAI_26_), 
        .B2(keyinput_f5), .ZN(n6952) );
  OAI221_X1 U7894 ( .B1(keyinput_f67), .B2(BE_N_REG_3__SCAN_IN), .C1(DATAI_26_), .C2(keyinput_f5), .A(n6952), .ZN(n6957) );
  AOI22_X1 U7895 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_f66), .B1(
        STATE_REG_1__SCAN_IN), .B2(keyinput_f102), .ZN(n6953) );
  OAI221_X1 U7896 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_f66), .C1(
        STATE_REG_1__SCAN_IN), .C2(keyinput_f102), .A(n6953), .ZN(n6956) );
  AOI22_X1 U7897 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_f44), .B1(
        REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .ZN(n6954) );
  OAI221_X1 U7898 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_f44), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_f57), .A(n6954), .ZN(n6955) );
  NOR4_X1 U7899 ( .A1(n6958), .A2(n6957), .A3(n6956), .A4(n6955), .ZN(n7111)
         );
  AOI22_X1 U7900 ( .A1(n6961), .A2(keyinput_f74), .B1(n6960), .B2(keyinput_f54), .ZN(n6959) );
  OAI221_X1 U7901 ( .B1(n6961), .B2(keyinput_f74), .C1(n6960), .C2(
        keyinput_f54), .A(n6959), .ZN(n7004) );
  OAI22_X1 U7902 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(keyinput_f106), .B2(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6962) );
  AOI221_X1 U7903 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(
        DATAWIDTH_REG_2__SCAN_IN), .C2(keyinput_f106), .A(n6962), .ZN(n6970)
         );
  OAI22_X1 U7904 ( .A1(n6964), .A2(keyinput_f29), .B1(keyinput_f45), .B2(
        FLUSH_REG_SCAN_IN), .ZN(n6963) );
  AOI221_X1 U7905 ( .B1(n6964), .B2(keyinput_f29), .C1(FLUSH_REG_SCAN_IN), 
        .C2(keyinput_f45), .A(n6963), .ZN(n6969) );
  OAI22_X1 U7906 ( .A1(keyinput_f122), .A2(n6967), .B1(n6966), .B2(
        keyinput_f100), .ZN(n6965) );
  AOI221_X1 U7907 ( .B1(n6967), .B2(keyinput_f122), .C1(n6966), .C2(
        keyinput_f100), .A(n6965), .ZN(n6968) );
  NAND3_X1 U7908 ( .A1(n6970), .A2(n6969), .A3(n6968), .ZN(n7003) );
  INV_X1 U7909 ( .A(DATAI_22_), .ZN(n6973) );
  OAI22_X1 U7910 ( .A1(n6973), .A2(keyinput_f9), .B1(n6972), .B2(keyinput_f123), .ZN(n6971) );
  AOI221_X1 U7911 ( .B1(n6973), .B2(keyinput_f9), .C1(keyinput_f123), .C2(
        n6972), .A(n6971), .ZN(n6985) );
  OAI22_X1 U7912 ( .A1(n4234), .A2(keyinput_f103), .B1(n6975), .B2(
        keyinput_f16), .ZN(n6974) );
  AOI221_X1 U7913 ( .B1(n4234), .B2(keyinput_f103), .C1(keyinput_f16), .C2(
        n6975), .A(n6974), .ZN(n6984) );
  OAI22_X1 U7914 ( .A1(keyinput_f119), .A2(n6978), .B1(n6977), .B2(
        keyinput_f40), .ZN(n6976) );
  AOI221_X1 U7915 ( .B1(n6978), .B2(keyinput_f119), .C1(n6977), .C2(
        keyinput_f40), .A(n6976), .ZN(n6983) );
  OAI22_X1 U7916 ( .A1(n6981), .A2(keyinput_f24), .B1(n6980), .B2(
        keyinput_f117), .ZN(n6979) );
  AOI221_X1 U7917 ( .B1(n6981), .B2(keyinput_f24), .C1(keyinput_f117), .C2(
        n6980), .A(n6979), .ZN(n6982) );
  NAND4_X1 U7918 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n7002)
         );
  OAI22_X1 U7919 ( .A1(keyinput_f36), .A2(n6988), .B1(n6987), .B2(keyinput_f69), .ZN(n6986) );
  AOI221_X1 U7920 ( .B1(n6988), .B2(keyinput_f36), .C1(n6987), .C2(
        keyinput_f69), .A(n6986), .ZN(n7000) );
  INV_X1 U7921 ( .A(keyinput_f115), .ZN(n6990) );
  OAI22_X1 U7922 ( .A1(n5683), .A2(keyinput_f59), .B1(n6990), .B2(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n6989) );
  AOI221_X1 U7923 ( .B1(n5683), .B2(keyinput_f59), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(n6990), .A(n6989), .ZN(n6999) );
  INV_X1 U7924 ( .A(DATAI_16_), .ZN(n6993) );
  OAI22_X1 U7925 ( .A1(n6993), .A2(keyinput_f15), .B1(n6992), .B2(keyinput_f82), .ZN(n6991) );
  AOI221_X1 U7926 ( .B1(n6993), .B2(keyinput_f15), .C1(keyinput_f82), .C2(
        n6992), .A(n6991), .ZN(n6998) );
  INV_X1 U7927 ( .A(keyinput_f108), .ZN(n6995) );
  OAI22_X1 U7928 ( .A1(keyinput_f33), .A2(n6996), .B1(n6995), .B2(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n6994) );
  AOI221_X1 U7929 ( .B1(n6996), .B2(keyinput_f33), .C1(n6995), .C2(
        DATAWIDTH_REG_4__SCAN_IN), .A(n6994), .ZN(n6997) );
  NAND4_X1 U7930 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), .ZN(n7001)
         );
  NOR4_X1 U7931 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), .ZN(n7110)
         );
  OAI22_X1 U7932 ( .A1(READY_N), .A2(keyinput_f35), .B1(keyinput_f104), .B2(
        DATAWIDTH_REG_0__SCAN_IN), .ZN(n7005) );
  AOI221_X1 U7933 ( .B1(READY_N), .B2(keyinput_f35), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput_f104), .A(n7005), .ZN(n7012)
         );
  OAI22_X1 U7934 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(keyinput_f113), .B2(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n7006) );
  AOI221_X1 U7935 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_f113), .A(n7006), .ZN(n7011)
         );
  OAI22_X1 U7936 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(
        BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_f50), .ZN(n7007) );
  AOI221_X1 U7937 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(keyinput_f50), .C2(
        BYTEENABLE_REG_3__SCAN_IN), .A(n7007), .ZN(n7010) );
  OAI22_X1 U7938 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(keyinput_f109), .B2(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n7008) );
  AOI221_X1 U7939 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(
        DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput_f109), .A(n7008), .ZN(n7009)
         );
  NAND4_X1 U7940 ( .A1(n7012), .A2(n7011), .A3(n7010), .A4(n7009), .ZN(n7108)
         );
  OAI22_X1 U7941 ( .A1(keyinput_f86), .A2(ADDRESS_REG_14__SCAN_IN), .B1(
        keyinput_f94), .B2(ADDRESS_REG_6__SCAN_IN), .ZN(n7013) );
  AOI221_X1 U7942 ( .B1(keyinput_f86), .B2(ADDRESS_REG_14__SCAN_IN), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput_f94), .A(n7013), .ZN(n7039) );
  INV_X1 U7943 ( .A(DATAI_20_), .ZN(n7019) );
  OAI22_X1 U7944 ( .A1(keyinput_f78), .A2(ADDRESS_REG_22__SCAN_IN), .B1(
        keyinput_f111), .B2(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7014) );
  AOI221_X1 U7945 ( .B1(keyinput_f78), .B2(ADDRESS_REG_22__SCAN_IN), .C1(
        DATAWIDTH_REG_7__SCAN_IN), .C2(keyinput_f111), .A(n7014), .ZN(n7017)
         );
  OAI22_X1 U7946 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(
        keyinput_f55), .B2(REIP_REG_27__SCAN_IN), .ZN(n7015) );
  AOI221_X1 U7947 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        REIP_REG_27__SCAN_IN), .C2(keyinput_f55), .A(n7015), .ZN(n7016) );
  OAI211_X1 U7948 ( .C1(n7019), .C2(keyinput_f11), .A(n7017), .B(n7016), .ZN(
        n7018) );
  AOI21_X1 U7949 ( .B1(n7019), .B2(keyinput_f11), .A(n7018), .ZN(n7038) );
  AOI22_X1 U7950 ( .A1(keyinput_f72), .A2(ADDRESS_REG_28__SCAN_IN), .B1(
        keyinput_f89), .B2(ADDRESS_REG_11__SCAN_IN), .ZN(n7020) );
  OAI221_X1 U7951 ( .B1(keyinput_f72), .B2(ADDRESS_REG_28__SCAN_IN), .C1(
        keyinput_f89), .C2(ADDRESS_REG_11__SCAN_IN), .A(n7020), .ZN(n7027) );
  AOI22_X1 U7952 ( .A1(keyinput_f80), .A2(ADDRESS_REG_20__SCAN_IN), .B1(
        DATAI_1_), .B2(keyinput_f30), .ZN(n7021) );
  OAI221_X1 U7953 ( .B1(keyinput_f80), .B2(ADDRESS_REG_20__SCAN_IN), .C1(
        DATAI_1_), .C2(keyinput_f30), .A(n7021), .ZN(n7026) );
  AOI22_X1 U7954 ( .A1(keyinput_f70), .A2(BE_N_REG_0__SCAN_IN), .B1(
        REIP_REG_18__SCAN_IN), .B2(keyinput_f64), .ZN(n7022) );
  OAI221_X1 U7955 ( .B1(keyinput_f70), .B2(BE_N_REG_0__SCAN_IN), .C1(
        REIP_REG_18__SCAN_IN), .C2(keyinput_f64), .A(n7022), .ZN(n7025) );
  AOI22_X1 U7956 ( .A1(keyinput_f47), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .ZN(n7023) );
  OAI221_X1 U7957 ( .B1(keyinput_f47), .B2(BYTEENABLE_REG_0__SCAN_IN), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_f61), .A(n7023), .ZN(n7024) );
  NOR4_X1 U7958 ( .A1(n7027), .A2(n7026), .A3(n7025), .A4(n7024), .ZN(n7037)
         );
  AOI22_X1 U7959 ( .A1(keyinput_f118), .A2(DATAWIDTH_REG_14__SCAN_IN), .B1(
        keyinput_f75), .B2(ADDRESS_REG_25__SCAN_IN), .ZN(n7028) );
  OAI221_X1 U7960 ( .B1(keyinput_f118), .B2(DATAWIDTH_REG_14__SCAN_IN), .C1(
        keyinput_f75), .C2(ADDRESS_REG_25__SCAN_IN), .A(n7028), .ZN(n7035) );
  AOI22_X1 U7961 ( .A1(keyinput_f97), .A2(ADDRESS_REG_3__SCAN_IN), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput_f63), .ZN(n7029) );
  OAI221_X1 U7962 ( .B1(keyinput_f97), .B2(ADDRESS_REG_3__SCAN_IN), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n7029), .ZN(n7034) );
  AOI22_X1 U7963 ( .A1(keyinput_f85), .A2(ADDRESS_REG_15__SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .ZN(n7030) );
  OAI221_X1 U7964 ( .B1(keyinput_f85), .B2(ADDRESS_REG_15__SCAN_IN), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_f58), .A(n7030), .ZN(n7033) );
  AOI22_X1 U7965 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(REIP_REG_30__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n7031) );
  OAI221_X1 U7966 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(REIP_REG_30__SCAN_IN), .C2(keyinput_f52), .A(n7031), .ZN(n7032) );
  NOR4_X1 U7967 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7036)
         );
  NAND4_X1 U7968 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7107)
         );
  OAI22_X1 U7969 ( .A1(n7042), .A2(keyinput_f13), .B1(n7041), .B2(keyinput_f98), .ZN(n7040) );
  AOI221_X1 U7970 ( .B1(n7042), .B2(keyinput_f13), .C1(keyinput_f98), .C2(
        n7041), .A(n7040), .ZN(n7055) );
  OAI22_X1 U7971 ( .A1(n7045), .A2(keyinput_f46), .B1(n7044), .B2(keyinput_f71), .ZN(n7043) );
  AOI221_X1 U7972 ( .B1(n7045), .B2(keyinput_f46), .C1(keyinput_f71), .C2(
        n7044), .A(n7043), .ZN(n7054) );
  OAI22_X1 U7973 ( .A1(n7048), .A2(keyinput_f62), .B1(n7047), .B2(
        keyinput_f120), .ZN(n7046) );
  AOI221_X1 U7974 ( .B1(n7048), .B2(keyinput_f62), .C1(keyinput_f120), .C2(
        n7047), .A(n7046), .ZN(n7053) );
  OAI22_X1 U7975 ( .A1(keyinput_f110), .A2(n7051), .B1(n7050), .B2(
        keyinput_f91), .ZN(n7049) );
  AOI221_X1 U7976 ( .B1(n7051), .B2(keyinput_f110), .C1(n7050), .C2(
        keyinput_f91), .A(n7049), .ZN(n7052) );
  NAND4_X1 U7977 ( .A1(n7055), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n7106)
         );
  AOI22_X1 U7978 ( .A1(n7058), .A2(keyinput_f93), .B1(n7057), .B2(keyinput_f51), .ZN(n7056) );
  OAI221_X1 U7979 ( .B1(n7058), .B2(keyinput_f93), .C1(n7057), .C2(
        keyinput_f51), .A(n7056), .ZN(n7071) );
  AOI22_X1 U7980 ( .A1(n7061), .A2(keyinput_f42), .B1(keyinput_f68), .B2(n7060), .ZN(n7059) );
  OAI221_X1 U7981 ( .B1(n7061), .B2(keyinput_f42), .C1(n7060), .C2(
        keyinput_f68), .A(n7059), .ZN(n7070) );
  AOI22_X1 U7982 ( .A1(n7064), .A2(keyinput_f48), .B1(n7063), .B2(keyinput_f31), .ZN(n7062) );
  OAI221_X1 U7983 ( .B1(n7064), .B2(keyinput_f48), .C1(n7063), .C2(
        keyinput_f31), .A(n7062), .ZN(n7069) );
  INV_X1 U7984 ( .A(keyinput_f127), .ZN(n7066) );
  AOI22_X1 U7985 ( .A1(n7067), .A2(keyinput_f23), .B1(
        DATAWIDTH_REG_23__SCAN_IN), .B2(n7066), .ZN(n7065) );
  OAI221_X1 U7986 ( .B1(n7067), .B2(keyinput_f23), .C1(n7066), .C2(
        DATAWIDTH_REG_23__SCAN_IN), .A(n7065), .ZN(n7068) );
  NOR4_X1 U7987 ( .A1(n7071), .A2(n7070), .A3(n7069), .A4(n7068), .ZN(n7104)
         );
  INV_X1 U7988 ( .A(DATAI_23_), .ZN(n7074) );
  AOI22_X1 U7989 ( .A1(n7074), .A2(keyinput_f8), .B1(keyinput_f116), .B2(n7073), .ZN(n7072) );
  OAI221_X1 U7990 ( .B1(n7074), .B2(keyinput_f8), .C1(n7073), .C2(
        keyinput_f116), .A(n7072), .ZN(n7087) );
  INV_X1 U7991 ( .A(DATAI_21_), .ZN(n7077) );
  AOI22_X1 U7992 ( .A1(n7077), .A2(keyinput_f10), .B1(keyinput_f83), .B2(n7076), .ZN(n7075) );
  OAI221_X1 U7993 ( .B1(n7077), .B2(keyinput_f10), .C1(n7076), .C2(
        keyinput_f83), .A(n7075), .ZN(n7086) );
  INV_X1 U7994 ( .A(DATAI_19_), .ZN(n7080) );
  AOI22_X1 U7995 ( .A1(n7080), .A2(keyinput_f12), .B1(n7079), .B2(keyinput_f19), .ZN(n7078) );
  OAI221_X1 U7996 ( .B1(n7080), .B2(keyinput_f12), .C1(n7079), .C2(
        keyinput_f19), .A(n7078), .ZN(n7085) );
  AOI22_X1 U7997 ( .A1(n7083), .A2(keyinput_f88), .B1(keyinput_f92), .B2(n7082), .ZN(n7081) );
  OAI221_X1 U7998 ( .B1(n7083), .B2(keyinput_f88), .C1(n7082), .C2(
        keyinput_f92), .A(n7081), .ZN(n7084) );
  NOR4_X1 U7999 ( .A1(n7087), .A2(n7086), .A3(n7085), .A4(n7084), .ZN(n7103)
         );
  OAI22_X1 U8000 ( .A1(n7090), .A2(keyinput_f27), .B1(n7089), .B2(keyinput_f28), .ZN(n7088) );
  AOI221_X1 U8001 ( .B1(n7090), .B2(keyinput_f27), .C1(keyinput_f28), .C2(
        n7089), .A(n7088), .ZN(n7102) );
  XOR2_X1 U8002 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_f41), .Z(n7100) );
  XOR2_X1 U8003 ( .A(keyinput_f107), .B(DATAWIDTH_REG_3__SCAN_IN), .Z(n7099)
         );
  AOI22_X1 U8004 ( .A1(n7093), .A2(keyinput_f60), .B1(n7092), .B2(keyinput_f43), .ZN(n7091) );
  OAI221_X1 U8005 ( .B1(n7093), .B2(keyinput_f60), .C1(n7092), .C2(
        keyinput_f43), .A(n7091), .ZN(n7098) );
  INV_X1 U8006 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7096) );
  INV_X1 U8007 ( .A(DATAI_31_), .ZN(n7095) );
  AOI22_X1 U8008 ( .A1(n7096), .A2(keyinput_f37), .B1(n7095), .B2(keyinput_f0), 
        .ZN(n7094) );
  OAI221_X1 U8009 ( .B1(n7096), .B2(keyinput_f37), .C1(n7095), .C2(keyinput_f0), .A(n7094), .ZN(n7097) );
  NOR4_X1 U8010 ( .A1(n7100), .A2(n7099), .A3(n7098), .A4(n7097), .ZN(n7101)
         );
  NAND4_X1 U8011 ( .A1(n7104), .A2(n7103), .A3(n7102), .A4(n7101), .ZN(n7105)
         );
  NOR4_X1 U8012 ( .A1(n7108), .A2(n7107), .A3(n7106), .A4(n7105), .ZN(n7109)
         );
  NAND4_X1 U8013 ( .A1(n7112), .A2(n7111), .A3(n7110), .A4(n7109), .ZN(n7114)
         );
  AOI21_X1 U8014 ( .B1(keyinput_f105), .B2(n7114), .A(n7116), .ZN(n7117) );
  INV_X1 U8015 ( .A(keyinput_f105), .ZN(n7113) );
  AOI21_X1 U8016 ( .B1(n7114), .B2(n7113), .A(keyinput_g105), .ZN(n7115) );
  AOI22_X1 U8017 ( .A1(keyinput_g105), .A2(n7117), .B1(n7116), .B2(n7115), 
        .ZN(n7118) );
  AOI21_X1 U8018 ( .B1(n7120), .B2(n7119), .A(n7118), .ZN(n7123) );
  AOI22_X1 U8019 ( .A1(n6716), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7121), .ZN(n7122) );
  XNOR2_X1 U8020 ( .A(n7123), .B(n7122), .ZN(U3445) );
  NOR2_X1 U3713 ( .A1(n4449), .A2(n5115), .ZN(n3489) );
  AND2_X1 U3933 ( .A1(n4092), .A2(n4091), .ZN(n5495) );
  OR2_X1 U3642 ( .A1(n3379), .A2(n4043), .ZN(n3356) );
  AND2_X2 U3650 ( .A1(n4528), .A2(n3209), .ZN(n3441) );
  NAND2_X1 U4031 ( .A1(n3402), .A2(n3401), .ZN(n3406) );
  CLKBUF_X1 U4071 ( .A(n3489), .Z(n4036) );
  CLKBUF_X1 U4075 ( .A(n4224), .Z(n5565) );
  AND2_X2 U4183 ( .A1(n4543), .A2(n4546), .ZN(n3316) );
  CLKBUF_X1 U4306 ( .A(n3480), .Z(n6609) );
endmodule

