

module b15_C_gen_AntiSAT_k_128_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2980, n2981, n2982, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794;

  NAND2_X1 U3428 ( .A1(n5609), .A2(n5608), .ZN(n5610) );
  CLKBUF_X1 U3429 ( .A(n4405), .Z(n3002) );
  AND2_X1 U3430 ( .A1(n5459), .A2(n5452), .ZN(n5523) );
  CLKBUF_X2 U3431 ( .A(n3545), .Z(n2990) );
  CLKBUF_X2 U3432 ( .A(n4230), .Z(n2997) );
  OAI211_X1 U3433 ( .C1(n3388), .C2(n3075), .A(n3073), .B(n3072), .ZN(n3429)
         );
  AND2_X1 U3434 ( .A1(n3098), .A2(n4276), .ZN(n3251) );
  CLKBUF_X2 U3435 ( .A(n3316), .Z(n3317) );
  CLKBUF_X1 U3436 ( .A(n3282), .Z(n4087) );
  CLKBUF_X2 U3437 ( .A(n3374), .Z(n3322) );
  BUF_X2 U3438 ( .A(n3276), .Z(n2985) );
  AND2_X1 U3439 ( .A1(n4430), .A2(n4445), .ZN(n3295) );
  CLKBUF_X1 U3440 ( .A(n4039), .Z(n2986) );
  AND2_X2 U3441 ( .A1(n3140), .A2(n3139), .ZN(n3969) );
  AND2_X2 U3442 ( .A1(n3140), .A2(n4404), .ZN(n3374) );
  BUF_X1 U3443 ( .A(n3290), .Z(n2988) );
  AND3_X1 U34450 ( .A1(n4286), .A2(n4272), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3580) );
  NAND2_X1 U34460 ( .A1(n4506), .A2(n4286), .ZN(n4168) );
  BUF_X1 U34470 ( .A(n5505), .Z(n5392) );
  NAND3_X1 U34480 ( .A1(n3018), .A2(n3181), .A3(n3009), .ZN(n4278) );
  NAND2_X1 U3449 ( .A1(n3407), .A2(n3406), .ZN(n4446) );
  NAND2_X1 U3450 ( .A1(n5482), .A2(n5483), .ZN(n5485) );
  OR2_X1 U34510 ( .A1(n5495), .A2(n5496), .ZN(n5498) );
  AND2_X1 U34520 ( .A1(n4384), .A2(n4383), .ZN(n4468) );
  INV_X1 U3454 ( .A(n6138), .ZN(n6201) );
  NAND2_X1 U34550 ( .A1(n4108), .A2(n3124), .ZN(n2980) );
  AND4_X1 U34560 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n2981)
         );
  NAND2_X2 U3457 ( .A1(n5619), .A2(n3539), .ZN(n5829) );
  NAND2_X2 U3458 ( .A1(n5990), .A2(n3130), .ZN(n5619) );
  AND2_X4 U34590 ( .A1(n3036), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3140) );
  NAND2_X4 U34600 ( .A1(n3289), .A2(n3288), .ZN(n3525) );
  NAND2_X2 U34610 ( .A1(n3531), .A2(n3530), .ZN(n5187) );
  AND2_X1 U34620 ( .A1(n3140), .A2(n4404), .ZN(n2982) );
  BUF_X4 U34640 ( .A(n3276), .Z(n2984) );
  BUF_X8 U3466 ( .A(n4039), .Z(n2987) );
  AND2_X2 U3467 ( .A1(n3145), .A2(n4430), .ZN(n4039) );
  BUF_X8 U34680 ( .A(n3290), .Z(n2989) );
  AND2_X2 U34690 ( .A1(n3139), .A2(n3145), .ZN(n3290) );
  AOI211_X1 U34700 ( .C1(n3097), .C2(n5359), .A(n5376), .B(n5370), .ZN(n5360)
         );
  NOR2_X1 U34710 ( .A1(n4525), .A2(n4489), .ZN(n6350) );
  NAND2_X1 U34720 ( .A1(n3055), .A2(n3054), .ZN(n5036) );
  NAND2_X1 U34730 ( .A1(n3097), .A2(n3096), .ZN(n4276) );
  INV_X2 U34740 ( .A(n5505), .ZN(n3097) );
  INV_X2 U3475 ( .A(n4278), .ZN(n3239) );
  CLKBUF_X2 U3476 ( .A(n3969), .Z(n4056) );
  BUF_X2 U3477 ( .A(n4086), .Z(n4034) );
  CLKBUF_X2 U3478 ( .A(n3379), .Z(n4079) );
  BUF_X2 U3479 ( .A(n3295), .Z(n4062) );
  CLKBUF_X2 U3480 ( .A(n3323), .Z(n4080) );
  AOI21_X1 U3481 ( .B1(n5564), .B2(n5563), .A(n5562), .ZN(n5565) );
  OR2_X1 U3482 ( .A1(n5610), .A2(n3090), .ZN(n3088) );
  AOI21_X1 U3483 ( .B1(n5569), .B2(n6266), .A(n5568), .ZN(n5570) );
  OAI21_X1 U3484 ( .B1(n3084), .B2(n3012), .A(n3083), .ZN(n5643) );
  OAI21_X1 U3485 ( .B1(n5408), .B2(n5410), .A(n5409), .ZN(n5583) );
  AOI21_X1 U3486 ( .B1(n5391), .B2(n5409), .A(n5390), .ZN(n5577) );
  OAI21_X1 U3487 ( .B1(n3016), .B2(n3026), .A(n2980), .ZN(n5902) );
  CLKBUF_X1 U3488 ( .A(n5389), .Z(n5409) );
  INV_X1 U3489 ( .A(n5648), .ZN(n5990) );
  OAI21_X1 U3490 ( .B1(n5735), .B2(n6335), .A(n5734), .ZN(n5736) );
  OR2_X1 U3491 ( .A1(n5989), .A2(n5238), .ZN(n5235) );
  INV_X2 U3492 ( .A(n5832), .ZN(n5989) );
  INV_X1 U3493 ( .A(n3545), .ZN(n5832) );
  XNOR2_X1 U3494 ( .A(n3521), .B(n3514), .ZN(n3678) );
  NAND2_X1 U3495 ( .A1(n3521), .A2(n3524), .ZN(n3545) );
  AND2_X1 U3496 ( .A1(n3661), .A2(n3660), .ZN(n4472) );
  NAND2_X1 U3497 ( .A1(n3500), .A2(n3499), .ZN(n3521) );
  NAND2_X1 U3498 ( .A1(n5523), .A2(n5522), .ZN(n6016) );
  OAI21_X1 U3499 ( .B1(n3649), .B2(n3522), .A(n3460), .ZN(n3461) );
  NAND2_X1 U3500 ( .A1(n4247), .A2(n3361), .ZN(n6264) );
  NAND2_X1 U3501 ( .A1(n3449), .A2(n3450), .ZN(n3479) );
  NAND2_X1 U3502 ( .A1(n3430), .A2(n4589), .ZN(n3431) );
  OR2_X1 U3503 ( .A1(n4525), .A2(n4496), .ZN(n6366) );
  XNOR2_X1 U3504 ( .A(n4446), .B(n4786), .ZN(n4429) );
  NAND2_X1 U3505 ( .A1(n3267), .A2(n3266), .ZN(n3268) );
  AND2_X1 U3506 ( .A1(n3345), .A2(n3346), .ZN(n3020) );
  AND2_X1 U3507 ( .A1(n3061), .A2(n3057), .ZN(n4384) );
  NAND4_X1 U3508 ( .A1(n3246), .A2(n3259), .A3(n4253), .A4(n3251), .ZN(n3103)
         );
  NAND2_X1 U3509 ( .A1(n3233), .A2(n4489), .ZN(n3259) );
  AND2_X1 U3510 ( .A1(n3236), .A2(n3235), .ZN(n3249) );
  AND2_X1 U3511 ( .A1(n3338), .A2(n3337), .ZN(n4417) );
  CLKBUF_X1 U3512 ( .A(n4230), .Z(n2996) );
  AND2_X1 U3513 ( .A1(n3242), .A2(n4305), .ZN(n3337) );
  NAND2_X1 U3514 ( .A1(n3253), .A2(n2993), .ZN(n5505) );
  OR2_X1 U3515 ( .A1(n3301), .A2(n3300), .ZN(n3353) );
  NOR2_X1 U3516 ( .A1(n4278), .A2(n3253), .ZN(n4304) );
  NAND2_X2 U3517 ( .A1(n3015), .A2(n2981), .ZN(n3253) );
  NAND2_X1 U3518 ( .A1(n3237), .A2(n3252), .ZN(n4305) );
  AND4_X2 U3519 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3260)
         );
  NAND2_X1 U3520 ( .A1(n3203), .A2(n3202), .ZN(n3553) );
  NAND2_X2 U3521 ( .A1(n3163), .A2(n3162), .ZN(n3252) );
  NAND2_X2 U3522 ( .A1(n3190), .A2(n3014), .ZN(n3622) );
  AND4_X1 U3523 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3162)
         );
  AND4_X1 U3524 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3150)
         );
  AND4_X1 U3525 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3202)
         );
  AND4_X1 U3526 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), .ZN(n3190)
         );
  AND4_X1 U3527 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3230)
         );
  AND4_X1 U3528 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3163)
         );
  AND4_X1 U3529 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3203)
         );
  AND4_X1 U3530 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), .ZN(n3014)
         );
  AND2_X1 U3531 ( .A1(n3037), .A2(n3035), .ZN(n3195) );
  AND4_X1 U3532 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3153)
         );
  NOR2_X1 U3533 ( .A1(n3128), .A2(n3129), .ZN(n3201) );
  AND4_X1 U3534 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3229)
         );
  AND4_X1 U3535 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3232)
         );
  AND4_X1 U3536 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3231)
         );
  AND4_X1 U3537 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3152)
         );
  AND4_X1 U3538 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3151)
         );
  NAND2_X1 U3539 ( .A1(n4103), .A2(n5872), .ZN(n6281) );
  AND2_X2 U3541 ( .A1(n3140), .A2(n4435), .ZN(n3316) );
  AND2_X2 U3542 ( .A1(n3139), .A2(n4445), .ZN(n4086) );
  AND2_X2 U3543 ( .A1(n3038), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4435)
         );
  AND2_X2 U3544 ( .A1(n4430), .A2(n4409), .ZN(n3271) );
  AND2_X2 U3545 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4409) );
  INV_X1 U3546 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3038) );
  NAND2_X2 U3548 ( .A1(n3264), .A2(n3265), .ZN(n3362) );
  INV_X2 U3549 ( .A(n2993), .ZN(n4496) );
  CLKBUF_X1 U3551 ( .A(n5187), .Z(n2992) );
  OR2_X4 U3552 ( .A1(n2994), .A2(n2995), .ZN(n2993) );
  NAND4_X1 U3553 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n2994)
         );
  NAND4_X1 U3554 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n2995)
         );
  NAND3_X1 U3555 ( .A1(n4459), .A2(n3076), .A3(n3429), .ZN(n3452) );
  OR2_X2 U3556 ( .A1(n4478), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U3557 ( .A1(n3342), .A2(n4112), .ZN(n6043) );
  NOR2_X2 U3558 ( .A1(n5361), .A2(n5360), .ZN(n5741) );
  AND2_X1 U3559 ( .A1(n3391), .A2(n3392), .ZN(n3081) );
  NOR2_X4 U3560 ( .A1(n3066), .A2(n3030), .ZN(n5411) );
  XNOR2_X1 U3561 ( .A(n3429), .B(n3394), .ZN(n3620) );
  AND2_X2 U3562 ( .A1(n5194), .A2(n5266), .ZN(n5264) );
  NOR2_X2 U3563 ( .A1(n5033), .A2(n3104), .ZN(n5194) );
  NAND2_X1 U3564 ( .A1(n5975), .A2(n3024), .ZN(n5572) );
  NAND2_X1 U3565 ( .A1(n5829), .A2(n3541), .ZN(n3034) );
  OR2_X1 U3566 ( .A1(n5973), .A2(n5580), .ZN(n5589) );
  OR2_X2 U3567 ( .A1(n5610), .A2(n3095), .ZN(n5617) );
  OAI21_X1 U3568 ( .B1(n5673), .B2(n3044), .A(n3042), .ZN(n5664) );
  NAND2_X1 U3569 ( .A1(n4286), .A2(n2993), .ZN(n4230) );
  NAND2_X2 U3570 ( .A1(n5975), .A2(n3544), .ZN(n5600) );
  OR2_X4 U3571 ( .A1(n5973), .A2(n5974), .ZN(n5975) );
  NAND2_X1 U3572 ( .A1(n4168), .A2(n5505), .ZN(n5369) );
  NAND2_X1 U3573 ( .A1(n4307), .A2(n5505), .ZN(n5345) );
  NAND2_X2 U3574 ( .A1(n5681), .A2(n3534), .ZN(n5673) );
  NAND2_X2 U3575 ( .A1(n5683), .A2(n5682), .ZN(n5681) );
  AND2_X2 U3576 ( .A1(n4106), .A2(n3950), .ZN(n4108) );
  NOR2_X2 U3577 ( .A1(n5432), .A2(n3109), .ZN(n4106) );
  AND2_X1 U3578 ( .A1(n3140), .A2(n4430), .ZN(n2999) );
  NAND2_X1 U3579 ( .A1(n3253), .A2(n2993), .ZN(n3000) );
  XNOR2_X1 U3580 ( .A(n3434), .B(n3433), .ZN(n5052) );
  NAND2_X2 U3581 ( .A1(n3362), .A2(n3268), .ZN(n3629) );
  NAND2_X2 U3582 ( .A1(n3452), .A2(n3431), .ZN(n3640) );
  AOI21_X2 U3583 ( .B1(n5233), .B2(n3048), .A(n3045), .ZN(n5687) );
  OAI21_X2 U3584 ( .B1(n5187), .B2(n3021), .A(n3532), .ZN(n5233) );
  BUF_X4 U3585 ( .A(n4457), .Z(n3001) );
  XNOR2_X1 U3586 ( .A(n3352), .B(n3393), .ZN(n4457) );
  AND2_X2 U3587 ( .A1(n3252), .A2(n3622), .ZN(n3339) );
  XNOR2_X1 U3588 ( .A(n3405), .B(n3406), .ZN(n4405) );
  AND2_X1 U3589 ( .A1(n4435), .A2(n4409), .ZN(n3004) );
  AND2_X4 U3590 ( .A1(n4435), .A2(n4409), .ZN(n3005) );
  AND2_X1 U3591 ( .A1(n4435), .A2(n4409), .ZN(n3373) );
  NOR2_X1 U3592 ( .A1(n4525), .A2(n4496), .ZN(n3006) );
  NOR2_X1 U3593 ( .A1(n4525), .A2(n4496), .ZN(n3007) );
  OR2_X1 U3594 ( .A1(n4272), .A2(n3053), .ZN(n3414) );
  OR2_X1 U3595 ( .A1(n6052), .A2(n6498), .ZN(n4264) );
  BUF_X1 U3596 ( .A(n3271), .Z(n4061) );
  NOR2_X1 U3597 ( .A1(n3355), .A2(n3553), .ZN(n3338) );
  NAND2_X1 U3598 ( .A1(n3027), .A2(n5487), .ZN(n3126) );
  AND2_X1 U3599 ( .A1(n3112), .A2(n5637), .ZN(n3111) );
  INV_X1 U3600 ( .A(n3113), .ZN(n3112) );
  NAND2_X1 U3601 ( .A1(n5318), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4073) );
  INV_X1 U3602 ( .A(n3657), .ZN(n4076) );
  NAND2_X1 U3603 ( .A1(n4641), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3760) );
  NOR2_X1 U3604 ( .A1(n3287), .A2(n3286), .ZN(n3288) );
  NOR2_X1 U3605 ( .A1(n3280), .A2(n3279), .ZN(n3289) );
  INV_X1 U3606 ( .A(n3525), .ZN(n3330) );
  INV_X1 U3607 ( .A(n3414), .ZN(n3387) );
  OR2_X1 U3608 ( .A1(n3347), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3348)
         );
  NAND2_X1 U3609 ( .A1(n3051), .A2(n3020), .ZN(n3364) );
  NOR2_X1 U3610 ( .A1(n3334), .A2(n3053), .ZN(n3052) );
  NAND2_X1 U3611 ( .A1(n3080), .A2(n3079), .ZN(n3078) );
  INV_X1 U3612 ( .A(n3392), .ZN(n3079) );
  INV_X1 U3613 ( .A(n3391), .ZN(n3080) );
  INV_X1 U3614 ( .A(n6498), .ZN(n4374) );
  NOR2_X2 U3615 ( .A1(n5389), .A2(n5391), .ZN(n5390) );
  INV_X1 U3616 ( .A(n4264), .ZN(n4232) );
  OR2_X1 U3617 ( .A1(n3608), .A2(n3607), .ZN(n6052) );
  AND2_X1 U3618 ( .A1(n4119), .A2(n3606), .ZN(n3607) );
  AND2_X1 U3619 ( .A1(n3260), .A2(n3622), .ZN(n3242) );
  AND2_X1 U3620 ( .A1(n3475), .A2(n3474), .ZN(n3478) );
  OR2_X1 U3621 ( .A1(n3496), .A2(n3495), .ZN(n3505) );
  OR2_X1 U3622 ( .A1(n3386), .A2(n3385), .ZN(n3395) );
  AOI21_X1 U3623 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6344), .A(n3594), 
        .ZN(n3601) );
  AND2_X1 U3624 ( .A1(n3592), .A2(n3591), .ZN(n3594) );
  NOR2_X1 U3625 ( .A1(n4168), .A2(n3060), .ZN(n3059) );
  NAND2_X1 U3626 ( .A1(n3697), .A2(n3107), .ZN(n3106) );
  INV_X1 U3627 ( .A(n5155), .ZN(n3107) );
  INV_X1 U3628 ( .A(n5034), .ZN(n3679) );
  CLKBUF_X1 U3629 ( .A(n3657), .Z(n4099) );
  NAND2_X1 U3630 ( .A1(n3101), .A2(n3100), .ZN(n4366) );
  NOR2_X1 U3631 ( .A1(n3252), .A2(n4641), .ZN(n3803) );
  OR2_X1 U3632 ( .A1(n5989), .A2(n3538), .ZN(n3539) );
  INV_X1 U3633 ( .A(n3043), .ZN(n3042) );
  OAI21_X1 U3634 ( .B1(n3535), .B2(n3044), .A(n5665), .ZN(n3043) );
  INV_X1 U3635 ( .A(n3536), .ZN(n3044) );
  INV_X1 U3636 ( .A(n3502), .ZN(n3499) );
  AND2_X1 U3637 ( .A1(n3249), .A2(n3611), .ZN(n4268) );
  NOR2_X1 U3638 ( .A1(n3390), .A2(n3017), .ZN(n3074) );
  OR2_X1 U3639 ( .A1(n6590), .A2(n4123), .ZN(n5447) );
  INV_X1 U3640 ( .A(n3760), .ZN(n5309) );
  NOR2_X1 U3641 ( .A1(n5420), .A2(n3126), .ZN(n3125) );
  INV_X1 U3642 ( .A(n3126), .ZN(n3124) );
  AND2_X1 U3643 ( .A1(n3905), .A2(n3904), .ZN(n5637) );
  AND2_X1 U3644 ( .A1(n3806), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3834)
         );
  NAND2_X1 U3645 ( .A1(n3834), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3850)
         );
  NOR2_X1 U3646 ( .A1(n3666), .A2(n5094), .ZN(n3674) );
  NAND2_X1 U3647 ( .A1(n3674), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3673)
         );
  NAND2_X1 U3648 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3642) );
  NOR2_X1 U3649 ( .A1(n5611), .A2(n3094), .ZN(n3092) );
  XNOR2_X1 U3650 ( .A(n3091), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3090)
         );
  NAND2_X1 U3651 ( .A1(n5627), .A2(n5793), .ZN(n3091) );
  OAI22_X1 U3652 ( .A1(n5643), .A2(n5642), .B1(n5606), .B2(n5989), .ZN(n5635)
         );
  XNOR2_X1 U3653 ( .A(n5989), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5665)
         );
  NOR2_X1 U3654 ( .A1(n3068), .A2(n5199), .ZN(n3067) );
  INV_X1 U3655 ( .A(n3069), .ZN(n3068) );
  AND2_X1 U3656 ( .A1(n4408), .A2(n4288), .ZN(n6472) );
  NAND2_X1 U3657 ( .A1(n3620), .A2(n3559), .ZN(n3402) );
  OAI21_X1 U3658 ( .B1(n4264), .B2(n4263), .A(n4262), .ZN(n4291) );
  OAI21_X1 U3659 ( .B1(n3313), .B2(n3312), .A(n3523), .ZN(n3314) );
  OAI211_X1 U3660 ( .C1(n3333), .C2(n3413), .A(n3332), .B(n3331), .ZN(n3392)
         );
  NAND2_X1 U3661 ( .A1(n3365), .A2(n3364), .ZN(n3405) );
  INV_X1 U3662 ( .A(n3620), .ZN(n4696) );
  INV_X1 U3663 ( .A(n4459), .ZN(n4589) );
  OR2_X1 U3664 ( .A1(n4746), .A2(n4964), .ZN(n4825) );
  NAND2_X1 U3665 ( .A1(n4377), .A2(n4376), .ZN(n6225) );
  XNOR2_X1 U3666 ( .A(n4126), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5567)
         );
  NOR2_X1 U3667 ( .A1(n4125), .A2(n4124), .ZN(n4126) );
  OR2_X1 U3668 ( .A1(n6262), .A2(n6275), .ZN(n6271) );
  NAND2_X1 U3669 ( .A1(n4232), .A2(n6476), .ZN(n6060) );
  OR2_X1 U3670 ( .A1(n3473), .A2(n3472), .ZN(n3481) );
  INV_X1 U3671 ( .A(n3478), .ZN(n3476) );
  AND2_X1 U3672 ( .A1(n3498), .A2(n3497), .ZN(n3502) );
  NAND2_X1 U3673 ( .A1(n3278), .A2(n3277), .ZN(n3279) );
  NAND2_X1 U3674 ( .A1(n2984), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3278) );
  AND2_X1 U3675 ( .A1(n3336), .A2(n3335), .ZN(n3346) );
  AOI22_X1 U3676 ( .A1(n2988), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U3677 ( .A1(n3969), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U3678 ( .A1(n3580), .A2(n3559), .ZN(n3600) );
  NAND2_X1 U3679 ( .A1(n4417), .A2(n4286), .ZN(n4110) );
  NAND2_X1 U3680 ( .A1(n3888), .A2(n3114), .ZN(n3113) );
  INV_X1 U3681 ( .A(n5511), .ZN(n3114) );
  NAND2_X1 U3682 ( .A1(n5291), .A2(n3121), .ZN(n3118) );
  NAND2_X1 U3683 ( .A1(n3123), .A2(n3122), .ZN(n3121) );
  INV_X1 U3684 ( .A(n5680), .ZN(n3122) );
  INV_X1 U3685 ( .A(n3774), .ZN(n3123) );
  NOR2_X1 U3686 ( .A1(n3119), .A2(n3117), .ZN(n3116) );
  INV_X1 U3687 ( .A(n5457), .ZN(n3117) );
  NOR2_X1 U3688 ( .A1(n5160), .A2(n3070), .ZN(n3069) );
  INV_X1 U3689 ( .A(n5150), .ZN(n3070) );
  NAND2_X1 U3690 ( .A1(n2990), .A2(n3528), .ZN(n3529) );
  NAND2_X1 U3691 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  NAND2_X1 U3692 ( .A1(n3243), .A2(n4254), .ZN(n3098) );
  OR2_X1 U3693 ( .A1(n4286), .A2(n3053), .ZN(n3413) );
  OR2_X1 U3694 ( .A1(n3329), .A2(n3328), .ZN(n3354) );
  AND2_X1 U3695 ( .A1(n3260), .A2(n4278), .ZN(n3192) );
  OR2_X1 U3696 ( .A1(n3002), .A2(n3350), .ZN(n4994) );
  INV_X1 U3697 ( .A(n3001), .ZN(n4961) );
  OR2_X1 U3698 ( .A1(n3640), .A2(n5877), .ZN(n4606) );
  NAND2_X1 U3699 ( .A1(n3379), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3700 ( .A1(n3316), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3035)
         );
  AOI22_X1 U3701 ( .A1(n3316), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U3702 ( .A1(n3380), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3169) );
  OR2_X1 U3703 ( .A1(n3425), .A2(n3424), .ZN(n3454) );
  AOI21_X1 U3704 ( .B1(n6504), .B2(n4453), .A(n5891), .ZN(n4488) );
  NOR2_X1 U3705 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4488), .ZN(n4916) );
  AND2_X1 U3706 ( .A1(n3002), .A2(n3350), .ZN(n4913) );
  INV_X1 U3707 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6455) );
  INV_X1 U3708 ( .A(n3600), .ZN(n3602) );
  OR2_X1 U3709 ( .A1(n3596), .A2(n3595), .ZN(n4114) );
  NAND2_X1 U3710 ( .A1(n3414), .A2(n3413), .ZN(n3606) );
  NAND2_X1 U3711 ( .A1(n4232), .A2(n6465), .ZN(n4224) );
  AND2_X1 U3712 ( .A1(n4171), .A2(n4170), .ZN(n5270) );
  INV_X1 U3713 ( .A(n6077), .ZN(n6188) );
  AND2_X1 U3714 ( .A1(n5447), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5380) );
  AND2_X1 U3715 ( .A1(n4192), .A2(n4191), .ZN(n5513) );
  NAND2_X1 U3716 ( .A1(n3063), .A2(n3062), .ZN(n5517) );
  INV_X1 U3717 ( .A(n5513), .ZN(n3062) );
  NAND2_X1 U3718 ( .A1(n4360), .A2(n4307), .ZN(n3057) );
  NAND2_X1 U3719 ( .A1(n4144), .A2(n3058), .ZN(n4383) );
  NOR2_X1 U3720 ( .A1(n4264), .A2(n4239), .ZN(n6227) );
  INV_X1 U3721 ( .A(n4110), .ZN(n6465) );
  AOI21_X1 U3722 ( .B1(n4102), .B2(n4101), .A(n4100), .ZN(n5308) );
  AND2_X1 U3723 ( .A1(n5334), .A2(n4099), .ZN(n4100) );
  OR2_X1 U3724 ( .A1(n4050), .A2(n5413), .ZN(n4054) );
  OR2_X1 U3725 ( .A1(n4054), .A2(n5400), .ZN(n4125) );
  AOI21_X1 U3726 ( .B1(n4053), .B2(n4052), .A(n4051), .ZN(n5410) );
  AND2_X1 U3727 ( .A1(n5412), .A2(n4099), .ZN(n4051) );
  AND2_X1 U3728 ( .A1(n4007), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4026)
         );
  OR2_X1 U3729 ( .A1(n5594), .A2(n4076), .ZN(n4030) );
  OR2_X1 U3730 ( .A1(n3963), .A2(n5612), .ZN(n3986) );
  NOR2_X1 U3731 ( .A1(n3986), .A2(n3985), .ZN(n4007) );
  AND2_X1 U3732 ( .A1(n3990), .A2(n3989), .ZN(n5478) );
  OR2_X1 U3733 ( .A1(n5623), .A2(n4076), .ZN(n3948) );
  NOR2_X1 U3734 ( .A1(n3919), .A2(n5631), .ZN(n3946) );
  NAND2_X1 U3735 ( .A1(n3946), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3963)
         );
  NAND2_X1 U3736 ( .A1(n3111), .A2(n3110), .ZN(n3109) );
  INV_X1 U3737 ( .A(n5501), .ZN(n3110) );
  AND2_X1 U3738 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3614), .ZN(n3903)
         );
  INV_X1 U3739 ( .A(n5432), .ZN(n3108) );
  NOR2_X1 U3740 ( .A1(n3850), .A2(n5653), .ZN(n3868) );
  NAND2_X1 U3741 ( .A1(n3868), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3885)
         );
  AND2_X1 U3742 ( .A1(n3836), .A2(n3835), .ZN(n5994) );
  NOR2_X1 U3743 ( .A1(n3790), .A2(n3791), .ZN(n3806) );
  NAND2_X1 U3744 ( .A1(n3785), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3790)
         );
  CLKBUF_X1 U3745 ( .A(n5444), .Z(n5445) );
  NOR2_X1 U3746 ( .A1(n3758), .A2(n3759), .ZN(n3785) );
  NAND2_X1 U3747 ( .A1(n3744), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3758)
         );
  INV_X1 U3748 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3759) );
  NOR2_X1 U3749 ( .A1(n3727), .A2(n5277), .ZN(n3744) );
  NAND2_X1 U3750 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3727)
         );
  INV_X1 U3751 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5277) );
  CLKBUF_X1 U3752 ( .A(n5264), .Z(n5265) );
  NAND2_X1 U3753 ( .A1(n3105), .A2(n5195), .ZN(n3104) );
  INV_X1 U3754 ( .A(n3106), .ZN(n3105) );
  NAND2_X1 U3755 ( .A1(n3681), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3698)
         );
  INV_X1 U3756 ( .A(n3673), .ZN(n3681) );
  AOI21_X1 U3757 ( .B1(n3678), .B2(n3803), .A(n3677), .ZN(n5034) );
  CLKBUF_X1 U3758 ( .A(n4681), .Z(n4682) );
  NAND2_X1 U3759 ( .A1(n3662), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3666)
         );
  AND2_X1 U3760 ( .A1(n3641), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3662)
         );
  OAI211_X1 U3761 ( .C1(n3653), .C2(n5305), .A(n3639), .B(n3638), .ZN(n4368)
         );
  NAND2_X1 U3762 ( .A1(n4362), .A2(n3637), .ZN(n4303) );
  NAND2_X1 U3763 ( .A1(n5393), .A2(n3065), .ZN(n3064) );
  NOR2_X1 U3764 ( .A1(n3030), .A2(n5474), .ZN(n3065) );
  AND2_X1 U3765 ( .A1(n4205), .A2(n4204), .ZN(n5496) );
  AND2_X1 U3766 ( .A1(n4201), .A2(n4200), .ZN(n5804) );
  NAND2_X1 U3767 ( .A1(n5989), .A2(n5839), .ZN(n3083) );
  AOI21_X1 U3768 ( .B1(n3042), .B2(n3044), .A(n3023), .ZN(n3039) );
  AND2_X1 U3769 ( .A1(n4183), .A2(n4182), .ZN(n5452) );
  AND2_X1 U3770 ( .A1(n4180), .A2(n4179), .ZN(n5460) );
  NOR2_X1 U3771 ( .A1(n5857), .A2(n5460), .ZN(n5459) );
  OR2_X1 U3772 ( .A1(n5859), .A2(n5860), .ZN(n5857) );
  AND2_X1 U3773 ( .A1(n5269), .A2(n5270), .ZN(n5294) );
  NAND2_X1 U3774 ( .A1(n5294), .A2(n5293), .ZN(n5859) );
  NOR2_X1 U3775 ( .A1(n3049), .A2(n3046), .ZN(n3048) );
  AOI21_X1 U3776 ( .B1(n5698), .B2(n3047), .A(n3046), .ZN(n3045) );
  INV_X1 U3777 ( .A(n5235), .ZN(n3049) );
  AND2_X1 U3778 ( .A1(n4167), .A2(n4166), .ZN(n5199) );
  NAND2_X1 U3779 ( .A1(n5151), .A2(n3069), .ZN(n5198) );
  NAND2_X1 U3780 ( .A1(n5151), .A2(n5150), .ZN(n5161) );
  INV_X1 U3781 ( .A(n4683), .ZN(n3054) );
  NAND2_X1 U3782 ( .A1(n3056), .A2(n4152), .ZN(n4622) );
  INV_X1 U3783 ( .A(n4474), .ZN(n4152) );
  INV_X1 U3784 ( .A(n4475), .ZN(n3056) );
  NOR2_X1 U3785 ( .A1(n6330), .A2(n6331), .ZN(n5725) );
  NOR2_X1 U3786 ( .A1(n4535), .A2(n4534), .ZN(n5708) );
  INV_X1 U3787 ( .A(n6341), .ZN(n4535) );
  OR2_X1 U3788 ( .A1(n5853), .A2(n4535), .ZN(n5823) );
  XNOR2_X1 U3789 ( .A(n3330), .B(n3353), .ZN(n3302) );
  NAND2_X1 U3790 ( .A1(n3364), .A2(n3363), .ZN(n3050) );
  NAND2_X1 U3791 ( .A1(n3390), .A2(n3017), .ZN(n3072) );
  INV_X1 U3792 ( .A(n3390), .ZN(n3075) );
  NAND2_X1 U3793 ( .A1(n3388), .A2(n3074), .ZN(n3073) );
  INV_X1 U3794 ( .A(n3077), .ZN(n3076) );
  OAI21_X1 U3795 ( .B1(n3393), .B2(n3081), .A(n3078), .ZN(n3077) );
  INV_X1 U3796 ( .A(n3081), .ZN(n3071) );
  NAND2_X1 U3797 ( .A1(n3393), .A2(n3078), .ZN(n3032) );
  INV_X1 U3798 ( .A(n5884), .ZN(n5318) );
  INV_X1 U3799 ( .A(n3405), .ZN(n3407) );
  INV_X1 U3800 ( .A(n3341), .ZN(n4112) );
  INV_X1 U3801 ( .A(n4440), .ZN(n6459) );
  NAND2_X1 U3802 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  INV_X1 U3803 ( .A(n4606), .ZN(n4962) );
  NAND2_X1 U3804 ( .A1(n4962), .A2(n4614), .ZN(n4826) );
  AND2_X1 U3805 ( .A1(n5877), .A2(n4458), .ZN(n4745) );
  AND2_X1 U3806 ( .A1(n3001), .A2(n4887), .ZN(n4695) );
  OR3_X1 U3807 ( .A1(n6580), .A2(STATE2_REG_0__SCAN_IN), .A3(n4488), .ZN(n4525) );
  INV_X1 U3808 ( .A(n4916), .ZN(n4790) );
  AND2_X1 U3809 ( .A1(n5447), .A2(n4127), .ZN(n6139) );
  INV_X1 U3810 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5159) );
  AND2_X1 U3811 ( .A1(n5447), .A2(n4134), .ZN(n6138) );
  INV_X1 U3812 ( .A(n6191), .ZN(n6170) );
  INV_X1 U3813 ( .A(n6178), .ZN(n6196) );
  INV_X1 U3814 ( .A(n6199), .ZN(n6181) );
  INV_X1 U3815 ( .A(n6210), .ZN(n5528) );
  AND2_X2 U3816 ( .A1(n4310), .A2(n4374), .ZN(n6210) );
  AND2_X1 U3817 ( .A1(n6225), .A2(n3339), .ZN(n6214) );
  AND2_X1 U3818 ( .A1(n6225), .A2(n4381), .ZN(n6217) );
  INV_X1 U3819 ( .A(n6225), .ZN(n6216) );
  OR2_X1 U3820 ( .A1(n6214), .A2(n6217), .ZN(n6220) );
  INV_X1 U3821 ( .A(n6220), .ZN(n6224) );
  BUF_X1 U3822 ( .A(n6258), .Z(n6251) );
  INV_X1 U3823 ( .A(n6484), .ZN(n6592) );
  OAI21_X1 U3824 ( .B1(n4254), .B2(n6485), .A(n4228), .ZN(n4299) );
  CLKBUF_X1 U3825 ( .A(n4351), .Z(n4359) );
  NAND2_X1 U3826 ( .A1(n4232), .A2(n4231), .ZN(n4376) );
  INV_X1 U3827 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5631) );
  AND2_X1 U3828 ( .A1(n3010), .A2(n5512), .ZN(n5982) );
  INV_X1 U3829 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5653) );
  INV_X1 U3830 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5094) );
  INV_X1 U3831 ( .A(n6281), .ZN(n6266) );
  INV_X1 U3832 ( .A(n6271), .ZN(n5695) );
  INV_X1 U3833 ( .A(n6060), .ZN(n6278) );
  XNOR2_X1 U3834 ( .A(n3552), .B(n3551), .ZN(n5746) );
  NAND2_X1 U3835 ( .A1(n5572), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3550) );
  AND2_X1 U3836 ( .A1(n5975), .A2(n3013), .ZN(n5591) );
  NAND2_X1 U3837 ( .A1(n5610), .A2(n3089), .ZN(n3087) );
  XNOR2_X1 U3838 ( .A(n3092), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3089)
         );
  NAND2_X1 U3839 ( .A1(n5664), .A2(n3537), .ZN(n5660) );
  NAND2_X1 U3840 ( .A1(n3041), .A2(n3536), .ZN(n5666) );
  NAND2_X1 U3841 ( .A1(n5673), .A2(n3535), .ZN(n3041) );
  NAND2_X1 U3842 ( .A1(n6032), .A2(n5865), .ZN(n6285) );
  AND2_X1 U3843 ( .A1(n4291), .A2(n4271), .ZN(n6337) );
  CLKBUF_X1 U3844 ( .A(n4478), .Z(n4479) );
  INV_X1 U3845 ( .A(n4696), .ZN(n5877) );
  INV_X1 U3846 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6344) );
  NOR2_X1 U3847 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6045) );
  INV_X1 U3848 ( .A(n4905), .ZN(n4865) );
  INV_X1 U3849 ( .A(n5120), .ZN(n5144) );
  INV_X1 U3850 ( .A(n5114), .ZN(n5143) );
  NOR2_X2 U3851 ( .A1(n4963), .A2(n4964), .ZN(n5026) );
  INV_X1 U3852 ( .A(n6448), .ZN(n5256) );
  NAND2_X1 U3853 ( .A1(n4745), .A2(n4964), .ZN(n4945) );
  NOR2_X1 U3854 ( .A1(n6689), .A2(n4790), .ZN(n6351) );
  NOR2_X1 U3855 ( .A1(n6675), .A2(n4790), .ZN(n6367) );
  NOR2_X1 U3856 ( .A1(n4505), .A2(n4790), .ZN(n6417) );
  NOR2_X1 U3857 ( .A1(n6694), .A2(n4790), .ZN(n6423) );
  NOR2_X1 U3858 ( .A1(n4625), .A2(n4790), .ZN(n6429) );
  NOR2_X1 U3859 ( .A1(n5035), .A2(n4790), .ZN(n6444) );
  OR2_X1 U3860 ( .A1(n6052), .A2(n6580), .ZN(n6492) );
  INV_X1 U3861 ( .A(n6595), .ZN(n6504) );
  INV_X1 U3862 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U3863 ( .C1(n6271), .C2(n5567), .A(n5730), .B(n5566), .ZN(n5568)
         );
  NAND2_X1 U3864 ( .A1(n5103), .A2(n3697), .ZN(n5102) );
  AOI21_X1 U3865 ( .B1(n3670), .B2(n3803), .A(n3669), .ZN(n4680) );
  INV_X1 U3866 ( .A(n4680), .ZN(n3671) );
  NAND2_X1 U3867 ( .A1(n3108), .A2(n3111), .ZN(n5499) );
  AND2_X1 U3868 ( .A1(n3103), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3008) );
  AND3_X1 U3869 ( .A1(n3180), .A2(n3179), .A3(n3178), .ZN(n3009) );
  OR2_X1 U3870 ( .A1(n5432), .A2(n5511), .ZN(n3010) );
  INV_X1 U3871 ( .A(n5422), .ZN(n3066) );
  AND2_X1 U3872 ( .A1(n3115), .A2(n3120), .ZN(n3011) );
  OR2_X1 U3873 ( .A1(n5989), .A2(n6289), .ZN(n5699) );
  INV_X1 U3874 ( .A(n5699), .ZN(n3046) );
  AND2_X1 U3875 ( .A1(n3086), .A2(n5832), .ZN(n3012) );
  AND2_X2 U3876 ( .A1(n3145), .A2(n4404), .ZN(n3380) );
  AND2_X2 U3877 ( .A1(n3139), .A2(n4409), .ZN(n3415) );
  AND2_X1 U3878 ( .A1(n3025), .A2(n3544), .ZN(n3013) );
  INV_X1 U3879 ( .A(n4286), .ZN(n4489) );
  AND4_X1 U3880 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3015)
         );
  AND2_X1 U3881 ( .A1(n5479), .A2(n5478), .ZN(n3016) );
  NAND2_X1 U3882 ( .A1(n3040), .A2(n3039), .ZN(n5648) );
  AND2_X1 U3883 ( .A1(n3387), .A2(n3395), .ZN(n3017) );
  NAND2_X1 U3884 ( .A1(n3372), .A2(n3371), .ZN(n3406) );
  AND2_X1 U3885 ( .A1(n4108), .A2(n5487), .ZN(n5479) );
  AND2_X1 U3886 ( .A1(n5339), .A2(n5489), .ZN(n5482) );
  AND4_X1 U3887 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n3018)
         );
  NAND2_X1 U3888 ( .A1(n5989), .A2(n5987), .ZN(n3019) );
  NOR2_X1 U3889 ( .A1(n5444), .A2(n5525), .ZN(n5526) );
  AND2_X1 U3890 ( .A1(n4108), .A2(n3125), .ZN(n5408) );
  NAND2_X1 U3891 ( .A1(n3071), .A2(n3032), .ZN(n3428) );
  INV_X1 U3892 ( .A(n3260), .ZN(n4272) );
  NOR2_X1 U3893 ( .A1(n5989), .A2(n5239), .ZN(n3021) );
  INV_X1 U3894 ( .A(n3337), .ZN(n3243) );
  OR2_X1 U3895 ( .A1(n5485), .A2(n5474), .ZN(n3022) );
  NOR2_X1 U3896 ( .A1(n5432), .A2(n3113), .ZN(n5503) );
  NAND2_X1 U3897 ( .A1(n3019), .A2(n3537), .ZN(n3023) );
  INV_X1 U3898 ( .A(n3086), .ZN(n3085) );
  NAND2_X1 U3899 ( .A1(n3539), .A2(n5839), .ZN(n3086) );
  INV_X1 U3900 ( .A(n3622), .ZN(n5314) );
  INV_X1 U3901 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5305) );
  INV_X1 U3902 ( .A(n3339), .ZN(n4378) );
  AND2_X1 U3903 ( .A1(n3115), .A2(n3116), .ZN(n5443) );
  NOR2_X1 U3904 ( .A1(n5033), .A2(n3106), .ZN(n5156) );
  XNOR2_X1 U3905 ( .A(n5291), .B(n3774), .ZN(n5679) );
  INV_X1 U3906 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U3907 ( .A1(n3243), .A2(n3245), .ZN(n4253) );
  INV_X1 U3908 ( .A(n3063), .ZN(n6015) );
  AND2_X1 U3909 ( .A1(n3013), .A2(n5757), .ZN(n3024) );
  AND2_X1 U3910 ( .A1(n2990), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3025)
         );
  INV_X1 U3911 ( .A(n3094), .ZN(n3093) );
  AND2_X1 U3912 ( .A1(n4009), .A2(n4008), .ZN(n3026) );
  NAND2_X1 U3913 ( .A1(n5805), .A2(n5804), .ZN(n5495) );
  AND2_X1 U3914 ( .A1(n3026), .A2(n5478), .ZN(n3027) );
  INV_X1 U3915 ( .A(n5627), .ZN(n3095) );
  NOR2_X1 U3916 ( .A1(n5989), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5627)
         );
  AND2_X1 U3917 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3028) );
  INV_X1 U3918 ( .A(n5530), .ZN(n6206) );
  INV_X1 U3919 ( .A(n3623), .ZN(n3761) );
  NOR2_X1 U3920 ( .A1(n4465), .A2(n4472), .ZN(n4471) );
  NAND3_X1 U3921 ( .A1(n3099), .A2(n3760), .A3(n3621), .ZN(n4367) );
  INV_X1 U3922 ( .A(n3559), .ZN(n3522) );
  AND2_X1 U3923 ( .A1(n3553), .A2(n2993), .ZN(n3559) );
  OR2_X1 U3924 ( .A1(n4622), .A2(n4623), .ZN(n4684) );
  INV_X1 U3925 ( .A(n4684), .ZN(n3055) );
  INV_X1 U3926 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3053) );
  INV_X1 U3927 ( .A(n3099), .ZN(n4302) );
  NAND2_X1 U3928 ( .A1(n4301), .A2(n4303), .ZN(n3099) );
  AND2_X1 U3929 ( .A1(n3116), .A2(n5446), .ZN(n3029) );
  XNOR2_X1 U3930 ( .A(n3061), .B(n4360), .ZN(n4274) );
  INV_X1 U3931 ( .A(n5101), .ZN(n3697) );
  AND2_X1 U3932 ( .A1(n5352), .A2(n5351), .ZN(n3030) );
  AND2_X1 U3933 ( .A1(n3852), .A2(n3851), .ZN(n3031) );
  INV_X1 U3934 ( .A(n3120), .ZN(n3119) );
  NAND2_X1 U3935 ( .A1(n3774), .A2(n5680), .ZN(n3120) );
  INV_X1 U3936 ( .A(n3612), .ZN(n3096) );
  NOR2_X2 U3937 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4445) );
  INV_X1 U3938 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3082) );
  INV_X1 U3939 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3060) );
  NAND2_X2 U3940 ( .A1(n3033), .A2(n3351), .ZN(n3393) );
  NAND2_X2 U3941 ( .A1(n3034), .A2(n3543), .ZN(n5973) );
  INV_X2 U3942 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3036) );
  AND2_X2 U3943 ( .A1(n3145), .A2(n4435), .ZN(n3379) );
  AND2_X2 U3944 ( .A1(n3334), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3145)
         );
  NAND2_X1 U3945 ( .A1(n5673), .A2(n3042), .ZN(n3040) );
  NAND2_X1 U3946 ( .A1(n5235), .A2(n5234), .ZN(n3047) );
  OAI21_X1 U3947 ( .B1(n5233), .B2(n5234), .A(n5235), .ZN(n5697) );
  OAI21_X2 U3948 ( .B1(n5687), .B2(n5690), .A(n5688), .ZN(n5683) );
  XNOR2_X1 U3949 ( .A(n3362), .B(n3050), .ZN(n4478) );
  NAND2_X1 U3950 ( .A1(n3103), .A2(n3052), .ZN(n3051) );
  INV_X1 U3951 ( .A(n5572), .ZN(n5564) );
  AND2_X2 U3952 ( .A1(n4496), .A2(n4286), .ZN(n4254) );
  NOR2_X4 U3953 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4430) );
  NOR2_X1 U3954 ( .A1(n2993), .A2(n3238), .ZN(n3343) );
  NOR2_X1 U3955 ( .A1(n4286), .A2(n2993), .ZN(n4267) );
  INV_X1 U3956 ( .A(n5372), .ZN(n5336) );
  AOI21_X1 U3957 ( .B1(n5372), .B2(n3060), .A(n3059), .ZN(n3058) );
  NAND2_X1 U3958 ( .A1(n4138), .A2(n4139), .ZN(n3061) );
  NOR2_X2 U3959 ( .A1(n5517), .A2(n4199), .ZN(n5805) );
  NOR2_X2 U3960 ( .A1(n6016), .A2(n6017), .ZN(n3063) );
  NOR3_X2 U3961 ( .A1(n5485), .A2(n5421), .A3(n3064), .ZN(n5370) );
  NOR3_X2 U3962 ( .A1(n5485), .A2(n5474), .A3(n5421), .ZN(n5422) );
  AND2_X2 U3963 ( .A1(n5151), .A2(n3067), .ZN(n5269) );
  AND2_X2 U3964 ( .A1(n3082), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3139)
         );
  INV_X1 U3965 ( .A(n5619), .ZN(n3084) );
  NAND2_X1 U3966 ( .A1(n5619), .A2(n3085), .ZN(n5830) );
  NAND2_X1 U3967 ( .A1(n3088), .A2(n3087), .ZN(n5787) );
  NAND2_X1 U3968 ( .A1(n5610), .A2(n3093), .ZN(n5629) );
  INV_X1 U3969 ( .A(n5610), .ZN(n5634) );
  NOR2_X1 U3970 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3094)
         );
  NAND4_X1 U3971 ( .A1(n3251), .A2(n3255), .A3(n3256), .A4(n4436), .ZN(n3257)
         );
  NAND2_X1 U3973 ( .A1(n3621), .A2(n3760), .ZN(n3102) );
  NAND2_X1 U3974 ( .A1(n3102), .A2(n4302), .ZN(n3100) );
  NAND2_X1 U3975 ( .A1(n4367), .A2(n4368), .ZN(n3101) );
  NAND2_X1 U3976 ( .A1(n3103), .A2(n3028), .ZN(n3248) );
  NAND2_X1 U3977 ( .A1(n3118), .A2(n3029), .ZN(n5444) );
  CLKBUF_X1 U3978 ( .A(n3118), .Z(n3115) );
  OR2_X1 U3979 ( .A1(n5327), .A2(n6281), .ZN(n4104) );
  AND2_X2 U3980 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U3981 ( .A1(n5408), .A2(n5410), .ZN(n5389) );
  AOI22_X1 U3982 ( .A1(n3969), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U3983 ( .A1(n3969), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3165) );
  AND2_X1 U3984 ( .A1(n2987), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U3985 ( .A1(n2986), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U3986 ( .A1(n3234), .A2(n3260), .ZN(n3236) );
  AND2_X1 U3987 ( .A1(n2985), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U3988 ( .A1(n3244), .A2(n3253), .ZN(n4111) );
  OR2_X1 U3989 ( .A1(n3244), .A2(n3610), .ZN(n5884) );
  XNOR2_X1 U3990 ( .A(n5390), .B(n5308), .ZN(n5327) );
  NAND2_X1 U3991 ( .A1(n5264), .A2(n5292), .ZN(n5291) );
  AOI22_X1 U3992 ( .A1(n2999), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U3993 ( .A1(n3283), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3284) );
  NOR2_X1 U3994 ( .A1(n6345), .A2(n4480), .ZN(n3127) );
  AND2_X1 U3995 ( .A1(n4291), .A2(n4273), .ZN(n6293) );
  INV_X1 U3996 ( .A(n6293), .ZN(n6335) );
  AND2_X1 U3997 ( .A1(n3004), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3128) );
  AND2_X1 U3998 ( .A1(n2982), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3129) );
  INV_X1 U3999 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3551) );
  INV_X1 U4000 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6049) );
  INV_X1 U4001 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4002 ( .A1(n5989), .A2(n5714), .ZN(n3130) );
  INV_X1 U4003 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3791) );
  AOI21_X1 U4004 ( .B1(n4951), .B2(STATE2_REG_3__SCAN_IN), .A(n4790), .ZN(
        n4957) );
  OR2_X1 U4005 ( .A1(n3571), .A2(n3570), .ZN(n3573) );
  NAND2_X1 U4006 ( .A1(n3285), .A2(n3284), .ZN(n3286) );
  AND2_X1 U4007 ( .A1(n3588), .A2(n3574), .ZN(n3577) );
  INV_X1 U4008 ( .A(n3314), .ZN(n3315) );
  AND2_X1 U4009 ( .A1(n4116), .A2(n4115), .ZN(n4117) );
  AOI22_X1 U4010 ( .A1(n3969), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3189) );
  INV_X1 U4011 ( .A(n5504), .ZN(n3888) );
  NOR2_X1 U4012 ( .A1(n3622), .A2(n4641), .ZN(n3623) );
  INV_X1 U4014 ( .A(n4107), .ZN(n3950) );
  INV_X1 U4015 ( .A(n3761), .ZN(n5310) );
  OR3_X1 U4016 ( .A1(n5989), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5755), 
        .ZN(n5559) );
  NAND2_X1 U4017 ( .A1(n3678), .A2(n3559), .ZN(n3517) );
  OR2_X1 U4018 ( .A1(n3446), .A2(n3445), .ZN(n3458) );
  AND4_X1 U4019 ( .A1(n5919), .A2(REIP_REG_25__SCAN_IN), .A3(
        REIP_REG_24__SCAN_IN), .A4(REIP_REG_26__SCAN_IN), .ZN(n5424) );
  INV_X1 U4020 ( .A(n3642), .ZN(n3613) );
  AND2_X1 U4021 ( .A1(n4157), .A2(n4156), .ZN(n4683) );
  NAND2_X1 U4022 ( .A1(n4026), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4050)
         );
  AND2_X1 U4023 ( .A1(n4151), .A2(n4150), .ZN(n4474) );
  OR2_X1 U4024 ( .A1(n4491), .A2(n6715), .ZN(n4483) );
  NAND2_X1 U4025 ( .A1(n4429), .A2(n3053), .ZN(n3427) );
  NAND2_X1 U4026 ( .A1(n3313), .A2(n3312), .ZN(n3308) );
  INV_X1 U4027 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6461) );
  AND2_X1 U4028 ( .A1(n4285), .A2(n4284), .ZN(n4408) );
  INV_X1 U4029 ( .A(n3885), .ZN(n3614) );
  NAND2_X1 U4030 ( .A1(n5380), .A2(n4129), .ZN(n6077) );
  NOR2_X1 U4031 ( .A1(n3698), .A2(n5159), .ZN(n3713) );
  INV_X1 U4032 ( .A(n5925), .ZN(n5438) );
  AND2_X1 U4033 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3613), .ZN(n3641)
         );
  AND2_X1 U4034 ( .A1(n5567), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4134) );
  INV_X1 U4035 ( .A(n3803), .ZN(n3789) );
  OR2_X1 U4036 ( .A1(n4229), .A2(n2997), .ZN(n4418) );
  NAND2_X1 U4037 ( .A1(n4031), .A2(n4030), .ZN(n5420) );
  AND2_X1 U4038 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  XNOR2_X1 U4039 ( .A(n3529), .B(n4159), .ZN(n5171) );
  INV_X1 U4040 ( .A(n2997), .ZN(n4307) );
  OR2_X1 U4041 ( .A1(n4836), .A2(n5877), .ZN(n4888) );
  INV_X1 U4042 ( .A(n4887), .ZN(n4964) );
  INV_X1 U4043 ( .A(n5206), .ZN(n5258) );
  NAND2_X1 U4044 ( .A1(n3412), .A2(n3411), .ZN(n4786) );
  OR2_X1 U4045 ( .A1(n4644), .A2(n4887), .ZN(n4864) );
  INV_X1 U4046 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5321) );
  INV_X1 U4047 ( .A(n4254), .ZN(n6594) );
  NAND2_X1 U4048 ( .A1(n4224), .A2(n4226), .ZN(n6590) );
  NOR2_X1 U4049 ( .A1(n5927), .A2(n5328), .ZN(n5919) );
  NAND2_X1 U4050 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3919)
         );
  AND2_X1 U4051 ( .A1(n5380), .A2(n4212), .ZN(n6178) );
  AND2_X1 U4052 ( .A1(n5447), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6191) );
  AND2_X1 U4053 ( .A1(n5380), .A2(n4217), .ZN(n6192) );
  INV_X1 U4054 ( .A(n6159), .ZN(n6173) );
  AOI21_X1 U4055 ( .B1(n5376), .B2(n5399), .A(n5375), .ZN(n5377) );
  NOR2_X1 U4056 ( .A1(n6592), .A2(n6227), .ZN(n6258) );
  INV_X1 U4057 ( .A(n4313), .ZN(n4356) );
  INV_X1 U4058 ( .A(n4376), .ZN(n4341) );
  INV_X1 U4059 ( .A(n5638), .ZN(n5965) );
  AND2_X1 U4060 ( .A1(n4268), .A2(n3096), .ZN(n6476) );
  AOI21_X1 U4061 ( .B1(n3628), .B2(n4887), .A(n4641), .ZN(n4364) );
  INV_X1 U4062 ( .A(n5823), .ZN(n5844) );
  INV_X1 U4063 ( .A(n6492), .ZN(n5891) );
  NAND2_X1 U4064 ( .A1(n4841), .A2(n4840), .ZN(n4863) );
  NOR2_X1 U4065 ( .A1(n4888), .A2(n4964), .ZN(n4905) );
  OAI21_X1 U4066 ( .B1(n5119), .B2(n5146), .A(n5212), .ZN(n5142) );
  OAI21_X1 U4067 ( .B1(n4703), .B2(n4702), .A(n4701), .ZN(n4727) );
  OAI21_X1 U4068 ( .B1(n4553), .B2(n4487), .A(n4486), .ZN(n4524) );
  INV_X1 U4069 ( .A(n6352), .ZN(n6394) );
  INV_X1 U4070 ( .A(n6407), .ZN(n6354) );
  INV_X1 U4071 ( .A(n4992), .ZN(n6401) );
  AND2_X1 U4072 ( .A1(n4965), .A2(n4964), .ZN(n5206) );
  AND2_X1 U4073 ( .A1(n5202), .A2(n5872), .ZN(n5210) );
  INV_X1 U4074 ( .A(n4826), .ZN(n6440) );
  INV_X1 U4075 ( .A(n5872), .ZN(n6353) );
  NOR2_X1 U4076 ( .A1(n6661), .A2(n4790), .ZN(n6411) );
  NOR2_X1 U4077 ( .A1(n6641), .A2(n4790), .ZN(n6435) );
  AND2_X1 U4078 ( .A1(n5321), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3609) );
  INV_X1 U4079 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6520) );
  INV_X1 U4080 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6715) );
  AND2_X1 U4081 ( .A1(n6520), .A2(STATE_REG_1__SCAN_IN), .ZN(n6791) );
  INV_X1 U4082 ( .A(n6192), .ZN(n6134) );
  INV_X1 U4083 ( .A(n6139), .ZN(n6150) );
  XOR2_X1 U4084 ( .A(n5378), .B(n5377), .Z(n5735) );
  NAND2_X1 U4085 ( .A1(n6210), .A2(n5314), .ZN(n5530) );
  INV_X1 U4086 ( .A(n6227), .ZN(n6260) );
  INV_X1 U4087 ( .A(n4299), .ZN(n4313) );
  INV_X1 U4088 ( .A(n6337), .ZN(n5870) );
  INV_X1 U4089 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4951) );
  NOR2_X1 U4090 ( .A1(n5001), .A2(n5000), .ZN(n5032) );
  AOI22_X1 U4091 ( .A1(n5210), .A2(n5207), .B1(n6345), .B2(n5204), .ZN(n5263)
         );
  NAND2_X1 U4092 ( .A1(n4962), .A2(n4695), .ZN(n6448) );
  NOR2_X1 U4093 ( .A1(n4792), .A2(n4791), .ZN(n4833) );
  INV_X1 U4094 ( .A(n6423), .ZN(n5250) );
  NAND2_X1 U4095 ( .A1(n3609), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6498) );
  INV_X1 U4096 ( .A(n6577), .ZN(n6508) );
  INV_X1 U4097 ( .A(n6570), .ZN(n6565) );
  NAND2_X1 U4098 ( .A1(n3415), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U4099 ( .A1(n2989), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4100 ( .A1(n4086), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U4101 ( .A1(n3295), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4102 ( .A1(n2985), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4103 ( .A1(n3316), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3137)
         );
  NAND2_X1 U4104 ( .A1(n3379), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U4105 ( .A1(n3283), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U4106 ( .A1(n3005), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3144)
         );
  NAND2_X1 U4107 ( .A1(n3969), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U4108 ( .A1(n3374), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3142)
         );
  NAND2_X1 U4109 ( .A1(n3271), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4110 ( .A1(n2987), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4111 ( .A1(n3380), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3148)
         );
  AND2_X2 U4112 ( .A1(n4409), .A2(n4404), .ZN(n3282) );
  NAND2_X1 U4113 ( .A1(n3282), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3147)
         );
  NAND2_X1 U4115 ( .A1(n3323), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3146)
         );
  AOI22_X1 U4116 ( .A1(n4086), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4117 ( .A1(n3415), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4118 ( .A1(n3374), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4119 ( .A1(n3316), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4120 ( .A1(n2986), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4121 ( .A1(n2988), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4122 ( .A1(n3379), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4123 ( .A1(n3005), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4124 ( .A1(n3415), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3164) );
  AND2_X2 U4125 ( .A1(n3202), .A2(n3203), .ZN(n3237) );
  OAI21_X1 U4126 ( .B1(n3260), .B2(n3252), .A(n4305), .ZN(n3191) );
  AOI22_X1 U4127 ( .A1(n3005), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4128 ( .A1(n3316), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4129 ( .A1(n4086), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4130 ( .A1(n2988), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3172) );
  NOR2_X1 U4131 ( .A1(n3177), .A2(n3176), .ZN(n3181) );
  AOI22_X1 U4132 ( .A1(n3374), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4133 ( .A1(n3380), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4134 ( .A1(n3969), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4135 ( .A1(n3380), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4136 ( .A1(n3316), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4137 ( .A1(n3373), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4138 ( .A1(n2986), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4139 ( .A1(n3379), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4140 ( .A1(n3374), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4141 ( .A1(n2988), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3186) );
  NAND3_X1 U4142 ( .A1(n3191), .A2(n3239), .A3(n3622), .ZN(n3193) );
  NAND3_X1 U4143 ( .A1(n3192), .A2(n4305), .A3(n3339), .ZN(n3341) );
  NAND2_X1 U4144 ( .A1(n3193), .A2(n3341), .ZN(n3212) );
  AOI22_X1 U4145 ( .A1(n4086), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4146 ( .A1(n2986), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4147 ( .A1(n2988), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4148 ( .A1(n3283), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4149 ( .A1(n3415), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3198) );
  INV_X1 U4150 ( .A(n3252), .ZN(n3628) );
  NAND2_X2 U4151 ( .A1(n3628), .A2(n3553), .ZN(n3244) );
  AOI22_X1 U4152 ( .A1(n2989), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4153 ( .A1(n3969), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4154 ( .A1(n3005), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4155 ( .A1(n3415), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4156 ( .A1(n3316), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4157 ( .A1(n2984), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4158 ( .A1(n3380), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4159 ( .A1(n2987), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3208) );
  NAND3_X1 U4160 ( .A1(n3212), .A2(n4496), .A3(n4111), .ZN(n3233) );
  NAND2_X1 U4161 ( .A1(n3415), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4162 ( .A1(n3969), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4163 ( .A1(n4086), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4164 ( .A1(n3295), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3213) );
  NAND2_X1 U4165 ( .A1(n3005), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4166 ( .A1(n3374), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3219)
         );
  NAND2_X1 U4167 ( .A1(n2989), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4168 ( .A1(n3271), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4169 ( .A1(n3316), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3224)
         );
  NAND2_X1 U4170 ( .A1(n3379), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4171 ( .A1(n2984), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4172 ( .A1(n3282), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3221)
         );
  NAND2_X1 U4173 ( .A1(n3380), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4174 ( .A1(n3283), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4175 ( .A1(n2986), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4176 ( .A1(n3323), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3225)
         );
  NAND4_X4 U4177 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n4286)
         );
  INV_X1 U4178 ( .A(n3244), .ZN(n3234) );
  AND2_X1 U4179 ( .A1(n4305), .A2(n3622), .ZN(n3235) );
  NAND2_X1 U4180 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6523) );
  OAI21_X1 U4181 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6523), .ZN(n4128) );
  INV_X1 U4182 ( .A(n4128), .ZN(n3238) );
  INV_X1 U4183 ( .A(n3343), .ZN(n3240) );
  NAND2_X1 U4184 ( .A1(n3239), .A2(n3253), .ZN(n3355) );
  AOI21_X1 U4185 ( .B1(n3237), .B2(n3240), .A(n3355), .ZN(n3241) );
  AND2_X1 U4186 ( .A1(n3249), .A2(n3241), .ZN(n3246) );
  NAND2_X1 U4187 ( .A1(n3260), .A2(n3553), .ZN(n3612) );
  AND2_X1 U4188 ( .A1(n3244), .A2(n4286), .ZN(n3245) );
  NAND2_X1 U4189 ( .A1(n6045), .A2(n3053), .ZN(n3615) );
  MUX2_X1 U4190 ( .A(n3615), .B(n3609), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3247) );
  NAND2_X1 U4191 ( .A1(n3248), .A2(n3247), .ZN(n3264) );
  INV_X1 U4192 ( .A(n3253), .ZN(n4506) );
  AOI21_X1 U4193 ( .B1(n3244), .B2(n4272), .A(n4506), .ZN(n3250) );
  AOI21_X1 U4194 ( .B1(n3249), .B2(n3250), .A(n4496), .ZN(n3258) );
  NAND2_X1 U4195 ( .A1(n6045), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6499) );
  AOI21_X1 U4196 ( .B1(n4278), .B2(n4286), .A(n6499), .ZN(n3256) );
  NAND2_X1 U4197 ( .A1(n3622), .A2(n4272), .ZN(n3610) );
  NOR2_X1 U4198 ( .A1(n3610), .A2(n3252), .ZN(n3254) );
  NAND2_X1 U4199 ( .A1(n3254), .A2(n4304), .ZN(n4436) );
  NAND2_X1 U4200 ( .A1(n4111), .A2(n4254), .ZN(n3255) );
  NOR2_X1 U4201 ( .A1(n3258), .A2(n3257), .ZN(n3263) );
  INV_X1 U4202 ( .A(n3259), .ZN(n3262) );
  NAND2_X1 U4203 ( .A1(n3559), .A2(n3260), .ZN(n3261) );
  NAND2_X1 U4204 ( .A1(n3262), .A2(n3261), .ZN(n4284) );
  NAND2_X1 U4205 ( .A1(n3263), .A2(n4284), .ZN(n3265) );
  INV_X1 U4206 ( .A(n3264), .ZN(n3267) );
  INV_X1 U4207 ( .A(n3265), .ZN(n3266) );
  AOI22_X1 U4208 ( .A1(n3317), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3275) );
  BUF_X1 U4209 ( .A(n3415), .Z(n3270) );
  BUF_X1 U4210 ( .A(n3380), .Z(n3269) );
  AOI22_X1 U4211 ( .A1(n3270), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4212 ( .A1(n3322), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4213 ( .A1(n2987), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3272) );
  NAND4_X1 U4214 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3280)
         );
  AOI22_X1 U4215 ( .A1(n4056), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4216 ( .A1(n2989), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3281) );
  INV_X1 U4217 ( .A(n3281), .ZN(n3287) );
  AOI22_X1 U4218 ( .A1(n4086), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4219 ( .A1(n4056), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4220 ( .A1(n3317), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4221 ( .A1(n3005), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4222 ( .A1(n2987), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3291) );
  NAND4_X1 U4223 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3301)
         );
  AOI22_X1 U4224 ( .A1(n3322), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4225 ( .A1(n3379), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4226 ( .A1(n4034), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4227 ( .A1(n3269), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3296) );
  NAND4_X1 U4228 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3300)
         );
  NAND2_X1 U4229 ( .A1(n3302), .A2(n3387), .ZN(n3312) );
  OAI21_X1 U4230 ( .B1(n3629), .B2(STATE2_REG_0__SCAN_IN), .A(n3312), .ZN(
        n3307) );
  INV_X1 U4231 ( .A(n3353), .ZN(n3305) );
  NAND2_X1 U4232 ( .A1(n3580), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3304) );
  AOI21_X1 U4233 ( .B1(n3260), .B2(n3525), .A(n3053), .ZN(n3303) );
  OAI211_X1 U4234 ( .C1(n3305), .C2(n4286), .A(n3304), .B(n3303), .ZN(n3306)
         );
  INV_X1 U4235 ( .A(n3306), .ZN(n3313) );
  NAND2_X1 U4236 ( .A1(n3307), .A2(n3306), .ZN(n3309) );
  NAND2_X2 U4237 ( .A1(n3309), .A2(n3308), .ZN(n4887) );
  NAND2_X1 U4238 ( .A1(n4489), .A2(n3253), .ZN(n3398) );
  OAI21_X1 U4239 ( .B1(n6594), .B2(n3353), .A(n3398), .ZN(n3310) );
  INV_X1 U4240 ( .A(n3310), .ZN(n3311) );
  OAI21_X1 U4241 ( .B1(n4887), .B2(n3522), .A(n3311), .ZN(n6273) );
  NAND2_X1 U4242 ( .A1(n6273), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6272)
         );
  XNOR2_X1 U4243 ( .A(n6272), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4249)
         );
  NAND2_X1 U4244 ( .A1(n3387), .A2(n3525), .ZN(n3523) );
  OAI21_X2 U4245 ( .B1(n3629), .B2(STATE2_REG_0__SCAN_IN), .A(n3315), .ZN(
        n3391) );
  AOI22_X1 U4246 ( .A1(n2989), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4247 ( .A1(n3317), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4248 ( .A1(n2987), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4249 ( .A1(n3005), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3318) );
  NAND4_X1 U4250 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3329)
         );
  AOI22_X1 U4251 ( .A1(n4056), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4252 ( .A1(n3322), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4253 ( .A1(n4085), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4254 ( .A1(n4034), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3324) );
  NAND4_X1 U4255 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3328)
         );
  INV_X1 U4256 ( .A(n3354), .ZN(n3333) );
  NAND2_X1 U4257 ( .A1(n3580), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4258 ( .A1(n3387), .A2(n3330), .ZN(n3331) );
  XNOR2_X1 U4259 ( .A(n3391), .B(n3392), .ZN(n3352) );
  INV_X1 U4260 ( .A(n3615), .ZN(n3370) );
  XNOR2_X1 U4261 ( .A(n6455), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6345)
         );
  NAND2_X1 U4262 ( .A1(n3370), .A2(n6345), .ZN(n3336) );
  INV_X1 U4263 ( .A(n3609), .ZN(n3369) );
  NAND2_X1 U4264 ( .A1(n3369), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3335) );
  NAND3_X1 U4265 ( .A1(n4267), .A2(n4304), .A3(n3237), .ZN(n4406) );
  AND2_X1 U4267 ( .A1(n4111), .A2(n4267), .ZN(n3342) );
  OAI211_X1 U4268 ( .C1(n4110), .C2(n3343), .A(n6794), .B(n6043), .ZN(n3344)
         );
  NAND2_X1 U4269 ( .A1(n3344), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3345) );
  INV_X1 U4270 ( .A(n3345), .ZN(n3349) );
  INV_X1 U4271 ( .A(n3346), .ZN(n3347) );
  NAND2_X1 U4272 ( .A1(n3349), .A2(n3348), .ZN(n3363) );
  INV_X1 U4273 ( .A(n4478), .ZN(n3350) );
  NAND2_X1 U4274 ( .A1(n3387), .A2(n3354), .ZN(n3351) );
  NAND2_X1 U4275 ( .A1(n3001), .A2(n3559), .ZN(n3359) );
  NAND2_X1 U4276 ( .A1(n3354), .A2(n3353), .ZN(n3396) );
  OAI21_X1 U4277 ( .B1(n3354), .B2(n3353), .A(n3396), .ZN(n3356) );
  INV_X1 U4278 ( .A(n3355), .ZN(n4279) );
  OAI211_X1 U4279 ( .C1(n3356), .C2(n6594), .A(n4279), .B(n3553), .ZN(n3357)
         );
  INV_X1 U4280 ( .A(n3357), .ZN(n3358) );
  NAND2_X1 U4281 ( .A1(n3359), .A2(n3358), .ZN(n4248) );
  NAND2_X1 U4282 ( .A1(n4249), .A2(n4248), .ZN(n4247) );
  INV_X1 U4283 ( .A(n6272), .ZN(n3360) );
  NAND2_X1 U4284 ( .A1(n3360), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3361)
         );
  NAND2_X1 U4285 ( .A1(n3363), .A2(n3362), .ZN(n3365) );
  NAND2_X1 U4286 ( .A1(n3008), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3372) );
  AND2_X1 U4287 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4288 ( .A1(n3366), .A2(n6461), .ZN(n4605) );
  INV_X1 U4289 ( .A(n3366), .ZN(n3367) );
  NAND2_X1 U4290 ( .A1(n3367), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3368) );
  NAND2_X1 U4291 ( .A1(n4605), .A2(n3368), .ZN(n4484) );
  AOI22_X1 U4292 ( .A1(n3370), .A2(n4484), .B1(n3369), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4293 ( .A1(n4405), .A2(n3053), .ZN(n3388) );
  AOI22_X1 U4294 ( .A1(n3005), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4295 ( .A1(n2989), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4296 ( .A1(n4056), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4297 ( .A1(n3270), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4298 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3386)
         );
  AOI22_X1 U4299 ( .A1(n3317), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4300 ( .A1(n2984), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4301 ( .A1(n3269), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4302 ( .A1(n2987), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4303 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3385)
         );
  INV_X1 U4304 ( .A(n3413), .ZN(n3389) );
  AOI22_X1 U4305 ( .A1(n3580), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3389), 
        .B2(n3395), .ZN(n3390) );
  INV_X1 U4306 ( .A(n3428), .ZN(n3394) );
  INV_X1 U4307 ( .A(n3395), .ZN(n3397) );
  NAND2_X1 U4308 ( .A1(n3396), .A2(n3397), .ZN(n3455) );
  OAI21_X1 U4309 ( .B1(n3397), .B2(n3396), .A(n3455), .ZN(n3400) );
  INV_X1 U4310 ( .A(n3398), .ZN(n3399) );
  AOI21_X1 U4311 ( .B1(n3400), .B2(n4254), .A(n3399), .ZN(n3401) );
  NAND2_X1 U4312 ( .A1(n3402), .A2(n3401), .ZN(n6263) );
  OAI21_X1 U4313 ( .B1(n6264), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6263), 
        .ZN(n3404) );
  NAND2_X1 U4314 ( .A1(n6264), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3403)
         );
  NAND2_X1 U4315 ( .A1(n3404), .A2(n3403), .ZN(n5051) );
  NAND2_X1 U4316 ( .A1(n3008), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3412) );
  NAND3_X1 U4317 ( .A1(n6344), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6349) );
  INV_X1 U4318 ( .A(n6349), .ZN(n3408) );
  NAND2_X1 U4319 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3408), .ZN(n6400) );
  NAND2_X1 U4320 ( .A1(n6344), .A2(n6400), .ZN(n3409) );
  NOR3_X1 U4321 ( .A1(n6344), .A2(n6461), .A3(n6455), .ZN(n4640) );
  NAND2_X1 U4322 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4640), .ZN(n4673) );
  NAND2_X1 U4323 ( .A1(n3409), .A2(n4673), .ZN(n4789) );
  OAI22_X1 U4324 ( .A1(n3615), .A2(n4789), .B1(n3609), .B2(n6344), .ZN(n3410)
         );
  INV_X1 U4325 ( .A(n3410), .ZN(n3411) );
  AOI22_X1 U4326 ( .A1(n3005), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4327 ( .A1(n2989), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4328 ( .A1(n4056), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4329 ( .A1(n3270), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3416) );
  NAND4_X1 U4330 ( .A1(n3419), .A2(n3418), .A3(n3417), .A4(n3416), .ZN(n3425)
         );
  AOI22_X1 U4331 ( .A1(n3317), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4332 ( .A1(n2985), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4333 ( .A1(n3269), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4334 ( .A1(n2987), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3420) );
  NAND4_X1 U4335 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3424)
         );
  AOI22_X1 U4336 ( .A1(n3606), .A2(n3454), .B1(n3580), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3426) );
  NAND2_X2 U4337 ( .A1(n3427), .A2(n3426), .ZN(n4459) );
  NAND2_X1 U4338 ( .A1(n3429), .A2(n3428), .ZN(n3430) );
  XNOR2_X1 U4339 ( .A(n3455), .B(n3454), .ZN(n3432) );
  OAI22_X2 U4340 ( .A1(n3640), .A2(n3522), .B1(n6594), .B2(n3432), .ZN(n3434)
         );
  INV_X1 U4341 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3433) );
  NAND2_X1 U4342 ( .A1(n5051), .A2(n5052), .ZN(n3436) );
  NAND2_X1 U4343 ( .A1(n3434), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3435)
         );
  NAND2_X1 U4344 ( .A1(n3436), .A2(n3435), .ZN(n4532) );
  INV_X1 U4345 ( .A(n3452), .ZN(n3449) );
  AOI22_X1 U4346 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n2989), .B1(n3270), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4347 ( .A1(n2987), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4348 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4079), .B1(n2984), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4349 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3269), .B1(n4080), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4350 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3446)
         );
  AOI22_X1 U4351 ( .A1(n3005), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4352 ( .A1(n4056), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4353 ( .A1(n4034), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4354 ( .A1(n3317), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4355 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  NAND2_X1 U4356 ( .A1(n3606), .A2(n3458), .ZN(n3448) );
  NAND2_X1 U4357 ( .A1(n3580), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4358 ( .A1(n3448), .A2(n3447), .ZN(n3450) );
  INV_X1 U4359 ( .A(n3450), .ZN(n3451) );
  NAND2_X1 U4360 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  NAND2_X1 U4361 ( .A1(n3479), .A2(n3453), .ZN(n3649) );
  NAND2_X1 U4362 ( .A1(n3455), .A2(n3454), .ZN(n3457) );
  INV_X1 U4363 ( .A(n3457), .ZN(n3459) );
  INV_X1 U4364 ( .A(n3458), .ZN(n3456) );
  OR2_X1 U4365 ( .A1(n3457), .A2(n3456), .ZN(n3504) );
  OAI211_X1 U4366 ( .C1(n3459), .C2(n3458), .A(n4254), .B(n3504), .ZN(n3460)
         );
  INV_X1 U4367 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4148) );
  XNOR2_X1 U4368 ( .A(n3461), .B(n4148), .ZN(n4533) );
  NAND2_X1 U4369 ( .A1(n4532), .A2(n4533), .ZN(n3463) );
  NAND2_X1 U4370 ( .A1(n3461), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3462)
         );
  NAND2_X1 U4371 ( .A1(n3463), .A2(n3462), .ZN(n4627) );
  INV_X1 U4372 ( .A(n3479), .ZN(n3477) );
  AOI22_X1 U4373 ( .A1(n3005), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4374 ( .A1(n2989), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4375 ( .A1(n4056), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4376 ( .A1(n3270), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3464) );
  NAND4_X1 U4377 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3473)
         );
  AOI22_X1 U4378 ( .A1(n3316), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4379 ( .A1(n2985), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4380 ( .A1(n3269), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4381 ( .A1(n2987), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4382 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3472)
         );
  NAND2_X1 U4383 ( .A1(n3606), .A2(n3481), .ZN(n3475) );
  NAND2_X1 U4384 ( .A1(n3580), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U4385 ( .A1(n3477), .A2(n3476), .ZN(n3501) );
  NAND2_X1 U4386 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  NAND2_X1 U4387 ( .A1(n3501), .A2(n3480), .ZN(n3665) );
  INV_X1 U4388 ( .A(n3481), .ZN(n3503) );
  XNOR2_X1 U4389 ( .A(n3504), .B(n3503), .ZN(n3482) );
  OAI22_X1 U4390 ( .A1(n3665), .A2(n3522), .B1(n3482), .B2(n6594), .ZN(n3484)
         );
  INV_X1 U4391 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3483) );
  XNOR2_X1 U4392 ( .A(n3484), .B(n3483), .ZN(n4628) );
  NAND2_X1 U4393 ( .A1(n4627), .A2(n4628), .ZN(n3486) );
  NAND2_X1 U4394 ( .A1(n3484), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3485)
         );
  NAND2_X1 U4395 ( .A1(n3486), .A2(n3485), .ZN(n4871) );
  INV_X1 U4396 ( .A(n3501), .ZN(n3500) );
  AOI22_X1 U4397 ( .A1(n4056), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4398 ( .A1(n2987), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4399 ( .A1(n4079), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4400 ( .A1(n4062), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3487) );
  NAND4_X1 U4401 ( .A1(n3490), .A2(n3489), .A3(n3488), .A4(n3487), .ZN(n3496)
         );
  AOI22_X1 U4402 ( .A1(n3005), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4403 ( .A1(n3316), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4404 ( .A1(n2989), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4405 ( .A1(n4034), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3491) );
  NAND4_X1 U4406 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3495)
         );
  NAND2_X1 U4407 ( .A1(n3606), .A2(n3505), .ZN(n3498) );
  NAND2_X1 U4408 ( .A1(n3580), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3497) );
  NAND2_X1 U4409 ( .A1(n3501), .A2(n3502), .ZN(n3670) );
  NAND3_X1 U4410 ( .A1(n3521), .A2(n3559), .A3(n3670), .ZN(n3508) );
  NOR2_X1 U4411 ( .A1(n3504), .A2(n3503), .ZN(n3506) );
  NAND2_X1 U4412 ( .A1(n3506), .A2(n3505), .ZN(n3527) );
  OAI211_X1 U4413 ( .C1(n3506), .C2(n3505), .A(n3527), .B(n4254), .ZN(n3507)
         );
  NAND2_X1 U4414 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  INV_X1 U4415 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4154) );
  XNOR2_X1 U4416 ( .A(n3509), .B(n4154), .ZN(n4872) );
  NAND2_X1 U4417 ( .A1(n4871), .A2(n4872), .ZN(n3511) );
  NAND2_X1 U4418 ( .A1(n3509), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3510)
         );
  NAND2_X1 U4419 ( .A1(n3511), .A2(n3510), .ZN(n5104) );
  NAND2_X1 U4420 ( .A1(n3606), .A2(n3525), .ZN(n3513) );
  NAND2_X1 U4421 ( .A1(n3580), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U4422 ( .A1(n3513), .A2(n3512), .ZN(n3514) );
  XNOR2_X1 U4423 ( .A(n3527), .B(n3525), .ZN(n3515) );
  NAND2_X1 U4424 ( .A1(n3515), .A2(n4254), .ZN(n3516) );
  INV_X1 U4425 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6301) );
  XNOR2_X1 U4426 ( .A(n3518), .B(n6301), .ZN(n5105) );
  NAND2_X1 U4427 ( .A1(n5104), .A2(n5105), .ZN(n3520) );
  NAND2_X1 U4428 ( .A1(n3518), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3519)
         );
  NAND2_X1 U4429 ( .A1(n3520), .A2(n3519), .ZN(n5170) );
  NOR2_X1 U4430 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  NAND2_X1 U4431 ( .A1(n3525), .A2(n4254), .ZN(n3526) );
  OR2_X1 U4432 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  INV_X1 U4433 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U4434 ( .A1(n5170), .A2(n5171), .ZN(n3531) );
  NAND2_X1 U4435 ( .A1(n3529), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3530)
         );
  INV_X1 U4436 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U4437 ( .A1(n2990), .A2(n5239), .ZN(n3532) );
  INV_X1 U4438 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5238) );
  AND2_X1 U4439 ( .A1(n5989), .A2(n5238), .ZN(n5234) );
  INV_X1 U4440 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U4441 ( .A1(n5989), .A2(n6289), .ZN(n5698) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3533) );
  NOR2_X1 U4443 ( .A1(n2990), .A2(n3533), .ZN(n5690) );
  NAND2_X1 U4444 ( .A1(n5989), .A2(n3533), .ZN(n5688) );
  XNOR2_X1 U4445 ( .A(n5989), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5682)
         );
  INV_X1 U4446 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U4447 ( .A1(n2990), .A2(n5711), .ZN(n3534) );
  INV_X1 U4448 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6041) );
  OR2_X1 U4449 ( .A1(n5989), .A2(n6041), .ZN(n3535) );
  NAND2_X1 U4450 ( .A1(n2990), .A2(n6041), .ZN(n3536) );
  INV_X1 U4451 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U4452 ( .A1(n2990), .A2(n5841), .ZN(n3537) );
  INV_X1 U4453 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U4454 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5714) );
  NOR2_X1 U4455 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5649) );
  INV_X1 U4456 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6007) );
  AND2_X1 U4457 ( .A1(n5649), .A2(n6007), .ZN(n3538) );
  NAND2_X1 U4458 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U4459 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U4460 ( .A1(n5782), .A2(n5719), .ZN(n5727) );
  AND2_X1 U4461 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U4462 ( .A1(n5727), .A2(n5814), .ZN(n3540) );
  NAND2_X1 U4463 ( .A1(n2990), .A2(n3540), .ZN(n3541) );
  NOR2_X1 U4464 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5813) );
  NOR2_X1 U4465 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5783) );
  NOR2_X1 U4466 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5798) );
  NAND3_X1 U4467 ( .A1(n5813), .A2(n5783), .A3(n5798), .ZN(n3542) );
  NAND2_X1 U4468 ( .A1(n5832), .A2(n3542), .ZN(n3543) );
  INV_X1 U4469 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6002) );
  XNOR2_X1 U4470 ( .A(n2990), .B(n6002), .ZN(n5974) );
  NAND2_X1 U4471 ( .A1(n2990), .A2(n6002), .ZN(n3544) );
  AND2_X1 U4472 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5757) );
  INV_X1 U4473 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3546) );
  INV_X1 U4474 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U4475 ( .A1(n3546), .A2(n5349), .ZN(n5755) );
  INV_X1 U4476 ( .A(n5559), .ZN(n3547) );
  NAND2_X1 U4477 ( .A1(n5600), .A2(n3547), .ZN(n5571) );
  NAND2_X1 U4478 ( .A1(n5571), .A2(n3548), .ZN(n3549) );
  NAND2_X1 U4479 ( .A1(n3550), .A2(n3549), .ZN(n3552) );
  NAND2_X1 U4480 ( .A1(n3606), .A2(n2993), .ZN(n3554) );
  NAND2_X1 U4481 ( .A1(n3554), .A2(n3553), .ZN(n3565) );
  INV_X1 U4482 ( .A(n3565), .ZN(n3569) );
  NAND2_X1 U4483 ( .A1(n6455), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3572) );
  NAND2_X1 U4484 ( .A1(n3334), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3555) );
  NAND2_X1 U4485 ( .A1(n3572), .A2(n3555), .ZN(n3571) );
  NAND2_X1 U4486 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n4951), .ZN(n3570) );
  INV_X1 U4487 ( .A(n3570), .ZN(n3556) );
  XNOR2_X1 U4488 ( .A(n3571), .B(n3556), .ZN(n4116) );
  AND2_X1 U4489 ( .A1(n4116), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3564) );
  INV_X1 U4490 ( .A(n3564), .ZN(n3568) );
  OAI21_X1 U4491 ( .B1(n4951), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3570), 
        .ZN(n3557) );
  INV_X1 U4492 ( .A(n3557), .ZN(n3560) );
  AOI21_X1 U4493 ( .B1(n3612), .B2(n3560), .A(n4489), .ZN(n3558) );
  AOI21_X1 U4494 ( .B1(n3237), .B2(n4286), .A(n2993), .ZN(n3585) );
  OR2_X1 U4495 ( .A1(n3558), .A2(n3585), .ZN(n3563) );
  NAND2_X1 U4496 ( .A1(n3560), .A2(n3606), .ZN(n3561) );
  NAND2_X1 U4497 ( .A1(n3600), .A2(n3561), .ZN(n3562) );
  OAI211_X1 U4498 ( .C1(n3565), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3567)
         );
  OR2_X1 U4499 ( .A1(n3600), .A2(n4116), .ZN(n3566) );
  OAI211_X1 U4500 ( .C1(n3569), .C2(n3568), .A(n3567), .B(n3566), .ZN(n3584)
         );
  NAND2_X1 U4501 ( .A1(n3573), .A2(n3572), .ZN(n3578) );
  INV_X1 U4502 ( .A(n3578), .ZN(n3576) );
  NAND2_X1 U4503 ( .A1(n6461), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3588) );
  NAND2_X1 U4504 ( .A1(n5305), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3574) );
  INV_X1 U4505 ( .A(n3577), .ZN(n3575) );
  NAND2_X1 U4506 ( .A1(n3576), .A2(n3575), .ZN(n3579) );
  NAND2_X1 U4507 ( .A1(n3578), .A2(n3577), .ZN(n3589) );
  AND2_X1 U4508 ( .A1(n3579), .A2(n3589), .ZN(n4118) );
  INV_X1 U4509 ( .A(n3580), .ZN(n3597) );
  NAND2_X1 U4510 ( .A1(n3606), .A2(n4118), .ZN(n3582) );
  INV_X1 U4511 ( .A(n3585), .ZN(n3581) );
  OAI211_X1 U4512 ( .C1(n4118), .C2(n3597), .A(n3582), .B(n3581), .ZN(n3583)
         );
  NAND2_X1 U4513 ( .A1(n3584), .A2(n3583), .ZN(n3587) );
  NAND3_X1 U4514 ( .A1(n3585), .A2(n4118), .A3(n3606), .ZN(n3586) );
  NAND2_X1 U4515 ( .A1(n3587), .A2(n3586), .ZN(n3599) );
  NAND2_X1 U4516 ( .A1(n3589), .A2(n3588), .ZN(n3592) );
  XNOR2_X1 U4517 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3591) );
  NAND2_X1 U4518 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3601), .ZN(n3590) );
  NOR2_X1 U4519 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3590), .ZN(n3596)
         );
  NOR2_X1 U4520 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  OR2_X1 U4521 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  NAND2_X1 U4522 ( .A1(n4114), .A2(n3597), .ZN(n3598) );
  NAND2_X1 U4523 ( .A1(n3599), .A2(n3598), .ZN(n3605) );
  AOI22_X1 U4524 ( .A1(n4114), .A2(n3602), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n3053), .ZN(n3604) );
  OAI222_X1 U4525 ( .A1(n6049), .A2(n3601), .B1(n6049), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3601), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4119) );
  AND2_X1 U4526 ( .A1(n4119), .A2(n3602), .ZN(n3603) );
  AOI21_X1 U4527 ( .B1(n3605), .B2(n3604), .A(n3603), .ZN(n3608) );
  AOI21_X1 U4528 ( .B1(n5884), .B2(n4489), .A(n3355), .ZN(n3611) );
  INV_X1 U4529 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5612) );
  INV_X1 U4530 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3985) );
  INV_X1 U4531 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5413) );
  INV_X1 U4532 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5400) );
  XNOR2_X1 U4533 ( .A(n4125), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5334)
         );
  NOR2_X2 U4534 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5872) );
  NAND2_X1 U4535 ( .A1(n6353), .A2(n3615), .ZN(n6591) );
  NAND2_X1 U4536 ( .A1(n6591), .A2(n3053), .ZN(n3616) );
  AND2_X2 U4537 ( .A1(n6060), .A2(n3616), .ZN(n6262) );
  NAND2_X1 U4538 ( .A1(n3053), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3618) );
  NAND2_X1 U4539 ( .A1(n6715), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3617) );
  AND2_X1 U4540 ( .A1(n3618), .A2(n3617), .ZN(n6275) );
  INV_X1 U4541 ( .A(n6262), .ZN(n6276) );
  INV_X1 U4542 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4124) );
  INV_X2 U4543 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U4544 ( .A1(n3053), .A2(n4641), .ZN(n6497) );
  INV_X1 U4545 ( .A(n6497), .ZN(n6507) );
  AND2_X2 U4546 ( .A1(n6045), .A2(n6507), .ZN(n6279) );
  NAND2_X1 U4547 ( .A1(n6279), .A2(REIP_REG_30__SCAN_IN), .ZN(n5740) );
  OAI21_X1 U4548 ( .B1(n6276), .B2(n4124), .A(n5740), .ZN(n3619) );
  AOI21_X1 U4549 ( .B1(n5334), .B2(n5695), .A(n3619), .ZN(n4105) );
  NAND2_X1 U4550 ( .A1(n3620), .A2(n3803), .ZN(n3621) );
  NAND2_X1 U4551 ( .A1(n3001), .A2(n3803), .ZN(n3627) );
  AOI22_X1 U4552 ( .A1(n5310), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4641), .ZN(n3625) );
  AND2_X1 U4553 ( .A1(n3339), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4554 ( .A1(n3630), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3624) );
  AND2_X1 U4555 ( .A1(n3625), .A2(n3624), .ZN(n3626) );
  NAND2_X1 U4556 ( .A1(n3627), .A2(n3626), .ZN(n4301) );
  OR2_X1 U4557 ( .A1(n3629), .A2(n3789), .ZN(n3635) );
  INV_X1 U4558 ( .A(n3630), .ZN(n3653) );
  NAND2_X1 U4559 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n4641), .ZN(n3632)
         );
  NAND2_X1 U4560 ( .A1(n5310), .A2(EAX_REG_0__SCAN_IN), .ZN(n3631) );
  OAI211_X1 U4561 ( .C1(n3653), .C2(n3036), .A(n3632), .B(n3631), .ZN(n3633)
         );
  INV_X1 U4562 ( .A(n3633), .ZN(n3634) );
  NAND2_X1 U4563 ( .A1(n3635), .A2(n3634), .ZN(n4363) );
  NAND2_X1 U4564 ( .A1(n4364), .A2(n4363), .ZN(n4362) );
  INV_X1 U4565 ( .A(n4363), .ZN(n3636) );
  NOR2_X2 U4566 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3657) );
  NAND2_X1 U4567 ( .A1(n3636), .A2(n3657), .ZN(n3637) );
  OAI21_X1 U4568 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3642), .ZN(n6270) );
  AOI22_X1 U4569 ( .A1(n4099), .A2(n6270), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4570 ( .A1(n5310), .A2(EAX_REG_2__SCAN_IN), .ZN(n3638) );
  INV_X1 U4571 ( .A(n3641), .ZN(n3654) );
  INV_X1 U4572 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3643) );
  NAND2_X1 U4573 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  NAND2_X1 U4574 ( .A1(n3654), .A2(n3644), .ZN(n5083) );
  AOI22_X1 U4575 ( .A1(n5083), .A2(n4099), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4576 ( .A1(n5310), .A2(EAX_REG_3__SCAN_IN), .ZN(n3645) );
  OAI211_X1 U4577 ( .C1(n3653), .C2(n3082), .A(n3646), .B(n3645), .ZN(n3647)
         );
  INV_X1 U4578 ( .A(n3647), .ZN(n3648) );
  OAI21_X1 U4579 ( .B1(n3640), .B2(n3789), .A(n3648), .ZN(n4466) );
  NAND2_X1 U4580 ( .A1(n4366), .A2(n4466), .ZN(n4465) );
  INV_X1 U4581 ( .A(n3649), .ZN(n3650) );
  NAND2_X1 U4582 ( .A1(n3650), .A2(n3803), .ZN(n3661) );
  NAND2_X1 U4583 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3652)
         );
  NAND2_X1 U4584 ( .A1(n5310), .A2(EAX_REG_4__SCAN_IN), .ZN(n3651) );
  OAI211_X1 U4585 ( .C1(n3653), .C2(n6049), .A(n3652), .B(n3651), .ZN(n3659)
         );
  INV_X1 U4586 ( .A(n3662), .ZN(n3656) );
  INV_X1 U4587 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U4588 ( .A1(n3654), .A2(n6171), .ZN(n3655) );
  NAND2_X1 U4589 ( .A1(n3656), .A2(n3655), .ZN(n6186) );
  AND2_X1 U4590 ( .A1(n6186), .A2(n3657), .ZN(n3658) );
  AOI21_X1 U4591 ( .B1(n3659), .B2(n4076), .A(n3658), .ZN(n3660) );
  OAI21_X1 U4592 ( .B1(n3662), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3666), 
        .ZN(n6167) );
  AOI22_X1 U4593 ( .A1(n6167), .A2(n3657), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3664) );
  NAND2_X1 U4594 ( .A1(n5310), .A2(EAX_REG_5__SCAN_IN), .ZN(n3663) );
  OAI211_X1 U4595 ( .C1(n3665), .C2(n3789), .A(n3664), .B(n3663), .ZN(n4620)
         );
  NAND2_X1 U4596 ( .A1(n4471), .A2(n4620), .ZN(n4619) );
  INV_X1 U4597 ( .A(n4619), .ZN(n3672) );
  NAND2_X1 U4598 ( .A1(n5310), .A2(EAX_REG_6__SCAN_IN), .ZN(n3668) );
  OAI21_X1 U4599 ( .B1(n6715), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4641), 
        .ZN(n3667) );
  XNOR2_X1 U4600 ( .A(n3666), .B(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5098) );
  AOI22_X1 U4601 ( .A1(n3668), .A2(n3667), .B1(n3657), .B2(n5098), .ZN(n3669)
         );
  NAND2_X1 U4602 ( .A1(n3672), .A2(n3671), .ZN(n4681) );
  INV_X1 U4603 ( .A(n4681), .ZN(n3680) );
  INV_X1 U4604 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3676) );
  OAI21_X1 U4605 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3674), .A(n3673), 
        .ZN(n6149) );
  AOI22_X1 U4606 ( .A1(n3657), .A2(n6149), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3675) );
  OAI21_X1 U4607 ( .B1(n3761), .B2(n3676), .A(n3675), .ZN(n3677) );
  NAND2_X1 U4608 ( .A1(n3680), .A2(n3679), .ZN(n5033) );
  XOR2_X1 U4609 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3681), .Z(n6137) );
  INV_X1 U4610 ( .A(n6137), .ZN(n3696) );
  AOI22_X1 U4611 ( .A1(n3322), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4612 ( .A1(n3316), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4613 ( .A1(n2985), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4614 ( .A1(n4034), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4615 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3691)
         );
  AOI22_X1 U4616 ( .A1(n2989), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4617 ( .A1(n3005), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4618 ( .A1(n3969), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4619 ( .A1(n2987), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4620 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3690)
         );
  NOR2_X1 U4621 ( .A1(n3691), .A2(n3690), .ZN(n3694) );
  NAND2_X1 U4622 ( .A1(n5310), .A2(EAX_REG_8__SCAN_IN), .ZN(n3693) );
  NAND2_X1 U4623 ( .A1(n5309), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3692)
         );
  OAI211_X1 U4624 ( .C1(n3789), .C2(n3694), .A(n3693), .B(n3692), .ZN(n3695)
         );
  AOI21_X1 U4625 ( .B1(n3696), .B2(n3657), .A(n3695), .ZN(n5101) );
  XNOR2_X1 U4626 ( .A(n3698), .B(n5159), .ZN(n5189) );
  AOI22_X1 U4627 ( .A1(n3969), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4628 ( .A1(n2987), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4629 ( .A1(n4079), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4630 ( .A1(n4034), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3699) );
  NAND4_X1 U4631 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n3708)
         );
  AOI22_X1 U4632 ( .A1(n3316), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4633 ( .A1(n3005), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4634 ( .A1(n3270), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4635 ( .A1(n2989), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4636 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3707)
         );
  NOR2_X1 U4637 ( .A1(n3708), .A2(n3707), .ZN(n3711) );
  NAND2_X1 U4638 ( .A1(n5310), .A2(EAX_REG_9__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4639 ( .A1(n5309), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3709)
         );
  OAI211_X1 U4640 ( .C1(n3789), .C2(n3711), .A(n3710), .B(n3709), .ZN(n3712)
         );
  AOI21_X1 U4641 ( .B1(n5189), .B2(n4099), .A(n3712), .ZN(n5155) );
  XOR2_X1 U4642 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3713), .Z(n6122) );
  AOI22_X1 U4643 ( .A1(n3005), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4644 ( .A1(n3270), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4645 ( .A1(n3316), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4646 ( .A1(n3969), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4647 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3723)
         );
  AOI22_X1 U4648 ( .A1(n4079), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4649 ( .A1(n2989), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4650 ( .A1(n4085), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4651 ( .A1(n3269), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3718) );
  NAND4_X1 U4652 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3722)
         );
  OR2_X1 U4653 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  AOI22_X1 U4654 ( .A1(n3803), .A2(n3724), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4655 ( .A1(n5310), .A2(EAX_REG_10__SCAN_IN), .ZN(n3725) );
  OAI211_X1 U4656 ( .C1(n6122), .C2(n4076), .A(n3726), .B(n3725), .ZN(n5195)
         );
  XNOR2_X1 U4657 ( .A(n3727), .B(n5277), .ZN(n5701) );
  NAND2_X1 U4658 ( .A1(n5701), .A2(n3657), .ZN(n3743) );
  AOI22_X1 U4659 ( .A1(n3005), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4660 ( .A1(n4034), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4661 ( .A1(n3316), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4662 ( .A1(n4056), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3728) );
  NAND4_X1 U4663 ( .A1(n3731), .A2(n3730), .A3(n3729), .A4(n3728), .ZN(n3737)
         );
  AOI22_X1 U4664 ( .A1(n4079), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4665 ( .A1(n3270), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4666 ( .A1(n4085), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4667 ( .A1(n2989), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4668 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3736)
         );
  NOR2_X1 U4669 ( .A1(n3737), .A2(n3736), .ZN(n3740) );
  NAND2_X1 U4670 ( .A1(n5310), .A2(EAX_REG_11__SCAN_IN), .ZN(n3739) );
  NAND2_X1 U4671 ( .A1(n5309), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3738)
         );
  OAI211_X1 U4672 ( .C1(n3789), .C2(n3740), .A(n3739), .B(n3738), .ZN(n3741)
         );
  INV_X1 U4673 ( .A(n3741), .ZN(n3742) );
  NAND2_X1 U4674 ( .A1(n3743), .A2(n3742), .ZN(n5266) );
  XOR2_X1 U4675 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3744), .Z(n6114) );
  INV_X1 U4676 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5297) );
  INV_X1 U4677 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5692) );
  OAI22_X1 U4678 ( .A1(n3761), .A2(n5297), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5692), .ZN(n3756) );
  AOI22_X1 U4679 ( .A1(n3969), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4680 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n2989), .B1(n3270), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4681 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4034), .B1(n3269), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4682 ( .A1(n4079), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4683 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3754)
         );
  AOI22_X1 U4684 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n2987), .B1(n4085), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4685 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3317), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4686 ( .A1(n3373), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4687 ( .A1(n4062), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4688 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3753)
         );
  OR2_X1 U4689 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  AOI22_X1 U4690 ( .A1(n3756), .A2(n4076), .B1(n3803), .B2(n3755), .ZN(n3757)
         );
  OAI21_X1 U4691 ( .B1(n6114), .B2(n4076), .A(n3757), .ZN(n5292) );
  XNOR2_X1 U4692 ( .A(n3758), .B(n3759), .ZN(n6100) );
  INV_X1 U4693 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6233) );
  OAI22_X1 U4694 ( .A1(n3761), .A2(n6233), .B1(n3760), .B2(n3759), .ZN(n3762)
         );
  AOI21_X1 U4695 ( .B1(n6100), .B2(n3657), .A(n3762), .ZN(n3774) );
  AOI22_X1 U4696 ( .A1(n3005), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4697 ( .A1(n2989), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4698 ( .A1(n3969), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4699 ( .A1(n3270), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4700 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3772)
         );
  AOI22_X1 U4701 ( .A1(n3316), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4702 ( .A1(n2984), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4703 ( .A1(n3269), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4704 ( .A1(n2987), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4705 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3771)
         );
  OR2_X1 U4706 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  NAND2_X1 U4707 ( .A1(n3803), .A2(n3773), .ZN(n5680) );
  AOI22_X1 U4708 ( .A1(n2989), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4709 ( .A1(n3317), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4710 ( .A1(n3270), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4711 ( .A1(n4085), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4712 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3784)
         );
  AOI22_X1 U4713 ( .A1(n3005), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4714 ( .A1(n4079), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4715 ( .A1(n4056), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4716 ( .A1(n3269), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3779) );
  NAND4_X1 U4717 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  NOR2_X1 U4718 ( .A1(n3784), .A2(n3783), .ZN(n3788) );
  XNOR2_X1 U4719 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3785), .ZN(n5675)
         );
  AOI22_X1 U4720 ( .A1(n4099), .A2(n5675), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U4721 ( .A1(n3623), .A2(EAX_REG_14__SCAN_IN), .ZN(n3786) );
  OAI211_X1 U4722 ( .C1(n3789), .C2(n3788), .A(n3787), .B(n3786), .ZN(n5457)
         );
  XOR2_X1 U4723 ( .A(n3791), .B(n3790), .Z(n5668) );
  AOI22_X1 U4724 ( .A1(n3005), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4725 ( .A1(n3316), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4726 ( .A1(n3269), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4727 ( .A1(n2989), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4728 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3801)
         );
  AOI22_X1 U4729 ( .A1(n4056), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4730 ( .A1(n2985), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4731 ( .A1(n4034), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4732 ( .A1(n4080), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4733 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3800)
         );
  OR2_X1 U4734 ( .A1(n3801), .A2(n3800), .ZN(n3802) );
  AOI22_X1 U4735 ( .A1(n3803), .A2(n3802), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U4736 ( .A1(n3623), .A2(EAX_REG_15__SCAN_IN), .ZN(n3804) );
  OAI211_X1 U4737 ( .C1(n5668), .C2(n4076), .A(n3805), .B(n3804), .ZN(n5446)
         );
  XNOR2_X1 U4738 ( .A(n3806), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6092)
         );
  AOI22_X1 U4739 ( .A1(n4056), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4740 ( .A1(n3317), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4741 ( .A1(n4034), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4742 ( .A1(n2987), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4743 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3816)
         );
  AOI22_X1 U4744 ( .A1(n2984), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4745 ( .A1(n3322), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4746 ( .A1(n3415), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4747 ( .A1(n2989), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4748 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3815)
         );
  NOR2_X1 U4749 ( .A1(n3816), .A2(n3815), .ZN(n3818) );
  AOI22_X1 U4750 ( .A1(n5310), .A2(EAX_REG_16__SCAN_IN), .B1(n5309), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3817) );
  OAI21_X1 U4751 ( .B1(n4073), .B2(n3818), .A(n3817), .ZN(n3819) );
  AOI21_X1 U4752 ( .B1(n6092), .B2(n3657), .A(n3819), .ZN(n5525) );
  AOI22_X1 U4753 ( .A1(n3380), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4754 ( .A1(n3317), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4755 ( .A1(n3270), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4756 ( .A1(n4034), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4757 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4758 ( .A1(n3373), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4759 ( .A1(n4079), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4760 ( .A1(n4056), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4761 ( .A1(n2989), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4762 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4763 ( .A1(n3829), .A2(n3828), .ZN(n3833) );
  NAND2_X1 U4764 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3830)
         );
  NAND2_X1 U4765 ( .A1(n4076), .A2(n3830), .ZN(n3831) );
  AOI21_X1 U4766 ( .B1(n3623), .B2(EAX_REG_17__SCAN_IN), .A(n3831), .ZN(n3832)
         );
  OAI21_X1 U4767 ( .B1(n4073), .B2(n3833), .A(n3832), .ZN(n3836) );
  OAI21_X1 U4768 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3834), .A(n3850), 
        .ZN(n6084) );
  OR2_X1 U4769 ( .A1(n4076), .A2(n6084), .ZN(n3835) );
  NAND2_X1 U4770 ( .A1(n5526), .A2(n5994), .ZN(n5431) );
  INV_X1 U4771 ( .A(n5431), .ZN(n3853) );
  AOI22_X1 U4772 ( .A1(n3373), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4773 ( .A1(n4056), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4774 ( .A1(n4079), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4775 ( .A1(n3380), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4776 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3846)
         );
  AOI22_X1 U4777 ( .A1(n3317), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4778 ( .A1(n3270), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4779 ( .A1(n2989), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4780 ( .A1(n2987), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4781 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3845)
         );
  NOR2_X1 U4782 ( .A1(n3846), .A2(n3845), .ZN(n3849) );
  OAI21_X1 U4783 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5653), .A(n4076), .ZN(
        n3847) );
  AOI21_X1 U4784 ( .B1(n3623), .B2(EAX_REG_18__SCAN_IN), .A(n3847), .ZN(n3848)
         );
  OAI21_X1 U4785 ( .B1(n4073), .B2(n3849), .A(n3848), .ZN(n3852) );
  XNOR2_X1 U4786 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3850), .ZN(n5655)
         );
  NAND2_X1 U4787 ( .A1(n3657), .A2(n5655), .ZN(n3851) );
  NAND2_X1 U4788 ( .A1(n3853), .A2(n3031), .ZN(n5432) );
  AOI22_X1 U4789 ( .A1(n4056), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4790 ( .A1(n2989), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4791 ( .A1(n4079), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4792 ( .A1(n2987), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4793 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3863)
         );
  AOI22_X1 U4794 ( .A1(n3317), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4795 ( .A1(n3373), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4796 ( .A1(n4034), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4797 ( .A1(n3269), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4798 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3862)
         );
  NOR2_X1 U4799 ( .A1(n3863), .A2(n3862), .ZN(n3867) );
  NAND2_X1 U4800 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3864)
         );
  NAND2_X1 U4801 ( .A1(n4076), .A2(n3864), .ZN(n3865) );
  AOI21_X1 U4802 ( .B1(n3623), .B2(EAX_REG_19__SCAN_IN), .A(n3865), .ZN(n3866)
         );
  OAI21_X1 U4803 ( .B1(n4073), .B2(n3867), .A(n3866), .ZN(n3870) );
  OAI21_X1 U4804 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3868), .A(n3885), 
        .ZN(n5986) );
  OR2_X1 U4805 ( .A1(n4076), .A2(n5986), .ZN(n3869) );
  NAND2_X1 U4806 ( .A1(n3870), .A2(n3869), .ZN(n5511) );
  AOI22_X1 U4807 ( .A1(n3322), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4808 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3317), .B1(n2985), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4809 ( .A1(n4034), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4810 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3380), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4811 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3880)
         );
  AOI22_X1 U4812 ( .A1(n2989), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4813 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4079), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4814 ( .A1(n3005), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4815 ( .A1(n4056), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4816 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3879)
         );
  NOR2_X1 U4817 ( .A1(n3880), .A2(n3879), .ZN(n3884) );
  NAND2_X1 U4818 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3881)
         );
  NAND2_X1 U4819 ( .A1(n4076), .A2(n3881), .ZN(n3882) );
  AOI21_X1 U4820 ( .B1(n3623), .B2(EAX_REG_20__SCAN_IN), .A(n3882), .ZN(n3883)
         );
  OAI21_X1 U4821 ( .B1(n4073), .B2(n3884), .A(n3883), .ZN(n3887) );
  XNOR2_X1 U4822 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3885), .ZN(n5944)
         );
  NAND2_X1 U4823 ( .A1(n3657), .A2(n5944), .ZN(n3886) );
  NAND2_X1 U4824 ( .A1(n3887), .A2(n3886), .ZN(n5504) );
  AOI22_X1 U4825 ( .A1(n3005), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4826 ( .A1(n2987), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4827 ( .A1(n4079), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4828 ( .A1(n4056), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4829 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4830 ( .A1(n3317), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4831 ( .A1(n3415), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4832 ( .A1(n2989), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4833 ( .A1(n4034), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4834 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  NOR2_X1 U4835 ( .A1(n3898), .A2(n3897), .ZN(n3902) );
  OAI21_X1 U4836 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6715), .A(n4641), 
        .ZN(n3899) );
  INV_X1 U4837 ( .A(n3899), .ZN(n3900) );
  AOI21_X1 U4838 ( .B1(n3623), .B2(EAX_REG_21__SCAN_IN), .A(n3900), .ZN(n3901)
         );
  OAI21_X1 U4839 ( .B1(n4073), .B2(n3902), .A(n3901), .ZN(n3905) );
  OAI21_X1 U4840 ( .B1(n3903), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3919), 
        .ZN(n5943) );
  OR2_X1 U4841 ( .A1(n5943), .A2(n4076), .ZN(n3904) );
  AOI22_X1 U4842 ( .A1(n3005), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4843 ( .A1(n2989), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4844 ( .A1(n4056), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4845 ( .A1(n3415), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4846 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3915)
         );
  AOI22_X1 U4847 ( .A1(n3317), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4848 ( .A1(n2985), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4849 ( .A1(n3269), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4850 ( .A1(n2987), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4851 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  NOR2_X1 U4852 ( .A1(n3915), .A2(n3914), .ZN(n3918) );
  AOI21_X1 U4853 ( .B1(n5631), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3916) );
  AOI21_X1 U4854 ( .B1(n3623), .B2(EAX_REG_22__SCAN_IN), .A(n3916), .ZN(n3917)
         );
  OAI21_X1 U4855 ( .B1(n4073), .B2(n3918), .A(n3917), .ZN(n3921) );
  XNOR2_X1 U4856 ( .A(n3919), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5929)
         );
  NAND2_X1 U4857 ( .A1(n5929), .A2(n3657), .ZN(n3920) );
  NAND2_X1 U4858 ( .A1(n3921), .A2(n3920), .ZN(n5501) );
  AOI22_X1 U4859 ( .A1(n3373), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4860 ( .A1(n4056), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4861 ( .A1(n4085), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4862 ( .A1(n4086), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4863 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3931)
         );
  AOI22_X1 U4864 ( .A1(n2989), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4865 ( .A1(n3317), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4866 ( .A1(n2987), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4867 ( .A1(n3415), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4868 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  NOR2_X1 U4869 ( .A1(n3931), .A2(n3930), .ZN(n3951) );
  AOI22_X1 U4870 ( .A1(n3969), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4871 ( .A1(n2984), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4872 ( .A1(n3322), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4873 ( .A1(n2987), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4874 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3941)
         );
  AOI22_X1 U4875 ( .A1(n3317), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4876 ( .A1(n3005), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4877 ( .A1(n2989), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4878 ( .A1(n3380), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4879 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3940)
         );
  NOR2_X1 U4880 ( .A1(n3941), .A2(n3940), .ZN(n3952) );
  XNOR2_X1 U4881 ( .A(n3951), .B(n3952), .ZN(n3945) );
  NAND2_X1 U4882 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3942)
         );
  NAND2_X1 U4883 ( .A1(n4076), .A2(n3942), .ZN(n3943) );
  AOI21_X1 U4884 ( .B1(n5310), .B2(EAX_REG_23__SCAN_IN), .A(n3943), .ZN(n3944)
         );
  OAI21_X1 U4885 ( .B1(n4073), .B2(n3945), .A(n3944), .ZN(n3949) );
  OR2_X1 U4886 ( .A1(n3946), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3947)
         );
  NAND2_X1 U4887 ( .A1(n3963), .A2(n3947), .ZN(n5623) );
  NAND2_X1 U4888 ( .A1(n3949), .A2(n3948), .ZN(n4107) );
  OR2_X1 U4889 ( .A1(n3952), .A2(n3951), .ZN(n3981) );
  AOI22_X1 U4890 ( .A1(n2987), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4891 ( .A1(n3317), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4892 ( .A1(n3005), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4893 ( .A1(n4085), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4894 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3962)
         );
  AOI22_X1 U4895 ( .A1(n4079), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4896 ( .A1(n3270), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4897 ( .A1(n4056), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4898 ( .A1(n2989), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4899 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3961)
         );
  NOR2_X1 U4900 ( .A1(n3962), .A2(n3961), .ZN(n3980) );
  XNOR2_X1 U4901 ( .A(n3981), .B(n3980), .ZN(n3968) );
  XNOR2_X1 U4902 ( .A(n3963), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5915)
         );
  NAND2_X1 U4903 ( .A1(n5310), .A2(EAX_REG_24__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U4904 ( .A1(n5309), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3964)
         );
  OAI211_X1 U4905 ( .C1(n5915), .C2(n4076), .A(n3965), .B(n3964), .ZN(n3966)
         );
  INV_X1 U4906 ( .A(n3966), .ZN(n3967) );
  OAI21_X1 U4907 ( .B1(n3968), .B2(n4073), .A(n3967), .ZN(n5487) );
  AOI22_X1 U4908 ( .A1(n3373), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4909 ( .A1(n3969), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4910 ( .A1(n2989), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4911 ( .A1(n3317), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4912 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3979)
         );
  AOI22_X1 U4913 ( .A1(n2987), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4914 ( .A1(n4079), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2985), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4915 ( .A1(n4062), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4916 ( .A1(n3269), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4917 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  NOR2_X1 U4918 ( .A1(n3979), .A2(n3978), .ZN(n3992) );
  OR2_X1 U4919 ( .A1(n3981), .A2(n3980), .ZN(n3991) );
  XNOR2_X1 U4920 ( .A(n3992), .B(n3991), .ZN(n3984) );
  OAI21_X1 U4921 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3985), .A(n4076), .ZN(
        n3982) );
  AOI21_X1 U4922 ( .B1(n3623), .B2(EAX_REG_25__SCAN_IN), .A(n3982), .ZN(n3983)
         );
  OAI21_X1 U4923 ( .B1(n3984), .B2(n4073), .A(n3983), .ZN(n3990) );
  AND2_X1 U4924 ( .A1(n3986), .A2(n3985), .ZN(n3987) );
  OR2_X1 U4925 ( .A1(n3987), .A2(n4007), .ZN(n5981) );
  INV_X1 U4926 ( .A(n5981), .ZN(n3988) );
  NAND2_X1 U4927 ( .A1(n3988), .A2(n3657), .ZN(n3989) );
  NOR2_X1 U4928 ( .A1(n3992), .A2(n3991), .ZN(n4021) );
  AOI22_X1 U4929 ( .A1(n3005), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4930 ( .A1(n2989), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4931 ( .A1(n4056), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4932 ( .A1(n3415), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4933 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4002)
         );
  AOI22_X1 U4934 ( .A1(n3317), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4935 ( .A1(n2985), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4936 ( .A1(n3269), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4937 ( .A1(n2987), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4938 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  OR2_X1 U4939 ( .A1(n4002), .A2(n4001), .ZN(n4020) );
  XNOR2_X1 U4940 ( .A(n4021), .B(n4020), .ZN(n4005) );
  INV_X1 U4941 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4006) );
  AOI21_X1 U4942 ( .B1(n4006), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4003) );
  AOI21_X1 U4943 ( .B1(n3623), .B2(EAX_REG_26__SCAN_IN), .A(n4003), .ZN(n4004)
         );
  OAI21_X1 U4944 ( .B1(n4005), .B2(n4073), .A(n4004), .ZN(n4009) );
  XNOR2_X1 U4945 ( .A(n4007), .B(n4006), .ZN(n5900) );
  NAND2_X1 U4946 ( .A1(n5900), .A2(n3657), .ZN(n4008) );
  AOI22_X1 U4947 ( .A1(n2989), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4948 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4079), .B1(n4085), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4949 ( .A1(n3373), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4950 ( .A1(n4056), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4951 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U4952 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3270), .B1(n3374), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4953 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3317), .B1(n2999), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4954 ( .A1(n4086), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4955 ( .A1(n2987), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4956 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  NOR2_X1 U4957 ( .A1(n4019), .A2(n4018), .ZN(n4033) );
  NAND2_X1 U4958 ( .A1(n4021), .A2(n4020), .ZN(n4032) );
  XNOR2_X1 U4959 ( .A(n4033), .B(n4032), .ZN(n4025) );
  NAND2_X1 U4960 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4022)
         );
  NAND2_X1 U4961 ( .A1(n4076), .A2(n4022), .ZN(n4023) );
  AOI21_X1 U4962 ( .B1(n5310), .B2(EAX_REG_27__SCAN_IN), .A(n4023), .ZN(n4024)
         );
  OAI21_X1 U4963 ( .B1(n4025), .B2(n4073), .A(n4024), .ZN(n4031) );
  INV_X1 U4964 ( .A(n4026), .ZN(n4028) );
  INV_X1 U4965 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4027) );
  NAND2_X1 U4966 ( .A1(n4028), .A2(n4027), .ZN(n4029) );
  NAND2_X1 U4967 ( .A1(n4050), .A2(n4029), .ZN(n5594) );
  NOR2_X1 U4968 ( .A1(n4033), .A2(n4032), .ZN(n4070) );
  AOI22_X1 U4969 ( .A1(n3373), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4970 ( .A1(n2989), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4971 ( .A1(n4056), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4972 ( .A1(n3415), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U4973 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4045)
         );
  AOI22_X1 U4974 ( .A1(n3317), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4975 ( .A1(n2984), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4976 ( .A1(n3269), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4977 ( .A1(n2987), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U4978 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  OR2_X1 U4979 ( .A1(n4045), .A2(n4044), .ZN(n4069) );
  INV_X1 U4980 ( .A(n4069), .ZN(n4046) );
  XNOR2_X1 U4981 ( .A(n4070), .B(n4046), .ZN(n4047) );
  INV_X1 U4982 ( .A(n4073), .ZN(n4096) );
  NAND2_X1 U4983 ( .A1(n4047), .A2(n4096), .ZN(n4053) );
  NAND2_X1 U4984 ( .A1(n4641), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U4985 ( .A1(n4076), .A2(n4048), .ZN(n4049) );
  AOI21_X1 U4986 ( .B1(n5310), .B2(EAX_REG_28__SCAN_IN), .A(n4049), .ZN(n4052)
         );
  XNOR2_X1 U4987 ( .A(n4050), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5412)
         );
  NAND2_X1 U4988 ( .A1(n4054), .A2(n5400), .ZN(n4055) );
  NAND2_X1 U4989 ( .A1(n4125), .A2(n4055), .ZN(n5575) );
  AOI22_X1 U4990 ( .A1(n4056), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4991 ( .A1(n3317), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U4992 ( .A1(n2989), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4993 ( .A1(n3380), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4057) );
  NAND4_X1 U4994 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4068)
         );
  AOI22_X1 U4995 ( .A1(n4086), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4996 ( .A1(n4079), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4997 ( .A1(n3005), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U4998 ( .A1(n3270), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U4999 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NOR2_X1 U5000 ( .A1(n4068), .A2(n4067), .ZN(n4078) );
  NAND2_X1 U5001 ( .A1(n4070), .A2(n4069), .ZN(n4077) );
  XNOR2_X1 U5002 ( .A(n4078), .B(n4077), .ZN(n4074) );
  AOI21_X1 U5003 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n4641), .A(n3657), 
        .ZN(n4072) );
  NAND2_X1 U5004 ( .A1(n5310), .A2(EAX_REG_29__SCAN_IN), .ZN(n4071) );
  OAI211_X1 U5005 ( .C1(n4074), .C2(n4073), .A(n4072), .B(n4071), .ZN(n4075)
         );
  OAI21_X1 U5006 ( .B1(n4076), .B2(n5575), .A(n4075), .ZN(n5391) );
  NOR2_X1 U5007 ( .A1(n4078), .A2(n4077), .ZN(n4095) );
  AOI22_X1 U5008 ( .A1(n3969), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5009 ( .A1(n3317), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5010 ( .A1(n2989), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5011 ( .A1(n2987), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4080), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4081) );
  NAND4_X1 U5012 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4093)
         );
  AOI22_X1 U5013 ( .A1(n2999), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5014 ( .A1(n3374), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5015 ( .A1(n4086), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5016 ( .A1(n3269), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5017 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  NOR2_X1 U5018 ( .A1(n4093), .A2(n4092), .ZN(n4094) );
  XNOR2_X1 U5019 ( .A(n4095), .B(n4094), .ZN(n4097) );
  NAND2_X1 U5020 ( .A1(n4097), .A2(n4096), .ZN(n4102) );
  AOI21_X1 U5021 ( .B1(n4124), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4098) );
  AOI21_X1 U5022 ( .B1(n5310), .B2(EAX_REG_30__SCAN_IN), .A(n4098), .ZN(n4101)
         );
  NAND3_X1 U5023 ( .A1(n3053), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6505) );
  INV_X1 U5024 ( .A(n6505), .ZN(n4103) );
  OAI211_X1 U5025 ( .C1(n5746), .C2(n6060), .A(n4105), .B(n4104), .ZN(U2956)
         );
  INV_X1 U5026 ( .A(n4106), .ZN(n5500) );
  AND2_X1 U5027 ( .A1(n5500), .A2(n4107), .ZN(n4109) );
  OR2_X1 U5028 ( .A1(n4109), .A2(n4108), .ZN(n5621) );
  AND2_X1 U5029 ( .A1(n4111), .A2(n4489), .ZN(n4113) );
  NAND2_X1 U5030 ( .A1(n4113), .A2(n4112), .ZN(n6468) );
  INV_X1 U5031 ( .A(n4114), .ZN(n4115) );
  NAND2_X1 U5032 ( .A1(n4118), .A2(n4117), .ZN(n4121) );
  INV_X1 U5033 ( .A(n4119), .ZN(n4120) );
  NAND2_X1 U5034 ( .A1(n4121), .A2(n4120), .ZN(n6467) );
  NOR2_X1 U5035 ( .A1(n6468), .A2(n6467), .ZN(n6053) );
  NAND2_X1 U5036 ( .A1(n6053), .A2(n4374), .ZN(n4226) );
  NOR2_X1 U5037 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6595) );
  NOR3_X1 U5038 ( .A1(n3053), .A2(n6580), .A3(n6504), .ZN(n6490) );
  NOR3_X1 U5039 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6497), .A3(n5321), .ZN(
        n6500) );
  OR2_X1 U5040 ( .A1(n6279), .A2(n6500), .ZN(n4122) );
  OR2_X1 U5041 ( .A1(n6490), .A2(n4122), .ZN(n4123) );
  NOR2_X1 U5042 ( .A1(n5567), .A2(n5321), .ZN(n4127) );
  NOR2_X1 U5043 ( .A1(n5621), .A2(n6150), .ZN(n4221) );
  NAND2_X1 U5044 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n4131) );
  NAND2_X1 U5045 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5952) );
  OR2_X1 U5046 ( .A1(n4128), .A2(STATE_REG_0__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U5047 ( .A1(n4496), .A2(n6514), .ZN(n4250) );
  INV_X1 U5048 ( .A(READY_N), .ZN(n6485) );
  NAND2_X1 U5049 ( .A1(n6715), .A2(n6485), .ZN(n4214) );
  INV_X1 U5050 ( .A(n4214), .ZN(n4213) );
  AND3_X1 U5051 ( .A1(n4250), .A2(n4213), .A3(n4286), .ZN(n4129) );
  INV_X1 U5052 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6075) );
  INV_X1 U5053 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6549) );
  INV_X1 U5054 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6544) );
  INV_X1 U5055 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6542) );
  INV_X1 U5056 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6532) );
  NAND3_X1 U5057 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6175) );
  INV_X1 U5058 ( .A(n6175), .ZN(n4130) );
  NAND2_X1 U5059 ( .A1(REIP_REG_4__SCAN_IN), .A2(n4130), .ZN(n4736) );
  NOR2_X1 U5060 ( .A1(n6532), .A2(n4736), .ZN(n4731) );
  NAND4_X1 U5061 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(n4731), .ZN(n5163) );
  INV_X1 U5062 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5276) );
  INV_X1 U5063 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6540) );
  INV_X1 U5064 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6537) );
  NOR3_X1 U5065 ( .A1(n5276), .A2(n6540), .A3(n6537), .ZN(n5274) );
  INV_X1 U5066 ( .A(n5274), .ZN(n6102) );
  NOR4_X1 U5067 ( .A1(n6544), .A2(n6542), .A3(n5163), .A4(n6102), .ZN(n5462)
         );
  NAND2_X1 U5068 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5462), .ZN(n5448) );
  NOR2_X1 U5069 ( .A1(n6549), .A2(n5448), .ZN(n6087) );
  NAND2_X1 U5070 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6087), .ZN(n6076) );
  NOR2_X1 U5071 ( .A1(n6075), .A2(n6076), .ZN(n4132) );
  NAND2_X1 U5072 ( .A1(n6188), .A2(n4132), .ZN(n5954) );
  NOR2_X1 U5073 ( .A1(n5952), .A2(n5954), .ZN(n5947) );
  NAND2_X1 U5074 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5947), .ZN(n5927) );
  INV_X1 U5075 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6560) );
  OAI21_X1 U5076 ( .B1(n4131), .B2(n5927), .A(n6560), .ZN(n4133) );
  NAND2_X1 U5077 ( .A1(n6077), .A2(n5447), .ZN(n5925) );
  AND2_X1 U5078 ( .A1(n5447), .A2(n4132), .ZN(n5437) );
  NAND4_X1 U5079 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5437), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5924) );
  NAND3_X1 U5080 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5328) );
  NOR2_X1 U5081 ( .A1(n5924), .A2(n5328), .ZN(n5330) );
  NOR2_X1 U5082 ( .A1(n5438), .A2(n5330), .ZN(n5916) );
  AND2_X1 U5083 ( .A1(n4133), .A2(n5916), .ZN(n4220) );
  INV_X1 U5084 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4135) );
  OAI22_X1 U5085 ( .A1(n4135), .A2(n6170), .B1(n5623), .B2(n6201), .ZN(n4219)
         );
  NOR2_X4 U5086 ( .A1(n3000), .A2(n2996), .ZN(n5372) );
  INV_X1 U5087 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4136) );
  NAND2_X1 U5088 ( .A1(n5372), .A2(n4136), .ZN(n4139) );
  INV_X1 U5089 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U5090 ( .A1(n4168), .A2(n5300), .ZN(n4137) );
  OAI211_X1 U5091 ( .C1(n2997), .C2(EBX_REG_1__SCAN_IN), .A(n4137), .B(n5505), 
        .ZN(n4138) );
  NAND2_X1 U5092 ( .A1(n4168), .A2(EBX_REG_0__SCAN_IN), .ZN(n4141) );
  INV_X1 U5093 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5094 ( .A1(n5505), .A2(n4365), .ZN(n4140) );
  NAND2_X1 U5095 ( .A1(n4141), .A2(n4140), .ZN(n4360) );
  INV_X1 U5096 ( .A(n4168), .ZN(n4142) );
  NAND2_X1 U5097 ( .A1(n4142), .A2(n2998), .ZN(n4203) );
  NAND2_X1 U5098 ( .A1(n2998), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4143)
         );
  AND2_X1 U5099 ( .A1(n4203), .A2(n4143), .ZN(n4144) );
  MUX2_X1 U5100 ( .A(n5345), .B(n5392), .S(EBX_REG_3__SCAN_IN), .Z(n4146) );
  OR2_X1 U5101 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4145)
         );
  AND2_X1 U5102 ( .A1(n4146), .A2(n4145), .ZN(n4467) );
  NAND2_X1 U5103 ( .A1(n4468), .A2(n4467), .ZN(n4475) );
  INV_X1 U5104 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4147) );
  NAND2_X1 U5105 ( .A1(n5372), .A2(n4147), .ZN(n4151) );
  NAND2_X1 U5106 ( .A1(n4168), .A2(n4148), .ZN(n4149) );
  OAI211_X1 U5107 ( .C1(n2997), .C2(EBX_REG_4__SCAN_IN), .A(n4149), .B(n5392), 
        .ZN(n4150) );
  MUX2_X1 U5108 ( .A(n5345), .B(n5392), .S(EBX_REG_5__SCAN_IN), .Z(n4153) );
  OAI21_X1 U5109 ( .B1(n5369), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4153), 
        .ZN(n4623) );
  INV_X1 U5110 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U5111 ( .A1(n5372), .A2(n4734), .ZN(n4157) );
  NAND2_X1 U5112 ( .A1(n4168), .A2(n4154), .ZN(n4155) );
  OAI211_X1 U5113 ( .C1(n2998), .C2(EBX_REG_6__SCAN_IN), .A(n4155), .B(n5392), 
        .ZN(n4156) );
  MUX2_X1 U5114 ( .A(n5345), .B(n5392), .S(EBX_REG_7__SCAN_IN), .Z(n4158) );
  OAI21_X1 U5115 ( .B1(n5369), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4158), 
        .ZN(n5037) );
  NOR2_X4 U5116 ( .A1(n5036), .A2(n5037), .ZN(n5151) );
  INV_X1 U5117 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U5118 ( .A1(n5372), .A2(n6135), .ZN(n4162) );
  NAND2_X1 U5119 ( .A1(n4168), .A2(n4159), .ZN(n4160) );
  OAI211_X1 U5120 ( .C1(n2998), .C2(EBX_REG_8__SCAN_IN), .A(n4160), .B(n5392), 
        .ZN(n4161) );
  NAND2_X1 U5121 ( .A1(n4162), .A2(n4161), .ZN(n5150) );
  MUX2_X1 U5122 ( .A(n5345), .B(n5392), .S(EBX_REG_9__SCAN_IN), .Z(n4164) );
  OR2_X1 U5123 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4163)
         );
  NAND2_X1 U5124 ( .A1(n4164), .A2(n4163), .ZN(n5160) );
  MUX2_X1 U5125 ( .A(n5336), .B(n4168), .S(EBX_REG_10__SCAN_IN), .Z(n4167) );
  NAND2_X1 U5126 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n2997), .ZN(n4165) );
  AND2_X1 U5127 ( .A1(n4203), .A2(n4165), .ZN(n4166) );
  OR2_X1 U5128 ( .A1(n5345), .A2(EBX_REG_11__SCAN_IN), .ZN(n4171) );
  NAND2_X1 U5129 ( .A1(n5392), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4169) );
  OAI211_X1 U5130 ( .C1(n2997), .C2(EBX_REG_11__SCAN_IN), .A(n4168), .B(n4169), 
        .ZN(n4170) );
  MUX2_X1 U5131 ( .A(n5336), .B(n4168), .S(EBX_REG_12__SCAN_IN), .Z(n4174) );
  NAND2_X1 U5132 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n2998), .ZN(n4172) );
  AND2_X1 U5133 ( .A1(n4203), .A2(n4172), .ZN(n4173) );
  NAND2_X1 U5134 ( .A1(n4174), .A2(n4173), .ZN(n5293) );
  OR2_X1 U5135 ( .A1(n5345), .A2(EBX_REG_13__SCAN_IN), .ZN(n4177) );
  NAND2_X1 U5136 ( .A1(n5392), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4175) );
  OAI211_X1 U5137 ( .C1(n2997), .C2(EBX_REG_13__SCAN_IN), .A(n4168), .B(n4175), 
        .ZN(n4176) );
  NAND2_X1 U5138 ( .A1(n4177), .A2(n4176), .ZN(n5860) );
  MUX2_X1 U5139 ( .A(n5336), .B(n4168), .S(EBX_REG_14__SCAN_IN), .Z(n4180) );
  NAND2_X1 U5140 ( .A1(n2998), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4178) );
  AND2_X1 U5141 ( .A1(n4203), .A2(n4178), .ZN(n4179) );
  OR2_X1 U5142 ( .A1(n5345), .A2(EBX_REG_15__SCAN_IN), .ZN(n4183) );
  NAND2_X1 U5143 ( .A1(n5392), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4181) );
  OAI211_X1 U5144 ( .C1(n2997), .C2(EBX_REG_15__SCAN_IN), .A(n4168), .B(n4181), 
        .ZN(n4182) );
  MUX2_X1 U5145 ( .A(n5336), .B(n4168), .S(EBX_REG_16__SCAN_IN), .Z(n4186) );
  NAND2_X1 U5146 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n2998), .ZN(n4184) );
  AND2_X1 U5147 ( .A1(n4203), .A2(n4184), .ZN(n4185) );
  NAND2_X1 U5148 ( .A1(n4186), .A2(n4185), .ZN(n5522) );
  OR2_X1 U5149 ( .A1(n5345), .A2(EBX_REG_17__SCAN_IN), .ZN(n4189) );
  NAND2_X1 U5150 ( .A1(n5392), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4187) );
  OAI211_X1 U5151 ( .C1(n2997), .C2(EBX_REG_17__SCAN_IN), .A(n4168), .B(n4187), 
        .ZN(n4188) );
  NAND2_X1 U5152 ( .A1(n4189), .A2(n4188), .ZN(n6017) );
  INV_X1 U5153 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U5154 ( .A1(n5372), .A2(n5961), .ZN(n4192) );
  INV_X1 U5155 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U5156 ( .A1(n4168), .A2(n5839), .ZN(n4190) );
  OAI211_X1 U5157 ( .C1(n2997), .C2(EBX_REG_19__SCAN_IN), .A(n4190), .B(n5392), 
        .ZN(n4191) );
  OR2_X1 U5158 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4195)
         );
  INV_X1 U5159 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4193) );
  NAND2_X1 U5160 ( .A1(n4307), .A2(n4193), .ZN(n4194) );
  AND2_X1 U5161 ( .A1(n4195), .A2(n4194), .ZN(n5507) );
  OR2_X1 U5162 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4197)
         );
  OR2_X1 U5163 ( .A1(n2998), .A2(EBX_REG_18__SCAN_IN), .ZN(n4196) );
  NAND2_X1 U5164 ( .A1(n4197), .A2(n4196), .ZN(n5506) );
  NAND2_X1 U5165 ( .A1(n5506), .A2(n5392), .ZN(n5434) );
  NAND2_X1 U5166 ( .A1(n3097), .A2(EBX_REG_20__SCAN_IN), .ZN(n4198) );
  OAI211_X1 U5167 ( .C1(n5507), .C2(n5506), .A(n5434), .B(n4198), .ZN(n4199)
         );
  MUX2_X1 U5168 ( .A(n5345), .B(n5392), .S(EBX_REG_21__SCAN_IN), .Z(n4201) );
  OR2_X1 U5169 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4200)
         );
  MUX2_X1 U5170 ( .A(n5336), .B(n4168), .S(EBX_REG_22__SCAN_IN), .Z(n4205) );
  NAND2_X1 U5171 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n2998), .ZN(n4202) );
  AND2_X1 U5172 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  OR2_X1 U5173 ( .A1(n5345), .A2(EBX_REG_23__SCAN_IN), .ZN(n4208) );
  NAND2_X1 U5174 ( .A1(n5392), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4206) );
  OAI211_X1 U5175 ( .C1(n2998), .C2(EBX_REG_23__SCAN_IN), .A(n4168), .B(n4206), 
        .ZN(n4207) );
  NAND2_X1 U5176 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  NOR2_X2 U5177 ( .A1(n5498), .A2(n4209), .ZN(n5339) );
  INV_X1 U5178 ( .A(n5339), .ZN(n5490) );
  NAND2_X1 U5179 ( .A1(n5498), .A2(n4209), .ZN(n4210) );
  NAND2_X1 U5180 ( .A1(n5490), .A2(n4210), .ZN(n5789) );
  NAND2_X1 U5181 ( .A1(n4214), .A2(EBX_REG_31__SCAN_IN), .ZN(n4211) );
  NOR2_X1 U5182 ( .A1(n2997), .A2(n4211), .ZN(n4212) );
  INV_X1 U5183 ( .A(n6514), .ZN(n4416) );
  NAND2_X1 U5184 ( .A1(n4416), .A2(n4213), .ZN(n6489) );
  AND2_X1 U5185 ( .A1(n4254), .A2(n6489), .ZN(n5379) );
  INV_X1 U5186 ( .A(n5379), .ZN(n4216) );
  INV_X1 U5187 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5469) );
  NAND3_X1 U5188 ( .A1(n4286), .A2(n5469), .A3(n4214), .ZN(n4215) );
  NAND2_X1 U5189 ( .A1(n4216), .A2(n4215), .ZN(n4217) );
  INV_X1 U5190 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5494) );
  OAI22_X1 U5191 ( .A1(n5789), .A2(n6196), .B1(n6134), .B2(n5494), .ZN(n4218)
         );
  OR4_X1 U5192 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(U2804) );
  INV_X1 U5193 ( .A(n6590), .ZN(n4223) );
  NAND2_X1 U5194 ( .A1(n4489), .A2(n2993), .ZN(n5060) );
  NAND2_X1 U5195 ( .A1(n6594), .A2(n5060), .ZN(n6058) );
  AND2_X1 U5196 ( .A1(n5872), .A2(n5321), .ZN(n4225) );
  OAI21_X1 U5197 ( .B1(n4225), .B2(READREQUEST_REG_SCAN_IN), .A(n4223), .ZN(
        n4222) );
  OAI21_X1 U5198 ( .B1(n4223), .B2(n6058), .A(n4222), .ZN(U3474) );
  INV_X1 U5199 ( .A(n4224), .ZN(n4228) );
  AOI211_X1 U5200 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4226), .A(n4225), .B(
        n4228), .ZN(n4227) );
  INV_X1 U5201 ( .A(n4227), .ZN(U2788) );
  NAND3_X1 U5202 ( .A1(n4232), .A2(n4496), .A3(n6465), .ZN(n4351) );
  NAND2_X1 U5203 ( .A1(n4299), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4233) );
  INV_X1 U5204 ( .A(n4417), .ZN(n4229) );
  NOR2_X1 U5205 ( .A1(n4418), .A2(READY_N), .ZN(n4231) );
  NAND2_X1 U5206 ( .A1(n4341), .A2(DATAI_13_), .ZN(n4320) );
  OAI211_X1 U5207 ( .C1(n4351), .C2(n6233), .A(n4233), .B(n4320), .ZN(U2952)
         );
  INV_X1 U5208 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5209 ( .A1(n4299), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U5210 ( .A1(n4341), .A2(DATAI_2_), .ZN(n4357) );
  OAI211_X1 U5211 ( .C1(n4396), .C2(n4351), .A(n4234), .B(n4357), .ZN(U2926)
         );
  INV_X1 U5212 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5213 ( .A1(n4299), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U5214 ( .A1(n4341), .A2(DATAI_3_), .ZN(n4347) );
  OAI211_X1 U5215 ( .C1(n4390), .C2(n4351), .A(n4235), .B(n4347), .ZN(U2927)
         );
  INV_X1 U5216 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U5217 ( .A1(n4299), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4236) );
  NAND2_X1 U5218 ( .A1(n4341), .A2(DATAI_1_), .ZN(n4354) );
  OAI211_X1 U5219 ( .C1(n4388), .C2(n4351), .A(n4236), .B(n4354), .ZN(U2925)
         );
  INV_X1 U5220 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4237) );
  INV_X1 U5221 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6229) );
  OAI222_X1 U5222 ( .A1(n6740), .A2(n4376), .B1(n4237), .B2(n4313), .C1(n4351), 
        .C2(n6229), .ZN(U2954) );
  INV_X1 U5223 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4346) );
  NOR2_X1 U5224 ( .A1(n6468), .A2(n4496), .ZN(n5324) );
  OR2_X1 U5225 ( .A1(n4229), .A2(n6594), .ZN(n6488) );
  INV_X1 U5226 ( .A(n6488), .ZN(n4238) );
  OAI21_X1 U5227 ( .B1(n5324), .B2(n4238), .A(n4416), .ZN(n4239) );
  NAND2_X1 U5228 ( .A1(n6227), .A2(n4286), .ZN(n4402) );
  NAND2_X1 U5229 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4453) );
  NOR2_X1 U5230 ( .A1(n4453), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6239) );
  INV_X1 U5231 ( .A(n6239), .ZN(n6484) );
  AOI22_X1 U5232 ( .A1(n6592), .A2(UWORD_REG_9__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4240) );
  OAI21_X1 U5233 ( .B1(n4346), .B2(n4402), .A(n4240), .ZN(U2898) );
  INV_X1 U5234 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U5235 ( .A1(n6592), .A2(UWORD_REG_10__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4241) );
  OAI21_X1 U5236 ( .B1(n4328), .B2(n4402), .A(n4241), .ZN(U2897) );
  INV_X1 U5237 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U5238 ( .A1(n6592), .A2(UWORD_REG_8__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4242) );
  OAI21_X1 U5239 ( .B1(n4343), .B2(n4402), .A(n4242), .ZN(U2899) );
  INV_X1 U5240 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U5241 ( .A1(n6592), .A2(UWORD_REG_12__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4243) );
  OAI21_X1 U5242 ( .B1(n4316), .B2(n4402), .A(n4243), .ZN(U2895) );
  INV_X1 U5243 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U5244 ( .A1(n6592), .A2(UWORD_REG_13__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4244) );
  OAI21_X1 U5245 ( .B1(n4322), .B2(n4402), .A(n4244), .ZN(U2894) );
  INV_X1 U5246 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U5247 ( .A1(n6592), .A2(UWORD_REG_11__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4245) );
  OAI21_X1 U5248 ( .B1(n4333), .B2(n4402), .A(n4245), .ZN(U2896) );
  INV_X1 U5249 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5250 ( .A1(n6592), .A2(UWORD_REG_14__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4246) );
  OAI21_X1 U5251 ( .B1(n4325), .B2(n4402), .A(n4246), .ZN(U2893) );
  OAI21_X1 U5252 ( .B1(n4249), .B2(n4248), .A(n4247), .ZN(n5077) );
  NAND2_X1 U5253 ( .A1(n4250), .A2(n6485), .ZN(n4251) );
  OAI211_X1 U5254 ( .C1(n4229), .C2(n4251), .A(n4286), .B(n4378), .ZN(n4252)
         );
  NAND2_X1 U5255 ( .A1(n4252), .A2(n3239), .ZN(n4263) );
  NOR2_X1 U5256 ( .A1(n5884), .A2(n4496), .ZN(n4288) );
  NAND2_X1 U5257 ( .A1(n6052), .A2(n4288), .ZN(n4260) );
  NAND2_X1 U5258 ( .A1(n3234), .A2(n4254), .ZN(n4255) );
  NAND2_X1 U5259 ( .A1(n4253), .A2(n4255), .ZN(n4280) );
  INV_X1 U5260 ( .A(n4280), .ZN(n4256) );
  NAND2_X1 U5261 ( .A1(n4268), .A2(n4256), .ZN(n4257) );
  NAND2_X1 U5262 ( .A1(n4257), .A2(n6468), .ZN(n4422) );
  NAND2_X1 U5263 ( .A1(n2993), .A2(n6514), .ZN(n4258) );
  NOR2_X1 U5264 ( .A1(READY_N), .A2(n6467), .ZN(n4370) );
  NAND3_X1 U5265 ( .A1(n4258), .A2(n4370), .A3(n4278), .ZN(n4259) );
  NAND3_X1 U5266 ( .A1(n4260), .A2(n4422), .A3(n4259), .ZN(n4261) );
  NAND2_X1 U5267 ( .A1(n4261), .A2(n4374), .ZN(n4262) );
  INV_X1 U5268 ( .A(n6476), .ZN(n4270) );
  OAI211_X1 U5269 ( .C1(n3260), .C2(n6794), .A(n4418), .B(n6043), .ZN(n4266)
         );
  INV_X1 U5270 ( .A(n4266), .ZN(n4269) );
  INV_X1 U5271 ( .A(n4267), .ZN(n4372) );
  INV_X1 U5272 ( .A(n4372), .ZN(n6054) );
  NAND2_X1 U5273 ( .A1(n4268), .A2(n6054), .ZN(n4412) );
  NAND3_X1 U5274 ( .A1(n4270), .A2(n4269), .A3(n4412), .ZN(n4271) );
  OAI21_X1 U5275 ( .B1(n6794), .B2(n4272), .A(n6488), .ZN(n4273) );
  XNOR2_X1 U5276 ( .A(n4274), .B(n4307), .ZN(n4311) );
  NAND2_X1 U5277 ( .A1(n6279), .A2(REIP_REG_1__SCAN_IN), .ZN(n5075) );
  INV_X1 U5278 ( .A(n5075), .ZN(n4290) );
  INV_X1 U5279 ( .A(n4291), .ZN(n4275) );
  INV_X1 U5280 ( .A(n6279), .ZN(n6323) );
  NAND2_X1 U5281 ( .A1(n4275), .A2(n6323), .ZN(n6340) );
  INV_X1 U5282 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6342) );
  AND2_X1 U5283 ( .A1(n3339), .A2(n4489), .ZN(n4277) );
  OAI22_X1 U5284 ( .A1(n3249), .A2(n5392), .B1(n3239), .B2(n4277), .ZN(n4283)
         );
  INV_X1 U5285 ( .A(n5369), .ZN(n5354) );
  OR2_X1 U5286 ( .A1(n5060), .A2(n4278), .ZN(n4421) );
  AOI21_X1 U5287 ( .B1(n5354), .B2(n4421), .A(n4279), .ZN(n4281) );
  OR2_X1 U5288 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  NOR2_X1 U5289 ( .A1(n4283), .A2(n4282), .ZN(n4285) );
  OAI211_X1 U5290 ( .C1(n4276), .C2(n4286), .A(n4408), .B(n4436), .ZN(n4287)
         );
  NAND2_X1 U5291 ( .A1(n4291), .A2(n4287), .ZN(n6033) );
  NAND2_X1 U5292 ( .A1(n4291), .A2(n6472), .ZN(n6322) );
  NAND2_X1 U5293 ( .A1(n6033), .A2(n6322), .ZN(n5853) );
  NAND2_X1 U5294 ( .A1(n6342), .A2(n5853), .ZN(n6333) );
  AOI21_X1 U5295 ( .B1(n6340), .B2(n6333), .A(n5300), .ZN(n4289) );
  AOI211_X1 U5296 ( .C1(n6293), .C2(n4311), .A(n4290), .B(n4289), .ZN(n4293)
         );
  NAND2_X1 U5297 ( .A1(n4291), .A2(n5324), .ZN(n6341) );
  NOR2_X1 U5298 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4535), .ZN(n4536)
         );
  OR3_X1 U5299 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4536), 
        .ZN(n4292) );
  OAI211_X1 U5300 ( .C1(n5077), .C2(n5870), .A(n4293), .B(n4292), .ZN(U3017)
         );
  INV_X1 U5301 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U5302 ( .A1(n4299), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4294) );
  NAND2_X1 U5303 ( .A1(n4341), .A2(DATAI_14_), .ZN(n4323) );
  OAI211_X1 U5304 ( .C1(n6231), .C2(n4359), .A(n4294), .B(n4323), .ZN(U2953)
         );
  INV_X1 U5305 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U5306 ( .A1(n4299), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4295) );
  NAND2_X1 U5307 ( .A1(n4341), .A2(DATAI_10_), .ZN(n4326) );
  OAI211_X1 U5308 ( .C1(n6238), .C2(n4359), .A(n4295), .B(n4326), .ZN(U2949)
         );
  NAND2_X1 U5309 ( .A1(n4299), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U5310 ( .A1(n4341), .A2(DATAI_12_), .ZN(n4314) );
  OAI211_X1 U5311 ( .C1(n5297), .C2(n4359), .A(n4296), .B(n4314), .ZN(U2951)
         );
  INV_X1 U5312 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U5313 ( .A1(n4299), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4297) );
  NAND2_X1 U5314 ( .A1(n4341), .A2(DATAI_9_), .ZN(n4344) );
  OAI211_X1 U5315 ( .C1(n6241), .C2(n4359), .A(n4297), .B(n4344), .ZN(U2948)
         );
  INV_X1 U5316 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5317 ( .A1(n4299), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U5318 ( .A1(n4341), .A2(DATAI_0_), .ZN(n4318) );
  OAI211_X1 U5319 ( .C1(n4394), .C2(n4359), .A(n4298), .B(n4318), .ZN(U2924)
         );
  INV_X1 U5320 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U5321 ( .A1(n4299), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U5322 ( .A1(n4341), .A2(DATAI_11_), .ZN(n4331) );
  OAI211_X1 U5323 ( .C1(n6236), .C2(n4359), .A(n4300), .B(n4331), .ZN(U2950)
         );
  OAI21_X1 U5324 ( .B1(n4303), .B2(n4301), .A(n3099), .ZN(n5081) );
  NAND2_X1 U5325 ( .A1(n6052), .A2(n6472), .ZN(n4424) );
  NAND3_X1 U5326 ( .A1(n4304), .A2(n3260), .A3(n5314), .ZN(n4306) );
  OR2_X1 U5327 ( .A1(n4306), .A2(n4305), .ZN(n4373) );
  INV_X1 U5328 ( .A(n4373), .ZN(n4308) );
  NAND2_X1 U5329 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  NAND2_X1 U5330 ( .A1(n4424), .A2(n4309), .ZN(n4310) );
  NAND2_X2 U5331 ( .A1(n6210), .A2(n3622), .ZN(n5533) );
  AOI22_X1 U5332 ( .A1(n6206), .A2(n4311), .B1(EBX_REG_1__SCAN_IN), .B2(n5528), 
        .ZN(n4312) );
  OAI21_X1 U5333 ( .B1(n5081), .B2(n5533), .A(n4312), .ZN(U2858) );
  NAND2_X1 U5334 ( .A1(n4356), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4315) );
  OAI211_X1 U5335 ( .C1(n4316), .C2(n4351), .A(n4315), .B(n4314), .ZN(U2936)
         );
  INV_X1 U5336 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U5337 ( .A1(n4356), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4317) );
  NAND2_X1 U5338 ( .A1(n4341), .A2(DATAI_6_), .ZN(n4337) );
  OAI211_X1 U5339 ( .C1(n6246), .C2(n4359), .A(n4317), .B(n4337), .ZN(U2945)
         );
  INV_X1 U5340 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U5341 ( .A1(n4356), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4319) );
  OAI211_X1 U5342 ( .C1(n6261), .C2(n4359), .A(n4319), .B(n4318), .ZN(U2939)
         );
  NAND2_X1 U5343 ( .A1(n4356), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4321) );
  OAI211_X1 U5344 ( .C1(n4322), .C2(n4359), .A(n4321), .B(n4320), .ZN(U2937)
         );
  NAND2_X1 U5345 ( .A1(n4356), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4324) );
  OAI211_X1 U5346 ( .C1(n4325), .C2(n4359), .A(n4324), .B(n4323), .ZN(U2938)
         );
  NAND2_X1 U5347 ( .A1(n4356), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4327) );
  OAI211_X1 U5348 ( .C1(n4328), .C2(n4351), .A(n4327), .B(n4326), .ZN(U2934)
         );
  INV_X1 U5349 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U5350 ( .A1(n4356), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4329) );
  NAND2_X1 U5351 ( .A1(n4341), .A2(DATAI_4_), .ZN(n4349) );
  OAI211_X1 U5352 ( .C1(n6250), .C2(n4359), .A(n4329), .B(n4349), .ZN(U2943)
         );
  INV_X1 U5353 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U5354 ( .A1(n4356), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4330) );
  NAND2_X1 U5355 ( .A1(n4341), .A2(DATAI_5_), .ZN(n4335) );
  OAI211_X1 U5356 ( .C1(n6248), .C2(n4359), .A(n4330), .B(n4335), .ZN(U2944)
         );
  NAND2_X1 U5357 ( .A1(n4356), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4332) );
  OAI211_X1 U5358 ( .C1(n4333), .C2(n4351), .A(n4332), .B(n4331), .ZN(U2935)
         );
  NAND2_X1 U5359 ( .A1(n4356), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4334) );
  NAND2_X1 U5360 ( .A1(n4341), .A2(DATAI_7_), .ZN(n4339) );
  OAI211_X1 U5361 ( .C1(n3676), .C2(n4359), .A(n4334), .B(n4339), .ZN(U2946)
         );
  INV_X1 U5362 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5363 ( .A1(n4356), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4336) );
  OAI211_X1 U5364 ( .C1(n4351), .C2(n4398), .A(n4336), .B(n4335), .ZN(U2929)
         );
  INV_X1 U5365 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5366 ( .A1(n4356), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U5367 ( .C1(n4400), .C2(n4359), .A(n4338), .B(n4337), .ZN(U2930)
         );
  INV_X1 U5368 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U5369 ( .A1(n4356), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4340) );
  OAI211_X1 U5370 ( .C1(n4403), .C2(n4351), .A(n4340), .B(n4339), .ZN(U2931)
         );
  NAND2_X1 U5371 ( .A1(n4356), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5372 ( .A1(n4341), .A2(DATAI_8_), .ZN(n4352) );
  OAI211_X1 U5373 ( .C1(n4343), .C2(n4351), .A(n4342), .B(n4352), .ZN(U2932)
         );
  NAND2_X1 U5374 ( .A1(n4356), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4345) );
  OAI211_X1 U5375 ( .C1(n4346), .C2(n4351), .A(n4345), .B(n4344), .ZN(U2933)
         );
  INV_X1 U5376 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U5377 ( .A1(n4356), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4348) );
  OAI211_X1 U5378 ( .C1(n6253), .C2(n4359), .A(n4348), .B(n4347), .ZN(U2942)
         );
  INV_X1 U5379 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U5380 ( .A1(n4356), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4350) );
  OAI211_X1 U5381 ( .C1(n4392), .C2(n4351), .A(n4350), .B(n4349), .ZN(U2928)
         );
  INV_X1 U5382 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U5383 ( .A1(n4356), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4353) );
  OAI211_X1 U5384 ( .C1(n6243), .C2(n4359), .A(n4353), .B(n4352), .ZN(U2947)
         );
  INV_X1 U5385 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U5386 ( .A1(n4356), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4355) );
  OAI211_X1 U5387 ( .C1(n6257), .C2(n4359), .A(n4355), .B(n4354), .ZN(U2940)
         );
  INV_X1 U5388 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U5389 ( .A1(n4356), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4358) );
  OAI211_X1 U5390 ( .C1(n6255), .C2(n4359), .A(n4358), .B(n4357), .ZN(U2941)
         );
  OR2_X1 U5391 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4361)
         );
  AND2_X1 U5392 ( .A1(n4361), .A2(n4360), .ZN(n5062) );
  INV_X1 U5393 ( .A(n5062), .ZN(n6334) );
  OAI21_X1 U5394 ( .B1(n4364), .B2(n4363), .A(n4362), .ZN(n6282) );
  OAI222_X1 U5395 ( .A1(n6334), .A2(n5530), .B1(n4365), .B2(n6210), .C1(n6282), 
        .C2(n5533), .ZN(U2859) );
  NOR2_X1 U5396 ( .A1(n4367), .A2(n4368), .ZN(n4369) );
  NOR2_X1 U5397 ( .A1(n4366), .A2(n4369), .ZN(n6267) );
  INV_X1 U5398 ( .A(n6267), .ZN(n4386) );
  INV_X1 U5399 ( .A(n4370), .ZN(n4371) );
  OAI22_X1 U5400 ( .A1(n6052), .A2(n4412), .B1(n6043), .B2(n4371), .ZN(n4427)
         );
  NOR2_X1 U5401 ( .A1(n4373), .A2(n4372), .ZN(n4375) );
  OAI21_X1 U5402 ( .B1(n4427), .B2(n4375), .A(n4374), .ZN(n4377) );
  NAND2_X1 U5403 ( .A1(n3237), .A2(n3622), .ZN(n4380) );
  AND2_X1 U5404 ( .A1(n4378), .A2(n4380), .ZN(n4379) );
  NAND2_X2 U5405 ( .A1(n6225), .A2(n4379), .ZN(n6226) );
  INV_X1 U5406 ( .A(n4380), .ZN(n4381) );
  AOI22_X1 U5407 ( .A1(n6220), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n6216), .ZN(n4382) );
  OAI21_X1 U5408 ( .B1(n4386), .B2(n6226), .A(n4382), .ZN(U2889) );
  NOR2_X1 U5409 ( .A1(n4384), .A2(n4383), .ZN(n4385) );
  OR2_X1 U5410 ( .A1(n4468), .A2(n4385), .ZN(n6324) );
  OAI222_X1 U5411 ( .A1(n4386), .A2(n5533), .B1(n3060), .B2(n6210), .C1(n5530), 
        .C2(n6324), .ZN(U2857) );
  INV_X1 U5412 ( .A(DATAI_1_), .ZN(n6675) );
  OAI222_X1 U5413 ( .A1(n5081), .A2(n6226), .B1(n6224), .B2(n6675), .C1(n6225), 
        .C2(n6257), .ZN(U2890) );
  AOI22_X1 U5414 ( .A1(n6239), .A2(UWORD_REG_1__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4387) );
  OAI21_X1 U5415 ( .B1(n4388), .B2(n4402), .A(n4387), .ZN(U2906) );
  AOI22_X1 U5416 ( .A1(n6239), .A2(UWORD_REG_3__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5417 ( .B1(n4390), .B2(n4402), .A(n4389), .ZN(U2904) );
  AOI22_X1 U5418 ( .A1(n6239), .A2(UWORD_REG_4__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4391) );
  OAI21_X1 U5419 ( .B1(n4392), .B2(n4402), .A(n4391), .ZN(U2903) );
  AOI22_X1 U5420 ( .A1(n6239), .A2(UWORD_REG_0__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4393) );
  OAI21_X1 U5421 ( .B1(n4394), .B2(n4402), .A(n4393), .ZN(U2907) );
  AOI22_X1 U5422 ( .A1(n6239), .A2(UWORD_REG_2__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4395) );
  OAI21_X1 U5423 ( .B1(n4396), .B2(n4402), .A(n4395), .ZN(U2905) );
  AOI22_X1 U5424 ( .A1(n6239), .A2(UWORD_REG_5__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4397) );
  OAI21_X1 U5425 ( .B1(n4398), .B2(n4402), .A(n4397), .ZN(U2902) );
  AOI22_X1 U5426 ( .A1(n6592), .A2(UWORD_REG_6__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4399) );
  OAI21_X1 U5427 ( .B1(n4400), .B2(n4402), .A(n4399), .ZN(U2901) );
  AOI22_X1 U5428 ( .A1(n6592), .A2(UWORD_REG_7__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4401) );
  OAI21_X1 U5429 ( .B1(n4403), .B2(n4402), .A(n4401), .ZN(U2900) );
  INV_X1 U5430 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6709) );
  NAND2_X1 U5431 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6709), .ZN(n4444) );
  INV_X1 U5432 ( .A(n4404), .ZN(n4443) );
  AND4_X1 U5433 ( .A1(n4276), .A2(n4229), .A3(n6043), .A4(n4406), .ZN(n4407)
         );
  NAND2_X1 U5434 ( .A1(n4408), .A2(n4407), .ZN(n5886) );
  INV_X1 U5435 ( .A(n5324), .ZN(n6452) );
  XNOR2_X1 U5436 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4411) );
  XNOR2_X1 U5437 ( .A(n4409), .B(n5305), .ZN(n4413) );
  INV_X1 U5438 ( .A(n4413), .ZN(n4410) );
  OAI22_X1 U5439 ( .A1(n6452), .A2(n4411), .B1(n4436), .B2(n4410), .ZN(n4415)
         );
  INV_X1 U5440 ( .A(n4412), .ZN(n6466) );
  NOR2_X1 U5441 ( .A1(n6472), .A2(n6466), .ZN(n4432) );
  NOR2_X1 U5442 ( .A1(n4432), .A2(n4413), .ZN(n4414) );
  AOI211_X1 U5443 ( .C1(n3002), .C2(n5886), .A(n4415), .B(n4414), .ZN(n5299)
         );
  OAI21_X1 U5444 ( .B1(n5324), .B2(n4417), .A(n4416), .ZN(n4419) );
  NAND2_X1 U5445 ( .A1(n4419), .A2(n4418), .ZN(n4420) );
  NAND2_X1 U5446 ( .A1(n4420), .A2(n6485), .ZN(n4425) );
  AND2_X1 U5447 ( .A1(n4422), .A2(n4421), .ZN(n4423) );
  OAI211_X1 U5448 ( .C1(n6052), .C2(n4425), .A(n4424), .B(n4423), .ZN(n4426)
         );
  OR2_X1 U5449 ( .A1(n4427), .A2(n4426), .ZN(n4440) );
  NOR2_X1 U5450 ( .A1(n4440), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4428)
         );
  AOI21_X1 U5451 ( .B1(n5299), .B2(n4440), .A(n4428), .ZN(n6462) );
  MUX2_X1 U5452 ( .A(n4430), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4409), 
        .Z(n4431) );
  NOR3_X1 U5453 ( .A1(n4432), .A2(n4404), .A3(n4431), .ZN(n4439) );
  NAND2_X1 U5454 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4434) );
  INV_X1 U5455 ( .A(n4434), .ZN(n4433) );
  MUX2_X1 U5456 ( .A(n4434), .B(n4433), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4437) );
  INV_X1 U5457 ( .A(n4409), .ZN(n5882) );
  AOI211_X1 U5458 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n5882), .A(n4435), .B(n3270), .ZN(n5895) );
  OAI22_X1 U5459 ( .A1(n6452), .A2(n4437), .B1(n5895), .B2(n4436), .ZN(n4438)
         );
  AOI211_X1 U5460 ( .C1(n3003), .C2(n5886), .A(n4439), .B(n4438), .ZN(n5897)
         );
  INV_X1 U5461 ( .A(n5897), .ZN(n4441) );
  MUX2_X1 U5462 ( .A(n4441), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6459), 
        .Z(n6450) );
  NAND3_X1 U5463 ( .A1(n6462), .A2(n6450), .A3(n5321), .ZN(n4442) );
  OAI21_X1 U5464 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(n6477) );
  INV_X1 U5465 ( .A(n6477), .ZN(n4451) );
  OAI21_X1 U5466 ( .B1(n6459), .B2(STATE2_REG_1__SCAN_IN), .A(n6709), .ZN(
        n4449) );
  INV_X1 U5467 ( .A(n4786), .ZN(n4582) );
  NOR2_X1 U5468 ( .A1(n4446), .A2(n4582), .ZN(n4447) );
  XNOR2_X1 U5469 ( .A(n4447), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6169)
         );
  OR3_X1 U5470 ( .A1(n6169), .A2(STATE2_REG_1__SCAN_IN), .A3(n6043), .ZN(n4448) );
  OAI21_X1 U5471 ( .B1(n4449), .B2(n6049), .A(n4448), .ZN(n6475) );
  INV_X1 U5472 ( .A(n6475), .ZN(n4450) );
  OAI21_X1 U5473 ( .B1(n4451), .B2(n4445), .A(n4450), .ZN(n4454) );
  NOR2_X1 U5474 ( .A1(n3053), .A2(n4453), .ZN(n5304) );
  OAI21_X1 U5475 ( .B1(n4454), .B2(FLUSH_REG_SCAN_IN), .A(n5304), .ZN(n4452)
         );
  NAND2_X1 U5476 ( .A1(n4452), .A2(n4790), .ZN(n6343) );
  NOR2_X1 U5477 ( .A1(n4454), .A2(n4453), .ZN(n6491) );
  AND2_X1 U5478 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6580), .ZN(n5878) );
  OAI22_X1 U5479 ( .A1(n4887), .A2(n6353), .B1(n3629), .B2(n5878), .ZN(n4455)
         );
  OAI21_X1 U5480 ( .B1(n6491), .B2(n4455), .A(n6343), .ZN(n4456) );
  OAI21_X1 U5481 ( .B1(n6343), .B2(n4951), .A(n4456), .ZN(U3465) );
  NOR2_X1 U5482 ( .A1(n3001), .A2(n4589), .ZN(n4458) );
  NAND2_X1 U5483 ( .A1(n4745), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4741) );
  NAND2_X1 U5484 ( .A1(n4741), .A2(n4606), .ZN(n4688) );
  INV_X1 U5485 ( .A(n4688), .ZN(n4461) );
  NAND2_X1 U5486 ( .A1(n3001), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5873) );
  NOR2_X1 U5487 ( .A1(n5873), .A2(n4459), .ZN(n4460) );
  NAND2_X1 U5488 ( .A1(n4460), .A2(n5877), .ZN(n4581) );
  AOI21_X1 U5489 ( .B1(n4461), .B2(n4581), .A(n6353), .ZN(n4463) );
  NAND2_X1 U5490 ( .A1(n5872), .A2(n6715), .ZN(n5113) );
  INV_X1 U5491 ( .A(n3003), .ZN(n4995) );
  OAI22_X1 U5492 ( .A1(n3640), .A2(n5113), .B1(n4995), .B2(n5878), .ZN(n4462)
         );
  OAI21_X1 U5493 ( .B1(n4463), .B2(n4462), .A(n6343), .ZN(n4464) );
  OAI21_X1 U5494 ( .B1(n6343), .B2(n6344), .A(n4464), .ZN(U3462) );
  OAI21_X1 U5495 ( .B1(n4366), .B2(n4466), .A(n4465), .ZN(n5093) );
  INV_X1 U5496 ( .A(DATAI_3_), .ZN(n4505) );
  OAI222_X1 U5497 ( .A1(n5093), .A2(n6226), .B1(n6224), .B2(n4505), .C1(n6225), 
        .C2(n6253), .ZN(U2888) );
  INV_X1 U5498 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4470) );
  OR2_X1 U5499 ( .A1(n4468), .A2(n4467), .ZN(n4469) );
  NAND2_X1 U5500 ( .A1(n4475), .A2(n4469), .ZN(n6310) );
  OAI222_X1 U5501 ( .A1(n5093), .A2(n5533), .B1(n4470), .B2(n6210), .C1(n6310), 
        .C2(n5530), .ZN(U2856) );
  AND2_X1 U5502 ( .A1(n4465), .A2(n4472), .ZN(n4473) );
  OR2_X1 U5503 ( .A1(n4471), .A2(n4473), .ZN(n6182) );
  NAND2_X1 U5504 ( .A1(n4475), .A2(n4474), .ZN(n4476) );
  AND2_X1 U5505 ( .A1(n4622), .A2(n4476), .ZN(n6177) );
  AOI22_X1 U5506 ( .A1(n6206), .A2(n6177), .B1(EBX_REG_4__SCAN_IN), .B2(n5528), 
        .ZN(n4477) );
  OAI21_X1 U5507 ( .B1(n6182), .B2(n5533), .A(n4477), .ZN(U2855) );
  INV_X1 U5508 ( .A(DATAI_4_), .ZN(n6694) );
  OAI222_X1 U5509 ( .A1(n6182), .A2(n6226), .B1(n6224), .B2(n6694), .C1(n6225), 
        .C2(n6250), .ZN(U2887) );
  AND2_X1 U5510 ( .A1(n4479), .A2(n3002), .ZN(n4787) );
  NAND2_X1 U5511 ( .A1(n4787), .A2(n5872), .ZN(n4794) );
  INV_X1 U5512 ( .A(n4794), .ZN(n4481) );
  AND2_X1 U5513 ( .A1(n4484), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6346) );
  INV_X1 U5514 ( .A(n4789), .ZN(n4480) );
  AOI22_X1 U5515 ( .A1(n4481), .A2(n4995), .B1(n6346), .B2(n3127), .ZN(n4531)
         );
  INV_X1 U5516 ( .A(DATAI_0_), .ZN(n6689) );
  INV_X1 U5517 ( .A(n6351), .ZN(n5218) );
  NOR2_X1 U5518 ( .A1(n4459), .A2(n3001), .ZN(n4482) );
  NAND2_X1 U5519 ( .A1(n5877), .A2(n4482), .ZN(n4491) );
  NAND2_X1 U5520 ( .A1(n4483), .A2(n5872), .ZN(n4553) );
  AND2_X1 U5521 ( .A1(n3001), .A2(n4964), .ZN(n4614) );
  NAND3_X1 U5522 ( .A1(n4696), .A2(n4614), .A3(n3640), .ZN(n4724) );
  INV_X1 U5523 ( .A(n5113), .ZN(n6356) );
  NAND2_X1 U5524 ( .A1(n4787), .A2(n4582), .ZN(n4543) );
  OAI21_X1 U5525 ( .B1(n4724), .B2(n6356), .A(n4543), .ZN(n4487) );
  NAND2_X1 U5526 ( .A1(n6455), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4748) );
  OR2_X1 U5527 ( .A1(n4748), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4550)
         );
  NOR2_X1 U5528 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4550), .ZN(n4528)
         );
  INV_X1 U5529 ( .A(n4528), .ZN(n4485) );
  NOR2_X1 U5530 ( .A1(n4484), .A2(n4641), .ZN(n4917) );
  OAI21_X1 U5531 ( .B1(n3127), .B2(n4641), .A(n4916), .ZN(n4834) );
  AOI211_X1 U5532 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4485), .A(n4917), .B(
        n4834), .ZN(n4486) );
  NAND2_X1 U5533 ( .A1(n4524), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4495) );
  INV_X1 U5534 ( .A(DATAI_24_), .ZN(n4490) );
  OR2_X1 U5535 ( .A1(n6281), .A2(n4490), .ZN(n5215) );
  INV_X1 U5536 ( .A(n4491), .ZN(n4548) );
  NAND2_X1 U5537 ( .A1(n4548), .A2(n4887), .ZN(n4574) );
  INV_X1 U5538 ( .A(DATAI_16_), .ZN(n4492) );
  OR2_X1 U5539 ( .A1(n6281), .A2(n4492), .ZN(n6365) );
  OAI22_X1 U5540 ( .A1(n5215), .A2(n4724), .B1(n4574), .B2(n6365), .ZN(n4493)
         );
  AOI21_X1 U5541 ( .B1(n6350), .B2(n4528), .A(n4493), .ZN(n4494) );
  OAI211_X1 U5542 ( .C1(n4531), .C2(n5218), .A(n4495), .B(n4494), .ZN(U3052)
         );
  INV_X1 U5543 ( .A(n6367), .ZN(n5224) );
  NAND2_X1 U5544 ( .A1(n4524), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4500) );
  INV_X1 U5545 ( .A(DATAI_25_), .ZN(n6733) );
  OR2_X1 U5546 ( .A1(n6281), .A2(n6733), .ZN(n5221) );
  INV_X1 U5547 ( .A(DATAI_17_), .ZN(n4497) );
  OR2_X1 U5548 ( .A1(n6281), .A2(n4497), .ZN(n6371) );
  OAI22_X1 U5549 ( .A1(n5221), .A2(n4724), .B1(n4574), .B2(n6371), .ZN(n4498)
         );
  AOI21_X1 U5550 ( .B1(n3006), .B2(n4528), .A(n4498), .ZN(n4499) );
  OAI211_X1 U5551 ( .C1(n4531), .C2(n5224), .A(n4500), .B(n4499), .ZN(U3053)
         );
  INV_X1 U5552 ( .A(DATAI_6_), .ZN(n6641) );
  INV_X1 U5553 ( .A(n6435), .ZN(n5246) );
  NAND2_X1 U5554 ( .A1(n4524), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4504) );
  NOR2_X2 U5555 ( .A1(n4525), .A2(n3628), .ZN(n6434) );
  INV_X1 U5556 ( .A(DATAI_30_), .ZN(n6703) );
  OR2_X1 U5557 ( .A1(n6281), .A2(n6703), .ZN(n6438) );
  INV_X1 U5558 ( .A(DATAI_22_), .ZN(n4501) );
  OR2_X1 U5559 ( .A1(n6281), .A2(n4501), .ZN(n6391) );
  OAI22_X1 U5560 ( .A1(n6438), .A2(n4724), .B1(n4574), .B2(n6391), .ZN(n4502)
         );
  AOI21_X1 U5561 ( .B1(n6434), .B2(n4528), .A(n4502), .ZN(n4503) );
  OAI211_X1 U5562 ( .C1(n4531), .C2(n5246), .A(n4504), .B(n4503), .ZN(U3058)
         );
  INV_X1 U5563 ( .A(n6417), .ZN(n5232) );
  NAND2_X1 U5564 ( .A1(n4524), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4511) );
  NOR2_X2 U5565 ( .A1(n4525), .A2(n4506), .ZN(n6416) );
  INV_X1 U5566 ( .A(DATAI_27_), .ZN(n4507) );
  OR2_X1 U5567 ( .A1(n6281), .A2(n4507), .ZN(n6420) );
  INV_X1 U5568 ( .A(DATAI_19_), .ZN(n4508) );
  OR2_X1 U5569 ( .A1(n6281), .A2(n4508), .ZN(n6379) );
  OAI22_X1 U5570 ( .A1(n6420), .A2(n4724), .B1(n4574), .B2(n6379), .ZN(n4509)
         );
  AOI21_X1 U5571 ( .B1(n6416), .B2(n4528), .A(n4509), .ZN(n4510) );
  OAI211_X1 U5572 ( .C1(n4531), .C2(n5232), .A(n4511), .B(n4510), .ZN(U3055)
         );
  INV_X1 U5573 ( .A(DATAI_2_), .ZN(n6661) );
  INV_X1 U5574 ( .A(n6411), .ZN(n5228) );
  NAND2_X1 U5575 ( .A1(n4524), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4515) );
  NOR2_X2 U5576 ( .A1(n4525), .A2(n3239), .ZN(n6410) );
  INV_X1 U5577 ( .A(DATAI_26_), .ZN(n6638) );
  OR2_X1 U5578 ( .A1(n6281), .A2(n6638), .ZN(n6414) );
  INV_X1 U5579 ( .A(DATAI_18_), .ZN(n4512) );
  OR2_X1 U5580 ( .A1(n6281), .A2(n4512), .ZN(n6375) );
  OAI22_X1 U5581 ( .A1(n6414), .A2(n4724), .B1(n4574), .B2(n6375), .ZN(n4513)
         );
  AOI21_X1 U5582 ( .B1(n6410), .B2(n4528), .A(n4513), .ZN(n4514) );
  OAI211_X1 U5583 ( .C1(n4531), .C2(n5228), .A(n4515), .B(n4514), .ZN(U3054)
         );
  INV_X1 U5584 ( .A(DATAI_5_), .ZN(n4625) );
  INV_X1 U5585 ( .A(n6429), .ZN(n5254) );
  NAND2_X1 U5586 ( .A1(n4524), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4519) );
  NOR2_X2 U5587 ( .A1(n4525), .A2(n3237), .ZN(n6428) );
  INV_X1 U5588 ( .A(DATAI_29_), .ZN(n6725) );
  OR2_X1 U5589 ( .A1(n6281), .A2(n6725), .ZN(n6432) );
  INV_X1 U5590 ( .A(DATAI_21_), .ZN(n4516) );
  OR2_X1 U5591 ( .A1(n6281), .A2(n4516), .ZN(n6387) );
  OAI22_X1 U5592 ( .A1(n6432), .A2(n4724), .B1(n4574), .B2(n6387), .ZN(n4517)
         );
  AOI21_X1 U5593 ( .B1(n6428), .B2(n4528), .A(n4517), .ZN(n4518) );
  OAI211_X1 U5594 ( .C1(n4531), .C2(n5254), .A(n4519), .B(n4518), .ZN(U3057)
         );
  NAND2_X1 U5595 ( .A1(n4524), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4523) );
  NOR2_X2 U5596 ( .A1(n4525), .A2(n3260), .ZN(n6422) );
  INV_X1 U5597 ( .A(DATAI_28_), .ZN(n4520) );
  OR2_X1 U5598 ( .A1(n6281), .A2(n4520), .ZN(n6426) );
  OR2_X1 U5599 ( .A1(n6281), .A2(n6716), .ZN(n6383) );
  OAI22_X1 U5600 ( .A1(n6426), .A2(n4724), .B1(n4574), .B2(n6383), .ZN(n4521)
         );
  AOI21_X1 U5601 ( .B1(n6422), .B2(n4528), .A(n4521), .ZN(n4522) );
  OAI211_X1 U5602 ( .C1(n4531), .C2(n5250), .A(n4523), .B(n4522), .ZN(U3056)
         );
  INV_X1 U5603 ( .A(DATAI_7_), .ZN(n5035) );
  INV_X1 U5604 ( .A(n6444), .ZN(n5262) );
  NAND2_X1 U5605 ( .A1(n4524), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4530) );
  NOR2_X2 U5606 ( .A1(n4525), .A2(n5314), .ZN(n6442) );
  INV_X1 U5607 ( .A(DATAI_31_), .ZN(n6650) );
  OR2_X1 U5608 ( .A1(n6281), .A2(n6650), .ZN(n6449) );
  INV_X1 U5609 ( .A(DATAI_23_), .ZN(n4526) );
  OR2_X1 U5610 ( .A1(n6281), .A2(n4526), .ZN(n6399) );
  OAI22_X1 U5611 ( .A1(n6449), .A2(n4724), .B1(n4574), .B2(n6399), .ZN(n4527)
         );
  AOI21_X1 U5612 ( .B1(n6442), .B2(n4528), .A(n4527), .ZN(n4529) );
  OAI211_X1 U5613 ( .C1(n4531), .C2(n5262), .A(n4530), .B(n4529), .ZN(U3059)
         );
  XNOR2_X1 U5614 ( .A(n4533), .B(n4532), .ZN(n5045) );
  INV_X1 U5615 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6330) );
  INV_X1 U5616 ( .A(n6033), .ZN(n4534) );
  NOR2_X1 U5617 ( .A1(n4536), .A2(n5708), .ZN(n5721) );
  NAND2_X1 U5618 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5721), .ZN(n6331)
         );
  INV_X1 U5619 ( .A(n6322), .ZN(n5720) );
  OR2_X1 U5620 ( .A1(n5725), .A2(n5720), .ZN(n4537) );
  OAI21_X1 U5621 ( .B1(n5300), .B2(n6342), .A(n6330), .ZN(n6318) );
  NAND2_X1 U5622 ( .A1(n4537), .A2(n6318), .ZN(n6311) );
  NAND2_X1 U5623 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4632) );
  INV_X1 U5624 ( .A(n4632), .ZN(n4538) );
  NOR2_X1 U5625 ( .A1(n6311), .A2(n4538), .ZN(n4629) );
  OAI21_X1 U5626 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4629), .ZN(n4542) );
  NOR2_X1 U5627 ( .A1(n6322), .A2(n6318), .ZN(n5177) );
  NOR2_X1 U5628 ( .A1(n6330), .A2(n5300), .ZN(n6320) );
  OAI21_X1 U5629 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6033), .A(n6340), 
        .ZN(n5709) );
  INV_X1 U5630 ( .A(n5709), .ZN(n4539) );
  OAI21_X1 U5631 ( .B1(n5708), .B2(n6320), .A(n4539), .ZN(n6317) );
  NOR2_X1 U5632 ( .A1(n5177), .A2(n6317), .ZN(n6316) );
  NAND2_X1 U5633 ( .A1(n6279), .A2(REIP_REG_4__SCAN_IN), .ZN(n5039) );
  OAI21_X1 U5634 ( .B1(n4148), .B2(n6316), .A(n5039), .ZN(n4540) );
  AOI21_X1 U5635 ( .B1(n6293), .B2(n6177), .A(n4540), .ZN(n4541) );
  OAI211_X1 U5636 ( .C1(n5870), .C2(n5045), .A(n4542), .B(n4541), .ZN(U3014)
         );
  INV_X1 U5637 ( .A(n4553), .ZN(n4547) );
  OR2_X1 U5638 ( .A1(n4543), .A2(n3629), .ZN(n4545) );
  NOR2_X1 U5639 ( .A1(n4951), .A2(n4550), .ZN(n4576) );
  INV_X1 U5640 ( .A(n4576), .ZN(n4544) );
  NAND2_X1 U5641 ( .A1(n4545), .A2(n4544), .ZN(n4552) );
  INV_X1 U5642 ( .A(n4550), .ZN(n4546) );
  AOI22_X1 U5643 ( .A1(n4547), .A2(n4552), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4546), .ZN(n4580) );
  NAND2_X1 U5644 ( .A1(n4548), .A2(n4964), .ZN(n6352) );
  OAI22_X1 U5645 ( .A1(n6352), .A2(n6391), .B1(n4574), .B2(n6438), .ZN(n4549)
         );
  AOI21_X1 U5646 ( .B1(n6434), .B2(n4576), .A(n4549), .ZN(n4555) );
  INV_X1 U5647 ( .A(n4957), .ZN(n4700) );
  AOI21_X1 U5648 ( .B1(n6353), .B2(n4550), .A(n4700), .ZN(n4551) );
  OAI21_X1 U5649 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n4577) );
  NAND2_X1 U5650 ( .A1(n4577), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4554) );
  OAI211_X1 U5651 ( .C1(n5246), .C2(n4580), .A(n4555), .B(n4554), .ZN(U3066)
         );
  OAI22_X1 U5652 ( .A1(n6352), .A2(n6371), .B1(n4574), .B2(n5221), .ZN(n4556)
         );
  AOI21_X1 U5653 ( .B1(n3006), .B2(n4576), .A(n4556), .ZN(n4558) );
  NAND2_X1 U5654 ( .A1(n4577), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4557) );
  OAI211_X1 U5655 ( .C1(n5224), .C2(n4580), .A(n4558), .B(n4557), .ZN(U3061)
         );
  OAI22_X1 U5656 ( .A1(n6352), .A2(n6375), .B1(n4574), .B2(n6414), .ZN(n4559)
         );
  AOI21_X1 U5657 ( .B1(n6410), .B2(n4576), .A(n4559), .ZN(n4561) );
  NAND2_X1 U5658 ( .A1(n4577), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4560) );
  OAI211_X1 U5659 ( .C1(n5228), .C2(n4580), .A(n4561), .B(n4560), .ZN(U3062)
         );
  OAI22_X1 U5660 ( .A1(n6352), .A2(n6383), .B1(n4574), .B2(n6426), .ZN(n4562)
         );
  AOI21_X1 U5661 ( .B1(n6422), .B2(n4576), .A(n4562), .ZN(n4564) );
  NAND2_X1 U5662 ( .A1(n4577), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4563) );
  OAI211_X1 U5663 ( .C1(n5250), .C2(n4580), .A(n4564), .B(n4563), .ZN(U3064)
         );
  OAI22_X1 U5664 ( .A1(n6352), .A2(n6365), .B1(n4574), .B2(n5215), .ZN(n4565)
         );
  AOI21_X1 U5665 ( .B1(n6350), .B2(n4576), .A(n4565), .ZN(n4567) );
  NAND2_X1 U5666 ( .A1(n4577), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4566) );
  OAI211_X1 U5667 ( .C1(n5218), .C2(n4580), .A(n4567), .B(n4566), .ZN(U3060)
         );
  OAI22_X1 U5668 ( .A1(n6352), .A2(n6387), .B1(n4574), .B2(n6432), .ZN(n4568)
         );
  AOI21_X1 U5669 ( .B1(n6428), .B2(n4576), .A(n4568), .ZN(n4570) );
  NAND2_X1 U5670 ( .A1(n4577), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4569) );
  OAI211_X1 U5671 ( .C1(n5254), .C2(n4580), .A(n4570), .B(n4569), .ZN(U3065)
         );
  OAI22_X1 U5672 ( .A1(n6352), .A2(n6379), .B1(n4574), .B2(n6420), .ZN(n4571)
         );
  AOI21_X1 U5673 ( .B1(n6416), .B2(n4576), .A(n4571), .ZN(n4573) );
  NAND2_X1 U5674 ( .A1(n4577), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4572) );
  OAI211_X1 U5675 ( .C1(n5232), .C2(n4580), .A(n4573), .B(n4572), .ZN(U3063)
         );
  OAI22_X1 U5676 ( .A1(n6352), .A2(n6399), .B1(n4574), .B2(n6449), .ZN(n4575)
         );
  AOI21_X1 U5677 ( .B1(n6442), .B2(n4576), .A(n4575), .ZN(n4579) );
  NAND2_X1 U5678 ( .A1(n4577), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4578) );
  OAI211_X1 U5679 ( .C1(n5262), .C2(n4580), .A(n4579), .B(n4578), .ZN(U3067)
         );
  NAND2_X1 U5680 ( .A1(n4581), .A2(n5872), .ZN(n4586) );
  NAND2_X1 U5681 ( .A1(n4913), .A2(n4582), .ZN(n6355) );
  OR2_X1 U5682 ( .A1(n6355), .A2(n3629), .ZN(n4583) );
  NAND2_X1 U5683 ( .A1(n4583), .A2(n6400), .ZN(n4585) );
  INV_X1 U5684 ( .A(n4585), .ZN(n4584) );
  OAI22_X1 U5685 ( .A1(n4586), .A2(n4584), .B1(n6349), .B2(n4641), .ZN(n6403)
         );
  OR2_X1 U5686 ( .A1(n4586), .A2(n4585), .ZN(n4588) );
  AOI21_X1 U5687 ( .B1(n6353), .B2(n6349), .A(n4700), .ZN(n4587) );
  NAND2_X1 U5688 ( .A1(n4588), .A2(n4587), .ZN(n6404) );
  AOI22_X1 U5689 ( .A1(n6367), .A2(n6403), .B1(INSTQUEUE_REG_7__1__SCAN_IN), 
        .B2(n6404), .ZN(n4592) );
  NAND3_X1 U5690 ( .A1(n5877), .A2(n4589), .A3(n4695), .ZN(n6407) );
  INV_X1 U5691 ( .A(n5221), .ZN(n6368) );
  AND3_X1 U5692 ( .A1(n3001), .A2(n4589), .A3(n4964), .ZN(n4590) );
  NAND2_X1 U5693 ( .A1(n5877), .A2(n4590), .ZN(n4992) );
  INV_X1 U5694 ( .A(n6371), .ZN(n5219) );
  AOI22_X1 U5695 ( .A1(n6354), .A2(n6368), .B1(n6401), .B2(n5219), .ZN(n4591)
         );
  OAI211_X1 U5696 ( .C1(n6400), .C2(n6366), .A(n4592), .B(n4591), .ZN(U3077)
         );
  INV_X1 U5697 ( .A(n6350), .ZN(n4990) );
  AOI22_X1 U5698 ( .A1(n6351), .A2(n6403), .B1(INSTQUEUE_REG_7__0__SCAN_IN), 
        .B2(n6404), .ZN(n4594) );
  INV_X1 U5699 ( .A(n5215), .ZN(n6362) );
  INV_X1 U5700 ( .A(n6365), .ZN(n5213) );
  AOI22_X1 U5701 ( .A1(n6354), .A2(n6362), .B1(n6401), .B2(n5213), .ZN(n4593)
         );
  OAI211_X1 U5702 ( .C1(n6400), .C2(n4990), .A(n4594), .B(n4593), .ZN(U3076)
         );
  INV_X1 U5703 ( .A(n6410), .ZN(n4983) );
  AOI22_X1 U5704 ( .A1(n6411), .A2(n6403), .B1(INSTQUEUE_REG_7__2__SCAN_IN), 
        .B2(n6404), .ZN(n4596) );
  INV_X1 U5705 ( .A(n6414), .ZN(n6372) );
  INV_X1 U5706 ( .A(n6375), .ZN(n6409) );
  AOI22_X1 U5707 ( .A1(n6354), .A2(n6372), .B1(n6401), .B2(n6409), .ZN(n4595)
         );
  OAI211_X1 U5708 ( .C1(n6400), .C2(n4983), .A(n4596), .B(n4595), .ZN(U3078)
         );
  INV_X1 U5709 ( .A(n6442), .ZN(n4971) );
  AOI22_X1 U5710 ( .A1(n6444), .A2(n6403), .B1(INSTQUEUE_REG_7__7__SCAN_IN), 
        .B2(n6404), .ZN(n4598) );
  INV_X1 U5711 ( .A(n6449), .ZN(n6395) );
  INV_X1 U5712 ( .A(n6399), .ZN(n6439) );
  AOI22_X1 U5713 ( .A1(n6354), .A2(n6395), .B1(n6401), .B2(n6439), .ZN(n4597)
         );
  OAI211_X1 U5714 ( .C1(n6400), .C2(n4971), .A(n4598), .B(n4597), .ZN(U3083)
         );
  INV_X1 U5715 ( .A(n6428), .ZN(n4974) );
  AOI22_X1 U5716 ( .A1(n6429), .A2(n6403), .B1(INSTQUEUE_REG_7__5__SCAN_IN), 
        .B2(n6404), .ZN(n4600) );
  INV_X1 U5717 ( .A(n6432), .ZN(n6384) );
  INV_X1 U5718 ( .A(n6387), .ZN(n6427) );
  AOI22_X1 U5719 ( .A1(n6354), .A2(n6384), .B1(n6401), .B2(n6427), .ZN(n4599)
         );
  OAI211_X1 U5720 ( .C1(n6400), .C2(n4974), .A(n4600), .B(n4599), .ZN(U3081)
         );
  INV_X1 U5721 ( .A(n6434), .ZN(n4977) );
  AOI22_X1 U5722 ( .A1(n6435), .A2(n6403), .B1(INSTQUEUE_REG_7__6__SCAN_IN), 
        .B2(n6404), .ZN(n4602) );
  INV_X1 U5723 ( .A(n6438), .ZN(n6388) );
  INV_X1 U5724 ( .A(n6391), .ZN(n6433) );
  AOI22_X1 U5725 ( .A1(n6354), .A2(n6388), .B1(n6401), .B2(n6433), .ZN(n4601)
         );
  OAI211_X1 U5726 ( .C1(n6400), .C2(n4977), .A(n4602), .B(n4601), .ZN(U3082)
         );
  INV_X1 U5727 ( .A(n6422), .ZN(n4980) );
  AOI22_X1 U5728 ( .A1(n6423), .A2(n6403), .B1(INSTQUEUE_REG_7__4__SCAN_IN), 
        .B2(n6404), .ZN(n4604) );
  INV_X1 U5729 ( .A(n6426), .ZN(n6380) );
  INV_X1 U5730 ( .A(n6383), .ZN(n6421) );
  AOI22_X1 U5731 ( .A1(n6354), .A2(n6380), .B1(n6401), .B2(n6421), .ZN(n4603)
         );
  OAI211_X1 U5732 ( .C1(n6400), .C2(n4980), .A(n4604), .B(n4603), .ZN(U3080)
         );
  INV_X1 U5733 ( .A(n4605), .ZN(n4691) );
  NAND2_X1 U5734 ( .A1(n4691), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6408) );
  NAND3_X1 U5735 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6461), .ZN(n5205) );
  INV_X1 U5736 ( .A(n5873), .ZN(n5876) );
  NAND2_X1 U5737 ( .A1(n4962), .A2(n5876), .ZN(n4611) );
  NOR2_X1 U5738 ( .A1(n3002), .A2(n4479), .ZN(n4690) );
  AND2_X1 U5739 ( .A1(n4690), .A2(n3003), .ZN(n5207) );
  INV_X1 U5740 ( .A(n3629), .ZN(n5063) );
  NAND2_X1 U5741 ( .A1(n5207), .A2(n5063), .ZN(n4607) );
  NAND2_X1 U5742 ( .A1(n4607), .A2(n6408), .ZN(n4609) );
  NAND3_X1 U5743 ( .A1(n4611), .A2(n5872), .A3(n4609), .ZN(n4608) );
  OAI21_X1 U5744 ( .B1(n5205), .B2(n4641), .A(n4608), .ZN(n6443) );
  NOR2_X1 U5745 ( .A1(n4609), .A2(n6353), .ZN(n4610) );
  NAND2_X1 U5746 ( .A1(n4611), .A2(n4610), .ZN(n4613) );
  AOI21_X1 U5747 ( .B1(n6353), .B2(n5205), .A(n4700), .ZN(n4612) );
  NAND2_X1 U5748 ( .A1(n4613), .A2(n4612), .ZN(n6445) );
  AOI22_X1 U5749 ( .A1(n6351), .A2(n6443), .B1(INSTQUEUE_REG_11__0__SCAN_IN), 
        .B2(n6445), .ZN(n4616) );
  AOI22_X1 U5750 ( .A1(n6362), .A2(n5256), .B1(n6440), .B2(n5213), .ZN(n4615)
         );
  OAI211_X1 U5751 ( .C1(n4990), .C2(n6408), .A(n4616), .B(n4615), .ZN(U3108)
         );
  AOI22_X1 U5752 ( .A1(n6367), .A2(n6443), .B1(INSTQUEUE_REG_11__1__SCAN_IN), 
        .B2(n6445), .ZN(n4618) );
  AOI22_X1 U5753 ( .A1(n6368), .A2(n5256), .B1(n6440), .B2(n5219), .ZN(n4617)
         );
  OAI211_X1 U5754 ( .C1(n6366), .C2(n6408), .A(n4618), .B(n4617), .ZN(U3109)
         );
  OR2_X1 U5755 ( .A1(n4471), .A2(n4620), .ZN(n4621) );
  AND2_X1 U5756 ( .A1(n4619), .A2(n4621), .ZN(n6165) );
  INV_X1 U5757 ( .A(n6165), .ZN(n4626) );
  AOI21_X1 U5758 ( .B1(n4623), .B2(n4622), .A(n3055), .ZN(n6157) );
  AOI22_X1 U5759 ( .A1(n6157), .A2(n6206), .B1(EBX_REG_5__SCAN_IN), .B2(n5528), 
        .ZN(n4624) );
  OAI21_X1 U5760 ( .B1(n4626), .B2(n5533), .A(n4624), .ZN(U2854) );
  OAI222_X1 U5761 ( .A1(n4626), .A2(n6226), .B1(n6224), .B2(n4625), .C1(n6225), 
        .C2(n6248), .ZN(U2886) );
  XNOR2_X1 U5762 ( .A(n4628), .B(n4627), .ZN(n5050) );
  NOR2_X1 U5763 ( .A1(n5720), .A2(n5725), .ZN(n4631) );
  INV_X1 U5764 ( .A(n4629), .ZN(n4630) );
  OAI211_X1 U5765 ( .C1(INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n4631), .A(n6316), 
        .B(n4630), .ZN(n4873) );
  OAI21_X1 U5766 ( .B1(n4632), .B2(n6311), .A(n3483), .ZN(n4633) );
  NAND2_X1 U5767 ( .A1(n4873), .A2(n4633), .ZN(n4635) );
  AND2_X1 U5768 ( .A1(n6279), .A2(REIP_REG_5__SCAN_IN), .ZN(n5046) );
  AOI21_X1 U5769 ( .B1(n6157), .B2(n6293), .A(n5046), .ZN(n4634) );
  OAI211_X1 U5770 ( .C1(n5050), .C2(n5870), .A(n4635), .B(n4634), .ZN(U3013)
         );
  AND2_X1 U5771 ( .A1(n3003), .A2(n5063), .ZN(n4954) );
  INV_X1 U5772 ( .A(n4673), .ZN(n4636) );
  AOI21_X1 U5773 ( .B1(n4954), .B2(n4913), .A(n4636), .ZN(n4642) );
  AND2_X1 U5774 ( .A1(n4459), .A2(n3001), .ZN(n4637) );
  AND2_X1 U5775 ( .A1(n5877), .A2(n4637), .ZN(n4643) );
  OAI21_X1 U5776 ( .B1(n4643), .B2(n6281), .A(n5113), .ZN(n4639) );
  NOR2_X1 U5777 ( .A1(n5872), .A2(n4640), .ZN(n4638) );
  AOI211_X2 U5778 ( .C1(n4642), .C2(n4639), .A(n4638), .B(n4700), .ZN(n4679)
         );
  INV_X1 U5779 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4648) );
  INV_X1 U5780 ( .A(n4640), .ZN(n4918) );
  OAI22_X1 U5781 ( .A1(n4642), .A2(n6353), .B1(n4641), .B2(n4918), .ZN(n4676)
         );
  INV_X1 U5782 ( .A(n4643), .ZN(n4644) );
  NAND3_X1 U5783 ( .A1(n5877), .A2(n4695), .A3(n4459), .ZN(n4944) );
  OAI22_X1 U5784 ( .A1(n4864), .A2(n6375), .B1(n4944), .B2(n6414), .ZN(n4646)
         );
  NOR2_X1 U5785 ( .A1(n4983), .A2(n4673), .ZN(n4645) );
  AOI211_X1 U5786 ( .C1(n6411), .C2(n4676), .A(n4646), .B(n4645), .ZN(n4647)
         );
  OAI21_X1 U5787 ( .B1(n4679), .B2(n4648), .A(n4647), .ZN(U3142) );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4652) );
  OAI22_X1 U5789 ( .A1(n4864), .A2(n6365), .B1(n4944), .B2(n5215), .ZN(n4650)
         );
  NOR2_X1 U5790 ( .A1(n4990), .A2(n4673), .ZN(n4649) );
  AOI211_X1 U5791 ( .C1(n6351), .C2(n4676), .A(n4650), .B(n4649), .ZN(n4651)
         );
  OAI21_X1 U5792 ( .B1(n4679), .B2(n4652), .A(n4651), .ZN(U3140) );
  INV_X1 U5793 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4656) );
  OAI22_X1 U5794 ( .A1(n4864), .A2(n6399), .B1(n4944), .B2(n6449), .ZN(n4654)
         );
  NOR2_X1 U5795 ( .A1(n4971), .A2(n4673), .ZN(n4653) );
  AOI211_X1 U5796 ( .C1(n6444), .C2(n4676), .A(n4654), .B(n4653), .ZN(n4655)
         );
  OAI21_X1 U5797 ( .B1(n4679), .B2(n4656), .A(n4655), .ZN(U3147) );
  INV_X1 U5798 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4660) );
  OAI22_X1 U5799 ( .A1(n4864), .A2(n6371), .B1(n4944), .B2(n5221), .ZN(n4658)
         );
  NOR2_X1 U5800 ( .A1(n6366), .A2(n4673), .ZN(n4657) );
  AOI211_X1 U5801 ( .C1(n6367), .C2(n4676), .A(n4658), .B(n4657), .ZN(n4659)
         );
  OAI21_X1 U5802 ( .B1(n4679), .B2(n4660), .A(n4659), .ZN(U3141) );
  INV_X1 U5803 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4664) );
  OAI22_X1 U5804 ( .A1(n4864), .A2(n6379), .B1(n4944), .B2(n6420), .ZN(n4662)
         );
  INV_X1 U5805 ( .A(n6416), .ZN(n4968) );
  NOR2_X1 U5806 ( .A1(n4968), .A2(n4673), .ZN(n4661) );
  AOI211_X1 U5807 ( .C1(n6417), .C2(n4676), .A(n4662), .B(n4661), .ZN(n4663)
         );
  OAI21_X1 U5808 ( .B1(n4679), .B2(n4664), .A(n4663), .ZN(U3143) );
  INV_X1 U5809 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4668) );
  OAI22_X1 U5810 ( .A1(n4864), .A2(n6383), .B1(n4944), .B2(n6426), .ZN(n4666)
         );
  NOR2_X1 U5811 ( .A1(n4980), .A2(n4673), .ZN(n4665) );
  AOI211_X1 U5812 ( .C1(n6423), .C2(n4676), .A(n4666), .B(n4665), .ZN(n4667)
         );
  OAI21_X1 U5813 ( .B1(n4679), .B2(n4668), .A(n4667), .ZN(U3144) );
  INV_X1 U5814 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4672) );
  OAI22_X1 U5815 ( .A1(n4864), .A2(n6391), .B1(n4944), .B2(n6438), .ZN(n4670)
         );
  NOR2_X1 U5816 ( .A1(n4977), .A2(n4673), .ZN(n4669) );
  AOI211_X1 U5817 ( .C1(n6435), .C2(n4676), .A(n4670), .B(n4669), .ZN(n4671)
         );
  OAI21_X1 U5818 ( .B1(n4679), .B2(n4672), .A(n4671), .ZN(U3146) );
  INV_X1 U5819 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4678) );
  OAI22_X1 U5820 ( .A1(n4864), .A2(n6387), .B1(n4944), .B2(n6432), .ZN(n4675)
         );
  NOR2_X1 U5821 ( .A1(n4974), .A2(n4673), .ZN(n4674) );
  AOI211_X1 U5822 ( .C1(n6429), .C2(n4676), .A(n4675), .B(n4674), .ZN(n4677)
         );
  OAI21_X1 U5823 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(U3145) );
  OAI21_X1 U5824 ( .B1(n3672), .B2(n3671), .A(n4682), .ZN(n5095) );
  NAND2_X1 U5825 ( .A1(n4684), .A2(n4683), .ZN(n4685) );
  NAND2_X1 U5826 ( .A1(n5036), .A2(n4685), .ZN(n4874) );
  OAI22_X1 U5827 ( .A1(n4874), .A2(n5530), .B1(n4734), .B2(n6210), .ZN(n4686)
         );
  INV_X1 U5828 ( .A(n4686), .ZN(n4687) );
  OAI21_X1 U5829 ( .B1(n5095), .B2(n5533), .A(n4687), .ZN(U2853) );
  NOR3_X1 U5830 ( .A1(n4688), .A2(n5877), .A3(n5873), .ZN(n4689) );
  NOR2_X1 U5831 ( .A1(n4689), .A2(n6353), .ZN(n4699) );
  NAND2_X1 U5832 ( .A1(n4995), .A2(n4690), .ZN(n5115) );
  OR2_X1 U5833 ( .A1(n5115), .A2(n3629), .ZN(n4692) );
  NAND2_X1 U5834 ( .A1(n4691), .A2(n6344), .ZN(n4694) );
  NAND2_X1 U5835 ( .A1(n4692), .A2(n4694), .ZN(n4702) );
  NAND3_X1 U5836 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6344), .A3(n6461), .ZN(n5117) );
  INV_X1 U5837 ( .A(n5117), .ZN(n4693) );
  AOI22_X1 U5838 ( .A1(n4699), .A2(n4702), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4693), .ZN(n4730) );
  INV_X1 U5839 ( .A(n4694), .ZN(n4726) );
  AND2_X1 U5840 ( .A1(n3640), .A2(n4695), .ZN(n4697) );
  AND2_X1 U5841 ( .A1(n4697), .A2(n4696), .ZN(n5114) );
  OAI22_X1 U5842 ( .A1(n5143), .A2(n6438), .B1(n6391), .B2(n4724), .ZN(n4698)
         );
  AOI21_X1 U5843 ( .B1(n6434), .B2(n4726), .A(n4698), .ZN(n4705) );
  INV_X1 U5844 ( .A(n4699), .ZN(n4703) );
  AOI21_X1 U5845 ( .B1(n6353), .B2(n5117), .A(n4700), .ZN(n4701) );
  NAND2_X1 U5846 ( .A1(n4727), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4704) );
  OAI211_X1 U5847 ( .C1(n4730), .C2(n5246), .A(n4705), .B(n4704), .ZN(U3050)
         );
  OAI22_X1 U5848 ( .A1(n5143), .A2(n6432), .B1(n6387), .B2(n4724), .ZN(n4706)
         );
  AOI21_X1 U5849 ( .B1(n6428), .B2(n4726), .A(n4706), .ZN(n4708) );
  NAND2_X1 U5850 ( .A1(n4727), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4707) );
  OAI211_X1 U5851 ( .C1(n4730), .C2(n5254), .A(n4708), .B(n4707), .ZN(U3049)
         );
  OAI22_X1 U5852 ( .A1(n5143), .A2(n5215), .B1(n6365), .B2(n4724), .ZN(n4709)
         );
  AOI21_X1 U5853 ( .B1(n6350), .B2(n4726), .A(n4709), .ZN(n4711) );
  NAND2_X1 U5854 ( .A1(n4727), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4710) );
  OAI211_X1 U5855 ( .C1(n4730), .C2(n5218), .A(n4711), .B(n4710), .ZN(U3044)
         );
  OAI22_X1 U5856 ( .A1(n5143), .A2(n6426), .B1(n6383), .B2(n4724), .ZN(n4712)
         );
  AOI21_X1 U5857 ( .B1(n6422), .B2(n4726), .A(n4712), .ZN(n4714) );
  NAND2_X1 U5858 ( .A1(n4727), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4713) );
  OAI211_X1 U5859 ( .C1(n4730), .C2(n5250), .A(n4714), .B(n4713), .ZN(U3048)
         );
  OAI22_X1 U5860 ( .A1(n5143), .A2(n6414), .B1(n6375), .B2(n4724), .ZN(n4715)
         );
  AOI21_X1 U5861 ( .B1(n6410), .B2(n4726), .A(n4715), .ZN(n4717) );
  NAND2_X1 U5862 ( .A1(n4727), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4716) );
  OAI211_X1 U5863 ( .C1(n4730), .C2(n5228), .A(n4717), .B(n4716), .ZN(U3046)
         );
  OAI22_X1 U5864 ( .A1(n5143), .A2(n5221), .B1(n6371), .B2(n4724), .ZN(n4718)
         );
  AOI21_X1 U5865 ( .B1(n3007), .B2(n4726), .A(n4718), .ZN(n4720) );
  NAND2_X1 U5866 ( .A1(n4727), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4719) );
  OAI211_X1 U5867 ( .C1(n4730), .C2(n5224), .A(n4720), .B(n4719), .ZN(U3045)
         );
  OAI22_X1 U5868 ( .A1(n5143), .A2(n6420), .B1(n6379), .B2(n4724), .ZN(n4721)
         );
  AOI21_X1 U5869 ( .B1(n6416), .B2(n4726), .A(n4721), .ZN(n4723) );
  NAND2_X1 U5870 ( .A1(n4727), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4722) );
  OAI211_X1 U5871 ( .C1(n4730), .C2(n5232), .A(n4723), .B(n4722), .ZN(U3047)
         );
  OAI22_X1 U5872 ( .A1(n5143), .A2(n6449), .B1(n6399), .B2(n4724), .ZN(n4725)
         );
  AOI21_X1 U5873 ( .B1(n6442), .B2(n4726), .A(n4725), .ZN(n4729) );
  NAND2_X1 U5874 ( .A1(n4727), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4728) );
  OAI211_X1 U5875 ( .C1(n4730), .C2(n5262), .A(n4729), .B(n4728), .ZN(U3051)
         );
  OAI222_X1 U5876 ( .A1(n5095), .A2(n6226), .B1(n6224), .B2(n6641), .C1(n6225), 
        .C2(n6246), .ZN(U2885) );
  INV_X1 U5877 ( .A(n4731), .ZN(n4732) );
  NAND2_X1 U5878 ( .A1(n6188), .A2(n4732), .ZN(n4733) );
  AND2_X1 U5879 ( .A1(n4733), .A2(n5447), .ZN(n6163) );
  INV_X1 U5880 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6130) );
  NAND3_X1 U5881 ( .A1(n5321), .A2(n5447), .A3(n5872), .ZN(n6159) );
  OAI22_X1 U5882 ( .A1(n4734), .A2(n6134), .B1(n6196), .B2(n4874), .ZN(n4735)
         );
  AOI211_X1 U5883 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6173), 
        .B(n4735), .ZN(n4738) );
  INV_X1 U5884 ( .A(n4736), .ZN(n4737) );
  NAND2_X1 U5885 ( .A1(n6188), .A2(n4737), .ZN(n6156) );
  NOR2_X1 U5886 ( .A1(n6156), .A2(n6532), .ZN(n6129) );
  NAND2_X1 U5887 ( .A1(n6129), .A2(n6130), .ZN(n6155) );
  OAI211_X1 U5888 ( .C1(n6163), .C2(n6130), .A(n4738), .B(n6155), .ZN(n4739)
         );
  AOI21_X1 U5889 ( .B1(n6138), .B2(n5098), .A(n4739), .ZN(n4740) );
  OAI21_X1 U5890 ( .B1(n6150), .B2(n5095), .A(n4740), .ZN(U2821) );
  NOR2_X1 U5891 ( .A1(n6344), .A2(n4748), .ZN(n4788) );
  INV_X1 U5892 ( .A(n4788), .ZN(n4744) );
  AND2_X1 U5893 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4788), .ZN(n4779)
         );
  AOI21_X1 U5894 ( .B1(n4954), .B2(n4787), .A(n4779), .ZN(n4750) );
  NAND2_X1 U5895 ( .A1(n4750), .A2(n4741), .ZN(n4742) );
  NOR2_X1 U5896 ( .A1(n6353), .A2(n4742), .ZN(n4743) );
  AOI211_X2 U5897 ( .C1(n6353), .C2(n4744), .A(n4743), .B(n4700), .ZN(n4784)
         );
  INV_X1 U5898 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4753) );
  INV_X1 U5899 ( .A(n4745), .ZN(n4746) );
  OAI22_X1 U5900 ( .A1(n6391), .A2(n4945), .B1(n4825), .B2(n6438), .ZN(n4747)
         );
  AOI21_X1 U5901 ( .B1(n6434), .B2(n4779), .A(n4747), .ZN(n4752) );
  NAND2_X1 U5902 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4749) );
  OAI22_X1 U5903 ( .A1(n4750), .A2(n6353), .B1(n4749), .B2(n4748), .ZN(n4780)
         );
  NAND2_X1 U5904 ( .A1(n6435), .A2(n4780), .ZN(n4751) );
  OAI211_X1 U5905 ( .C1(n4784), .C2(n4753), .A(n4752), .B(n4751), .ZN(U3130)
         );
  INV_X1 U5906 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4757) );
  OAI22_X1 U5907 ( .A1(n6365), .A2(n4945), .B1(n4825), .B2(n5215), .ZN(n4754)
         );
  AOI21_X1 U5908 ( .B1(n6350), .B2(n4779), .A(n4754), .ZN(n4756) );
  NAND2_X1 U5909 ( .A1(n6351), .A2(n4780), .ZN(n4755) );
  OAI211_X1 U5910 ( .C1(n4784), .C2(n4757), .A(n4756), .B(n4755), .ZN(U3124)
         );
  INV_X1 U5911 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4761) );
  OAI22_X1 U5912 ( .A1(n6375), .A2(n4945), .B1(n4825), .B2(n6414), .ZN(n4758)
         );
  AOI21_X1 U5913 ( .B1(n6410), .B2(n4779), .A(n4758), .ZN(n4760) );
  NAND2_X1 U5914 ( .A1(n6411), .A2(n4780), .ZN(n4759) );
  OAI211_X1 U5915 ( .C1(n4784), .C2(n4761), .A(n4760), .B(n4759), .ZN(U3126)
         );
  INV_X1 U5916 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4765) );
  OAI22_X1 U5917 ( .A1(n6387), .A2(n4945), .B1(n4825), .B2(n6432), .ZN(n4762)
         );
  AOI21_X1 U5918 ( .B1(n6428), .B2(n4779), .A(n4762), .ZN(n4764) );
  NAND2_X1 U5919 ( .A1(n6429), .A2(n4780), .ZN(n4763) );
  OAI211_X1 U5920 ( .C1(n4784), .C2(n4765), .A(n4764), .B(n4763), .ZN(U3129)
         );
  INV_X1 U5921 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4769) );
  OAI22_X1 U5922 ( .A1(n6379), .A2(n4945), .B1(n4825), .B2(n6420), .ZN(n4766)
         );
  AOI21_X1 U5923 ( .B1(n6416), .B2(n4779), .A(n4766), .ZN(n4768) );
  NAND2_X1 U5924 ( .A1(n6417), .A2(n4780), .ZN(n4767) );
  OAI211_X1 U5925 ( .C1(n4784), .C2(n4769), .A(n4768), .B(n4767), .ZN(U3127)
         );
  INV_X1 U5926 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4773) );
  OAI22_X1 U5927 ( .A1(n6399), .A2(n4945), .B1(n4825), .B2(n6449), .ZN(n4770)
         );
  AOI21_X1 U5928 ( .B1(n6442), .B2(n4779), .A(n4770), .ZN(n4772) );
  NAND2_X1 U5929 ( .A1(n6444), .A2(n4780), .ZN(n4771) );
  OAI211_X1 U5930 ( .C1(n4784), .C2(n4773), .A(n4772), .B(n4771), .ZN(U3131)
         );
  INV_X1 U5931 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4777) );
  OAI22_X1 U5932 ( .A1(n6371), .A2(n4945), .B1(n4825), .B2(n5221), .ZN(n4774)
         );
  AOI21_X1 U5933 ( .B1(n3006), .B2(n4779), .A(n4774), .ZN(n4776) );
  NAND2_X1 U5934 ( .A1(n6367), .A2(n4780), .ZN(n4775) );
  OAI211_X1 U5935 ( .C1(n4784), .C2(n4777), .A(n4776), .B(n4775), .ZN(U3125)
         );
  INV_X1 U5936 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4783) );
  OAI22_X1 U5937 ( .A1(n6383), .A2(n4945), .B1(n4825), .B2(n6426), .ZN(n4778)
         );
  AOI21_X1 U5938 ( .B1(n6422), .B2(n4779), .A(n4778), .ZN(n4782) );
  NAND2_X1 U5939 ( .A1(n6423), .A2(n4780), .ZN(n4781) );
  OAI211_X1 U5940 ( .C1(n4784), .C2(n4783), .A(n4782), .B(n4781), .ZN(U3128)
         );
  AOI21_X1 U5941 ( .B1(n4826), .B2(n4825), .A(n6715), .ZN(n4785) );
  AOI211_X1 U5942 ( .C1(n4787), .C2(n4786), .A(n6353), .B(n4785), .ZN(n4792)
         );
  AND2_X1 U5943 ( .A1(n4951), .A2(n4788), .ZN(n4828) );
  INV_X1 U5944 ( .A(n4917), .ZN(n5203) );
  OR2_X1 U5945 ( .A1(n6345), .A2(n4789), .ZN(n5003) );
  AOI21_X1 U5946 ( .B1(n5003), .B2(STATE2_REG_2__SCAN_IN), .A(n4790), .ZN(
        n4998) );
  OAI211_X1 U5947 ( .C1(n6580), .C2(n4828), .A(n5203), .B(n4998), .ZN(n4791)
         );
  INV_X1 U5948 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4800) );
  OAI22_X1 U5949 ( .A1(n4826), .A2(n6426), .B1(n4825), .B2(n6383), .ZN(n4793)
         );
  AOI21_X1 U5950 ( .B1(n6422), .B2(n4828), .A(n4793), .ZN(n4799) );
  OR2_X1 U5951 ( .A1(n4794), .A2(n4995), .ZN(n4797) );
  INV_X1 U5952 ( .A(n5003), .ZN(n4795) );
  NAND2_X1 U5953 ( .A1(n4795), .A2(n6346), .ZN(n4796) );
  NAND2_X1 U5954 ( .A1(n4797), .A2(n4796), .ZN(n4829) );
  NAND2_X1 U5955 ( .A1(n6423), .A2(n4829), .ZN(n4798) );
  OAI211_X1 U5956 ( .C1(n4833), .C2(n4800), .A(n4799), .B(n4798), .ZN(U3120)
         );
  INV_X1 U5957 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4804) );
  OAI22_X1 U5958 ( .A1(n4826), .A2(n5221), .B1(n4825), .B2(n6371), .ZN(n4801)
         );
  AOI21_X1 U5959 ( .B1(n3007), .B2(n4828), .A(n4801), .ZN(n4803) );
  NAND2_X1 U5960 ( .A1(n6367), .A2(n4829), .ZN(n4802) );
  OAI211_X1 U5961 ( .C1(n4833), .C2(n4804), .A(n4803), .B(n4802), .ZN(U3117)
         );
  INV_X1 U5962 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4808) );
  OAI22_X1 U5963 ( .A1(n4826), .A2(n6449), .B1(n4825), .B2(n6399), .ZN(n4805)
         );
  AOI21_X1 U5964 ( .B1(n6442), .B2(n4828), .A(n4805), .ZN(n4807) );
  NAND2_X1 U5965 ( .A1(n6444), .A2(n4829), .ZN(n4806) );
  OAI211_X1 U5966 ( .C1(n4833), .C2(n4808), .A(n4807), .B(n4806), .ZN(U3123)
         );
  INV_X1 U5967 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4812) );
  OAI22_X1 U5968 ( .A1(n4826), .A2(n6420), .B1(n4825), .B2(n6379), .ZN(n4809)
         );
  AOI21_X1 U5969 ( .B1(n6416), .B2(n4828), .A(n4809), .ZN(n4811) );
  NAND2_X1 U5970 ( .A1(n6417), .A2(n4829), .ZN(n4810) );
  OAI211_X1 U5971 ( .C1(n4833), .C2(n4812), .A(n4811), .B(n4810), .ZN(U3119)
         );
  INV_X1 U5972 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4816) );
  OAI22_X1 U5973 ( .A1(n4826), .A2(n6432), .B1(n4825), .B2(n6387), .ZN(n4813)
         );
  AOI21_X1 U5974 ( .B1(n6428), .B2(n4828), .A(n4813), .ZN(n4815) );
  NAND2_X1 U5975 ( .A1(n6429), .A2(n4829), .ZN(n4814) );
  OAI211_X1 U5976 ( .C1(n4833), .C2(n4816), .A(n4815), .B(n4814), .ZN(U3121)
         );
  INV_X1 U5977 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4820) );
  OAI22_X1 U5978 ( .A1(n4826), .A2(n5215), .B1(n4825), .B2(n6365), .ZN(n4817)
         );
  AOI21_X1 U5979 ( .B1(n6350), .B2(n4828), .A(n4817), .ZN(n4819) );
  NAND2_X1 U5980 ( .A1(n6351), .A2(n4829), .ZN(n4818) );
  OAI211_X1 U5981 ( .C1(n4833), .C2(n4820), .A(n4819), .B(n4818), .ZN(U3116)
         );
  INV_X1 U5982 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4824) );
  OAI22_X1 U5983 ( .A1(n4826), .A2(n6438), .B1(n4825), .B2(n6391), .ZN(n4821)
         );
  AOI21_X1 U5984 ( .B1(n6434), .B2(n4828), .A(n4821), .ZN(n4823) );
  NAND2_X1 U5985 ( .A1(n6435), .A2(n4829), .ZN(n4822) );
  OAI211_X1 U5986 ( .C1(n4833), .C2(n4824), .A(n4823), .B(n4822), .ZN(U3122)
         );
  INV_X1 U5987 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4832) );
  OAI22_X1 U5988 ( .A1(n4826), .A2(n6414), .B1(n4825), .B2(n6375), .ZN(n4827)
         );
  AOI21_X1 U5989 ( .B1(n6410), .B2(n4828), .A(n4827), .ZN(n4831) );
  NAND2_X1 U5990 ( .A1(n6411), .A2(n4829), .ZN(n4830) );
  OAI211_X1 U5991 ( .C1(n4833), .C2(n4832), .A(n4831), .B(n4830), .ZN(U3118)
         );
  OR2_X1 U5992 ( .A1(n4994), .A2(n3003), .ZN(n4838) );
  INV_X1 U5993 ( .A(n4838), .ZN(n4880) );
  AOI22_X1 U5994 ( .A1(n4880), .A2(n5872), .B1(n4917), .B2(n3127), .ZN(n4870)
         );
  NAND3_X1 U5995 ( .A1(n6344), .A2(n6461), .A3(n6455), .ZN(n4884) );
  NOR2_X1 U5996 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4884), .ZN(n4867)
         );
  INV_X1 U5997 ( .A(n4867), .ZN(n4835) );
  AOI211_X1 U5998 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4835), .A(n6346), .B(
        n4834), .ZN(n4841) );
  NAND2_X1 U5999 ( .A1(n3640), .A2(n4961), .ZN(n4836) );
  INV_X1 U6000 ( .A(n4864), .ZN(n4837) );
  OAI21_X1 U6001 ( .B1(n4905), .B2(n4837), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4839) );
  NAND3_X1 U6002 ( .A1(n4839), .A2(n5872), .A3(n4838), .ZN(n4840) );
  NAND2_X1 U6003 ( .A1(n4863), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4844) );
  OAI22_X1 U6004 ( .A1(n4865), .A2(n6365), .B1(n5215), .B2(n4864), .ZN(n4842)
         );
  AOI21_X1 U6005 ( .B1(n6350), .B2(n4867), .A(n4842), .ZN(n4843) );
  OAI211_X1 U6006 ( .C1(n4870), .C2(n5218), .A(n4844), .B(n4843), .ZN(U3020)
         );
  NAND2_X1 U6007 ( .A1(n4863), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4847) );
  OAI22_X1 U6008 ( .A1(n4865), .A2(n6391), .B1(n6438), .B2(n4864), .ZN(n4845)
         );
  AOI21_X1 U6009 ( .B1(n6434), .B2(n4867), .A(n4845), .ZN(n4846) );
  OAI211_X1 U6010 ( .C1(n4870), .C2(n5246), .A(n4847), .B(n4846), .ZN(U3026)
         );
  NAND2_X1 U6011 ( .A1(n4863), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4850) );
  OAI22_X1 U6012 ( .A1(n4865), .A2(n6399), .B1(n6449), .B2(n4864), .ZN(n4848)
         );
  AOI21_X1 U6013 ( .B1(n6442), .B2(n4867), .A(n4848), .ZN(n4849) );
  OAI211_X1 U6014 ( .C1(n4870), .C2(n5262), .A(n4850), .B(n4849), .ZN(U3027)
         );
  NAND2_X1 U6015 ( .A1(n4863), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4853) );
  OAI22_X1 U6016 ( .A1(n4865), .A2(n6379), .B1(n6420), .B2(n4864), .ZN(n4851)
         );
  AOI21_X1 U6017 ( .B1(n6416), .B2(n4867), .A(n4851), .ZN(n4852) );
  OAI211_X1 U6018 ( .C1(n4870), .C2(n5232), .A(n4853), .B(n4852), .ZN(U3023)
         );
  NAND2_X1 U6019 ( .A1(n4863), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4856) );
  OAI22_X1 U6020 ( .A1(n4865), .A2(n6371), .B1(n5221), .B2(n4864), .ZN(n4854)
         );
  AOI21_X1 U6021 ( .B1(n3006), .B2(n4867), .A(n4854), .ZN(n4855) );
  OAI211_X1 U6022 ( .C1(n4870), .C2(n5224), .A(n4856), .B(n4855), .ZN(U3021)
         );
  NAND2_X1 U6023 ( .A1(n4863), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4859) );
  OAI22_X1 U6024 ( .A1(n4865), .A2(n6387), .B1(n6432), .B2(n4864), .ZN(n4857)
         );
  AOI21_X1 U6025 ( .B1(n6428), .B2(n4867), .A(n4857), .ZN(n4858) );
  OAI211_X1 U6026 ( .C1(n4870), .C2(n5254), .A(n4859), .B(n4858), .ZN(U3025)
         );
  NAND2_X1 U6027 ( .A1(n4863), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4862) );
  OAI22_X1 U6028 ( .A1(n4865), .A2(n6383), .B1(n6426), .B2(n4864), .ZN(n4860)
         );
  AOI21_X1 U6029 ( .B1(n6422), .B2(n4867), .A(n4860), .ZN(n4861) );
  OAI211_X1 U6030 ( .C1(n4870), .C2(n5250), .A(n4862), .B(n4861), .ZN(U3024)
         );
  NAND2_X1 U6031 ( .A1(n4863), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4869) );
  OAI22_X1 U6032 ( .A1(n4865), .A2(n6375), .B1(n6414), .B2(n4864), .ZN(n4866)
         );
  AOI21_X1 U6033 ( .B1(n6410), .B2(n4867), .A(n4866), .ZN(n4868) );
  OAI211_X1 U6034 ( .C1(n4870), .C2(n5228), .A(n4869), .B(n4868), .ZN(U3022)
         );
  XNOR2_X1 U6035 ( .A(n4871), .B(n4872), .ZN(n5100) );
  NAND2_X1 U6036 ( .A1(n4873), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4878)
         );
  NAND3_X1 U6037 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n5176) );
  NOR2_X1 U6038 ( .A1(n5176), .A2(n6311), .ZN(n4876) );
  OAI22_X1 U6039 ( .A1(n6335), .A2(n4874), .B1(n6130), .B2(n6323), .ZN(n4875)
         );
  AOI21_X1 U6040 ( .B1(n4876), .B2(n4154), .A(n4875), .ZN(n4877) );
  OAI211_X1 U6041 ( .C1(n5100), .C2(n5870), .A(n4878), .B(n4877), .ZN(U3012)
         );
  NOR2_X1 U6042 ( .A1(n4951), .A2(n4884), .ZN(n4879) );
  INV_X1 U6043 ( .A(n4879), .ZN(n4908) );
  AOI21_X1 U6044 ( .B1(n4880), .B2(n5063), .A(n4879), .ZN(n4886) );
  INV_X1 U6045 ( .A(n4888), .ZN(n4881) );
  AOI21_X1 U6046 ( .B1(n4881), .B2(STATEBS16_REG_SCAN_IN), .A(n6353), .ZN(
        n4883) );
  AOI22_X1 U6047 ( .A1(n4886), .A2(n4883), .B1(n6353), .B2(n4884), .ZN(n4882)
         );
  NAND2_X1 U6048 ( .A1(n4957), .A2(n4882), .ZN(n4904) );
  INV_X1 U6049 ( .A(n4883), .ZN(n4885) );
  OAI22_X1 U6050 ( .A1(n4886), .A2(n4885), .B1(n4641), .B2(n4884), .ZN(n4903)
         );
  AOI22_X1 U6051 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4904), .B1(n6367), 
        .B2(n4903), .ZN(n4890) );
  NOR2_X1 U6052 ( .A1(n4888), .A2(n4887), .ZN(n5120) );
  AOI22_X1 U6053 ( .A1(n5219), .A2(n5120), .B1(n4905), .B2(n6368), .ZN(n4889)
         );
  OAI211_X1 U6054 ( .C1(n6366), .C2(n4908), .A(n4890), .B(n4889), .ZN(U3029)
         );
  AOI22_X1 U6055 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4904), .B1(n6417), 
        .B2(n4903), .ZN(n4892) );
  INV_X1 U6056 ( .A(n6379), .ZN(n6415) );
  INV_X1 U6057 ( .A(n6420), .ZN(n6376) );
  AOI22_X1 U6058 ( .A1(n6415), .A2(n5120), .B1(n4905), .B2(n6376), .ZN(n4891)
         );
  OAI211_X1 U6059 ( .C1(n4968), .C2(n4908), .A(n4892), .B(n4891), .ZN(U3031)
         );
  AOI22_X1 U6060 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4904), .B1(n6444), 
        .B2(n4903), .ZN(n4894) );
  AOI22_X1 U6061 ( .A1(n6439), .A2(n5120), .B1(n4905), .B2(n6395), .ZN(n4893)
         );
  OAI211_X1 U6062 ( .C1(n4971), .C2(n4908), .A(n4894), .B(n4893), .ZN(U3035)
         );
  AOI22_X1 U6063 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4904), .B1(n6423), 
        .B2(n4903), .ZN(n4896) );
  AOI22_X1 U6064 ( .A1(n6421), .A2(n5120), .B1(n4905), .B2(n6380), .ZN(n4895)
         );
  OAI211_X1 U6065 ( .C1(n4980), .C2(n4908), .A(n4896), .B(n4895), .ZN(U3032)
         );
  AOI22_X1 U6066 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4904), .B1(n6429), 
        .B2(n4903), .ZN(n4898) );
  AOI22_X1 U6067 ( .A1(n6427), .A2(n5120), .B1(n4905), .B2(n6384), .ZN(n4897)
         );
  OAI211_X1 U6068 ( .C1(n4974), .C2(n4908), .A(n4898), .B(n4897), .ZN(U3033)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4904), .B1(n6435), 
        .B2(n4903), .ZN(n4900) );
  AOI22_X1 U6070 ( .A1(n6433), .A2(n5120), .B1(n4905), .B2(n6388), .ZN(n4899)
         );
  OAI211_X1 U6071 ( .C1(n4977), .C2(n4908), .A(n4900), .B(n4899), .ZN(U3034)
         );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4904), .B1(n6351), 
        .B2(n4903), .ZN(n4902) );
  AOI22_X1 U6073 ( .A1(n5213), .A2(n5120), .B1(n4905), .B2(n6362), .ZN(n4901)
         );
  OAI211_X1 U6074 ( .C1(n4990), .C2(n4908), .A(n4902), .B(n4901), .ZN(U3028)
         );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4904), .B1(n6411), 
        .B2(n4903), .ZN(n4907) );
  AOI22_X1 U6076 ( .A1(n6409), .A2(n5120), .B1(n4905), .B2(n6372), .ZN(n4906)
         );
  OAI211_X1 U6077 ( .C1(n4983), .C2(n4908), .A(n4907), .B(n4906), .ZN(U3030)
         );
  NAND2_X1 U6078 ( .A1(n4913), .A2(n5872), .ZN(n6348) );
  INV_X1 U6079 ( .A(n6348), .ZN(n4910) );
  INV_X1 U6080 ( .A(n6346), .ZN(n4999) );
  NOR2_X1 U6081 ( .A1(n4999), .A2(n6344), .ZN(n4909) );
  AOI22_X1 U6082 ( .A1(n4910), .A2(n3003), .B1(n6345), .B2(n4909), .ZN(n4950)
         );
  INV_X1 U6083 ( .A(n4945), .ZN(n4912) );
  INV_X1 U6084 ( .A(n4944), .ZN(n4911) );
  NOR3_X1 U6085 ( .A1(n4912), .A2(n4911), .A3(n6353), .ZN(n4915) );
  INV_X1 U6086 ( .A(n4913), .ZN(n4914) );
  OAI21_X1 U6087 ( .B1(n4915), .B2(n6356), .A(n4914), .ZN(n4921) );
  OAI21_X1 U6088 ( .B1(n6345), .B2(n4641), .A(n4916), .ZN(n5118) );
  NOR2_X1 U6089 ( .A1(n4917), .A2(n5118), .ZN(n6360) );
  NOR2_X1 U6090 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4918), .ZN(n4947)
         );
  INV_X1 U6091 ( .A(n4947), .ZN(n4919) );
  AOI21_X1 U6092 ( .B1(n4919), .B2(STATE2_REG_3__SCAN_IN), .A(n6344), .ZN(
        n4920) );
  NAND3_X1 U6093 ( .A1(n4921), .A2(n6360), .A3(n4920), .ZN(n4943) );
  NAND2_X1 U6094 ( .A1(n4943), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4924)
         );
  OAI22_X1 U6095 ( .A1(n4945), .A2(n6426), .B1(n6383), .B2(n4944), .ZN(n4922)
         );
  AOI21_X1 U6096 ( .B1(n6422), .B2(n4947), .A(n4922), .ZN(n4923) );
  OAI211_X1 U6097 ( .C1(n5250), .C2(n4950), .A(n4924), .B(n4923), .ZN(U3136)
         );
  NAND2_X1 U6098 ( .A1(n4943), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4927)
         );
  OAI22_X1 U6099 ( .A1(n4945), .A2(n6432), .B1(n6387), .B2(n4944), .ZN(n4925)
         );
  AOI21_X1 U6100 ( .B1(n6428), .B2(n4947), .A(n4925), .ZN(n4926) );
  OAI211_X1 U6101 ( .C1(n5254), .C2(n4950), .A(n4927), .B(n4926), .ZN(U3137)
         );
  NAND2_X1 U6102 ( .A1(n4943), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4930)
         );
  OAI22_X1 U6103 ( .A1(n4945), .A2(n6438), .B1(n6391), .B2(n4944), .ZN(n4928)
         );
  AOI21_X1 U6104 ( .B1(n6434), .B2(n4947), .A(n4928), .ZN(n4929) );
  OAI211_X1 U6105 ( .C1(n5246), .C2(n4950), .A(n4930), .B(n4929), .ZN(U3138)
         );
  NAND2_X1 U6106 ( .A1(n4943), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4933)
         );
  OAI22_X1 U6107 ( .A1(n4945), .A2(n5215), .B1(n6365), .B2(n4944), .ZN(n4931)
         );
  AOI21_X1 U6108 ( .B1(n6350), .B2(n4947), .A(n4931), .ZN(n4932) );
  OAI211_X1 U6109 ( .C1(n5218), .C2(n4950), .A(n4933), .B(n4932), .ZN(U3132)
         );
  NAND2_X1 U6110 ( .A1(n4943), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4936)
         );
  OAI22_X1 U6111 ( .A1(n4945), .A2(n5221), .B1(n6371), .B2(n4944), .ZN(n4934)
         );
  AOI21_X1 U6112 ( .B1(n3007), .B2(n4947), .A(n4934), .ZN(n4935) );
  OAI211_X1 U6113 ( .C1(n5224), .C2(n4950), .A(n4936), .B(n4935), .ZN(U3133)
         );
  NAND2_X1 U6114 ( .A1(n4943), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4939)
         );
  OAI22_X1 U6115 ( .A1(n4945), .A2(n6414), .B1(n6375), .B2(n4944), .ZN(n4937)
         );
  AOI21_X1 U6116 ( .B1(n6410), .B2(n4947), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6117 ( .C1(n5228), .C2(n4950), .A(n4939), .B(n4938), .ZN(U3134)
         );
  NAND2_X1 U6118 ( .A1(n4943), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4942)
         );
  OAI22_X1 U6119 ( .A1(n4945), .A2(n6420), .B1(n6379), .B2(n4944), .ZN(n4940)
         );
  AOI21_X1 U6120 ( .B1(n6416), .B2(n4947), .A(n4940), .ZN(n4941) );
  OAI211_X1 U6121 ( .C1(n5232), .C2(n4950), .A(n4942), .B(n4941), .ZN(U3135)
         );
  NAND2_X1 U6122 ( .A1(n4943), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4949)
         );
  OAI22_X1 U6123 ( .A1(n4945), .A2(n6449), .B1(n6399), .B2(n4944), .ZN(n4946)
         );
  AOI21_X1 U6124 ( .B1(n6442), .B2(n4947), .A(n4946), .ZN(n4948) );
  OAI211_X1 U6125 ( .C1(n5262), .C2(n4950), .A(n4949), .B(n4948), .ZN(U3139)
         );
  NAND3_X1 U6126 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6461), .A3(n6455), .ZN(n4997) );
  NOR2_X1 U6127 ( .A1(n4951), .A2(n4997), .ZN(n4952) );
  INV_X1 U6128 ( .A(n4952), .ZN(n4991) );
  INV_X1 U6129 ( .A(n4994), .ZN(n4953) );
  AOI21_X1 U6130 ( .B1(n4954), .B2(n4953), .A(n4952), .ZN(n4960) );
  NOR2_X1 U6131 ( .A1(n3001), .A2(n6715), .ZN(n4955) );
  AOI21_X1 U6132 ( .B1(n4962), .B2(n4955), .A(n6353), .ZN(n4958) );
  AOI22_X1 U6133 ( .A1(n4960), .A2(n4958), .B1(n6353), .B2(n4997), .ZN(n4956)
         );
  NAND2_X1 U6134 ( .A1(n4957), .A2(n4956), .ZN(n4987) );
  INV_X1 U6135 ( .A(n4958), .ZN(n4959) );
  OAI22_X1 U6136 ( .A1(n4960), .A2(n4959), .B1(n4641), .B2(n4997), .ZN(n4986)
         );
  AOI22_X1 U6137 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4987), .B1(n6417), 
        .B2(n4986), .ZN(n4967) );
  INV_X1 U6138 ( .A(n4963), .ZN(n4965) );
  AOI22_X1 U6139 ( .A1(n5026), .A2(n6376), .B1(n5206), .B2(n6415), .ZN(n4966)
         );
  OAI211_X1 U6140 ( .C1(n4991), .C2(n4968), .A(n4967), .B(n4966), .ZN(U3095)
         );
  AOI22_X1 U6141 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4987), .B1(n6444), 
        .B2(n4986), .ZN(n4970) );
  AOI22_X1 U6142 ( .A1(n5026), .A2(n6395), .B1(n5206), .B2(n6439), .ZN(n4969)
         );
  OAI211_X1 U6143 ( .C1(n4991), .C2(n4971), .A(n4970), .B(n4969), .ZN(U3099)
         );
  AOI22_X1 U6144 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4987), .B1(n6429), 
        .B2(n4986), .ZN(n4973) );
  AOI22_X1 U6145 ( .A1(n5026), .A2(n6384), .B1(n5206), .B2(n6427), .ZN(n4972)
         );
  OAI211_X1 U6146 ( .C1(n4991), .C2(n4974), .A(n4973), .B(n4972), .ZN(U3097)
         );
  AOI22_X1 U6147 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4987), .B1(n6435), 
        .B2(n4986), .ZN(n4976) );
  AOI22_X1 U6148 ( .A1(n5026), .A2(n6388), .B1(n5206), .B2(n6433), .ZN(n4975)
         );
  OAI211_X1 U6149 ( .C1(n4991), .C2(n4977), .A(n4976), .B(n4975), .ZN(U3098)
         );
  AOI22_X1 U6150 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4987), .B1(n6423), 
        .B2(n4986), .ZN(n4979) );
  AOI22_X1 U6151 ( .A1(n5026), .A2(n6380), .B1(n5206), .B2(n6421), .ZN(n4978)
         );
  OAI211_X1 U6152 ( .C1(n4991), .C2(n4980), .A(n4979), .B(n4978), .ZN(U3096)
         );
  AOI22_X1 U6153 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4987), .B1(n6411), 
        .B2(n4986), .ZN(n4982) );
  AOI22_X1 U6154 ( .A1(n5026), .A2(n6372), .B1(n5206), .B2(n6409), .ZN(n4981)
         );
  OAI211_X1 U6155 ( .C1(n4991), .C2(n4983), .A(n4982), .B(n4981), .ZN(U3094)
         );
  AOI22_X1 U6156 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4987), .B1(n6367), 
        .B2(n4986), .ZN(n4985) );
  AOI22_X1 U6157 ( .A1(n5026), .A2(n6368), .B1(n5206), .B2(n5219), .ZN(n4984)
         );
  OAI211_X1 U6158 ( .C1(n4991), .C2(n6366), .A(n4985), .B(n4984), .ZN(U3093)
         );
  AOI22_X1 U6159 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4987), .B1(n6351), 
        .B2(n4986), .ZN(n4989) );
  AOI22_X1 U6160 ( .A1(n5026), .A2(n6362), .B1(n5206), .B2(n5213), .ZN(n4988)
         );
  OAI211_X1 U6161 ( .C1(n4991), .C2(n4990), .A(n4989), .B(n4988), .ZN(U3092)
         );
  INV_X1 U6162 ( .A(n5026), .ZN(n4993) );
  NAND3_X1 U6163 ( .A1(n4993), .A2(n5872), .A3(n4992), .ZN(n4996) );
  NOR2_X1 U6164 ( .A1(n4995), .A2(n4994), .ZN(n5002) );
  AOI21_X1 U6165 ( .B1(n4996), .B2(n5113), .A(n5002), .ZN(n5001) );
  NOR2_X1 U6166 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4997), .ZN(n5027)
         );
  OAI211_X1 U6167 ( .C1(n6580), .C2(n5027), .A(n4999), .B(n4998), .ZN(n5000)
         );
  INV_X1 U6168 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U6169 ( .A1(n5026), .A2(n6433), .B1(n6388), .B2(n6401), .ZN(n5006)
         );
  INV_X1 U6170 ( .A(n5002), .ZN(n5004) );
  OAI22_X1 U6171 ( .A1(n5004), .A2(n6353), .B1(n5203), .B2(n5003), .ZN(n5028)
         );
  AOI22_X1 U6172 ( .A1(n6435), .A2(n5028), .B1(n6434), .B2(n5027), .ZN(n5005)
         );
  OAI211_X1 U6173 ( .C1(n5032), .C2(n5007), .A(n5006), .B(n5005), .ZN(U3090)
         );
  INV_X1 U6174 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U6175 ( .A1(n5026), .A2(n6409), .B1(n6372), .B2(n6401), .ZN(n5009)
         );
  AOI22_X1 U6176 ( .A1(n6411), .A2(n5028), .B1(n6410), .B2(n5027), .ZN(n5008)
         );
  OAI211_X1 U6177 ( .C1(n5032), .C2(n5010), .A(n5009), .B(n5008), .ZN(U3086)
         );
  INV_X1 U6178 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5013) );
  AOI22_X1 U6179 ( .A1(n5026), .A2(n6415), .B1(n6376), .B2(n6401), .ZN(n5012)
         );
  AOI22_X1 U6180 ( .A1(n6417), .A2(n5028), .B1(n6416), .B2(n5027), .ZN(n5011)
         );
  OAI211_X1 U6181 ( .C1(n5032), .C2(n5013), .A(n5012), .B(n5011), .ZN(U3087)
         );
  INV_X1 U6182 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5016) );
  AOI22_X1 U6183 ( .A1(n5026), .A2(n6439), .B1(n6395), .B2(n6401), .ZN(n5015)
         );
  AOI22_X1 U6184 ( .A1(n6444), .A2(n5028), .B1(n6442), .B2(n5027), .ZN(n5014)
         );
  OAI211_X1 U6185 ( .C1(n5032), .C2(n5016), .A(n5015), .B(n5014), .ZN(U3091)
         );
  INV_X1 U6186 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5019) );
  AOI22_X1 U6187 ( .A1(n5026), .A2(n6427), .B1(n6384), .B2(n6401), .ZN(n5018)
         );
  AOI22_X1 U6188 ( .A1(n6429), .A2(n5028), .B1(n6428), .B2(n5027), .ZN(n5017)
         );
  OAI211_X1 U6189 ( .C1(n5032), .C2(n5019), .A(n5018), .B(n5017), .ZN(U3089)
         );
  INV_X1 U6190 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5022) );
  AOI22_X1 U6191 ( .A1(n5026), .A2(n6421), .B1(n6380), .B2(n6401), .ZN(n5021)
         );
  AOI22_X1 U6192 ( .A1(n6423), .A2(n5028), .B1(n6422), .B2(n5027), .ZN(n5020)
         );
  OAI211_X1 U6193 ( .C1(n5032), .C2(n5022), .A(n5021), .B(n5020), .ZN(U3088)
         );
  INV_X1 U6194 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5025) );
  AOI22_X1 U6195 ( .A1(n5026), .A2(n5213), .B1(n6362), .B2(n6401), .ZN(n5024)
         );
  AOI22_X1 U6196 ( .A1(n6351), .A2(n5028), .B1(n6350), .B2(n5027), .ZN(n5023)
         );
  OAI211_X1 U6197 ( .C1(n5032), .C2(n5025), .A(n5024), .B(n5023), .ZN(U3084)
         );
  INV_X1 U6198 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6199 ( .A1(n5026), .A2(n5219), .B1(n6368), .B2(n6401), .ZN(n5030)
         );
  AOI22_X1 U6200 ( .A1(n6367), .A2(n5028), .B1(n3007), .B2(n5027), .ZN(n5029)
         );
  OAI211_X1 U6201 ( .C1(n5032), .C2(n5031), .A(n5030), .B(n5029), .ZN(U3085)
         );
  INV_X1 U6202 ( .A(n5033), .ZN(n5103) );
  AOI21_X1 U6203 ( .B1(n5034), .B2(n4682), .A(n5103), .ZN(n5108) );
  INV_X1 U6204 ( .A(n5108), .ZN(n6151) );
  OAI222_X1 U6205 ( .A1(n6151), .A2(n6226), .B1(n6224), .B2(n5035), .C1(n6225), 
        .C2(n3676), .ZN(U2884) );
  INV_X1 U6206 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5038) );
  AOI21_X1 U6207 ( .B1(n5037), .B2(n5036), .A(n5151), .ZN(n6146) );
  INV_X1 U6208 ( .A(n6146), .ZN(n6304) );
  OAI222_X1 U6209 ( .A1(n6151), .A2(n5533), .B1(n5038), .B2(n6210), .C1(n5530), 
        .C2(n6304), .ZN(U2852) );
  INV_X1 U6210 ( .A(n6182), .ZN(n5043) );
  INV_X1 U6211 ( .A(n5039), .ZN(n5040) );
  AOI21_X1 U6212 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5040), 
        .ZN(n5041) );
  OAI21_X1 U6213 ( .B1(n6271), .B2(n6186), .A(n5041), .ZN(n5042) );
  AOI21_X1 U6214 ( .B1(n5043), .B2(n6266), .A(n5042), .ZN(n5044) );
  OAI21_X1 U6215 ( .B1(n6060), .B2(n5045), .A(n5044), .ZN(U2982) );
  AOI21_X1 U6216 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5046), 
        .ZN(n5047) );
  OAI21_X1 U6217 ( .B1(n6271), .B2(n6167), .A(n5047), .ZN(n5048) );
  AOI21_X1 U6218 ( .B1(n6165), .B2(n6266), .A(n5048), .ZN(n5049) );
  OAI21_X1 U6219 ( .B1(n6060), .B2(n5050), .A(n5049), .ZN(U2981) );
  XOR2_X1 U6220 ( .A(n5051), .B(n5052), .Z(n6314) );
  INV_X1 U6221 ( .A(n6314), .ZN(n5058) );
  INV_X1 U6222 ( .A(n5093), .ZN(n5056) );
  NAND2_X1 U6223 ( .A1(n6279), .A2(REIP_REG_3__SCAN_IN), .ZN(n6309) );
  INV_X1 U6224 ( .A(n6309), .ZN(n5053) );
  AOI21_X1 U6225 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5053), 
        .ZN(n5054) );
  OAI21_X1 U6226 ( .B1(n6271), .B2(n5083), .A(n5054), .ZN(n5055) );
  AOI21_X1 U6227 ( .B1(n5056), .B2(n6266), .A(n5055), .ZN(n5057) );
  OAI21_X1 U6228 ( .B1(n5058), .B2(n6060), .A(n5057), .ZN(U2983) );
  NAND2_X1 U6229 ( .A1(n5380), .A2(n6054), .ZN(n5059) );
  NAND2_X1 U6230 ( .A1(n6150), .A2(n5059), .ZN(n6199) );
  INV_X1 U6231 ( .A(n5060), .ZN(n5061) );
  NAND2_X1 U6232 ( .A1(n5380), .A2(n5061), .ZN(n6168) );
  INV_X1 U6233 ( .A(n6168), .ZN(n6193) );
  AOI22_X1 U6234 ( .A1(n6193), .A2(n5063), .B1(n6178), .B2(n5062), .ZN(n5067)
         );
  NAND2_X1 U6235 ( .A1(n5925), .A2(REIP_REG_0__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6236 ( .A1(n6192), .A2(EBX_REG_0__SCAN_IN), .ZN(n5065) );
  OAI21_X1 U6237 ( .B1(n6191), .B2(n6138), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5064) );
  AND4_X1 U6238 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n5068)
         );
  OAI21_X1 U6239 ( .B1(n6181), .B2(n6282), .A(n5068), .ZN(U2827) );
  AOI22_X1 U6240 ( .A1(n6193), .A2(n3350), .B1(n6178), .B2(n4274), .ZN(n5073)
         );
  INV_X1 U6241 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5069) );
  AOI22_X1 U6242 ( .A1(n6188), .A2(n5069), .B1(n6192), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5072) );
  INV_X1 U6243 ( .A(n5447), .ZN(n6187) );
  AOI22_X1 U6244 ( .A1(n6191), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6187), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5071) );
  INV_X1 U6245 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6246 ( .A1(n6138), .A2(n5076), .ZN(n5070) );
  AND4_X1 U6247 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(n5074)
         );
  OAI21_X1 U6248 ( .B1(n5081), .B2(n6181), .A(n5074), .ZN(U2826) );
  OAI21_X1 U6249 ( .B1(n6276), .B2(n5076), .A(n5075), .ZN(n5079) );
  NOR2_X1 U6250 ( .A1(n5077), .A2(n6060), .ZN(n5078) );
  AOI211_X1 U6251 ( .C1(n5695), .C2(n5076), .A(n5079), .B(n5078), .ZN(n5080)
         );
  OAI21_X1 U6252 ( .B1(n6281), .B2(n5081), .A(n5080), .ZN(U2985) );
  NAND2_X1 U6253 ( .A1(n6188), .A2(n6175), .ZN(n5090) );
  NAND2_X1 U6254 ( .A1(n5090), .A2(n5447), .ZN(n6174) );
  NAND2_X1 U6255 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .ZN(
        n5089) );
  INV_X1 U6256 ( .A(n6310), .ZN(n5082) );
  AOI22_X1 U6257 ( .A1(n6193), .A2(n3003), .B1(n6178), .B2(n5082), .ZN(n5088)
         );
  INV_X1 U6258 ( .A(n5083), .ZN(n5084) );
  AOI22_X1 U6259 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6191), .B1(n6138), 
        .B2(n5084), .ZN(n5086) );
  NAND2_X1 U6260 ( .A1(n6192), .A2(EBX_REG_3__SCAN_IN), .ZN(n5085) );
  AND2_X1 U6261 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  OAI211_X1 U6262 ( .C1(n5090), .C2(n5089), .A(n5088), .B(n5087), .ZN(n5091)
         );
  AOI21_X1 U6263 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6174), .A(n5091), .ZN(n5092)
         );
  OAI21_X1 U6264 ( .B1(n5093), .B2(n6181), .A(n5092), .ZN(U2824) );
  OAI22_X1 U6265 ( .A1(n6276), .A2(n5094), .B1(n6323), .B2(n6130), .ZN(n5097)
         );
  NOR2_X1 U6266 ( .A1(n5095), .A2(n6281), .ZN(n5096) );
  AOI211_X1 U6267 ( .C1(n5695), .C2(n5098), .A(n5097), .B(n5096), .ZN(n5099)
         );
  OAI21_X1 U6268 ( .B1(n6060), .B2(n5100), .A(n5099), .ZN(U2980) );
  OAI21_X1 U6269 ( .B1(n5103), .B2(n3697), .A(n5102), .ZN(n5175) );
  INV_X1 U6270 ( .A(DATAI_8_), .ZN(n6636) );
  OAI222_X1 U6271 ( .A1(n5175), .A2(n6226), .B1(n6224), .B2(n6636), .C1(n6225), 
        .C2(n6243), .ZN(U2883) );
  XOR2_X1 U6272 ( .A(n5104), .B(n5105), .Z(n6306) );
  INV_X1 U6273 ( .A(n6306), .ZN(n5110) );
  NAND2_X1 U6274 ( .A1(n6279), .A2(REIP_REG_7__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U6275 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5106)
         );
  OAI211_X1 U6276 ( .C1(n6271), .C2(n6149), .A(n6303), .B(n5106), .ZN(n5107)
         );
  AOI21_X1 U6277 ( .B1(n5108), .B2(n6266), .A(n5107), .ZN(n5109) );
  OAI21_X1 U6278 ( .B1(n5110), .B2(n6060), .A(n5109), .ZN(U2979) );
  INV_X1 U6279 ( .A(n5115), .ZN(n5112) );
  NOR2_X1 U6280 ( .A1(n5203), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5111)
         );
  AOI22_X1 U6281 ( .A1(n5112), .A2(n5872), .B1(n6345), .B2(n5111), .ZN(n5149)
         );
  OAI21_X1 U6282 ( .B1(n5120), .B2(n5114), .A(n5113), .ZN(n5116) );
  AOI21_X1 U6283 ( .B1(n5116), .B2(n5115), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5119) );
  NOR2_X1 U6284 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5117), .ZN(n5146)
         );
  NOR2_X1 U6285 ( .A1(n6346), .A2(n5118), .ZN(n5212) );
  NAND2_X1 U6286 ( .A1(n5142), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5123) );
  OAI22_X1 U6287 ( .A1(n5144), .A2(n5221), .B1(n6371), .B2(n5143), .ZN(n5121)
         );
  AOI21_X1 U6288 ( .B1(n3007), .B2(n5146), .A(n5121), .ZN(n5122) );
  OAI211_X1 U6289 ( .C1(n5149), .C2(n5224), .A(n5123), .B(n5122), .ZN(U3037)
         );
  NAND2_X1 U6290 ( .A1(n5142), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5126) );
  OAI22_X1 U6291 ( .A1(n5144), .A2(n6432), .B1(n6387), .B2(n5143), .ZN(n5124)
         );
  AOI21_X1 U6292 ( .B1(n6428), .B2(n5146), .A(n5124), .ZN(n5125) );
  OAI211_X1 U6293 ( .C1(n5149), .C2(n5254), .A(n5126), .B(n5125), .ZN(U3041)
         );
  NAND2_X1 U6294 ( .A1(n5142), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5129) );
  OAI22_X1 U6295 ( .A1(n5144), .A2(n5215), .B1(n6365), .B2(n5143), .ZN(n5127)
         );
  AOI21_X1 U6296 ( .B1(n6350), .B2(n5146), .A(n5127), .ZN(n5128) );
  OAI211_X1 U6297 ( .C1(n5149), .C2(n5218), .A(n5129), .B(n5128), .ZN(U3036)
         );
  NAND2_X1 U6298 ( .A1(n5142), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5132) );
  OAI22_X1 U6299 ( .A1(n5144), .A2(n6426), .B1(n6383), .B2(n5143), .ZN(n5130)
         );
  AOI21_X1 U6300 ( .B1(n6422), .B2(n5146), .A(n5130), .ZN(n5131) );
  OAI211_X1 U6301 ( .C1(n5149), .C2(n5250), .A(n5132), .B(n5131), .ZN(U3040)
         );
  NAND2_X1 U6302 ( .A1(n5142), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5135) );
  OAI22_X1 U6303 ( .A1(n5144), .A2(n6449), .B1(n6399), .B2(n5143), .ZN(n5133)
         );
  AOI21_X1 U6304 ( .B1(n6442), .B2(n5146), .A(n5133), .ZN(n5134) );
  OAI211_X1 U6305 ( .C1(n5149), .C2(n5262), .A(n5135), .B(n5134), .ZN(U3043)
         );
  NAND2_X1 U6306 ( .A1(n5142), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5138) );
  OAI22_X1 U6307 ( .A1(n5144), .A2(n6438), .B1(n6391), .B2(n5143), .ZN(n5136)
         );
  AOI21_X1 U6308 ( .B1(n6434), .B2(n5146), .A(n5136), .ZN(n5137) );
  OAI211_X1 U6309 ( .C1(n5149), .C2(n5246), .A(n5138), .B(n5137), .ZN(U3042)
         );
  NAND2_X1 U6310 ( .A1(n5142), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5141) );
  OAI22_X1 U6311 ( .A1(n5144), .A2(n6420), .B1(n6379), .B2(n5143), .ZN(n5139)
         );
  AOI21_X1 U6312 ( .B1(n6416), .B2(n5146), .A(n5139), .ZN(n5140) );
  OAI211_X1 U6313 ( .C1(n5149), .C2(n5232), .A(n5141), .B(n5140), .ZN(U3039)
         );
  NAND2_X1 U6314 ( .A1(n5142), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5148) );
  OAI22_X1 U6315 ( .A1(n5144), .A2(n6414), .B1(n6375), .B2(n5143), .ZN(n5145)
         );
  AOI21_X1 U6316 ( .B1(n6410), .B2(n5146), .A(n5145), .ZN(n5147) );
  OAI211_X1 U6317 ( .C1(n5149), .C2(n5228), .A(n5148), .B(n5147), .ZN(U3038)
         );
  INV_X1 U6318 ( .A(n5175), .ZN(n6140) );
  INV_X1 U6319 ( .A(n5533), .ZN(n6207) );
  OR2_X1 U6320 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U6321 ( .A1(n5161), .A2(n5152), .ZN(n6133) );
  OAI22_X1 U6322 ( .A1(n6133), .A2(n5530), .B1(n6135), .B2(n6210), .ZN(n5153)
         );
  AOI21_X1 U6323 ( .B1(n6140), .B2(n6207), .A(n5153), .ZN(n5154) );
  INV_X1 U6324 ( .A(n5154), .ZN(U2851) );
  AND2_X1 U6325 ( .A1(n5102), .A2(n5155), .ZN(n5157) );
  OR2_X1 U6326 ( .A1(n5157), .A2(n5156), .ZN(n5193) );
  NOR2_X1 U6327 ( .A1(n6187), .A2(n5163), .ZN(n5273) );
  NOR2_X1 U6328 ( .A1(n5438), .A2(n5273), .ZN(n6132) );
  AOI22_X1 U6329 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6192), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6132), .ZN(n5158) );
  OAI211_X1 U6330 ( .C1(n6170), .C2(n5159), .A(n5158), .B(n6159), .ZN(n5167)
         );
  NAND2_X1 U6331 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  NAND2_X1 U6332 ( .A1(n5198), .A2(n5162), .ZN(n6291) );
  INV_X1 U6333 ( .A(n5189), .ZN(n5164) );
  NOR2_X1 U6334 ( .A1(n6077), .A2(n5163), .ZN(n5275) );
  INV_X1 U6335 ( .A(n5275), .ZN(n6103) );
  NOR2_X1 U6336 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6103), .ZN(n6124) );
  AOI21_X1 U6337 ( .B1(n6138), .B2(n5164), .A(n6124), .ZN(n5165) );
  OAI21_X1 U6338 ( .B1(n6196), .B2(n6291), .A(n5165), .ZN(n5166) );
  NOR2_X1 U6339 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  OAI21_X1 U6340 ( .B1(n6150), .B2(n5193), .A(n5168), .ZN(U2818) );
  INV_X1 U6341 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5169) );
  OAI222_X1 U6342 ( .A1(n5193), .A2(n5533), .B1(n5169), .B2(n6210), .C1(n5530), 
        .C2(n6291), .ZN(U2850) );
  INV_X1 U6343 ( .A(DATAI_9_), .ZN(n6722) );
  OAI222_X1 U6344 ( .A1(n5193), .A2(n6226), .B1(n6224), .B2(n6722), .C1(n6225), 
        .C2(n6241), .ZN(U2882) );
  XOR2_X1 U6345 ( .A(n5170), .B(n5171), .Z(n5180) );
  NAND2_X1 U6346 ( .A1(n5180), .A2(n6278), .ZN(n5174) );
  AND2_X1 U6347 ( .A1(n6279), .A2(REIP_REG_8__SCAN_IN), .ZN(n5183) );
  AND2_X1 U6348 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5172)
         );
  AOI211_X1 U6349 ( .C1(n5695), .C2(n6137), .A(n5183), .B(n5172), .ZN(n5173)
         );
  OAI211_X1 U6350 ( .C1(n6281), .C2(n5175), .A(n5174), .B(n5173), .ZN(U2978)
         );
  NOR2_X1 U6351 ( .A1(n4154), .A2(n5176), .ZN(n5707) );
  INV_X1 U6352 ( .A(n5707), .ZN(n5181) );
  OAI21_X1 U6353 ( .B1(n5181), .B2(n5177), .A(n5823), .ZN(n5178) );
  INV_X1 U6354 ( .A(n5178), .ZN(n5179) );
  NOR2_X1 U6355 ( .A1(n6317), .A2(n5179), .ZN(n6308) );
  NAND2_X1 U6356 ( .A1(n5180), .A2(n6337), .ZN(n5186) );
  NOR2_X1 U6357 ( .A1(n5181), .A2(n6311), .ZN(n6300) );
  NOR2_X1 U6358 ( .A1(n6301), .A2(n4159), .ZN(n5706) );
  AOI21_X1 U6359 ( .B1(n6301), .B2(n4159), .A(n5706), .ZN(n5184) );
  NOR2_X1 U6360 ( .A1(n6133), .A2(n6335), .ZN(n5182) );
  AOI211_X1 U6361 ( .C1(n6300), .C2(n5184), .A(n5183), .B(n5182), .ZN(n5185)
         );
  OAI211_X1 U6362 ( .C1(n6308), .C2(n4159), .A(n5186), .B(n5185), .ZN(U3010)
         );
  XNOR2_X1 U6363 ( .A(n2990), .B(n5239), .ZN(n5188) );
  XNOR2_X1 U6364 ( .A(n2992), .B(n5188), .ZN(n6296) );
  NAND2_X1 U6365 ( .A1(n6296), .A2(n6278), .ZN(n5192) );
  NOR2_X1 U6366 ( .A1(n6323), .A2(n6537), .ZN(n6292) );
  NOR2_X1 U6367 ( .A1(n6271), .A2(n5189), .ZN(n5190) );
  AOI211_X1 U6368 ( .C1(n6262), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6292), 
        .B(n5190), .ZN(n5191) );
  OAI211_X1 U6369 ( .C1(n6281), .C2(n5193), .A(n5192), .B(n5191), .ZN(U2977)
         );
  NOR2_X1 U6370 ( .A1(n5156), .A2(n5195), .ZN(n5196) );
  OR2_X1 U6371 ( .A1(n5194), .A2(n5196), .ZN(n6121) );
  AOI22_X1 U6372 ( .A1(n6220), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6216), .ZN(n5197) );
  OAI21_X1 U6373 ( .B1(n6121), .B2(n6226), .A(n5197), .ZN(U2881) );
  INV_X1 U6374 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5201) );
  AOI21_X1 U6375 ( .B1(n5199), .B2(n5198), .A(n5269), .ZN(n5200) );
  INV_X1 U6376 ( .A(n5200), .ZN(n6118) );
  OAI222_X1 U6377 ( .A1(n6121), .A2(n5533), .B1(n5201), .B2(n6210), .C1(n5530), 
        .C2(n6118), .ZN(U2849) );
  OAI21_X1 U6378 ( .B1(n5206), .B2(n5256), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5202) );
  NOR2_X1 U6379 ( .A1(n5203), .A2(n6344), .ZN(n5204) );
  NOR2_X1 U6380 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5205), .ZN(n5260)
         );
  INV_X1 U6381 ( .A(n5207), .ZN(n5209) );
  INV_X1 U6382 ( .A(n5260), .ZN(n5208) );
  AOI22_X1 U6383 ( .A1(n5210), .A2(n5209), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5208), .ZN(n5211) );
  OAI211_X1 U6384 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4641), .A(n5212), .B(n5211), .ZN(n5255) );
  AOI22_X1 U6385 ( .A1(n5256), .A2(n5213), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5255), .ZN(n5214) );
  OAI21_X1 U6386 ( .B1(n5258), .B2(n5215), .A(n5214), .ZN(n5216) );
  AOI21_X1 U6387 ( .B1(n6350), .B2(n5260), .A(n5216), .ZN(n5217) );
  OAI21_X1 U6388 ( .B1(n5263), .B2(n5218), .A(n5217), .ZN(U3100) );
  AOI22_X1 U6389 ( .A1(n5256), .A2(n5219), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5255), .ZN(n5220) );
  OAI21_X1 U6390 ( .B1(n5258), .B2(n5221), .A(n5220), .ZN(n5222) );
  AOI21_X1 U6391 ( .B1(n3006), .B2(n5260), .A(n5222), .ZN(n5223) );
  OAI21_X1 U6392 ( .B1(n5263), .B2(n5224), .A(n5223), .ZN(U3101) );
  AOI22_X1 U6393 ( .A1(n5256), .A2(n6409), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5255), .ZN(n5225) );
  OAI21_X1 U6394 ( .B1(n5258), .B2(n6414), .A(n5225), .ZN(n5226) );
  AOI21_X1 U6395 ( .B1(n6410), .B2(n5260), .A(n5226), .ZN(n5227) );
  OAI21_X1 U6396 ( .B1(n5263), .B2(n5228), .A(n5227), .ZN(U3102) );
  AOI22_X1 U6397 ( .A1(n5256), .A2(n6415), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5255), .ZN(n5229) );
  OAI21_X1 U6398 ( .B1(n5258), .B2(n6420), .A(n5229), .ZN(n5230) );
  AOI21_X1 U6399 ( .B1(n6416), .B2(n5260), .A(n5230), .ZN(n5231) );
  OAI21_X1 U6400 ( .B1(n5263), .B2(n5232), .A(n5231), .ZN(U3103) );
  INV_X1 U6401 ( .A(n5234), .ZN(n5236) );
  NAND2_X1 U6402 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  XNOR2_X1 U6403 ( .A(n5233), .B(n5237), .ZN(n5290) );
  OAI21_X1 U6404 ( .B1(n5844), .B2(n5706), .A(n6308), .ZN(n6295) );
  OAI22_X1 U6405 ( .A1(n6118), .A2(n6335), .B1(n6540), .B2(n6323), .ZN(n5241)
         );
  NAND2_X1 U6406 ( .A1(n5706), .A2(n6300), .ZN(n6299) );
  AOI221_X1 U6407 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5239), .C2(n5238), .A(n6299), 
        .ZN(n5240) );
  AOI211_X1 U6408 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6295), .A(n5241), .B(n5240), .ZN(n5242) );
  OAI21_X1 U6409 ( .B1(n5870), .B2(n5290), .A(n5242), .ZN(U3008) );
  AOI22_X1 U6410 ( .A1(n5256), .A2(n6433), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5255), .ZN(n5243) );
  OAI21_X1 U6411 ( .B1(n5258), .B2(n6438), .A(n5243), .ZN(n5244) );
  AOI21_X1 U6412 ( .B1(n6434), .B2(n5260), .A(n5244), .ZN(n5245) );
  OAI21_X1 U6413 ( .B1(n5263), .B2(n5246), .A(n5245), .ZN(U3106) );
  AOI22_X1 U6414 ( .A1(n5256), .A2(n6421), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5255), .ZN(n5247) );
  OAI21_X1 U6415 ( .B1(n5258), .B2(n6426), .A(n5247), .ZN(n5248) );
  AOI21_X1 U6416 ( .B1(n6422), .B2(n5260), .A(n5248), .ZN(n5249) );
  OAI21_X1 U6417 ( .B1(n5263), .B2(n5250), .A(n5249), .ZN(U3104) );
  AOI22_X1 U6418 ( .A1(n5256), .A2(n6427), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5255), .ZN(n5251) );
  OAI21_X1 U6419 ( .B1(n5258), .B2(n6432), .A(n5251), .ZN(n5252) );
  AOI21_X1 U6420 ( .B1(n6428), .B2(n5260), .A(n5252), .ZN(n5253) );
  OAI21_X1 U6421 ( .B1(n5263), .B2(n5254), .A(n5253), .ZN(U3105) );
  AOI22_X1 U6422 ( .A1(n5256), .A2(n6439), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5255), .ZN(n5257) );
  OAI21_X1 U6423 ( .B1(n5258), .B2(n6449), .A(n5257), .ZN(n5259) );
  AOI21_X1 U6424 ( .B1(n6442), .B2(n5260), .A(n5259), .ZN(n5261) );
  OAI21_X1 U6425 ( .B1(n5263), .B2(n5262), .A(n5261), .ZN(U3107) );
  NOR2_X1 U6426 ( .A1(n5194), .A2(n5266), .ZN(n5267) );
  OR2_X1 U6427 ( .A1(n5265), .A2(n5267), .ZN(n5705) );
  INV_X1 U6428 ( .A(n5294), .ZN(n5268) );
  OAI21_X1 U6429 ( .B1(n5270), .B2(n5269), .A(n5268), .ZN(n5282) );
  INV_X1 U6430 ( .A(n5282), .ZN(n6284) );
  AOI22_X1 U6431 ( .A1(n6284), .A2(n6206), .B1(EBX_REG_11__SCAN_IN), .B2(n5528), .ZN(n5271) );
  OAI21_X1 U6432 ( .B1(n5705), .B2(n5533), .A(n5271), .ZN(U2848) );
  AOI22_X1 U6433 ( .A1(n6220), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6216), .ZN(n5272) );
  OAI21_X1 U6434 ( .B1(n5705), .B2(n6226), .A(n5272), .ZN(U2880) );
  AOI21_X1 U6435 ( .B1(n5274), .B2(n5273), .A(n5438), .ZN(n6112) );
  NAND2_X1 U6436 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5275), .ZN(n6119) );
  OAI21_X1 U6437 ( .B1(n6540), .B2(n6119), .A(n5276), .ZN(n5284) );
  INV_X1 U6438 ( .A(n5701), .ZN(n5280) );
  INV_X1 U6439 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5278) );
  OAI22_X1 U6440 ( .A1(n5278), .A2(n6134), .B1(n5277), .B2(n6170), .ZN(n5279)
         );
  AOI211_X1 U6441 ( .C1(n6138), .C2(n5280), .A(n5279), .B(n6173), .ZN(n5281)
         );
  OAI21_X1 U6442 ( .B1(n5282), .B2(n6196), .A(n5281), .ZN(n5283) );
  AOI21_X1 U6443 ( .B1(n6112), .B2(n5284), .A(n5283), .ZN(n5285) );
  OAI21_X1 U6444 ( .B1(n5705), .B2(n6150), .A(n5285), .ZN(U2816) );
  AOI22_X1 U6445 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6279), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6446 ( .A1(n5695), .A2(n6122), .ZN(n5286) );
  OAI211_X1 U6447 ( .C1(n6121), .C2(n6281), .A(n5287), .B(n5286), .ZN(n5288)
         );
  INV_X1 U6448 ( .A(n5288), .ZN(n5289) );
  OAI21_X1 U6449 ( .B1(n5290), .B2(n6060), .A(n5289), .ZN(U2976) );
  OAI21_X1 U6450 ( .B1(n5265), .B2(n5292), .A(n5291), .ZN(n6113) );
  INV_X1 U6451 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5296) );
  OR2_X1 U6452 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  NAND2_X1 U6453 ( .A1(n5859), .A2(n5295), .ZN(n6109) );
  OAI222_X1 U6454 ( .A1(n6113), .A2(n5533), .B1(n5296), .B2(n6210), .C1(n5530), 
        .C2(n6109), .ZN(U2847) );
  INV_X1 U6455 ( .A(DATAI_12_), .ZN(n5298) );
  OAI222_X1 U6456 ( .A1(n6113), .A2(n6226), .B1(n5298), .B2(n6224), .C1(n5297), 
        .C2(n6225), .ZN(U2879) );
  INV_X1 U6457 ( .A(n5299), .ZN(n5303) );
  INV_X1 U6458 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5731) );
  AOI22_X1 U6459 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5731), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5300), .ZN(n5889) );
  NOR2_X1 U6460 ( .A1(n5321), .A2(n6342), .ZN(n5888) );
  INV_X1 U6461 ( .A(n5888), .ZN(n5322) );
  NAND3_X1 U6462 ( .A1(n5891), .A2(n4409), .A3(n5305), .ZN(n5301) );
  OAI21_X1 U6463 ( .B1(n5889), .B2(n5322), .A(n5301), .ZN(n5302) );
  AOI21_X1 U6464 ( .B1(n5303), .B2(n6045), .A(n5302), .ZN(n5307) );
  INV_X1 U6465 ( .A(n5304), .ZN(n6578) );
  OAI22_X1 U6466 ( .A1(n6459), .A2(n6498), .B1(n6578), .B2(n6709), .ZN(n6044)
         );
  AOI21_X1 U6467 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n3053), .A(n6044), .ZN(
        n5893) );
  AOI21_X1 U6468 ( .B1(n5891), .B2(n5882), .A(n5893), .ZN(n5306) );
  OAI22_X1 U6469 ( .A1(n5307), .A2(n5893), .B1(n5306), .B2(n5305), .ZN(U3459)
         );
  NAND2_X1 U6470 ( .A1(n5390), .A2(n5308), .ZN(n5313) );
  AOI22_X1 U6471 ( .A1(n5310), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5309), .ZN(n5311) );
  INV_X1 U6472 ( .A(n5311), .ZN(n5312) );
  XNOR2_X2 U6473 ( .A(n5313), .B(n5312), .ZN(n5569) );
  NAND3_X1 U6474 ( .A1(n5569), .A2(n5314), .A3(n6225), .ZN(n5316) );
  AOI22_X1 U6475 ( .A1(n6214), .A2(DATAI_31_), .B1(n6216), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6476 ( .A1(n5316), .A2(n5315), .ZN(U2860) );
  INV_X1 U6477 ( .A(n5886), .ZN(n5317) );
  OR2_X1 U6478 ( .A1(n3629), .A2(n5317), .ZN(n5320) );
  NAND2_X1 U6479 ( .A1(n5318), .A2(n3036), .ZN(n5319) );
  AND2_X1 U6480 ( .A1(n5320), .A2(n5319), .ZN(n6451) );
  OAI21_X1 U6481 ( .B1(n6451), .B2(STATE2_REG_3__SCAN_IN), .A(n5321), .ZN(
        n5323) );
  AOI22_X1 U6482 ( .A1(n5323), .A2(n5322), .B1(n5891), .B2(n3036), .ZN(n5326)
         );
  AOI21_X1 U6483 ( .B1(n5324), .B2(n6045), .A(n5893), .ZN(n5325) );
  OAI22_X1 U6484 ( .A1(n5326), .A2(n5893), .B1(n5325), .B2(n3036), .ZN(U3461)
         );
  NAND3_X1 U6485 ( .A1(n5424), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6486 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5383) );
  INV_X1 U6487 ( .A(n5383), .ZN(n5333) );
  INV_X1 U6488 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6669) );
  INV_X1 U6489 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6731) );
  INV_X1 U6490 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6653) );
  NOR3_X1 U6491 ( .A1(n6669), .A2(n6731), .A3(n6653), .ZN(n5329) );
  AOI21_X1 U6492 ( .B1(n5330), .B2(n5329), .A(n5438), .ZN(n5905) );
  AND2_X1 U6493 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5331) );
  NOR2_X1 U6494 ( .A1(n6077), .A2(n5331), .ZN(n5332) );
  OR2_X1 U6495 ( .A1(n5905), .A2(n5332), .ZN(n5402) );
  INV_X1 U6496 ( .A(n5402), .ZN(n5417) );
  OAI21_X1 U6497 ( .B1(n5405), .B2(n5333), .A(n5417), .ZN(n5386) );
  INV_X1 U6498 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6719) );
  INV_X1 U6499 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6573) );
  OAI21_X1 U6500 ( .B1(n5405), .B2(n6719), .A(n6573), .ZN(n5364) );
  INV_X1 U6501 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5368) );
  AOI22_X1 U6502 ( .A1(n5334), .A2(n6138), .B1(n6191), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5335) );
  OAI21_X1 U6503 ( .B1(n6134), .B2(n5368), .A(n5335), .ZN(n5363) );
  MUX2_X1 U6504 ( .A(n5336), .B(n4168), .S(EBX_REG_24__SCAN_IN), .Z(n5338) );
  NAND2_X1 U6505 ( .A1(n2997), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6506 ( .A1(n5338), .A2(n5337), .ZN(n5489) );
  MUX2_X1 U6507 ( .A(n5345), .B(n5392), .S(EBX_REG_25__SCAN_IN), .Z(n5341) );
  OR2_X1 U6508 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5340)
         );
  AND2_X1 U6509 ( .A1(n5341), .A2(n5340), .ZN(n5483) );
  INV_X1 U6510 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U6511 ( .A1(n5372), .A2(n5908), .ZN(n5344) );
  INV_X1 U6512 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6513 ( .A1(n4168), .A2(n5598), .ZN(n5342) );
  OAI211_X1 U6514 ( .C1(n2997), .C2(EBX_REG_26__SCAN_IN), .A(n5342), .B(n5392), 
        .ZN(n5343) );
  AND2_X1 U6515 ( .A1(n5344), .A2(n5343), .ZN(n5474) );
  MUX2_X1 U6516 ( .A(n5345), .B(n5392), .S(EBX_REG_27__SCAN_IN), .Z(n5347) );
  OR2_X1 U6517 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5346)
         );
  NAND2_X1 U6518 ( .A1(n5347), .A2(n5346), .ZN(n5421) );
  INV_X1 U6519 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6520 ( .A1(n5372), .A2(n5348), .ZN(n5352) );
  NAND2_X1 U6521 ( .A1(n4168), .A2(n5349), .ZN(n5350) );
  OAI211_X1 U6522 ( .C1(n2998), .C2(EBX_REG_28__SCAN_IN), .A(n5350), .B(n5392), 
        .ZN(n5351) );
  NOR2_X1 U6523 ( .A1(n2998), .A2(EBX_REG_29__SCAN_IN), .ZN(n5353) );
  AOI21_X1 U6524 ( .B1(n5354), .B2(n3548), .A(n5353), .ZN(n5393) );
  INV_X1 U6525 ( .A(n5370), .ZN(n5358) );
  NAND2_X1 U6526 ( .A1(n5369), .A2(EBX_REG_30__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6527 ( .A1(n2998), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5355) );
  AND2_X1 U6528 ( .A1(n5356), .A2(n5355), .ZN(n5376) );
  INV_X1 U6529 ( .A(n5376), .ZN(n5357) );
  NOR2_X1 U6530 ( .A1(n5370), .A2(n3097), .ZN(n5375) );
  AOI211_X1 U6531 ( .C1(n5411), .C2(n5358), .A(n5357), .B(n5375), .ZN(n5361)
         );
  INV_X1 U6532 ( .A(n5411), .ZN(n5359) );
  NOR2_X1 U6533 ( .A1(n5741), .A2(n6196), .ZN(n5362) );
  AOI211_X1 U6534 ( .C1(n5386), .C2(n5364), .A(n5363), .B(n5362), .ZN(n5365)
         );
  OAI21_X1 U6535 ( .B1(n5327), .B2(n6150), .A(n5365), .ZN(U2797) );
  AOI22_X1 U6536 ( .A1(n6214), .A2(DATAI_30_), .B1(n6216), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6537 ( .A1(n6217), .A2(DATAI_14_), .ZN(n5366) );
  OAI211_X1 U6538 ( .C1(n5327), .C2(n6226), .A(n5367), .B(n5366), .ZN(U2861)
         );
  OAI222_X1 U6539 ( .A1(n5533), .A2(n5327), .B1(n5530), .B2(n5741), .C1(n5368), 
        .C2(n6210), .ZN(U2829) );
  OAI22_X1 U6540 ( .A1(n5369), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n2997), .ZN(n5378) );
  NAND2_X1 U6541 ( .A1(n5370), .A2(n5392), .ZN(n5374) );
  INV_X1 U6542 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5371) );
  AND2_X1 U6543 ( .A1(n5372), .A2(n5371), .ZN(n5394) );
  NAND2_X1 U6544 ( .A1(n5411), .A2(n5394), .ZN(n5373) );
  NAND2_X1 U6545 ( .A1(n5374), .A2(n5373), .ZN(n5399) );
  NAND2_X1 U6546 ( .A1(n5569), .A2(n6139), .ZN(n5388) );
  INV_X1 U6547 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5382) );
  NAND3_X1 U6548 ( .A1(n5380), .A2(EBX_REG_31__SCAN_IN), .A3(n5379), .ZN(n5381) );
  OAI21_X1 U6549 ( .B1(n6170), .B2(n5382), .A(n5381), .ZN(n5385) );
  NOR3_X1 U6550 ( .A1(n5405), .A2(REIP_REG_31__SCAN_IN), .A3(n5383), .ZN(n5384) );
  AOI211_X1 U6551 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5386), .A(n5385), .B(n5384), .ZN(n5387) );
  OAI211_X1 U6552 ( .C1(n5735), .C2(n6196), .A(n5388), .B(n5387), .ZN(U2796)
         );
  INV_X1 U6553 ( .A(n5577), .ZN(n5536) );
  NAND2_X1 U6554 ( .A1(n5393), .A2(n5392), .ZN(n5396) );
  INV_X1 U6555 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U6556 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NOR2_X1 U6557 ( .A1(n5411), .A2(n5397), .ZN(n5398) );
  NOR2_X1 U6558 ( .A1(n5399), .A2(n5398), .ZN(n5750) );
  OAI22_X1 U6559 ( .A1(n5400), .A2(n6170), .B1(n6201), .B2(n5575), .ZN(n5401)
         );
  AOI21_X1 U6560 ( .B1(n6192), .B2(EBX_REG_29__SCAN_IN), .A(n5401), .ZN(n5404)
         );
  NAND2_X1 U6561 ( .A1(n5402), .A2(REIP_REG_29__SCAN_IN), .ZN(n5403) );
  OAI211_X1 U6562 ( .C1(n5405), .C2(REIP_REG_29__SCAN_IN), .A(n5404), .B(n5403), .ZN(n5406) );
  AOI21_X1 U6563 ( .B1(n5750), .B2(n6178), .A(n5406), .ZN(n5407) );
  OAI21_X1 U6564 ( .B1(n5536), .B2(n6150), .A(n5407), .ZN(U2798) );
  AOI21_X1 U6565 ( .B1(n3030), .B2(n3066), .A(n5411), .ZN(n5760) );
  INV_X1 U6566 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6706) );
  NAND3_X1 U6567 ( .A1(n5424), .A2(REIP_REG_27__SCAN_IN), .A3(n6706), .ZN(
        n5416) );
  INV_X1 U6568 ( .A(n5412), .ZN(n5585) );
  OAI22_X1 U6569 ( .A1(n5413), .A2(n6170), .B1(n6201), .B2(n5585), .ZN(n5414)
         );
  AOI21_X1 U6570 ( .B1(n6192), .B2(EBX_REG_28__SCAN_IN), .A(n5414), .ZN(n5415)
         );
  OAI211_X1 U6571 ( .C1(n5417), .C2(n6706), .A(n5416), .B(n5415), .ZN(n5418)
         );
  AOI21_X1 U6572 ( .B1(n5760), .B2(n6178), .A(n5418), .ZN(n5419) );
  OAI21_X1 U6573 ( .B1(n5583), .B2(n6150), .A(n5419), .ZN(U2799) );
  AOI21_X1 U6574 ( .B1(n5420), .B2(n2980), .A(n5408), .ZN(n5596) );
  INV_X1 U6575 ( .A(n5596), .ZN(n5541) );
  AND2_X1 U6576 ( .A1(n3022), .A2(n5421), .ZN(n5423) );
  OR2_X1 U6577 ( .A1(n5423), .A2(n5422), .ZN(n5472) );
  INV_X1 U6578 ( .A(n5472), .ZN(n5765) );
  INV_X1 U6579 ( .A(n5424), .ZN(n5428) );
  AOI22_X1 U6580 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6191), .ZN(n5425) );
  OAI21_X1 U6581 ( .B1(n5594), .B2(n6201), .A(n5425), .ZN(n5426) );
  AOI21_X1 U6582 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5905), .A(n5426), .ZN(n5427) );
  OAI21_X1 U6583 ( .B1(n5428), .B2(REIP_REG_27__SCAN_IN), .A(n5427), .ZN(n5429) );
  AOI21_X1 U6584 ( .B1(n5765), .B2(n6178), .A(n5429), .ZN(n5430) );
  OAI21_X1 U6585 ( .B1(n5541), .B2(n6150), .A(n5430), .ZN(U2800) );
  OAI21_X1 U6586 ( .B1(n3853), .B2(n3031), .A(n5432), .ZN(n5658) );
  NAND2_X1 U6587 ( .A1(n3097), .A2(EBX_REG_18__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6588 ( .A1(n5434), .A2(n5433), .ZN(n5516) );
  OR2_X1 U6589 ( .A1(n6015), .A2(n5516), .ZN(n5514) );
  NAND2_X1 U6590 ( .A1(n6015), .A2(n5516), .ZN(n5435) );
  NAND2_X1 U6591 ( .A1(n5514), .A2(n5435), .ZN(n5520) );
  INV_X1 U6592 ( .A(n5520), .ZN(n6009) );
  INV_X1 U6593 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5521) );
  INV_X1 U6594 ( .A(n5655), .ZN(n5436) );
  OAI22_X1 U6595 ( .A1(n6134), .A2(n5521), .B1(n5436), .B2(n6201), .ZN(n5441)
         );
  INV_X1 U6596 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6554) );
  NOR2_X1 U6597 ( .A1(n5438), .A2(n5437), .ZN(n6081) );
  INV_X1 U6598 ( .A(n6081), .ZN(n5955) );
  AOI21_X1 U6599 ( .B1(n6191), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6173), 
        .ZN(n5439) );
  OAI221_X1 U6600 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5954), .C1(n6554), .C2(
        n5955), .A(n5439), .ZN(n5440) );
  AOI211_X1 U6601 ( .C1(n6009), .C2(n6178), .A(n5441), .B(n5440), .ZN(n5442)
         );
  OAI21_X1 U6602 ( .B1(n5658), .B2(n6150), .A(n5442), .ZN(U2809) );
  OAI21_X1 U6603 ( .B1(n5443), .B2(n5446), .A(n5445), .ZN(n5671) );
  NAND2_X1 U6604 ( .A1(n6188), .A2(n5448), .ZN(n5464) );
  NAND2_X1 U6605 ( .A1(n5447), .A2(n5464), .ZN(n6085) );
  INV_X1 U6606 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5450) );
  NOR3_X1 U6607 ( .A1(n6077), .A2(REIP_REG_15__SCAN_IN), .A3(n5448), .ZN(n6086) );
  AOI211_X1 U6608 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6173), 
        .B(n6086), .ZN(n5449) );
  OAI21_X1 U6609 ( .B1(n5450), .B2(n6134), .A(n5449), .ZN(n5451) );
  AOI21_X1 U6610 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6085), .A(n5451), .ZN(n5456) );
  INV_X1 U6611 ( .A(n5452), .ZN(n5454) );
  INV_X1 U6612 ( .A(n5459), .ZN(n5453) );
  AOI21_X1 U6613 ( .B1(n5454), .B2(n5453), .A(n5523), .ZN(n6025) );
  AOI22_X1 U6614 ( .A1(n6025), .A2(n6178), .B1(n6138), .B2(n5668), .ZN(n5455)
         );
  OAI211_X1 U6615 ( .C1(n5671), .C2(n6150), .A(n5456), .B(n5455), .ZN(U2812)
         );
  NOR2_X1 U6616 ( .A1(n3011), .A2(n5457), .ZN(n5458) );
  NOR2_X1 U6617 ( .A1(n5443), .A2(n5458), .ZN(n5677) );
  INV_X1 U6618 ( .A(n5677), .ZN(n5558) );
  AOI21_X1 U6619 ( .B1(n5460), .B2(n5857), .A(n5459), .ZN(n6038) );
  AOI21_X1 U6620 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6085), .A(n6173), .ZN(n5461) );
  OAI21_X1 U6621 ( .B1(n6201), .B2(n5675), .A(n5461), .ZN(n5467) );
  INV_X1 U6622 ( .A(n5462), .ZN(n5465) );
  AOI22_X1 U6623 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6191), .ZN(n5463) );
  OAI21_X1 U6624 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5466) );
  AOI211_X1 U6625 ( .C1(n6038), .C2(n6178), .A(n5467), .B(n5466), .ZN(n5468)
         );
  OAI21_X1 U6626 ( .B1(n5558), .B2(n6150), .A(n5468), .ZN(U2813) );
  OAI22_X1 U6627 ( .A1(n5735), .A2(n5530), .B1(n6210), .B2(n5469), .ZN(U2828)
         );
  AOI22_X1 U6628 ( .A1(n5750), .A2(n6206), .B1(EBX_REG_29__SCAN_IN), .B2(n5528), .ZN(n5470) );
  OAI21_X1 U6629 ( .B1(n5536), .B2(n5533), .A(n5470), .ZN(U2830) );
  AOI22_X1 U6630 ( .A1(n5760), .A2(n6206), .B1(EBX_REG_28__SCAN_IN), .B2(n5528), .ZN(n5471) );
  OAI21_X1 U6631 ( .B1(n5583), .B2(n5533), .A(n5471), .ZN(U2831) );
  INV_X1 U6632 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5473) );
  OAI222_X1 U6633 ( .A1(n5541), .A2(n5533), .B1(n5473), .B2(n6210), .C1(n5530), 
        .C2(n5472), .ZN(U2832) );
  NAND2_X1 U6634 ( .A1(n5485), .A2(n5474), .ZN(n5475) );
  NAND2_X1 U6635 ( .A1(n3022), .A2(n5475), .ZN(n5901) );
  OAI22_X1 U6636 ( .A1(n5901), .A2(n5530), .B1(n5908), .B2(n6210), .ZN(n5476)
         );
  INV_X1 U6637 ( .A(n5476), .ZN(n5477) );
  OAI21_X1 U6638 ( .B1(n5902), .B2(n5533), .A(n5477), .ZN(U2833) );
  INV_X1 U6639 ( .A(n5478), .ZN(n5481) );
  INV_X1 U6640 ( .A(n5479), .ZN(n5480) );
  AOI21_X1 U6641 ( .B1(n5481), .B2(n5480), .A(n3016), .ZN(n5978) );
  INV_X1 U6642 ( .A(n5978), .ZN(n5546) );
  OR2_X1 U6643 ( .A1(n5482), .A2(n5483), .ZN(n5484) );
  AND2_X1 U6644 ( .A1(n5485), .A2(n5484), .ZN(n5998) );
  AOI22_X1 U6645 ( .A1(n5998), .A2(n6206), .B1(EBX_REG_25__SCAN_IN), .B2(n5528), .ZN(n5486) );
  OAI21_X1 U6646 ( .B1(n5546), .B2(n5533), .A(n5486), .ZN(U2834) );
  NOR2_X1 U6647 ( .A1(n4108), .A2(n5487), .ZN(n5488) );
  OR2_X1 U6648 ( .A1(n5479), .A2(n5488), .ZN(n5614) );
  INV_X1 U6649 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5493) );
  INV_X1 U6650 ( .A(n5489), .ZN(n5491) );
  AOI21_X1 U6651 ( .B1(n5491), .B2(n5490), .A(n5482), .ZN(n5917) );
  INV_X1 U6652 ( .A(n5917), .ZN(n5492) );
  OAI222_X1 U6653 ( .A1(n5533), .A2(n5614), .B1(n6210), .B2(n5493), .C1(n5492), 
        .C2(n5530), .ZN(U2835) );
  OAI222_X1 U6654 ( .A1(n5621), .A2(n5533), .B1(n5494), .B2(n6210), .C1(n5789), 
        .C2(n5530), .ZN(U2836) );
  NAND2_X1 U6655 ( .A1(n5495), .A2(n5496), .ZN(n5497) );
  NAND2_X1 U6656 ( .A1(n5498), .A2(n5497), .ZN(n5936) );
  INV_X1 U6657 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5502) );
  AOI21_X1 U6658 ( .B1(n5501), .B2(n5499), .A(n4106), .ZN(n5926) );
  INV_X1 U6659 ( .A(n5926), .ZN(n5553) );
  OAI222_X1 U6660 ( .A1(n5936), .A2(n5530), .B1(n6210), .B2(n5502), .C1(n5553), 
        .C2(n5533), .ZN(U2837) );
  AOI21_X1 U6661 ( .B1(n5504), .B2(n3010), .A(n5503), .ZN(n5968) );
  INV_X1 U6662 ( .A(n5968), .ZN(n5510) );
  MUX2_X1 U6663 ( .A(n5506), .B(n5392), .S(n5517), .Z(n5508) );
  XNOR2_X1 U6664 ( .A(n5508), .B(n5507), .ZN(n5945) );
  AOI22_X1 U6665 ( .A1(n5945), .A2(n6206), .B1(EBX_REG_20__SCAN_IN), .B2(n5528), .ZN(n5509) );
  OAI21_X1 U6666 ( .B1(n5510), .B2(n5533), .A(n5509), .ZN(U2839) );
  NAND2_X1 U6667 ( .A1(n5432), .A2(n5511), .ZN(n5512) );
  NAND2_X1 U6668 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  OAI21_X1 U6669 ( .B1(n5517), .B2(n5516), .A(n5515), .ZN(n5957) );
  OAI22_X1 U6670 ( .A1(n5957), .A2(n5530), .B1(n5961), .B2(n6210), .ZN(n5518)
         );
  AOI21_X1 U6671 ( .B1(n5982), .B2(n6207), .A(n5518), .ZN(n5519) );
  INV_X1 U6672 ( .A(n5519), .ZN(U2840) );
  OAI222_X1 U6673 ( .A1(n5658), .A2(n5533), .B1(n5521), .B2(n6210), .C1(n5520), 
        .C2(n5530), .ZN(U2841) );
  OR2_X1 U6674 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  NAND2_X1 U6675 ( .A1(n6016), .A2(n5524), .ZN(n6097) );
  INV_X1 U6676 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6090) );
  AND2_X1 U6677 ( .A1(n5445), .A2(n5525), .ZN(n5527) );
  OR2_X1 U6678 ( .A1(n5527), .A2(n5526), .ZN(n6093) );
  OAI222_X1 U6679 ( .A1(n6097), .A2(n5530), .B1(n6210), .B2(n6090), .C1(n6093), 
        .C2(n5533), .ZN(U2843) );
  AOI22_X1 U6680 ( .A1(n6025), .A2(n6206), .B1(EBX_REG_15__SCAN_IN), .B2(n5528), .ZN(n5529) );
  OAI21_X1 U6681 ( .B1(n5671), .B2(n5533), .A(n5529), .ZN(U2844) );
  INV_X1 U6682 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5532) );
  INV_X1 U6683 ( .A(n6038), .ZN(n5531) );
  OAI222_X1 U6684 ( .A1(n5558), .A2(n5533), .B1(n6210), .B2(n5532), .C1(n5531), 
        .C2(n5530), .ZN(U2845) );
  AOI22_X1 U6685 ( .A1(n6214), .A2(DATAI_29_), .B1(n6216), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6686 ( .A1(n6217), .A2(DATAI_13_), .ZN(n5534) );
  OAI211_X1 U6687 ( .C1(n5536), .C2(n6226), .A(n5535), .B(n5534), .ZN(U2862)
         );
  AOI22_X1 U6688 ( .A1(n6214), .A2(DATAI_28_), .B1(n6216), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6689 ( .A1(n6217), .A2(DATAI_12_), .ZN(n5537) );
  OAI211_X1 U6690 ( .C1(n5583), .C2(n6226), .A(n5538), .B(n5537), .ZN(U2863)
         );
  AOI22_X1 U6691 ( .A1(n6214), .A2(DATAI_27_), .B1(n6216), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U6692 ( .A1(n6217), .A2(DATAI_11_), .ZN(n5539) );
  OAI211_X1 U6693 ( .C1(n5541), .C2(n6226), .A(n5540), .B(n5539), .ZN(U2864)
         );
  AOI22_X1 U6694 ( .A1(n6217), .A2(DATAI_10_), .B1(n6216), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U6695 ( .A1(n6214), .A2(DATAI_26_), .ZN(n5542) );
  OAI211_X1 U6696 ( .C1(n5902), .C2(n6226), .A(n5543), .B(n5542), .ZN(U2865)
         );
  AOI22_X1 U6697 ( .A1(n6217), .A2(DATAI_9_), .B1(n6216), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6698 ( .A1(n6214), .A2(DATAI_25_), .ZN(n5544) );
  OAI211_X1 U6699 ( .C1(n5546), .C2(n6226), .A(n5545), .B(n5544), .ZN(U2866)
         );
  AOI22_X1 U6700 ( .A1(n6217), .A2(DATAI_8_), .B1(n6216), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6701 ( .A1(n6214), .A2(DATAI_24_), .ZN(n5547) );
  OAI211_X1 U6702 ( .C1(n5614), .C2(n6226), .A(n5548), .B(n5547), .ZN(U2867)
         );
  AOI22_X1 U6703 ( .A1(n6214), .A2(DATAI_23_), .B1(n6216), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6704 ( .A1(n6217), .A2(DATAI_7_), .ZN(n5549) );
  OAI211_X1 U6705 ( .C1(n5621), .C2(n6226), .A(n5550), .B(n5549), .ZN(U2868)
         );
  AOI22_X1 U6706 ( .A1(n6217), .A2(DATAI_6_), .B1(n6216), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6707 ( .A1(n6214), .A2(DATAI_22_), .ZN(n5551) );
  OAI211_X1 U6708 ( .C1(n5553), .C2(n6226), .A(n5552), .B(n5551), .ZN(U2869)
         );
  AOI22_X1 U6709 ( .A1(n6214), .A2(DATAI_18_), .B1(n6216), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6710 ( .A1(n6217), .A2(DATAI_2_), .ZN(n5554) );
  OAI211_X1 U6711 ( .C1(n5658), .C2(n6226), .A(n5555), .B(n5554), .ZN(U2873)
         );
  AOI22_X1 U6712 ( .A1(n6220), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6216), .ZN(n5556) );
  OAI21_X1 U6713 ( .B1(n5671), .B2(n6226), .A(n5556), .ZN(U2876) );
  AOI22_X1 U6714 ( .A1(n6220), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6216), .ZN(n5557) );
  OAI21_X1 U6715 ( .B1(n5558), .B2(n6226), .A(n5557), .ZN(U2877) );
  NOR2_X1 U6716 ( .A1(n3548), .A2(n3551), .ZN(n5563) );
  INV_X1 U6717 ( .A(n5975), .ZN(n5561) );
  NOR3_X1 U6718 ( .A1(n5559), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5560) );
  XNOR2_X1 U6719 ( .A(n5565), .B(n5731), .ZN(n5738) );
  NAND2_X1 U6720 ( .A1(n6279), .A2(REIP_REG_31__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6721 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5566)
         );
  OAI21_X1 U6722 ( .B1(n5738), .B2(n6060), .A(n5570), .ZN(U2955) );
  NAND2_X1 U6723 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  XNOR2_X1 U6724 ( .A(n5573), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5754)
         );
  AND2_X1 U6725 ( .A1(n6279), .A2(REIP_REG_29__SCAN_IN), .ZN(n5749) );
  AOI21_X1 U6726 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5749), 
        .ZN(n5574) );
  OAI21_X1 U6727 ( .B1(n6271), .B2(n5575), .A(n5574), .ZN(n5576) );
  AOI21_X1 U6728 ( .B1(n5577), .B2(n6266), .A(n5576), .ZN(n5578) );
  OAI21_X1 U6729 ( .B1(n5754), .B2(n6060), .A(n5578), .ZN(U2957) );
  INV_X1 U6730 ( .A(n5600), .ZN(n5579) );
  NAND3_X1 U6731 ( .A1(n5579), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5989), .ZN(n5581) );
  NAND2_X1 U6732 ( .A1(n6002), .A2(n5598), .ZN(n5774) );
  OR2_X1 U6733 ( .A1(n5989), .A2(n5774), .ZN(n5580) );
  AOI22_X2 U6734 ( .A1(n5581), .A2(n5589), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5598), .ZN(n5582) );
  XNOR2_X1 U6735 ( .A(n5582), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5763)
         );
  INV_X1 U6736 ( .A(n5583), .ZN(n5587) );
  AND2_X1 U6737 ( .A1(n6279), .A2(REIP_REG_28__SCAN_IN), .ZN(n5759) );
  AOI21_X1 U6738 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5759), 
        .ZN(n5584) );
  OAI21_X1 U6739 ( .B1(n6271), .B2(n5585), .A(n5584), .ZN(n5586) );
  AOI21_X1 U6740 ( .B1(n5587), .B2(n6266), .A(n5586), .ZN(n5588) );
  OAI21_X1 U6741 ( .B1(n6060), .B2(n5763), .A(n5588), .ZN(U2958) );
  INV_X1 U6742 ( .A(n5589), .ZN(n5590) );
  OR2_X1 U6743 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  XNOR2_X1 U6744 ( .A(n5592), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5771)
         );
  AND2_X1 U6745 ( .A1(n6279), .A2(REIP_REG_27__SCAN_IN), .ZN(n5764) );
  AOI21_X1 U6746 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5764), 
        .ZN(n5593) );
  OAI21_X1 U6747 ( .B1(n6271), .B2(n5594), .A(n5593), .ZN(n5595) );
  AOI21_X1 U6748 ( .B1(n5596), .B2(n6266), .A(n5595), .ZN(n5597) );
  OAI21_X1 U6749 ( .B1(n5771), .B2(n6060), .A(n5597), .ZN(U2959) );
  XNOR2_X1 U6750 ( .A(n2990), .B(n5598), .ZN(n5599) );
  XNOR2_X1 U6751 ( .A(n5600), .B(n5599), .ZN(n5780) );
  INV_X1 U6752 ( .A(n5902), .ZN(n5604) );
  INV_X1 U6753 ( .A(n5900), .ZN(n5602) );
  AND2_X1 U6754 ( .A1(n6279), .A2(REIP_REG_26__SCAN_IN), .ZN(n5772) );
  AOI21_X1 U6755 ( .B1(n6262), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5772), 
        .ZN(n5601) );
  OAI21_X1 U6756 ( .B1(n6271), .B2(n5602), .A(n5601), .ZN(n5603) );
  AOI21_X1 U6757 ( .B1(n5604), .B2(n6266), .A(n5603), .ZN(n5605) );
  OAI21_X1 U6758 ( .B1(n6060), .B2(n5780), .A(n5605), .ZN(U2960) );
  INV_X1 U6759 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5606) );
  XNOR2_X1 U6760 ( .A(n2990), .B(n5606), .ZN(n5642) );
  INV_X1 U6761 ( .A(n5635), .ZN(n5609) );
  INV_X1 U6762 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U6763 ( .A(n2990), .B(n5607), .ZN(n5636) );
  INV_X1 U6764 ( .A(n5636), .ZN(n5608) );
  NAND3_X1 U6765 ( .A1(n5989), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5611) );
  AND2_X1 U6766 ( .A1(n6279), .A2(REIP_REG_24__SCAN_IN), .ZN(n5781) );
  NOR2_X1 U6767 ( .A1(n6276), .A2(n5612), .ZN(n5613) );
  AOI211_X1 U6768 ( .C1(n5695), .C2(n5915), .A(n5781), .B(n5613), .ZN(n5616)
         );
  INV_X1 U6769 ( .A(n5614), .ZN(n5918) );
  NAND2_X1 U6770 ( .A1(n5918), .A2(n6266), .ZN(n5615) );
  OAI211_X1 U6771 ( .C1(n5787), .C2(n6060), .A(n5616), .B(n5615), .ZN(U2962)
         );
  INV_X1 U6772 ( .A(n5782), .ZN(n5799) );
  NAND3_X1 U6773 ( .A1(n5989), .A2(n5814), .A3(n5799), .ZN(n5618) );
  OAI21_X1 U6774 ( .B1(n5619), .B2(n5618), .A(n5617), .ZN(n5620) );
  XNOR2_X1 U6775 ( .A(n5620), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5796)
         );
  INV_X1 U6776 ( .A(n5621), .ZN(n5625) );
  NAND2_X1 U6777 ( .A1(n6279), .A2(REIP_REG_23__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6778 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5622)
         );
  OAI211_X1 U6779 ( .C1(n6271), .C2(n5623), .A(n5788), .B(n5622), .ZN(n5624)
         );
  AOI21_X1 U6780 ( .B1(n5625), .B2(n6266), .A(n5624), .ZN(n5626) );
  OAI21_X1 U6781 ( .B1(n5796), .B2(n6060), .A(n5626), .ZN(U2963) );
  AOI21_X1 U6782 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5989), .A(n5627), 
        .ZN(n5628) );
  XNOR2_X1 U6783 ( .A(n5629), .B(n5628), .ZN(n5803) );
  NAND2_X1 U6784 ( .A1(n5695), .A2(n5929), .ZN(n5630) );
  NAND2_X1 U6785 ( .A1(n6279), .A2(REIP_REG_22__SCAN_IN), .ZN(n5797) );
  OAI211_X1 U6786 ( .C1(n6276), .C2(n5631), .A(n5630), .B(n5797), .ZN(n5632)
         );
  AOI21_X1 U6787 ( .B1(n5926), .B2(n6266), .A(n5632), .ZN(n5633) );
  OAI21_X1 U6788 ( .B1(n5803), .B2(n6060), .A(n5633), .ZN(U2964) );
  AOI21_X1 U6789 ( .B1(n5636), .B2(n5635), .A(n5634), .ZN(n5812) );
  OAI21_X1 U6790 ( .B1(n5503), .B2(n5637), .A(n5499), .ZN(n5638) );
  NAND2_X1 U6791 ( .A1(n6279), .A2(REIP_REG_21__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U6792 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5639)
         );
  OAI211_X1 U6793 ( .C1(n6271), .C2(n5943), .A(n5806), .B(n5639), .ZN(n5640)
         );
  AOI21_X1 U6794 ( .B1(n5965), .B2(n6266), .A(n5640), .ZN(n5641) );
  OAI21_X1 U6795 ( .B1(n5812), .B2(n6060), .A(n5641), .ZN(U2965) );
  XNOR2_X1 U6796 ( .A(n5643), .B(n5642), .ZN(n5827) );
  INV_X1 U6797 ( .A(n5944), .ZN(n5645) );
  NAND2_X1 U6798 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5644)
         );
  NAND2_X1 U6799 ( .A1(n6279), .A2(REIP_REG_20__SCAN_IN), .ZN(n5816) );
  OAI211_X1 U6800 ( .C1(n6271), .C2(n5645), .A(n5644), .B(n5816), .ZN(n5646)
         );
  AOI21_X1 U6801 ( .B1(n5968), .B2(n6266), .A(n5646), .ZN(n5647) );
  OAI21_X1 U6802 ( .B1(n6060), .B2(n5827), .A(n5647), .ZN(U2966) );
  INV_X1 U6803 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5820) );
  NOR3_X1 U6804 ( .A1(n5648), .A2(n5832), .A3(n5820), .ZN(n5992) );
  INV_X1 U6805 ( .A(n5664), .ZN(n5650) );
  NAND3_X1 U6806 ( .A1(n5650), .A2(n5832), .A3(n5649), .ZN(n5991) );
  INV_X1 U6807 ( .A(n5991), .ZN(n5651) );
  NOR2_X1 U6808 ( .A1(n5992), .A2(n5651), .ZN(n5652) );
  XNOR2_X1 U6809 ( .A(n5652), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6010)
         );
  NAND2_X1 U6810 ( .A1(n6010), .A2(n6278), .ZN(n5657) );
  OAI22_X1 U6811 ( .A1(n6276), .A2(n5653), .B1(n6323), .B2(n6554), .ZN(n5654)
         );
  AOI21_X1 U6812 ( .B1(n5695), .B2(n5655), .A(n5654), .ZN(n5656) );
  OAI211_X1 U6813 ( .C1(n6281), .C2(n5658), .A(n5657), .B(n5656), .ZN(U2968)
         );
  XNOR2_X1 U6814 ( .A(n2990), .B(n5987), .ZN(n5659) );
  XNOR2_X1 U6815 ( .A(n5660), .B(n5659), .ZN(n5851) );
  INV_X1 U6816 ( .A(n6093), .ZN(n6215) );
  NAND2_X1 U6817 ( .A1(n6279), .A2(REIP_REG_16__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6818 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5661)
         );
  OAI211_X1 U6819 ( .C1(n6271), .C2(n6092), .A(n5845), .B(n5661), .ZN(n5662)
         );
  AOI21_X1 U6820 ( .B1(n6215), .B2(n6266), .A(n5662), .ZN(n5663) );
  OAI21_X1 U6821 ( .B1(n5851), .B2(n6060), .A(n5663), .ZN(U2970) );
  OAI21_X1 U6822 ( .B1(n5666), .B2(n5665), .A(n5664), .ZN(n6027) );
  NAND2_X1 U6823 ( .A1(n6027), .A2(n6278), .ZN(n5670) );
  NAND2_X1 U6824 ( .A1(n6279), .A2(REIP_REG_15__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U6825 ( .B1(n6276), .B2(n3791), .A(n6023), .ZN(n5667) );
  AOI21_X1 U6826 ( .B1(n5695), .B2(n5668), .A(n5667), .ZN(n5669) );
  OAI211_X1 U6827 ( .C1(n6281), .C2(n5671), .A(n5670), .B(n5669), .ZN(U2971)
         );
  XNOR2_X1 U6828 ( .A(n5989), .B(n6041), .ZN(n5672) );
  XNOR2_X1 U6829 ( .A(n5673), .B(n5672), .ZN(n6036) );
  AOI22_X1 U6830 ( .A1(n6262), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6279), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5674) );
  OAI21_X1 U6831 ( .B1(n6271), .B2(n5675), .A(n5674), .ZN(n5676) );
  AOI21_X1 U6832 ( .B1(n5677), .B2(n6266), .A(n5676), .ZN(n5678) );
  OAI21_X1 U6833 ( .B1(n6060), .B2(n6036), .A(n5678), .ZN(U2972) );
  XNOR2_X1 U6834 ( .A(n5679), .B(n5680), .ZN(n6099) );
  OAI21_X1 U6835 ( .B1(n5683), .B2(n5682), .A(n2991), .ZN(n5852) );
  NAND2_X1 U6836 ( .A1(n5852), .A2(n6278), .ZN(n5686) );
  NOR2_X1 U6837 ( .A1(n6323), .A2(n6544), .ZN(n5861) );
  NOR2_X1 U6838 ( .A1(n6271), .A2(n6100), .ZN(n5684) );
  AOI211_X1 U6839 ( .C1(n6262), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5861), 
        .B(n5684), .ZN(n5685) );
  OAI211_X1 U6840 ( .C1(n6099), .C2(n6281), .A(n5686), .B(n5685), .ZN(U2973)
         );
  INV_X1 U6841 ( .A(n5688), .ZN(n5689) );
  NOR2_X1 U6842 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  XNOR2_X1 U6843 ( .A(n5687), .B(n5691), .ZN(n5871) );
  OAI22_X1 U6844 ( .A1(n6276), .A2(n5692), .B1(n6323), .B2(n6542), .ZN(n5694)
         );
  NOR2_X1 U6845 ( .A1(n6113), .A2(n6281), .ZN(n5693) );
  AOI211_X1 U6846 ( .C1(n5695), .C2(n6114), .A(n5694), .B(n5693), .ZN(n5696)
         );
  OAI21_X1 U6847 ( .B1(n5871), .B2(n6060), .A(n5696), .ZN(U2974) );
  NAND2_X1 U6848 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  XNOR2_X1 U6849 ( .A(n5697), .B(n5700), .ZN(n6286) );
  NAND2_X1 U6850 ( .A1(n6286), .A2(n6278), .ZN(n5704) );
  NOR2_X1 U6851 ( .A1(n6323), .A2(n5276), .ZN(n6283) );
  NOR2_X1 U6852 ( .A1(n6271), .A2(n5701), .ZN(n5702) );
  AOI211_X1 U6853 ( .C1(n6262), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6283), 
        .B(n5702), .ZN(n5703) );
  OAI211_X1 U6854 ( .C1(n6281), .C2(n5705), .A(n5704), .B(n5703), .ZN(U2975)
         );
  INV_X1 U6855 ( .A(n5757), .ZN(n5747) );
  AND2_X1 U6856 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5773) );
  AND4_X1 U6857 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5707), .A4(n5706), .ZN(n5726)
         );
  NAND2_X1 U6858 ( .A1(n6318), .A2(n5726), .ZN(n5724) );
  AOI21_X1 U6859 ( .B1(n5726), .B2(n6320), .A(n5708), .ZN(n5710) );
  AOI211_X1 U6860 ( .C1(n5720), .C2(n5724), .A(n5710), .B(n5709), .ZN(n6290)
         );
  NAND2_X1 U6861 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5855) );
  NOR2_X1 U6862 ( .A1(n5711), .A2(n5855), .ZN(n6031) );
  NAND2_X1 U6863 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6031), .ZN(n5842) );
  NAND2_X1 U6864 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5848) );
  NOR2_X1 U6865 ( .A1(n5842), .A2(n5848), .ZN(n5821) );
  INV_X1 U6866 ( .A(n5821), .ZN(n5712) );
  NAND2_X1 U6867 ( .A1(n5823), .A2(n5712), .ZN(n5713) );
  NAND2_X1 U6868 ( .A1(n6290), .A2(n5713), .ZN(n6014) );
  INV_X1 U6869 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U6870 ( .A1(n5715), .A2(n5814), .ZN(n5716) );
  AND2_X1 U6871 ( .A1(n5823), .A2(n5716), .ZN(n5717) );
  OR2_X1 U6872 ( .A1(n6014), .A2(n5717), .ZN(n5810) );
  AND2_X1 U6873 ( .A1(n5823), .A2(n5782), .ZN(n5718) );
  NOR2_X1 U6874 ( .A1(n5810), .A2(n5718), .ZN(n5790) );
  OAI21_X1 U6875 ( .B1(n5721), .B2(n5720), .A(n5719), .ZN(n5722) );
  NAND2_X1 U6876 ( .A1(n5790), .A2(n5722), .ZN(n6001) );
  INV_X1 U6877 ( .A(n6001), .ZN(n5723) );
  OAI21_X1 U6878 ( .B1(n5844), .B2(n5773), .A(n5723), .ZN(n5769) );
  AOI21_X1 U6879 ( .B1(n5747), .B2(n5823), .A(n5769), .ZN(n5751) );
  OAI21_X1 U6880 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5844), .A(n5751), 
        .ZN(n5744) );
  AOI21_X1 U6881 ( .B1(n3551), .B2(n5823), .A(n5744), .ZN(n5732) );
  OR2_X1 U6882 ( .A1(n6322), .A2(n5724), .ZN(n6032) );
  NAND2_X1 U6883 ( .A1(n5726), .A2(n5725), .ZN(n5865) );
  NAND3_X1 U6884 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5821), .A3(n6285), .ZN(n6013) );
  NOR2_X1 U6885 ( .A1(n6007), .A2(n6013), .ZN(n5836) );
  NAND2_X1 U6886 ( .A1(n5836), .A2(n5814), .ZN(n5807) );
  INV_X1 U6887 ( .A(n5727), .ZN(n5728) );
  NOR2_X1 U6888 ( .A1(n5807), .A2(n5728), .ZN(n6003) );
  NAND2_X1 U6889 ( .A1(n6003), .A2(n5773), .ZN(n5767) );
  OR3_X1 U6890 ( .A1(n5767), .A2(n5747), .A3(n3548), .ZN(n5739) );
  OR3_X1 U6891 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n3551), 
        .ZN(n5729) );
  OAI211_X1 U6892 ( .C1(n5732), .C2(n5731), .A(n5730), .B(n5729), .ZN(n5733)
         );
  INV_X1 U6893 ( .A(n5733), .ZN(n5734) );
  INV_X1 U6894 ( .A(n5736), .ZN(n5737) );
  OAI21_X1 U6895 ( .B1(n5738), .B2(n5870), .A(n5737), .ZN(U2987) );
  NOR2_X1 U6896 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5743)
         );
  OAI21_X1 U6897 ( .B1(n5741), .B2(n6335), .A(n5740), .ZN(n5742) );
  AOI211_X1 U6898 ( .C1(INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n5744), .A(n5743), .B(n5742), .ZN(n5745) );
  OAI21_X1 U6899 ( .B1(n5746), .B2(n5870), .A(n5745), .ZN(U2988) );
  NOR3_X1 U6900 ( .A1(n5767), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5747), 
        .ZN(n5748) );
  AOI211_X1 U6901 ( .C1(n5750), .C2(n6293), .A(n5749), .B(n5748), .ZN(n5753)
         );
  OR2_X1 U6902 ( .A1(n5751), .A2(n3548), .ZN(n5752) );
  OAI211_X1 U6903 ( .C1(n5754), .C2(n5870), .A(n5753), .B(n5752), .ZN(U2989)
         );
  INV_X1 U6904 ( .A(n5755), .ZN(n5756) );
  NOR3_X1 U6905 ( .A1(n5767), .A2(n5757), .A3(n5756), .ZN(n5758) );
  AOI211_X1 U6906 ( .C1(n5760), .C2(n6293), .A(n5759), .B(n5758), .ZN(n5762)
         );
  NAND2_X1 U6907 ( .A1(n5769), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5761) );
  OAI211_X1 U6908 ( .C1(n5763), .C2(n5870), .A(n5762), .B(n5761), .ZN(U2990)
         );
  AOI21_X1 U6909 ( .B1(n5765), .B2(n6293), .A(n5764), .ZN(n5766) );
  OAI21_X1 U6910 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5767), .A(n5766), 
        .ZN(n5768) );
  AOI21_X1 U6911 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5769), .A(n5768), 
        .ZN(n5770) );
  OAI21_X1 U6912 ( .B1(n5771), .B2(n5870), .A(n5770), .ZN(U2991) );
  INV_X1 U6913 ( .A(n5772), .ZN(n5777) );
  INV_X1 U6914 ( .A(n5773), .ZN(n5775) );
  NAND3_X1 U6915 ( .A1(n6003), .A2(n5775), .A3(n5774), .ZN(n5776) );
  OAI211_X1 U6916 ( .C1(n5901), .C2(n6335), .A(n5777), .B(n5776), .ZN(n5778)
         );
  AOI21_X1 U6917 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6001), .A(n5778), 
        .ZN(n5779) );
  OAI21_X1 U6918 ( .B1(n5780), .B2(n5870), .A(n5779), .ZN(U2992) );
  AOI21_X1 U6919 ( .B1(n5917), .B2(n6293), .A(n5781), .ZN(n5786) );
  NOR2_X1 U6920 ( .A1(n5807), .A2(n5782), .ZN(n5794) );
  INV_X1 U6921 ( .A(n5783), .ZN(n5784) );
  OAI211_X1 U6922 ( .C1(n5794), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n6001), .B(n5784), .ZN(n5785) );
  OAI211_X1 U6923 ( .C1(n5787), .C2(n5870), .A(n5786), .B(n5785), .ZN(U2994)
         );
  INV_X1 U6924 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U6925 ( .B1(n5789), .B2(n6335), .A(n5788), .ZN(n5792) );
  NOR2_X1 U6926 ( .A1(n5790), .A2(n5793), .ZN(n5791) );
  AOI211_X1 U6927 ( .C1(n5794), .C2(n5793), .A(n5792), .B(n5791), .ZN(n5795)
         );
  OAI21_X1 U6928 ( .B1(n5796), .B2(n5870), .A(n5795), .ZN(U2995) );
  OAI21_X1 U6929 ( .B1(n5936), .B2(n6335), .A(n5797), .ZN(n5801) );
  NOR3_X1 U6930 ( .A1(n5807), .A2(n5799), .A3(n5798), .ZN(n5800) );
  AOI211_X1 U6931 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5810), .A(n5801), .B(n5800), .ZN(n5802) );
  OAI21_X1 U6932 ( .B1(n5803), .B2(n5870), .A(n5802), .ZN(U2996) );
  OAI21_X1 U6933 ( .B1(n5805), .B2(n5804), .A(n5495), .ZN(n5940) );
  OAI21_X1 U6934 ( .B1(n5940), .B2(n6335), .A(n5806), .ZN(n5809) );
  NOR2_X1 U6935 ( .A1(n5807), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5808)
         );
  AOI211_X1 U6936 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5810), .A(n5809), .B(n5808), .ZN(n5811) );
  OAI21_X1 U6937 ( .B1(n5812), .B2(n5870), .A(n5811), .ZN(U2997) );
  NOR2_X1 U6938 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  NAND2_X1 U6939 ( .A1(n5836), .A2(n5815), .ZN(n5819) );
  INV_X1 U6940 ( .A(n5816), .ZN(n5817) );
  AOI21_X1 U6941 ( .B1(n5945), .B2(n6293), .A(n5817), .ZN(n5818) );
  AND2_X1 U6942 ( .A1(n5819), .A2(n5818), .ZN(n5826) );
  NAND2_X1 U6943 ( .A1(n5821), .A2(n5820), .ZN(n6021) );
  OAI22_X1 U6944 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6322), .B1(n6021), .B2(n5865), .ZN(n5822) );
  NOR2_X1 U6945 ( .A1(n6014), .A2(n5822), .ZN(n6006) );
  NAND2_X1 U6946 ( .A1(n5823), .A2(n6007), .ZN(n5824) );
  NAND2_X1 U6947 ( .A1(n6006), .A2(n5824), .ZN(n5828) );
  NAND2_X1 U6948 ( .A1(n5828), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5825) );
  OAI211_X1 U6949 ( .C1(n5827), .C2(n5870), .A(n5826), .B(n5825), .ZN(U2998)
         );
  INV_X1 U6950 ( .A(n5828), .ZN(n5840) );
  INV_X1 U6951 ( .A(n5829), .ZN(n5831) );
  OAI21_X1 U6952 ( .B1(n5831), .B2(n5839), .A(n5830), .ZN(n5833) );
  XNOR2_X1 U6953 ( .A(n5833), .B(n5832), .ZN(n5983) );
  NAND2_X1 U6954 ( .A1(n5983), .A2(n6337), .ZN(n5838) );
  INV_X1 U6955 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5834) );
  OAI22_X1 U6956 ( .A1(n5957), .A2(n6335), .B1(n6323), .B2(n5834), .ZN(n5835)
         );
  AOI21_X1 U6957 ( .B1(n5836), .B2(n5839), .A(n5835), .ZN(n5837) );
  OAI211_X1 U6958 ( .C1(n5840), .C2(n5839), .A(n5838), .B(n5837), .ZN(U2999)
         );
  NAND3_X1 U6959 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6031), .A3(n6285), .ZN(n6030) );
  AOI21_X1 U6960 ( .B1(n5841), .B2(n5987), .A(n6030), .ZN(n5849) );
  INV_X1 U6961 ( .A(n5842), .ZN(n5843) );
  OAI21_X1 U6962 ( .B1(n5844), .B2(n5843), .A(n6290), .ZN(n6026) );
  NAND2_X1 U6963 ( .A1(n6026), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5846) );
  OAI211_X1 U6964 ( .C1(n6335), .C2(n6097), .A(n5846), .B(n5845), .ZN(n5847)
         );
  AOI21_X1 U6965 ( .B1(n5849), .B2(n5848), .A(n5847), .ZN(n5850) );
  OAI21_X1 U6966 ( .B1(n5851), .B2(n5870), .A(n5850), .ZN(U3002) );
  INV_X1 U6967 ( .A(n5852), .ZN(n5864) );
  NAND2_X1 U6968 ( .A1(n5855), .A2(n5853), .ZN(n5854) );
  OAI211_X1 U6969 ( .C1(n6031), .C2(n6341), .A(n6290), .B(n5854), .ZN(n6034)
         );
  NOR2_X1 U6970 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5855), .ZN(n5856)
         );
  AOI22_X1 U6971 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6034), .B1(n5856), .B2(n6285), .ZN(n5863) );
  INV_X1 U6972 ( .A(n5857), .ZN(n5858) );
  AOI21_X1 U6973 ( .B1(n5860), .B2(n5859), .A(n5858), .ZN(n6205) );
  AOI21_X1 U6974 ( .B1(n6205), .B2(n6293), .A(n5861), .ZN(n5862) );
  OAI211_X1 U6975 ( .C1(n5864), .C2(n5870), .A(n5863), .B(n5862), .ZN(U3005)
         );
  OAI221_X1 U6976 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6322), .C1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5865), .A(n6290), .ZN(n5868) );
  OAI22_X1 U6977 ( .A1(n6109), .A2(n6335), .B1(n6542), .B2(n6323), .ZN(n5867)
         );
  INV_X1 U6978 ( .A(n6285), .ZN(n6022) );
  NOR3_X1 U6979 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6022), .A3(n6289), 
        .ZN(n5866) );
  AOI211_X1 U6980 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n5868), .A(n5867), .B(n5866), .ZN(n5869) );
  OAI21_X1 U6981 ( .B1(n5871), .B2(n5870), .A(n5869), .ZN(U3006) );
  OAI211_X1 U6982 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3001), .A(n5873), .B(
        n5872), .ZN(n5874) );
  OAI21_X1 U6983 ( .B1(n5878), .B2(n4479), .A(n5874), .ZN(n5875) );
  MUX2_X1 U6984 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5875), .S(n6343), 
        .Z(U3464) );
  XNOR2_X1 U6985 ( .A(n5877), .B(n5876), .ZN(n5880) );
  INV_X1 U6986 ( .A(n3002), .ZN(n5879) );
  OAI22_X1 U6987 ( .A1(n5880), .A2(n6353), .B1(n5879), .B2(n5878), .ZN(n5881)
         );
  MUX2_X1 U6988 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5881), .S(n6343), 
        .Z(U3463) );
  INV_X1 U6989 ( .A(n4445), .ZN(n5883) );
  NAND2_X1 U6990 ( .A1(n5883), .A2(n5882), .ZN(n5887) );
  OAI22_X1 U6991 ( .A1(n6452), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n5887), .B2(n5884), .ZN(n5885) );
  AOI21_X1 U6992 ( .B1(n3350), .B2(n5886), .A(n5885), .ZN(n6453) );
  INV_X1 U6993 ( .A(n6045), .ZN(n5896) );
  INV_X1 U6994 ( .A(n5887), .ZN(n5890) );
  AOI22_X1 U6995 ( .A1(n5891), .A2(n5890), .B1(n5889), .B2(n5888), .ZN(n5892)
         );
  OAI21_X1 U6996 ( .B1(n6453), .B2(n5896), .A(n5892), .ZN(n5894) );
  INV_X1 U6997 ( .A(n5893), .ZN(n6050) );
  MUX2_X1 U6998 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n5894), .S(n6050), 
        .Z(U3460) );
  OAI22_X1 U6999 ( .A1(n5897), .A2(n5896), .B1(n5895), .B2(n6492), .ZN(n5898)
         );
  MUX2_X1 U7000 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5898), .S(n6050), 
        .Z(U3456) );
  AND2_X1 U7001 ( .A1(n6251), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7002 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6191), .B1(n5900), 
        .B2(n6138), .ZN(n5907) );
  NAND2_X1 U7003 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5919), .ZN(n5909) );
  OAI21_X1 U7004 ( .B1(n6653), .B2(n5909), .A(n6731), .ZN(n5904) );
  OAI22_X1 U7005 ( .A1(n5902), .A2(n6150), .B1(n6196), .B2(n5901), .ZN(n5903)
         );
  AOI21_X1 U7006 ( .B1(n5905), .B2(n5904), .A(n5903), .ZN(n5906) );
  OAI211_X1 U7007 ( .C1(n5908), .C2(n6134), .A(n5907), .B(n5906), .ZN(U2801)
         );
  AOI21_X1 U7008 ( .B1(n5919), .B2(n6669), .A(n5916), .ZN(n5914) );
  NOR2_X1 U7009 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5909), .ZN(n5911) );
  OAI22_X1 U7010 ( .A1(n3985), .A2(n6170), .B1(n5981), .B2(n6201), .ZN(n5910)
         );
  AOI211_X1 U7011 ( .C1(n6192), .C2(EBX_REG_25__SCAN_IN), .A(n5911), .B(n5910), 
        .ZN(n5913) );
  AOI22_X1 U7012 ( .A1(n5978), .A2(n6139), .B1(n6178), .B2(n5998), .ZN(n5912)
         );
  OAI211_X1 U7013 ( .C1(n5914), .C2(n6653), .A(n5913), .B(n5912), .ZN(U2802)
         );
  AOI22_X1 U7014 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6191), .ZN(n5923) );
  AOI22_X1 U7015 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5916), .B1(n5915), .B2(
        n6138), .ZN(n5922) );
  AOI22_X1 U7016 ( .A1(n5918), .A2(n6139), .B1(n6178), .B2(n5917), .ZN(n5921)
         );
  NAND2_X1 U7017 ( .A1(n5919), .A2(n6669), .ZN(n5920) );
  NAND4_X1 U7018 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(U2803)
         );
  AND2_X1 U7019 ( .A1(n5925), .A2(n5924), .ZN(n5946) );
  NOR2_X1 U7020 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5927), .ZN(n5939) );
  NAND2_X1 U7021 ( .A1(n5926), .A2(n6139), .ZN(n5933) );
  NOR2_X1 U7022 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5927), .ZN(n5928) );
  AOI22_X1 U7023 ( .A1(n6191), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5928), .ZN(n5932) );
  NAND2_X1 U7024 ( .A1(n6192), .A2(EBX_REG_22__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7025 ( .A1(n6138), .A2(n5929), .ZN(n5930) );
  NAND4_X1 U7026 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n5934)
         );
  AOI221_X1 U7027 ( .B1(n5946), .B2(REIP_REG_22__SCAN_IN), .C1(n5939), .C2(
        REIP_REG_22__SCAN_IN), .A(n5934), .ZN(n5935) );
  OAI21_X1 U7028 ( .B1(n5936), .B2(n6196), .A(n5935), .ZN(U2805) );
  INV_X1 U7029 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5964) );
  INV_X1 U7030 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5937) );
  OAI22_X1 U7031 ( .A1(n5964), .A2(n6134), .B1(n5937), .B2(n6170), .ZN(n5938)
         );
  AOI211_X1 U7032 ( .C1(n5946), .C2(REIP_REG_21__SCAN_IN), .A(n5939), .B(n5938), .ZN(n5942) );
  INV_X1 U7033 ( .A(n5940), .ZN(n5962) );
  AOI22_X1 U7034 ( .A1(n5965), .A2(n6139), .B1(n6178), .B2(n5962), .ZN(n5941)
         );
  OAI211_X1 U7035 ( .C1(n5943), .C2(n6201), .A(n5942), .B(n5941), .ZN(U2806)
         );
  AOI22_X1 U7036 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6191), .ZN(n5951) );
  AOI22_X1 U7037 ( .A1(n5968), .A2(n6139), .B1(n6138), .B2(n5944), .ZN(n5950)
         );
  NAND2_X1 U7038 ( .A1(n6178), .A2(n5945), .ZN(n5949) );
  OAI21_X1 U7039 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5947), .A(n5946), .ZN(n5948) );
  NAND4_X1 U7040 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(U2807)
         );
  OAI21_X1 U7041 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5952), .ZN(n5953) );
  OAI22_X1 U7042 ( .A1(n5834), .A2(n5955), .B1(n5954), .B2(n5953), .ZN(n5956)
         );
  AOI211_X1 U7043 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6173), 
        .B(n5956), .ZN(n5960) );
  OAI22_X1 U7044 ( .A1(n5957), .A2(n6196), .B1(n5986), .B2(n6201), .ZN(n5958)
         );
  AOI21_X1 U7045 ( .B1(n5982), .B2(n6139), .A(n5958), .ZN(n5959) );
  OAI211_X1 U7046 ( .C1(n5961), .C2(n6134), .A(n5960), .B(n5959), .ZN(U2808)
         );
  AOI22_X1 U7047 ( .A1(n5965), .A2(n6207), .B1(n6206), .B2(n5962), .ZN(n5963)
         );
  OAI21_X1 U7048 ( .B1(n6210), .B2(n5964), .A(n5963), .ZN(U2838) );
  INV_X1 U7049 ( .A(n6226), .ZN(n6221) );
  AOI22_X1 U7050 ( .A1(n5965), .A2(n6221), .B1(n6214), .B2(DATAI_21_), .ZN(
        n5967) );
  AOI22_X1 U7051 ( .A1(n6217), .A2(DATAI_5_), .B1(n6216), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7052 ( .A1(n5967), .A2(n5966), .ZN(U2870) );
  AOI22_X1 U7053 ( .A1(n5968), .A2(n6221), .B1(n6214), .B2(DATAI_20_), .ZN(
        n5970) );
  AOI22_X1 U7054 ( .A1(n6217), .A2(DATAI_4_), .B1(n6216), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7055 ( .A1(n5970), .A2(n5969), .ZN(U2871) );
  AOI22_X1 U7056 ( .A1(n5982), .A2(n6221), .B1(n6214), .B2(DATAI_19_), .ZN(
        n5972) );
  AOI22_X1 U7057 ( .A1(n6217), .A2(DATAI_3_), .B1(n6216), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7058 ( .A1(n5972), .A2(n5971), .ZN(U2872) );
  AOI22_X1 U7059 ( .A1(n6279), .A2(REIP_REG_25__SCAN_IN), .B1(n6262), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5980) );
  INV_X1 U7060 ( .A(n5973), .ZN(n5977) );
  INV_X1 U7061 ( .A(n5974), .ZN(n5976) );
  OAI21_X1 U7062 ( .B1(n5977), .B2(n5976), .A(n5975), .ZN(n5999) );
  AOI22_X1 U7063 ( .A1(n5978), .A2(n6266), .B1(n6278), .B2(n5999), .ZN(n5979)
         );
  OAI211_X1 U7064 ( .C1(n6271), .C2(n5981), .A(n5980), .B(n5979), .ZN(U2961)
         );
  AOI22_X1 U7065 ( .A1(n6279), .A2(REIP_REG_19__SCAN_IN), .B1(n6262), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5985) );
  AOI22_X1 U7066 ( .A1(n5983), .A2(n6278), .B1(n6266), .B2(n5982), .ZN(n5984)
         );
  OAI211_X1 U7067 ( .C1(n6271), .C2(n5986), .A(n5985), .B(n5984), .ZN(U2967)
         );
  AOI22_X1 U7068 ( .A1(n6279), .A2(REIP_REG_17__SCAN_IN), .B1(n6262), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5997) );
  NAND3_X1 U7069 ( .A1(n5648), .A2(n5832), .A3(n5987), .ZN(n5988) );
  AOI22_X1 U7070 ( .A1(n5990), .A2(n5989), .B1(n5988), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5993) );
  OAI21_X1 U7071 ( .B1(n5993), .B2(n5992), .A(n5991), .ZN(n6018) );
  OR2_X1 U7072 ( .A1(n5526), .A2(n5994), .ZN(n5995) );
  AND2_X1 U7073 ( .A1(n5431), .A2(n5995), .ZN(n6211) );
  AOI22_X1 U7074 ( .A1(n6018), .A2(n6278), .B1(n6266), .B2(n6211), .ZN(n5996)
         );
  OAI211_X1 U7075 ( .C1(n6271), .C2(n6084), .A(n5997), .B(n5996), .ZN(U2969)
         );
  AOI22_X1 U7076 ( .A1(n5999), .A2(n6337), .B1(n6293), .B2(n5998), .ZN(n6005)
         );
  NOR2_X1 U7077 ( .A1(n6323), .A2(n6653), .ZN(n6000) );
  AOI221_X1 U7078 ( .B1(n6003), .B2(n6002), .C1(n6001), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6000), .ZN(n6004) );
  NAND2_X1 U7079 ( .A1(n6005), .A2(n6004), .ZN(U2993) );
  OAI22_X1 U7080 ( .A1(n6007), .A2(n6006), .B1(n6323), .B2(n6554), .ZN(n6008)
         );
  INV_X1 U7081 ( .A(n6008), .ZN(n6012) );
  AOI22_X1 U7082 ( .A1(n6010), .A2(n6337), .B1(n6293), .B2(n6009), .ZN(n6011)
         );
  OAI211_X1 U7083 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n6013), .A(n6012), .B(n6011), .ZN(U3000) );
  AOI22_X1 U7084 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6014), .B1(n6279), .B2(REIP_REG_17__SCAN_IN), .ZN(n6020) );
  AOI21_X1 U7085 ( .B1(n6017), .B2(n6016), .A(n3063), .ZN(n6202) );
  AOI22_X1 U7086 ( .A1(n6018), .A2(n6337), .B1(n6293), .B2(n6202), .ZN(n6019)
         );
  OAI211_X1 U7087 ( .C1(n6022), .C2(n6021), .A(n6020), .B(n6019), .ZN(U3001)
         );
  INV_X1 U7088 ( .A(n6023), .ZN(n6024) );
  AOI21_X1 U7089 ( .B1(n6025), .B2(n6293), .A(n6024), .ZN(n6029) );
  AOI22_X1 U7090 ( .A1(n6027), .A2(n6337), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6026), .ZN(n6028) );
  OAI211_X1 U7091 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6030), .A(n6029), .B(n6028), .ZN(U3003) );
  NAND2_X1 U7092 ( .A1(n6031), .A2(n6285), .ZN(n6042) );
  AOI21_X1 U7093 ( .B1(n6033), .B2(n6032), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n6035) );
  NOR2_X1 U7094 ( .A1(n6035), .A2(n6034), .ZN(n6040) );
  INV_X1 U7095 ( .A(n6036), .ZN(n6037) );
  AOI222_X1 U7096 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6279), .B1(n6293), .B2(
        n6038), .C1(n6337), .C2(n6037), .ZN(n6039) );
  OAI221_X1 U7097 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6042), .C1(
        n6041), .C2(n6040), .A(n6039), .ZN(U3004) );
  INV_X1 U7098 ( .A(n6169), .ZN(n6047) );
  INV_X1 U7099 ( .A(n6043), .ZN(n6046) );
  NAND4_X1 U7100 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n6048)
         );
  OAI21_X1 U7101 ( .B1(n6050), .B2(n6049), .A(n6048), .ZN(U3455) );
  INV_X1 U7102 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6697) );
  INV_X1 U7103 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U7104 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6515), .ZN(n6051) );
  AOI21_X1 U7105 ( .B1(STATE_REG_0__SCAN_IN), .B2(n6051), .A(n6791), .ZN(n6577) );
  OAI21_X1 U7106 ( .B1(n6791), .B2(n6697), .A(n6508), .ZN(U2789) );
  INV_X1 U7107 ( .A(n6052), .ZN(n6473) );
  OAI22_X1 U7108 ( .A1(n6473), .A2(n6054), .B1(n6465), .B2(n6053), .ZN(n6059)
         );
  OAI21_X1 U7109 ( .B1(n6059), .B2(n6498), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6055) );
  OAI21_X1 U7110 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6499), .A(n6055), .ZN(
        U2790) );
  INV_X2 U7111 ( .A(n6791), .ZN(n6790) );
  NOR2_X1 U7112 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6057) );
  OAI21_X1 U7113 ( .B1(n6057), .B2(D_C_N_REG_SCAN_IN), .A(n6790), .ZN(n6056)
         );
  OAI21_X1 U7114 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6790), .A(n6056), .ZN(
        U2791) );
  OAI21_X1 U7115 ( .B1(BS16_N), .B2(n6057), .A(n6577), .ZN(n6575) );
  OAI21_X1 U7116 ( .B1(n6577), .B2(n6715), .A(n6575), .ZN(U2792) );
  AOI21_X1 U7117 ( .B1(n6058), .B2(n6514), .A(READY_N), .ZN(n6593) );
  NOR2_X1 U7118 ( .A1(n6059), .A2(n6593), .ZN(n6478) );
  NOR2_X1 U7119 ( .A1(n6478), .A2(n6498), .ZN(n6589) );
  OAI21_X1 U7120 ( .B1(n6589), .B2(n6709), .A(n6060), .ZN(U2793) );
  NOR4_X1 U7121 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6064) );
  NOR4_X1 U7122 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6063) );
  NOR4_X1 U7123 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6062) );
  NOR4_X1 U7124 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6061) );
  NAND4_X1 U7125 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n6070)
         );
  NOR4_X1 U7126 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n6068) );
  AOI211_X1 U7127 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6067) );
  NOR4_X1 U7128 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6066) );
  NOR4_X1 U7129 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6065) );
  NAND4_X1 U7130 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(n6069)
         );
  NOR2_X1 U7131 ( .A1(n6070), .A2(n6069), .ZN(n6586) );
  INV_X1 U7132 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6072) );
  NOR3_X1 U7133 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6073) );
  OAI21_X1 U7134 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6073), .A(n6586), .ZN(n6071)
         );
  OAI21_X1 U7135 ( .B1(n6586), .B2(n6072), .A(n6071), .ZN(U2794) );
  INV_X1 U7136 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6576) );
  AOI21_X1 U7137 ( .B1(n5069), .B2(n6576), .A(n6073), .ZN(n6074) );
  INV_X1 U7138 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6724) );
  INV_X1 U7139 ( .A(n6586), .ZN(n6582) );
  AOI22_X1 U7140 ( .A1(n6586), .A2(n6074), .B1(n6724), .B2(n6582), .ZN(U2795)
         );
  OAI21_X1 U7141 ( .B1(n6077), .B2(n6076), .A(n6075), .ZN(n6080) );
  AOI22_X1 U7142 ( .A1(EBX_REG_17__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6191), .ZN(n6078) );
  INV_X1 U7143 ( .A(n6078), .ZN(n6079) );
  AOI211_X1 U7144 ( .C1(n6081), .C2(n6080), .A(n6173), .B(n6079), .ZN(n6083)
         );
  AOI22_X1 U7145 ( .A1(n6211), .A2(n6139), .B1(n6178), .B2(n6202), .ZN(n6082)
         );
  OAI211_X1 U7146 ( .C1(n6084), .C2(n6201), .A(n6083), .B(n6082), .ZN(U2810)
         );
  OAI21_X1 U7147 ( .B1(n6086), .B2(n6085), .A(REIP_REG_16__SCAN_IN), .ZN(n6089) );
  INV_X1 U7148 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6551) );
  NAND3_X1 U7149 ( .A1(n6188), .A2(n6551), .A3(n6087), .ZN(n6088) );
  OAI211_X1 U7150 ( .C1(n6134), .C2(n6090), .A(n6089), .B(n6088), .ZN(n6091)
         );
  AOI211_X1 U7151 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6173), 
        .B(n6091), .ZN(n6096) );
  OAI22_X1 U7152 ( .A1(n6093), .A2(n6150), .B1(n6092), .B2(n6201), .ZN(n6094)
         );
  INV_X1 U7153 ( .A(n6094), .ZN(n6095) );
  OAI211_X1 U7154 ( .C1(n6196), .C2(n6097), .A(n6096), .B(n6095), .ZN(U2811)
         );
  AOI22_X1 U7155 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6192), .B1(n6178), .B2(n6205), .ZN(n6107) );
  NOR4_X1 U7156 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6542), .A3(n6102), .A4(n6103), .ZN(n6098) );
  AOI211_X1 U7157 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6173), 
        .B(n6098), .ZN(n6106) );
  INV_X1 U7158 ( .A(n6099), .ZN(n6222) );
  INV_X1 U7159 ( .A(n6100), .ZN(n6101) );
  AOI22_X1 U7160 ( .A1(n6222), .A2(n6139), .B1(n6138), .B2(n6101), .ZN(n6105)
         );
  NOR3_X1 U7161 ( .A1(n6103), .A2(REIP_REG_12__SCAN_IN), .A3(n6102), .ZN(n6111) );
  OAI21_X1 U7162 ( .B1(n6112), .B2(n6111), .A(REIP_REG_13__SCAN_IN), .ZN(n6104) );
  NAND4_X1 U7163 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(U2814)
         );
  AOI22_X1 U7164 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6191), .ZN(n6108) );
  OAI211_X1 U7165 ( .C1(n6196), .C2(n6109), .A(n6108), .B(n6159), .ZN(n6110)
         );
  AOI211_X1 U7166 ( .C1(n6112), .C2(REIP_REG_12__SCAN_IN), .A(n6111), .B(n6110), .ZN(n6117) );
  INV_X1 U7167 ( .A(n6113), .ZN(n6115) );
  AOI22_X1 U7168 ( .A1(n6115), .A2(n6139), .B1(n6114), .B2(n6138), .ZN(n6116)
         );
  NAND2_X1 U7169 ( .A1(n6117), .A2(n6116), .ZN(U2815) );
  OAI22_X1 U7170 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6119), .B1(n6196), .B2(
        n6118), .ZN(n6120) );
  AOI211_X1 U7171 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6173), 
        .B(n6120), .ZN(n6128) );
  INV_X1 U7172 ( .A(n6121), .ZN(n6123) );
  AOI22_X1 U7173 ( .A1(n6123), .A2(n6139), .B1(n6138), .B2(n6122), .ZN(n6127)
         );
  OAI21_X1 U7174 ( .B1(n6132), .B2(n6124), .A(REIP_REG_10__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7175 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6192), .ZN(n6125) );
  NAND4_X1 U7176 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(U2817)
         );
  INV_X1 U7177 ( .A(n6129), .ZN(n6131) );
  NOR2_X1 U7178 ( .A1(n6131), .A2(n6130), .ZN(n6145) );
  AOI21_X1 U7179 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6145), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6144) );
  INV_X1 U7180 ( .A(n6132), .ZN(n6143) );
  OAI22_X1 U7181 ( .A1(n6135), .A2(n6134), .B1(n6196), .B2(n6133), .ZN(n6136)
         );
  AOI211_X1 U7182 ( .C1(n6191), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6173), 
        .B(n6136), .ZN(n6142) );
  AOI22_X1 U7183 ( .A1(n6140), .A2(n6139), .B1(n6138), .B2(n6137), .ZN(n6141)
         );
  OAI211_X1 U7184 ( .C1(n6144), .C2(n6143), .A(n6142), .B(n6141), .ZN(U2819)
         );
  INV_X1 U7185 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6535) );
  INV_X1 U7186 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6148) );
  AOI22_X1 U7187 ( .A1(n6178), .A2(n6146), .B1(n6145), .B2(n6535), .ZN(n6147)
         );
  OAI211_X1 U7188 ( .C1(n6170), .C2(n6148), .A(n6147), .B(n6159), .ZN(n6153)
         );
  OAI22_X1 U7189 ( .A1(n6151), .A2(n6150), .B1(n6149), .B2(n6201), .ZN(n6152)
         );
  AOI211_X1 U7190 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6192), .A(n6153), .B(n6152), 
        .ZN(n6154) );
  OAI221_X1 U7191 ( .B1(n6535), .B2(n6163), .C1(n6535), .C2(n6155), .A(n6154), 
        .ZN(U2820) );
  AND2_X1 U7192 ( .A1(n6156), .A2(n6532), .ZN(n6162) );
  AOI22_X1 U7193 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6192), .B1(n6178), .B2(n6157), 
        .ZN(n6158) );
  NAND2_X1 U7194 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  AOI21_X1 U7195 ( .B1(n6191), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6160), 
        .ZN(n6161) );
  OAI21_X1 U7196 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6164) );
  AOI21_X1 U7197 ( .B1(n6165), .B2(n6199), .A(n6164), .ZN(n6166) );
  OAI21_X1 U7198 ( .B1(n6167), .B2(n6201), .A(n6166), .ZN(U2822) );
  OAI22_X1 U7199 ( .A1(n6171), .A2(n6170), .B1(n6169), .B2(n6168), .ZN(n6172)
         );
  AOI211_X1 U7200 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6174), .A(n6173), .B(n6172), 
        .ZN(n6185) );
  NOR2_X1 U7201 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6175), .ZN(n6176) );
  AOI22_X1 U7202 ( .A1(n6176), .A2(n6188), .B1(n6192), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n6180) );
  NAND2_X1 U7203 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  OAI211_X1 U7204 ( .C1(n6182), .C2(n6181), .A(n6180), .B(n6179), .ZN(n6183)
         );
  INV_X1 U7205 ( .A(n6183), .ZN(n6184) );
  OAI211_X1 U7206 ( .C1(n6186), .C2(n6201), .A(n6185), .B(n6184), .ZN(U2823)
         );
  INV_X1 U7207 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6526) );
  AOI211_X1 U7208 ( .C1(n6188), .C2(n5069), .A(n6187), .B(n6526), .ZN(n6190)
         );
  AOI21_X1 U7209 ( .B1(n6188), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6189) );
  NOR2_X1 U7210 ( .A1(n6190), .A2(n6189), .ZN(n6198) );
  AOI22_X1 U7211 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6192), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6191), .ZN(n6195) );
  NAND2_X1 U7212 ( .A1(n6193), .A2(n3002), .ZN(n6194) );
  OAI211_X1 U7213 ( .C1(n6196), .C2(n6324), .A(n6195), .B(n6194), .ZN(n6197)
         );
  AOI211_X1 U7214 ( .C1(n6267), .C2(n6199), .A(n6198), .B(n6197), .ZN(n6200)
         );
  OAI21_X1 U7215 ( .B1(n6270), .B2(n6201), .A(n6200), .ZN(U2825) );
  INV_X1 U7216 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6204) );
  AOI22_X1 U7217 ( .A1(n6211), .A2(n6207), .B1(n6206), .B2(n6202), .ZN(n6203)
         );
  OAI21_X1 U7218 ( .B1(n6210), .B2(n6204), .A(n6203), .ZN(U2842) );
  INV_X1 U7219 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6209) );
  AOI22_X1 U7220 ( .A1(n6222), .A2(n6207), .B1(n6206), .B2(n6205), .ZN(n6208)
         );
  OAI21_X1 U7221 ( .B1(n6210), .B2(n6209), .A(n6208), .ZN(U2846) );
  AOI22_X1 U7222 ( .A1(n6211), .A2(n6221), .B1(n6214), .B2(DATAI_17_), .ZN(
        n6213) );
  AOI22_X1 U7223 ( .A1(n6217), .A2(DATAI_1_), .B1(n6216), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7224 ( .A1(n6213), .A2(n6212), .ZN(U2874) );
  AOI22_X1 U7225 ( .A1(n6215), .A2(n6221), .B1(n6214), .B2(DATAI_16_), .ZN(
        n6219) );
  AOI22_X1 U7226 ( .A1(n6217), .A2(DATAI_0_), .B1(n6216), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7227 ( .A1(n6219), .A2(n6218), .ZN(U2875) );
  AOI22_X1 U7228 ( .A1(n6222), .A2(n6221), .B1(DATAI_13_), .B2(n6220), .ZN(
        n6223) );
  OAI21_X1 U7229 ( .B1(n6233), .B2(n6225), .A(n6223), .ZN(U2878) );
  OAI222_X1 U7230 ( .A1(n6282), .A2(n6226), .B1(n6225), .B2(n6261), .C1(n6224), 
        .C2(n6689), .ZN(U2891) );
  AOI22_X1 U7231 ( .A1(n6592), .A2(LWORD_REG_15__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7232 ( .B1(n6229), .B2(n6260), .A(n6228), .ZN(U2908) );
  AOI22_X1 U7233 ( .A1(n6592), .A2(LWORD_REG_14__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7234 ( .B1(n6231), .B2(n6260), .A(n6230), .ZN(U2909) );
  AOI22_X1 U7235 ( .A1(n6592), .A2(LWORD_REG_13__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7236 ( .B1(n6233), .B2(n6260), .A(n6232), .ZN(U2910) );
  AOI22_X1 U7237 ( .A1(n6239), .A2(LWORD_REG_12__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6234) );
  OAI21_X1 U7238 ( .B1(n5297), .B2(n6260), .A(n6234), .ZN(U2911) );
  AOI22_X1 U7239 ( .A1(n6239), .A2(LWORD_REG_11__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7240 ( .B1(n6236), .B2(n6260), .A(n6235), .ZN(U2912) );
  AOI22_X1 U7241 ( .A1(n6239), .A2(LWORD_REG_10__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6237) );
  OAI21_X1 U7242 ( .B1(n6238), .B2(n6260), .A(n6237), .ZN(U2913) );
  AOI22_X1 U7243 ( .A1(n6239), .A2(LWORD_REG_9__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U7244 ( .B1(n6241), .B2(n6260), .A(n6240), .ZN(U2914) );
  AOI22_X1 U7245 ( .A1(n6592), .A2(LWORD_REG_8__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6242) );
  OAI21_X1 U7246 ( .B1(n6243), .B2(n6260), .A(n6242), .ZN(U2915) );
  AOI22_X1 U7247 ( .A1(n6592), .A2(LWORD_REG_7__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6244) );
  OAI21_X1 U7248 ( .B1(n3676), .B2(n6260), .A(n6244), .ZN(U2916) );
  AOI22_X1 U7249 ( .A1(n6592), .A2(LWORD_REG_6__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6245) );
  OAI21_X1 U7250 ( .B1(n6246), .B2(n6260), .A(n6245), .ZN(U2917) );
  AOI22_X1 U7251 ( .A1(n6592), .A2(LWORD_REG_5__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U7252 ( .B1(n6248), .B2(n6260), .A(n6247), .ZN(U2918) );
  AOI22_X1 U7253 ( .A1(n6592), .A2(LWORD_REG_4__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6249) );
  OAI21_X1 U7254 ( .B1(n6250), .B2(n6260), .A(n6249), .ZN(U2919) );
  AOI22_X1 U7255 ( .A1(n6592), .A2(LWORD_REG_3__SCAN_IN), .B1(n6251), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U7256 ( .B1(n6253), .B2(n6260), .A(n6252), .ZN(U2920) );
  AOI22_X1 U7257 ( .A1(n6592), .A2(LWORD_REG_2__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U7258 ( .B1(n6255), .B2(n6260), .A(n6254), .ZN(U2921) );
  AOI22_X1 U7259 ( .A1(n6592), .A2(LWORD_REG_1__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6256) );
  OAI21_X1 U7260 ( .B1(n6257), .B2(n6260), .A(n6256), .ZN(U2922) );
  AOI22_X1 U7261 ( .A1(n6592), .A2(LWORD_REG_0__SCAN_IN), .B1(n6258), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7262 ( .B1(n6261), .B2(n6260), .A(n6259), .ZN(U2923) );
  AOI22_X1 U7263 ( .A1(n6279), .A2(REIP_REG_2__SCAN_IN), .B1(n6262), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6269) );
  XNOR2_X1 U7264 ( .A(n6264), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6265)
         );
  XNOR2_X1 U7265 ( .A(n6263), .B(n6265), .ZN(n6327) );
  AOI22_X1 U7266 ( .A1(n6267), .A2(n6266), .B1(n6327), .B2(n6278), .ZN(n6268)
         );
  OAI211_X1 U7267 ( .C1(n6271), .C2(n6270), .A(n6269), .B(n6268), .ZN(U2984)
         );
  OAI21_X1 U7268 ( .B1(n6273), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6272), 
        .ZN(n6274) );
  INV_X1 U7269 ( .A(n6274), .ZN(n6338) );
  NAND2_X1 U7270 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  AOI22_X1 U7271 ( .A1(n6338), .A2(n6278), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6277), .ZN(n6280) );
  NAND2_X1 U7272 ( .A1(n6279), .A2(REIP_REG_0__SCAN_IN), .ZN(n6332) );
  OAI211_X1 U7273 ( .C1(n6282), .C2(n6281), .A(n6280), .B(n6332), .ZN(U2986)
         );
  AOI21_X1 U7274 ( .B1(n6284), .B2(n6293), .A(n6283), .ZN(n6288) );
  AOI22_X1 U7275 ( .A1(n6337), .A2(n6286), .B1(n6289), .B2(n6285), .ZN(n6287)
         );
  OAI211_X1 U7276 ( .C1(n6290), .C2(n6289), .A(n6288), .B(n6287), .ZN(U3007)
         );
  INV_X1 U7277 ( .A(n6291), .ZN(n6294) );
  AOI21_X1 U7278 ( .B1(n6294), .B2(n6293), .A(n6292), .ZN(n6298) );
  AOI22_X1 U7279 ( .A1(n6296), .A2(n6337), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6295), .ZN(n6297) );
  OAI211_X1 U7280 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6299), .A(n6298), 
        .B(n6297), .ZN(U3009) );
  NAND2_X1 U7281 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  OAI211_X1 U7282 ( .C1(n6304), .C2(n6335), .A(n6303), .B(n6302), .ZN(n6305)
         );
  AOI21_X1 U7283 ( .B1(n6306), .B2(n6337), .A(n6305), .ZN(n6307) );
  OAI21_X1 U7284 ( .B1(n6308), .B2(n6301), .A(n6307), .ZN(U3011) );
  OAI21_X1 U7285 ( .B1(n6335), .B2(n6310), .A(n6309), .ZN(n6313) );
  NOR2_X1 U7286 ( .A1(n6311), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6312)
         );
  AOI211_X1 U7287 ( .C1(n6337), .C2(n6314), .A(n6313), .B(n6312), .ZN(n6315)
         );
  OAI21_X1 U7288 ( .B1(n6316), .B2(n3433), .A(n6315), .ZN(U3015) );
  INV_X1 U7289 ( .A(n6317), .ZN(n6329) );
  INV_X1 U7290 ( .A(n6318), .ZN(n6319) );
  AOI21_X1 U7291 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6320), .A(n6319), 
        .ZN(n6321) );
  NOR2_X1 U7292 ( .A1(n6322), .A2(n6321), .ZN(n6326) );
  OAI22_X1 U7293 ( .A1(n6335), .A2(n6324), .B1(n6526), .B2(n6323), .ZN(n6325)
         );
  AOI211_X1 U7294 ( .C1(n6327), .C2(n6337), .A(n6326), .B(n6325), .ZN(n6328)
         );
  OAI221_X1 U7295 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6331), .C1(n6330), .C2(n6329), .A(n6328), .ZN(U3016) );
  OAI211_X1 U7296 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n6332), .ZN(n6336)
         );
  AOI21_X1 U7297 ( .B1(n6338), .B2(n6337), .A(n6336), .ZN(n6339) );
  OAI221_X1 U7298 ( .B1(n6342), .B2(n6341), .C1(n6342), .C2(n6340), .A(n6339), 
        .ZN(U3018) );
  INV_X1 U7299 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6482) );
  NOR2_X1 U7300 ( .A1(n6482), .A2(n6343), .ZN(U3019) );
  NAND3_X1 U7301 ( .A1(n6346), .A2(n6345), .A3(n6344), .ZN(n6347) );
  OAI21_X1 U7302 ( .B1(n6348), .B2(n3003), .A(n6347), .ZN(n6393) );
  NOR2_X1 U7303 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6349), .ZN(n6392)
         );
  AOI22_X1 U7304 ( .A1(n6351), .A2(n6393), .B1(n6350), .B2(n6392), .ZN(n6364)
         );
  NOR3_X1 U7305 ( .A1(n6394), .A2(n6354), .A3(n6353), .ZN(n6357) );
  OAI21_X1 U7306 ( .B1(n6357), .B2(n6356), .A(n6355), .ZN(n6361) );
  INV_X1 U7307 ( .A(n6392), .ZN(n6358) );
  AOI21_X1 U7308 ( .B1(n6358), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6359) );
  NAND3_X1 U7309 ( .A1(n6361), .A2(n6360), .A3(n6359), .ZN(n6396) );
  AOI22_X1 U7310 ( .A1(n6396), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6362), 
        .B2(n6394), .ZN(n6363) );
  OAI211_X1 U7311 ( .C1(n6365), .C2(n6407), .A(n6364), .B(n6363), .ZN(U3068)
         );
  AOI22_X1 U7312 ( .A1(n6367), .A2(n6393), .B1(n3006), .B2(n6392), .ZN(n6370)
         );
  AOI22_X1 U7313 ( .A1(n6396), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6368), 
        .B2(n6394), .ZN(n6369) );
  OAI211_X1 U7314 ( .C1(n6371), .C2(n6407), .A(n6370), .B(n6369), .ZN(U3069)
         );
  AOI22_X1 U7315 ( .A1(n6411), .A2(n6393), .B1(n6410), .B2(n6392), .ZN(n6374)
         );
  AOI22_X1 U7316 ( .A1(n6396), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6372), 
        .B2(n6394), .ZN(n6373) );
  OAI211_X1 U7317 ( .C1(n6375), .C2(n6407), .A(n6374), .B(n6373), .ZN(U3070)
         );
  AOI22_X1 U7318 ( .A1(n6417), .A2(n6393), .B1(n6416), .B2(n6392), .ZN(n6378)
         );
  AOI22_X1 U7319 ( .A1(n6396), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6376), 
        .B2(n6394), .ZN(n6377) );
  OAI211_X1 U7320 ( .C1(n6379), .C2(n6407), .A(n6378), .B(n6377), .ZN(U3071)
         );
  AOI22_X1 U7321 ( .A1(n6423), .A2(n6393), .B1(n6422), .B2(n6392), .ZN(n6382)
         );
  AOI22_X1 U7322 ( .A1(n6396), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6380), 
        .B2(n6394), .ZN(n6381) );
  OAI211_X1 U7323 ( .C1(n6383), .C2(n6407), .A(n6382), .B(n6381), .ZN(U3072)
         );
  AOI22_X1 U7324 ( .A1(n6429), .A2(n6393), .B1(n6428), .B2(n6392), .ZN(n6386)
         );
  AOI22_X1 U7325 ( .A1(n6396), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6384), 
        .B2(n6394), .ZN(n6385) );
  OAI211_X1 U7326 ( .C1(n6387), .C2(n6407), .A(n6386), .B(n6385), .ZN(U3073)
         );
  AOI22_X1 U7327 ( .A1(n6435), .A2(n6393), .B1(n6434), .B2(n6392), .ZN(n6390)
         );
  AOI22_X1 U7328 ( .A1(n6396), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6388), 
        .B2(n6394), .ZN(n6389) );
  OAI211_X1 U7329 ( .C1(n6391), .C2(n6407), .A(n6390), .B(n6389), .ZN(U3074)
         );
  AOI22_X1 U7330 ( .A1(n6444), .A2(n6393), .B1(n6442), .B2(n6392), .ZN(n6398)
         );
  AOI22_X1 U7331 ( .A1(n6396), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6395), 
        .B2(n6394), .ZN(n6397) );
  OAI211_X1 U7332 ( .C1(n6399), .C2(n6407), .A(n6398), .B(n6397), .ZN(U3075)
         );
  INV_X1 U7333 ( .A(n6400), .ZN(n6402) );
  AOI22_X1 U7334 ( .A1(n6416), .A2(n6402), .B1(n6415), .B2(n6401), .ZN(n6406)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6404), .B1(n6417), 
        .B2(n6403), .ZN(n6405) );
  OAI211_X1 U7336 ( .C1(n6420), .C2(n6407), .A(n6406), .B(n6405), .ZN(U3079)
         );
  INV_X1 U7337 ( .A(n6408), .ZN(n6441) );
  AOI22_X1 U7338 ( .A1(n6410), .A2(n6441), .B1(n6440), .B2(n6409), .ZN(n6413)
         );
  AOI22_X1 U7339 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6445), .B1(n6411), 
        .B2(n6443), .ZN(n6412) );
  OAI211_X1 U7340 ( .C1(n6414), .C2(n6448), .A(n6413), .B(n6412), .ZN(U3110)
         );
  AOI22_X1 U7341 ( .A1(n6416), .A2(n6441), .B1(n6440), .B2(n6415), .ZN(n6419)
         );
  AOI22_X1 U7342 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6445), .B1(n6417), 
        .B2(n6443), .ZN(n6418) );
  OAI211_X1 U7343 ( .C1(n6420), .C2(n6448), .A(n6419), .B(n6418), .ZN(U3111)
         );
  AOI22_X1 U7344 ( .A1(n6422), .A2(n6441), .B1(n6440), .B2(n6421), .ZN(n6425)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6445), .B1(n6423), 
        .B2(n6443), .ZN(n6424) );
  OAI211_X1 U7346 ( .C1(n6426), .C2(n6448), .A(n6425), .B(n6424), .ZN(U3112)
         );
  AOI22_X1 U7347 ( .A1(n6428), .A2(n6441), .B1(n6440), .B2(n6427), .ZN(n6431)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6445), .B1(n6429), 
        .B2(n6443), .ZN(n6430) );
  OAI211_X1 U7349 ( .C1(n6432), .C2(n6448), .A(n6431), .B(n6430), .ZN(U3113)
         );
  AOI22_X1 U7350 ( .A1(n6434), .A2(n6441), .B1(n6440), .B2(n6433), .ZN(n6437)
         );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6445), .B1(n6435), 
        .B2(n6443), .ZN(n6436) );
  OAI211_X1 U7352 ( .C1(n6438), .C2(n6448), .A(n6437), .B(n6436), .ZN(U3114)
         );
  AOI22_X1 U7353 ( .A1(n6442), .A2(n6441), .B1(n6440), .B2(n6439), .ZN(n6447)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6445), .B1(n6444), 
        .B2(n6443), .ZN(n6446) );
  OAI211_X1 U7355 ( .C1(n6449), .C2(n6448), .A(n6447), .B(n6446), .ZN(U3115)
         );
  INV_X1 U7356 ( .A(n6450), .ZN(n6464) );
  OAI211_X1 U7357 ( .C1(n3036), .C2(n6452), .A(n6451), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6456) );
  INV_X1 U7358 ( .A(n6453), .ZN(n6454) );
  OAI21_X1 U7359 ( .B1(n6455), .B2(n6456), .A(n6454), .ZN(n6458) );
  NAND2_X1 U7360 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  OAI21_X1 U7361 ( .B1(n6459), .B2(n6458), .A(n6457), .ZN(n6460) );
  AOI222_X1 U7362 ( .A1(n6462), .A2(n6461), .B1(n6462), .B2(n6460), .C1(n6461), 
        .C2(n6460), .ZN(n6463) );
  AOI222_X1 U7363 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6464), .B1(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6463), .C1(n6464), .C2(n6463), 
        .ZN(n6483) );
  NOR3_X1 U7364 ( .A1(n6466), .A2(n6476), .A3(n6465), .ZN(n6470) );
  INV_X1 U7365 ( .A(n6467), .ZN(n6469) );
  OAI22_X1 U7366 ( .A1(n6473), .A2(n6470), .B1(n6469), .B2(n6468), .ZN(n6471)
         );
  AOI21_X1 U7367 ( .B1(n6473), .B2(n6472), .A(n6471), .ZN(n6588) );
  INV_X1 U7368 ( .A(n6588), .ZN(n6474) );
  NOR4_X1 U7369 ( .A1(n6477), .A2(n6476), .A3(n6475), .A4(n6474), .ZN(n6480)
         );
  OAI21_X1 U7370 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6478), 
        .ZN(n6479) );
  NAND2_X1 U7371 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  AOI21_X1 U7372 ( .B1(n6483), .B2(n6482), .A(n6481), .ZN(n6495) );
  INV_X1 U7373 ( .A(n6495), .ZN(n6486) );
  OAI22_X1 U7374 ( .A1(n6486), .A2(n6498), .B1(n6485), .B2(n6484), .ZN(n6487)
         );
  OAI21_X1 U7375 ( .B1(n6489), .B2(n6488), .A(n6487), .ZN(n6579) );
  OAI21_X1 U7376 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6485), .A(n6579), .ZN(
        n6496) );
  AOI221_X1 U7377 ( .B1(n6491), .B2(STATE2_REG_0__SCAN_IN), .C1(n6496), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6490), .ZN(n6494) );
  OAI211_X1 U7378 ( .C1(n6504), .C2(n6492), .A(n3053), .B(n6579), .ZN(n6493)
         );
  OAI211_X1 U7379 ( .C1(n6495), .C2(n6498), .A(n6494), .B(n6493), .ZN(U3148)
         );
  NAND3_X1 U7380 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6497), .A3(n6496), .ZN(
        n6503) );
  OAI21_X1 U7381 ( .B1(READY_N), .B2(n6499), .A(n6498), .ZN(n6501) );
  AOI21_X1 U7382 ( .B1(n6501), .B2(n6579), .A(n6500), .ZN(n6502) );
  NAND2_X1 U7383 ( .A1(n6503), .A2(n6502), .ZN(U3149) );
  OAI211_X1 U7384 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6485), .A(n6578), .B(
        n6504), .ZN(n6506) );
  OAI21_X1 U7385 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(U3150) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6508), .ZN(U3151) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6508), .ZN(U3152) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6508), .ZN(U3153) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6508), .ZN(U3154) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6508), .ZN(U3155) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6508), .ZN(U3156) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6508), .ZN(U3157) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6508), .ZN(U3158) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6508), .ZN(U3159) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6508), .ZN(U3160) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6508), .ZN(U3161) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6508), .ZN(U3162) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6508), .ZN(U3163) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6508), .ZN(U3164) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6508), .ZN(U3165) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6508), .ZN(U3166) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6508), .ZN(U3167) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6508), .ZN(U3168) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6508), .ZN(U3169) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6508), .ZN(U3170) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6508), .ZN(U3171) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6508), .ZN(U3172) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6508), .ZN(U3173) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6508), .ZN(U3174) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6508), .ZN(U3175) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6508), .ZN(U3176) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6508), .ZN(U3177) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6508), .ZN(U3178) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6508), .ZN(U3179) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6508), .ZN(U3180) );
  INV_X1 U7416 ( .A(n6523), .ZN(n6510) );
  AOI22_X1 U7417 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6524) );
  INV_X1 U7418 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6519) );
  INV_X1 U7419 ( .A(HOLD), .ZN(n6652) );
  NOR2_X1 U7420 ( .A1(n6519), .A2(n6652), .ZN(n6511) );
  INV_X1 U7421 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6739) );
  OAI21_X1 U7422 ( .B1(n6511), .B2(n6739), .A(n6790), .ZN(n6509) );
  OAI211_X1 U7423 ( .C1(NA_N), .C2(n6515), .A(n6520), .B(n6523), .ZN(n6516) );
  OAI211_X1 U7424 ( .C1(n6510), .C2(n6524), .A(n6509), .B(n6516), .ZN(U3181)
         );
  NOR2_X1 U7425 ( .A1(n6520), .A2(n6739), .ZN(n6512) );
  OAI22_X1 U7426 ( .A1(n6512), .A2(n6511), .B1(n6515), .B2(n6652), .ZN(n6513)
         );
  OAI211_X1 U7427 ( .C1(n6519), .C2(n6485), .A(n6514), .B(n6513), .ZN(U3182)
         );
  INV_X1 U7428 ( .A(NA_N), .ZN(n6707) );
  NAND2_X1 U7429 ( .A1(READY_N), .A2(n6707), .ZN(n6518) );
  OAI221_X1 U7430 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_1__SCAN_IN), 
        .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6518), .A(n6515), .ZN(n6517) );
  OAI211_X1 U7431 ( .C1(n6520), .C2(HOLD), .A(n6517), .B(n6516), .ZN(n6522) );
  OR4_X1 U7432 ( .A1(n6520), .A2(n6519), .A3(n6739), .A4(n6518), .ZN(n6521) );
  OAI211_X1 U7433 ( .C1(n6524), .C2(n6523), .A(n6522), .B(n6521), .ZN(U3183)
         );
  NOR2_X2 U7434 ( .A1(n6790), .A2(STATE_REG_2__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7435 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6791), .ZN(n6572) );
  INV_X1 U7436 ( .A(n6572), .ZN(n6563) );
  AOI22_X1 U7437 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6790), .ZN(n6525) );
  OAI21_X1 U7438 ( .B1(n6526), .B2(n6565), .A(n6525), .ZN(U3184) );
  INV_X1 U7439 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6529) );
  AOI22_X1 U7440 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6790), .ZN(n6527) );
  OAI21_X1 U7441 ( .B1(n6529), .B2(n6565), .A(n6527), .ZN(U3185) );
  AOI22_X1 U7442 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6790), .ZN(n6528) );
  OAI21_X1 U7443 ( .B1(n6529), .B2(n6572), .A(n6528), .ZN(U3186) );
  AOI22_X1 U7444 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6790), .ZN(n6530) );
  OAI21_X1 U7445 ( .B1(n6532), .B2(n6565), .A(n6530), .ZN(U3187) );
  AOI22_X1 U7446 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6790), .ZN(n6531) );
  OAI21_X1 U7447 ( .B1(n6532), .B2(n6572), .A(n6531), .ZN(U3188) );
  AOI22_X1 U7448 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6790), .ZN(n6533) );
  OAI21_X1 U7449 ( .B1(n6535), .B2(n6565), .A(n6533), .ZN(U3189) );
  AOI22_X1 U7450 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6790), .ZN(n6534) );
  OAI21_X1 U7451 ( .B1(n6535), .B2(n6572), .A(n6534), .ZN(U3190) );
  AOI22_X1 U7452 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6790), .ZN(n6536) );
  OAI21_X1 U7453 ( .B1(n6537), .B2(n6565), .A(n6536), .ZN(U3191) );
  AOI22_X1 U7454 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6790), .ZN(n6538) );
  OAI21_X1 U7455 ( .B1(n6540), .B2(n6565), .A(n6538), .ZN(U3192) );
  AOI22_X1 U7456 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6790), .ZN(n6539) );
  OAI21_X1 U7457 ( .B1(n6540), .B2(n6572), .A(n6539), .ZN(U3193) );
  AOI22_X1 U7458 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6790), .ZN(n6541) );
  OAI21_X1 U7459 ( .B1(n6542), .B2(n6565), .A(n6541), .ZN(U3194) );
  AOI22_X1 U7460 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6790), .ZN(n6543) );
  OAI21_X1 U7461 ( .B1(n6544), .B2(n6565), .A(n6543), .ZN(U3195) );
  INV_X1 U7462 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6547) );
  AOI22_X1 U7463 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6790), .ZN(n6545) );
  OAI21_X1 U7464 ( .B1(n6547), .B2(n6565), .A(n6545), .ZN(U3196) );
  AOI22_X1 U7465 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6790), .ZN(n6546) );
  OAI21_X1 U7466 ( .B1(n6547), .B2(n6572), .A(n6546), .ZN(U3197) );
  AOI22_X1 U7467 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6790), .ZN(n6548) );
  OAI21_X1 U7468 ( .B1(n6549), .B2(n6572), .A(n6548), .ZN(U3198) );
  AOI22_X1 U7469 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6790), .ZN(n6550) );
  OAI21_X1 U7470 ( .B1(n6551), .B2(n6572), .A(n6550), .ZN(U3199) );
  AOI22_X1 U7471 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6790), .ZN(n6552) );
  OAI21_X1 U7472 ( .B1(n6554), .B2(n6565), .A(n6552), .ZN(U3200) );
  AOI22_X1 U7473 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6790), .ZN(n6553) );
  OAI21_X1 U7474 ( .B1(n6554), .B2(n6572), .A(n6553), .ZN(U3201) );
  INV_X1 U7475 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6673) );
  AOI22_X1 U7476 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6790), .ZN(n6555) );
  OAI21_X1 U7477 ( .B1(n6673), .B2(n6565), .A(n6555), .ZN(U3202) );
  AOI22_X1 U7478 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6790), .ZN(n6556) );
  OAI21_X1 U7479 ( .B1(n6673), .B2(n6572), .A(n6556), .ZN(U3203) );
  INV_X1 U7480 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6757) );
  AOI22_X1 U7481 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6790), .ZN(n6557) );
  OAI21_X1 U7482 ( .B1(n6757), .B2(n6572), .A(n6557), .ZN(U3204) );
  AOI22_X1 U7483 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6790), .ZN(n6558) );
  OAI21_X1 U7484 ( .B1(n6560), .B2(n6565), .A(n6558), .ZN(U3205) );
  AOI22_X1 U7485 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6790), .ZN(n6559) );
  OAI21_X1 U7486 ( .B1(n6560), .B2(n6572), .A(n6559), .ZN(U3206) );
  AOI22_X1 U7487 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6790), .ZN(n6561) );
  OAI21_X1 U7488 ( .B1(n6653), .B2(n6565), .A(n6561), .ZN(U3207) );
  AOI22_X1 U7489 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6790), .ZN(n6562) );
  OAI21_X1 U7490 ( .B1(n6731), .B2(n6565), .A(n6562), .ZN(U3208) );
  INV_X1 U7491 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6567) );
  AOI22_X1 U7492 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6563), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6790), .ZN(n6564) );
  OAI21_X1 U7493 ( .B1(n6567), .B2(n6565), .A(n6564), .ZN(U3209) );
  AOI22_X1 U7494 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6790), .ZN(n6566) );
  OAI21_X1 U7495 ( .B1(n6567), .B2(n6572), .A(n6566), .ZN(U3210) );
  AOI22_X1 U7496 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6790), .ZN(n6568) );
  OAI21_X1 U7497 ( .B1(n6706), .B2(n6572), .A(n6568), .ZN(U3211) );
  AOI22_X1 U7498 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6790), .ZN(n6569) );
  OAI21_X1 U7499 ( .B1(n6719), .B2(n6572), .A(n6569), .ZN(U3212) );
  AOI22_X1 U7500 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6790), .ZN(n6571) );
  OAI21_X1 U7501 ( .B1(n6573), .B2(n6572), .A(n6571), .ZN(U3213) );
  MUX2_X1 U7502 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6790), .Z(U3446) );
  MUX2_X1 U7503 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6790), .Z(U3447) );
  MUX2_X1 U7504 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6790), .Z(U3448) );
  OAI21_X1 U7505 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6577), .A(n6575), .ZN(
        n6574) );
  INV_X1 U7506 ( .A(n6574), .ZN(U3451) );
  OAI21_X1 U7507 ( .B1(n6577), .B2(n6576), .A(n6575), .ZN(U3452) );
  OAI221_X1 U7508 ( .B1(n6580), .B2(STATE2_REG_0__SCAN_IN), .C1(n6580), .C2(
        n6579), .A(n6578), .ZN(U3453) );
  AOI21_X1 U7509 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6581) );
  AOI22_X1 U7510 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6581), .B2(n5069), .ZN(n6584) );
  INV_X1 U7511 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6583) );
  AOI22_X1 U7512 ( .A1(n6586), .A2(n6584), .B1(n6583), .B2(n6582), .ZN(U3468)
         );
  INV_X1 U7513 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6718) );
  OAI21_X1 U7514 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6586), .ZN(n6585) );
  OAI21_X1 U7515 ( .B1(n6586), .B2(n6718), .A(n6585), .ZN(U3469) );
  INV_X1 U7516 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6737) );
  AOI22_X1 U7517 ( .A1(n6791), .A2(READREQUEST_REG_SCAN_IN), .B1(n6737), .B2(
        n6790), .ZN(U3470) );
  INV_X1 U7518 ( .A(MORE_REG_SCAN_IN), .ZN(n6691) );
  INV_X1 U7519 ( .A(n6589), .ZN(n6587) );
  AOI22_X1 U7520 ( .A1(n6589), .A2(n6588), .B1(n6691), .B2(n6587), .ZN(U3471)
         );
  AOI211_X1 U7521 ( .C1(n6592), .C2(n6485), .A(n6591), .B(n6590), .ZN(n6599)
         );
  OAI211_X1 U7522 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6594), .A(n6593), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6596) );
  AOI21_X1 U7523 ( .B1(n6596), .B2(STATE2_REG_0__SCAN_IN), .A(n6595), .ZN(
        n6598) );
  NAND2_X1 U7524 ( .A1(n6599), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6597) );
  OAI21_X1 U7525 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(U3472) );
  INV_X1 U7526 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6642) );
  INV_X1 U7527 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7528 ( .A1(n6791), .A2(n6642), .B1(n6668), .B2(n6790), .ZN(U3473)
         );
  INV_X1 U7529 ( .A(DATAI_10_), .ZN(n6789) );
  AOI22_X1 U7530 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_f55), .ZN(n6600) );
  OAI221_X1 U7531 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(REIP_REG_27__SCAN_IN), .C2(keyinput_f55), .A(n6600), .ZN(n6607) );
  AOI22_X1 U7532 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_9_), .B2(
        keyinput_f22), .ZN(n6601) );
  OAI221_X1 U7533 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(DATAI_9_), .C2(
        keyinput_f22), .A(n6601), .ZN(n6606) );
  AOI22_X1 U7534 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(DATAI_30_), .B2(
        keyinput_f1), .ZN(n6602) );
  OAI221_X1 U7535 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(DATAI_30_), .C2(
        keyinput_f1), .A(n6602), .ZN(n6605) );
  AOI22_X1 U7536 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(DATAI_3_), .B2(
        keyinput_f28), .ZN(n6603) );
  OAI221_X1 U7537 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(DATAI_3_), .C2(
        keyinput_f28), .A(n6603), .ZN(n6604) );
  NOR4_X1 U7538 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n6634)
         );
  XNOR2_X1 U7539 ( .A(DATAI_22_), .B(keyinput_f9), .ZN(n6614) );
  AOI22_X1 U7540 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(n5834), .B2(
        keyinput_f63), .ZN(n6608) );
  OAI221_X1 U7541 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(n5834), .C2(
        keyinput_f63), .A(n6608), .ZN(n6613) );
  AOI22_X1 U7542 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .ZN(n6609) );
  OAI221_X1 U7543 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_f51), .A(n6609), .ZN(n6612) );
  AOI22_X1 U7544 ( .A1(keyinput_f49), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        DATAI_20_), .B2(keyinput_f11), .ZN(n6610) );
  OAI221_X1 U7545 ( .B1(keyinput_f49), .B2(BYTEENABLE_REG_2__SCAN_IN), .C1(
        DATAI_20_), .C2(keyinput_f11), .A(n6610), .ZN(n6611) );
  NOR4_X1 U7546 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n6633)
         );
  AOI22_X1 U7547 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .ZN(n6615) );
  OAI221_X1 U7548 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_f60), .A(n6615), .ZN(n6622) );
  AOI22_X1 U7549 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_f45), .B1(DATAI_16_), 
        .B2(keyinput_f15), .ZN(n6616) );
  OAI221_X1 U7550 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_f45), .C1(DATAI_16_), 
        .C2(keyinput_f15), .A(n6616), .ZN(n6621) );
  AOI22_X1 U7551 ( .A1(keyinput_f47), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_f59), .ZN(n6617) );
  OAI221_X1 U7552 ( .B1(keyinput_f47), .B2(BYTEENABLE_REG_0__SCAN_IN), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_f59), .A(n6617), .ZN(n6620) );
  AOI22_X1 U7553 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .ZN(n6618) );
  OAI221_X1 U7554 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_f53), .A(n6618), .ZN(n6619) );
  NOR4_X1 U7555 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6632)
         );
  AOI22_X1 U7556 ( .A1(keyinput_f48), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .ZN(n6623) );
  OAI221_X1 U7557 ( .B1(keyinput_f48), .B2(BYTEENABLE_REG_1__SCAN_IN), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_f52), .A(n6623), .ZN(n6630) );
  AOI22_X1 U7558 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(keyinput_f34), .B2(BS16_N), .ZN(n6624) );
  OAI221_X1 U7559 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(
        keyinput_f34), .C2(BS16_N), .A(n6624), .ZN(n6629) );
  AOI22_X1 U7560 ( .A1(keyinput_f50), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        DATAI_7_), .B2(keyinput_f24), .ZN(n6625) );
  OAI221_X1 U7561 ( .B1(keyinput_f50), .B2(BYTEENABLE_REG_3__SCAN_IN), .C1(
        DATAI_7_), .C2(keyinput_f24), .A(n6625), .ZN(n6628) );
  AOI22_X1 U7562 ( .A1(keyinput_f41), .A2(D_C_N_REG_SCAN_IN), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .ZN(n6626) );
  OAI221_X1 U7563 ( .B1(keyinput_f41), .B2(D_C_N_REG_SCAN_IN), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_f54), .A(n6626), .ZN(n6627) );
  NOR4_X1 U7564 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n6631)
         );
  NAND4_X1 U7565 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6685)
         );
  AOI22_X1 U7566 ( .A1(n6636), .A2(keyinput_f23), .B1(n6731), .B2(keyinput_f56), .ZN(n6635) );
  OAI221_X1 U7567 ( .B1(n6636), .B2(keyinput_f23), .C1(n6731), .C2(
        keyinput_f56), .A(n6635), .ZN(n6646) );
  INV_X1 U7568 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7569 ( .A1(n6736), .A2(keyinput_f39), .B1(n6638), .B2(keyinput_f5), 
        .ZN(n6637) );
  OAI221_X1 U7570 ( .B1(n6736), .B2(keyinput_f39), .C1(n6638), .C2(keyinput_f5), .A(n6637), .ZN(n6645) );
  AOI22_X1 U7571 ( .A1(n6697), .A2(keyinput_f38), .B1(n5298), .B2(keyinput_f19), .ZN(n6639) );
  OAI221_X1 U7572 ( .B1(n6697), .B2(keyinput_f38), .C1(n5298), .C2(
        keyinput_f19), .A(n6639), .ZN(n6644) );
  AOI22_X1 U7573 ( .A1(n6642), .A2(keyinput_f32), .B1(n6641), .B2(keyinput_f25), .ZN(n6640) );
  OAI221_X1 U7574 ( .B1(n6642), .B2(keyinput_f32), .C1(n6641), .C2(
        keyinput_f25), .A(n6640), .ZN(n6643) );
  NOR4_X1 U7575 ( .A1(n6646), .A2(n6645), .A3(n6644), .A4(n6643), .ZN(n6683)
         );
  AOI22_X1 U7576 ( .A1(n6757), .A2(keyinput_f61), .B1(keyinput_f33), .B2(n6707), .ZN(n6647) );
  OAI221_X1 U7577 ( .B1(n6757), .B2(keyinput_f61), .C1(n6707), .C2(
        keyinput_f33), .A(n6647), .ZN(n6657) );
  AOI22_X1 U7578 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(n6733), .B2(
        keyinput_f6), .ZN(n6648) );
  OAI221_X1 U7579 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(n6733), .C2(
        keyinput_f6), .A(n6648), .ZN(n6656) );
  AOI22_X1 U7580 ( .A1(n6739), .A2(keyinput_f42), .B1(n6650), .B2(keyinput_f0), 
        .ZN(n6649) );
  OAI221_X1 U7581 ( .B1(n6739), .B2(keyinput_f42), .C1(n6650), .C2(keyinput_f0), .A(n6649), .ZN(n6655) );
  AOI22_X1 U7582 ( .A1(n6653), .A2(keyinput_f57), .B1(keyinput_f36), .B2(n6652), .ZN(n6651) );
  OAI221_X1 U7583 ( .B1(n6653), .B2(keyinput_f57), .C1(n6652), .C2(
        keyinput_f36), .A(n6651), .ZN(n6654) );
  NOR4_X1 U7584 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6682)
         );
  AOI22_X1 U7585 ( .A1(n6691), .A2(keyinput_f44), .B1(n6715), .B2(keyinput_f43), .ZN(n6658) );
  OAI221_X1 U7586 ( .B1(n6691), .B2(keyinput_f44), .C1(n6715), .C2(
        keyinput_f43), .A(n6658), .ZN(n6666) );
  INV_X1 U7587 ( .A(DATAI_13_), .ZN(n6734) );
  INV_X1 U7588 ( .A(DATAI_15_), .ZN(n6740) );
  AOI22_X1 U7589 ( .A1(n6734), .A2(keyinput_f18), .B1(keyinput_f16), .B2(n6740), .ZN(n6659) );
  OAI221_X1 U7590 ( .B1(n6734), .B2(keyinput_f18), .C1(n6740), .C2(
        keyinput_f16), .A(n6659), .ZN(n6665) );
  INV_X1 U7591 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6696) );
  AOI22_X1 U7592 ( .A1(n6696), .A2(keyinput_f37), .B1(n6661), .B2(keyinput_f29), .ZN(n6660) );
  OAI221_X1 U7593 ( .B1(n6696), .B2(keyinput_f37), .C1(n6661), .C2(
        keyinput_f29), .A(n6660), .ZN(n6664) );
  AOI22_X1 U7594 ( .A1(n6485), .A2(keyinput_f35), .B1(keyinput_f2), .B2(n6725), 
        .ZN(n6662) );
  OAI221_X1 U7595 ( .B1(n6485), .B2(keyinput_f35), .C1(n6725), .C2(keyinput_f2), .A(n6662), .ZN(n6663) );
  NOR4_X1 U7596 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6681)
         );
  AOI22_X1 U7597 ( .A1(n6669), .A2(keyinput_f58), .B1(keyinput_f40), .B2(n6668), .ZN(n6667) );
  OAI221_X1 U7598 ( .B1(n6669), .B2(keyinput_f58), .C1(n6668), .C2(
        keyinput_f40), .A(n6667), .ZN(n6679) );
  INV_X1 U7599 ( .A(DATAI_14_), .ZN(n6671) );
  AOI22_X1 U7600 ( .A1(n6671), .A2(keyinput_f17), .B1(keyinput_f12), .B2(n4508), .ZN(n6670) );
  OAI221_X1 U7601 ( .B1(n6671), .B2(keyinput_f17), .C1(n4508), .C2(
        keyinput_f12), .A(n6670), .ZN(n6678) );
  AOI22_X1 U7602 ( .A1(n6673), .A2(keyinput_f62), .B1(keyinput_f14), .B2(n4497), .ZN(n6672) );
  OAI221_X1 U7603 ( .B1(n6673), .B2(keyinput_f62), .C1(n4497), .C2(
        keyinput_f14), .A(n6672), .ZN(n6677) );
  AOI22_X1 U7604 ( .A1(n6675), .A2(keyinput_f30), .B1(n6694), .B2(keyinput_f27), .ZN(n6674) );
  OAI221_X1 U7605 ( .B1(n6675), .B2(keyinput_f30), .C1(n6694), .C2(
        keyinput_f27), .A(n6674), .ZN(n6676) );
  NOR4_X1 U7606 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6680)
         );
  NAND4_X1 U7607 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  OAI22_X1 U7608 ( .A1(keyinput_f21), .A2(n6789), .B1(n6685), .B2(n6684), .ZN(
        n6686) );
  AOI21_X1 U7609 ( .B1(keyinput_f21), .B2(n6789), .A(n6686), .ZN(n6788) );
  INV_X1 U7610 ( .A(BS16_N), .ZN(n6688) );
  AOI22_X1 U7611 ( .A1(n6689), .A2(keyinput_g31), .B1(keyinput_g34), .B2(n6688), .ZN(n6687) );
  OAI221_X1 U7612 ( .B1(n6689), .B2(keyinput_g31), .C1(n6688), .C2(
        keyinput_g34), .A(n6687), .ZN(n6701) );
  AOI22_X1 U7613 ( .A1(n4526), .A2(keyinput_g8), .B1(keyinput_g44), .B2(n6691), 
        .ZN(n6690) );
  OAI221_X1 U7614 ( .B1(n4526), .B2(keyinput_g8), .C1(n6691), .C2(keyinput_g44), .A(n6690), .ZN(n6700) );
  INV_X1 U7615 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6693) );
  AOI22_X1 U7616 ( .A1(n6694), .A2(keyinput_g27), .B1(n6693), .B2(keyinput_g51), .ZN(n6692) );
  OAI221_X1 U7617 ( .B1(n6694), .B2(keyinput_g27), .C1(n6693), .C2(
        keyinput_g51), .A(n6692), .ZN(n6699) );
  AOI22_X1 U7618 ( .A1(n6697), .A2(keyinput_g38), .B1(n6696), .B2(keyinput_g37), .ZN(n6695) );
  OAI221_X1 U7619 ( .B1(n6697), .B2(keyinput_g38), .C1(n6696), .C2(
        keyinput_g37), .A(n6695), .ZN(n6698) );
  NOR4_X1 U7620 ( .A1(n6701), .A2(n6700), .A3(n6699), .A4(n6698), .ZN(n6748)
         );
  AOI22_X1 U7621 ( .A1(n6485), .A2(keyinput_g35), .B1(keyinput_g1), .B2(n6703), 
        .ZN(n6702) );
  OAI221_X1 U7622 ( .B1(n6485), .B2(keyinput_g35), .C1(n6703), .C2(keyinput_g1), .A(n6702), .ZN(n6713) );
  AOI22_X1 U7623 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6704) );
  OAI221_X1 U7624 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6704), .ZN(n6712) );
  AOI22_X1 U7625 ( .A1(n6707), .A2(keyinput_g33), .B1(n6706), .B2(keyinput_g54), .ZN(n6705) );
  OAI221_X1 U7626 ( .B1(n6707), .B2(keyinput_g33), .C1(n6706), .C2(
        keyinput_g54), .A(n6705), .ZN(n6711) );
  AOI22_X1 U7627 ( .A1(n5298), .A2(keyinput_g19), .B1(keyinput_g45), .B2(n6709), .ZN(n6708) );
  OAI221_X1 U7628 ( .B1(n5298), .B2(keyinput_g19), .C1(n6709), .C2(
        keyinput_g45), .A(n6708), .ZN(n6710) );
  NOR4_X1 U7629 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6747)
         );
  INV_X1 U7630 ( .A(DATAI_20_), .ZN(n6716) );
  AOI22_X1 U7631 ( .A1(n6716), .A2(keyinput_g11), .B1(n6715), .B2(keyinput_g43), .ZN(n6714) );
  OAI221_X1 U7632 ( .B1(n6716), .B2(keyinput_g11), .C1(n6715), .C2(
        keyinput_g43), .A(n6714), .ZN(n6729) );
  AOI22_X1 U7633 ( .A1(n6719), .A2(keyinput_g53), .B1(keyinput_g47), .B2(n6718), .ZN(n6717) );
  OAI221_X1 U7634 ( .B1(n6719), .B2(keyinput_g53), .C1(n6718), .C2(
        keyinput_g47), .A(n6717), .ZN(n6728) );
  INV_X1 U7635 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7636 ( .A1(n6722), .A2(keyinput_g22), .B1(n6721), .B2(keyinput_g60), .ZN(n6720) );
  OAI221_X1 U7637 ( .B1(n6722), .B2(keyinput_g22), .C1(n6721), .C2(
        keyinput_g60), .A(n6720), .ZN(n6727) );
  AOI22_X1 U7638 ( .A1(n6725), .A2(keyinput_g2), .B1(keyinput_g50), .B2(n6724), 
        .ZN(n6723) );
  OAI221_X1 U7639 ( .B1(n6725), .B2(keyinput_g2), .C1(n6724), .C2(keyinput_g50), .A(n6723), .ZN(n6726) );
  NOR4_X1 U7640 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6746)
         );
  AOI22_X1 U7641 ( .A1(n6731), .A2(keyinput_g56), .B1(keyinput_g14), .B2(n4497), .ZN(n6730) );
  OAI221_X1 U7642 ( .B1(n6731), .B2(keyinput_g56), .C1(n4497), .C2(
        keyinput_g14), .A(n6730), .ZN(n6744) );
  AOI22_X1 U7643 ( .A1(n6734), .A2(keyinput_g18), .B1(keyinput_g6), .B2(n6733), 
        .ZN(n6732) );
  OAI221_X1 U7644 ( .B1(n6734), .B2(keyinput_g18), .C1(n6733), .C2(keyinput_g6), .A(n6732), .ZN(n6743) );
  AOI22_X1 U7645 ( .A1(n6737), .A2(keyinput_g46), .B1(n6736), .B2(keyinput_g39), .ZN(n6735) );
  OAI221_X1 U7646 ( .B1(n6737), .B2(keyinput_g46), .C1(n6736), .C2(
        keyinput_g39), .A(n6735), .ZN(n6742) );
  AOI22_X1 U7647 ( .A1(n6740), .A2(keyinput_g16), .B1(keyinput_g42), .B2(n6739), .ZN(n6738) );
  OAI221_X1 U7648 ( .B1(n6740), .B2(keyinput_g16), .C1(n6739), .C2(
        keyinput_g42), .A(n6738), .ZN(n6741) );
  NOR4_X1 U7649 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6745)
         );
  NAND4_X1 U7650 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6786)
         );
  AOI22_X1 U7651 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_24_), .B2(
        keyinput_g7), .ZN(n6749) );
  OAI221_X1 U7652 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_24_), .C2(
        keyinput_g7), .A(n6749), .ZN(n6756) );
  AOI22_X1 U7653 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(DATAI_22_), .B2(
        keyinput_g9), .ZN(n6750) );
  OAI221_X1 U7654 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_22_), .C2(
        keyinput_g9), .A(n6750), .ZN(n6755) );
  AOI22_X1 U7655 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n6751) );
  OAI221_X1 U7656 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n6751), .ZN(n6754) );
  AOI22_X1 U7657 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n6752) );
  OAI221_X1 U7658 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(DATAI_11_), .C2(
        keyinput_g20), .A(n6752), .ZN(n6753) );
  NOR4_X1 U7659 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6784)
         );
  XNOR2_X1 U7660 ( .A(n6757), .B(keyinput_g61), .ZN(n6764) );
  AOI22_X1 U7661 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n6758) );
  OAI221_X1 U7662 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(REIP_REG_19__SCAN_IN), .C2(keyinput_g63), .A(n6758), .ZN(n6763) );
  AOI22_X1 U7663 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_7_), .B2(
        keyinput_g24), .ZN(n6759) );
  OAI221_X1 U7664 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_7_), .C2(
        keyinput_g24), .A(n6759), .ZN(n6762) );
  AOI22_X1 U7665 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_g40), .B1(DATAI_1_), 
        .B2(keyinput_g30), .ZN(n6760) );
  OAI221_X1 U7666 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .C1(DATAI_1_), 
        .C2(keyinput_g30), .A(n6760), .ZN(n6761) );
  NOR4_X1 U7667 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6783)
         );
  AOI22_X1 U7668 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g49), .ZN(n6765) );
  OAI221_X1 U7669 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_g49), .A(n6765), .ZN(n6772)
         );
  AOI22_X1 U7670 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_g62), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6766) );
  OAI221_X1 U7671 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6766), .ZN(n6771) );
  AOI22_X1 U7672 ( .A1(HOLD), .A2(keyinput_g36), .B1(DATAI_8_), .B2(
        keyinput_g23), .ZN(n6767) );
  OAI221_X1 U7673 ( .B1(HOLD), .B2(keyinput_g36), .C1(DATAI_8_), .C2(
        keyinput_g23), .A(n6767), .ZN(n6770) );
  AOI22_X1 U7674 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6768) );
  OAI221_X1 U7675 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6768), .ZN(n6769) );
  NOR4_X1 U7676 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6782)
         );
  AOI22_X1 U7677 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(DATAI_27_), .B2(
        keyinput_g4), .ZN(n6773) );
  OAI221_X1 U7678 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(DATAI_27_), .C2(
        keyinput_g4), .A(n6773), .ZN(n6780) );
  AOI22_X1 U7679 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        DATAI_26_), .B2(keyinput_g5), .ZN(n6774) );
  OAI221_X1 U7680 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        DATAI_26_), .C2(keyinput_g5), .A(n6774), .ZN(n6779) );
  AOI22_X1 U7681 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_g55), .ZN(n6775) );
  OAI221_X1 U7682 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6775), .ZN(n6778) );
  AOI22_X1 U7683 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(REIP_REG_30__SCAN_IN), 
        .B2(keyinput_g52), .ZN(n6776) );
  OAI221_X1 U7684 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(REIP_REG_30__SCAN_IN), .C2(keyinput_g52), .A(n6776), .ZN(n6777) );
  NOR4_X1 U7685 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6781)
         );
  NAND4_X1 U7686 ( .A1(n6784), .A2(n6783), .A3(n6782), .A4(n6781), .ZN(n6785)
         );
  OAI22_X1 U7687 ( .A1(keyinput_g21), .A2(n6789), .B1(n6786), .B2(n6785), .ZN(
        n6787) );
  AOI211_X1 U7688 ( .C1(keyinput_g21), .C2(n6789), .A(n6788), .B(n6787), .ZN(
        n6793) );
  AOI22_X1 U7689 ( .A1(n6791), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6790), .ZN(n6792) );
  XNOR2_X1 U7690 ( .A(n6793), .B(n6792), .ZN(U3445) );
  AND2_X1 U3972 ( .A1(n4435), .A2(n4445), .ZN(n3283) );
  AND2_X1 U4114 ( .A1(n4445), .A2(n4404), .ZN(n3323) );
  CLKBUF_X2 U3444 ( .A(n3283), .Z(n4085) );
  CLKBUF_X1 U34530 ( .A(n4230), .Z(n2998) );
  CLKBUF_X1 U34630 ( .A(n5681), .Z(n2991) );
  CLKBUF_X1 U34650 ( .A(n4429), .Z(n3003) );
  OR2_X1 U3540 ( .A1(n4406), .A2(n4378), .ZN(n6794) );
  AND2_X1 U3547 ( .A1(n3140), .A2(n4430), .ZN(n3276) );
endmodule

