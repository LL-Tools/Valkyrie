

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3426, n3427, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211;

  CLKBUF_X2 U34600 ( .A(n5105), .Z(n5162) );
  AND2_X1 U34610 ( .A1(n4001), .A2(n4000), .ZN(n5985) );
  OR2_X1 U34620 ( .A1(n3768), .A2(n3767), .ZN(n3769) );
  CLKBUF_X2 U34630 ( .A(n5829), .Z(n5850) );
  CLKBUF_X2 U34640 ( .A(n3702), .Z(n5860) );
  CLKBUF_X2 U34650 ( .A(n3720), .Z(n5966) );
  CLKBUF_X2 U3466 ( .A(n3639), .Z(n5859) );
  NAND2_X1 U3467 ( .A1(n4519), .A2(n3675), .ZN(n5145) );
  CLKBUF_X2 U34680 ( .A(n3661), .Z(n4680) );
  AND2_X1 U34690 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5124) );
  INV_X2 U34700 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3513) );
  CLKBUF_X1 U34710 ( .A(n5876), .Z(n3426) );
  NOR2_X1 U34720 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), 
        .ZN(n5876) );
  INV_X2 U34740 ( .A(n3677), .ZN(n4528) );
  INV_X1 U3475 ( .A(n5805), .ZN(n5819) );
  INV_X1 U3476 ( .A(n3661), .ZN(n3675) );
  AND2_X1 U3477 ( .A1(n3675), .A2(n3677), .ZN(n3836) );
  NOR2_X1 U3478 ( .A1(n6050), .A2(n6031), .ZN(n6030) );
  NAND2_X1 U3479 ( .A1(n3913), .A2(n3924), .ZN(n5895) );
  AND3_X1 U3480 ( .A1(n3576), .A2(n3575), .A3(n3574), .ZN(n3582) );
  INV_X1 U3481 ( .A(n7061), .ZN(n7101) );
  NAND2_X1 U3483 ( .A1(n4485), .A2(n7136), .ZN(n7108) );
  CLKBUF_X3 U3484 ( .A(n3640), .Z(n3433) );
  INV_X1 U3485 ( .A(n4639), .ZN(n4863) );
  INV_X2 U3486 ( .A(n3830), .ZN(n3508) );
  NAND2_X2 U3487 ( .A1(n3793), .A2(n3792), .ZN(n3830) );
  AND4_X2 U3488 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3559)
         );
  NAND2_X4 U3489 ( .A1(n3582), .A2(n3581), .ZN(n4006) );
  AND2_X4 U3490 ( .A1(n3502), .A2(n3501), .ZN(n4462) );
  BUF_X4 U3491 ( .A(n3645), .Z(n4363) );
  NAND2_X4 U3492 ( .A1(n4503), .A2(n3427), .ZN(n4965) );
  NAND4_X2 U3494 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3427)
         );
  XNOR2_X2 U3497 ( .A(n3768), .B(n3766), .ZN(n3490) );
  NAND2_X2 U3498 ( .A1(n3712), .A2(n3711), .ZN(n3768) );
  XNOR2_X2 U3499 ( .A(n5143), .B(n5141), .ZN(n4636) );
  NAND2_X2 U3500 ( .A1(n3809), .A2(n3808), .ZN(n5143) );
  NAND2_X1 U3501 ( .A1(n5607), .A2(n5606), .ZN(n5605) );
  NAND2_X1 U3502 ( .A1(n3903), .A2(n3902), .ZN(n3913) );
  NAND2_X1 U3503 ( .A1(n3861), .A2(n3831), .ZN(n4869) );
  CLKBUF_X2 U3504 ( .A(n4144), .Z(n5855) );
  BUF_X2 U3505 ( .A(n3820), .Z(n5858) );
  BUF_X2 U3506 ( .A(n3713), .Z(n5845) );
  BUF_X2 U3507 ( .A(n3719), .Z(n4436) );
  BUF_X2 U3508 ( .A(n4096), .Z(n5856) );
  BUF_X2 U3509 ( .A(n3714), .Z(n5849) );
  BUF_X2 U3510 ( .A(n3866), .Z(n5848) );
  AND2_X2 U3511 ( .A1(n3531), .A2(n5124), .ZN(n3702) );
  NOR2_X2 U3512 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3530) );
  AND2_X2 U3513 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4535) );
  OAI21_X1 U3514 ( .B1(n6191), .B2(n5898), .A(n6182), .ZN(n5936) );
  AND2_X1 U3515 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  OR2_X1 U3516 ( .A1(n6168), .A2(n6291), .ZN(n4458) );
  OAI21_X1 U3517 ( .B1(n4448), .B2(n4449), .A(n5842), .ZN(n6168) );
  NOR2_X2 U3518 ( .A1(n6060), .A2(n3482), .ZN(n6046) );
  AND2_X1 U3519 ( .A1(n5622), .A2(n3447), .ZN(n5680) );
  NAND2_X1 U3520 ( .A1(n5574), .A2(n4165), .ZN(n5622) );
  OR2_X1 U3521 ( .A1(n3909), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6793)
         );
  XNOR2_X1 U3522 ( .A(n3913), .B(n3912), .ZN(n4059) );
  AND2_X1 U3523 ( .A1(n3471), .A2(n4023), .ZN(n4599) );
  INV_X1 U3524 ( .A(n4869), .ZN(n5156) );
  CLKBUF_X1 U3525 ( .A(n4639), .Z(n5222) );
  XNOR2_X1 U3526 ( .A(n3807), .B(n3808), .ZN(n5223) );
  XNOR2_X1 U3527 ( .A(n3772), .B(n3773), .ZN(n4637) );
  NAND2_X1 U3528 ( .A1(n3736), .A2(n3735), .ZN(n5934) );
  NOR2_X1 U3529 ( .A1(n4603), .A2(n4585), .ZN(n4631) );
  AND2_X1 U3530 ( .A1(n4558), .A2(n4507), .ZN(n5165) );
  INV_X1 U3531 ( .A(n4003), .ZN(n5892) );
  AND2_X1 U3532 ( .A1(n4528), .A2(n3672), .ZN(n3673) );
  NAND2_X1 U3533 ( .A1(n3655), .A2(n4680), .ZN(n4488) );
  NOR2_X1 U3534 ( .A1(n3661), .A2(n7170), .ZN(n3678) );
  CLKBUF_X1 U3535 ( .A(n3657), .Z(n4662) );
  NAND2_X1 U3536 ( .A1(n3560), .A2(n3559), .ZN(n3657) );
  AND4_X2 U3537 ( .A1(n3540), .A2(n3539), .A3(n3538), .A4(n3537), .ZN(n3688)
         );
  AND4_X1 U3538 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3576)
         );
  AND4_X1 U3539 ( .A1(n3536), .A2(n3535), .A3(n3534), .A4(n3533), .ZN(n3537)
         );
  AND4_X1 U3540 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3602)
         );
  AND4_X1 U3541 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3600)
         );
  AND4_X1 U3542 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3539)
         );
  AND4_X1 U3543 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3603)
         );
  AND4_X1 U3544 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3560)
         );
  AND4_X1 U3545 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3538)
         );
  AND4_X1 U3546 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(n3575)
         );
  AND4_X1 U3547 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3620)
         );
  AND4_X1 U3548 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3540)
         );
  AND4_X1 U3549 ( .A1(n3573), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n3574)
         );
  AND2_X2 U3550 ( .A1(n3531), .A2(n3530), .ZN(n3719) );
  OR2_X2 U3551 ( .A1(n7183), .A2(n6456), .ZN(n6453) );
  AND2_X2 U3552 ( .A1(n3532), .A2(n5124), .ZN(n4096) );
  BUF_X2 U3553 ( .A(n3704), .Z(n5846) );
  AND2_X2 U3554 ( .A1(n3449), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5964)
         );
  AND2_X2 U3555 ( .A1(n5124), .A2(n4535), .ZN(n5829) );
  AND2_X1 U3556 ( .A1(n3519), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3524)
         );
  NAND2_X1 U3558 ( .A1(n3940), .A2(n3437), .ZN(n3430) );
  NAND2_X1 U3559 ( .A1(n3757), .A2(n3756), .ZN(n3431) );
  NAND2_X1 U3560 ( .A1(n3771), .A2(n3685), .ZN(n3432) );
  NAND2_X1 U3561 ( .A1(n3940), .A2(n3437), .ZN(n6257) );
  NAND2_X1 U3562 ( .A1(n3757), .A2(n3756), .ZN(n4605) );
  NAND2_X1 U3563 ( .A1(n3771), .A2(n3685), .ZN(n3772) );
  OAI21_X1 U3564 ( .B1(n4605), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4606), 
        .ZN(n3764) );
  NAND2_X1 U3565 ( .A1(n3804), .A2(n3803), .ZN(n6663) );
  NAND2_X2 U3566 ( .A1(n3508), .A2(n3829), .ZN(n3861) );
  NAND2_X2 U3567 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  OAI21_X2 U3568 ( .B1(n3938), .B2(n6388), .A(n6217), .ZN(n6243) );
  AND2_X1 U3569 ( .A1(n5124), .A2(n4535), .ZN(n3434) );
  OR2_X4 U3570 ( .A1(n3634), .A2(n3633), .ZN(n3671) );
  NAND2_X2 U3571 ( .A1(n6283), .A2(n3505), .ZN(n6225) );
  NAND2_X2 U3572 ( .A1(n6285), .A2(n6284), .ZN(n6283) );
  NAND4_X1 U3573 ( .A1(n3659), .A2(n3636), .A3(n4652), .A4(n4006), .ZN(n4551)
         );
  NAND2_X2 U3574 ( .A1(n3680), .A2(n3679), .ZN(n3771) );
  NAND2_X2 U3575 ( .A1(n5605), .A2(n3931), .ZN(n5641) );
  AND2_X4 U3576 ( .A1(n3531), .A2(n5964), .ZN(n3714) );
  NAND2_X2 U3577 ( .A1(n3857), .A2(n3856), .ZN(n3858) );
  OAI21_X2 U3578 ( .B1(n4797), .B2(n4796), .A(n3859), .ZN(n4801) );
  XNOR2_X2 U3579 ( .A(n3858), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4796)
         );
  NAND2_X1 U3580 ( .A1(n3508), .A2(n3507), .ZN(n3877) );
  AND2_X1 U3581 ( .A1(n3829), .A2(n3860), .ZN(n3507) );
  NAND2_X1 U3582 ( .A1(n3637), .A2(n4006), .ZN(n4463) );
  NAND2_X1 U3583 ( .A1(n4468), .A2(n4463), .ZN(n3502) );
  INV_X1 U3584 ( .A(n3877), .ZN(n3874) );
  AND2_X1 U3585 ( .A1(n3489), .A2(n3488), .ZN(n3487) );
  INV_X1 U3586 ( .A(n5995), .ZN(n3488) );
  AOI21_X1 U3587 ( .B1(n5223), .B2(n7159), .A(n3791), .ZN(n3794) );
  AND2_X1 U3588 ( .A1(n6020), .A2(n3487), .ZN(n5994) );
  INV_X1 U3589 ( .A(n4775), .ZN(n4485) );
  NOR2_X1 U3590 ( .A1(n4503), .A2(n3503), .ZN(n3501) );
  AND3_X2 U3591 ( .A1(n3674), .A2(n3673), .A3(n5892), .ZN(n4519) );
  AND2_X1 U3592 ( .A1(n4503), .A2(n4675), .ZN(n3674) );
  AND2_X1 U3593 ( .A1(n3667), .A2(n3666), .ZN(n3681) );
  OR2_X1 U3594 ( .A1(n3872), .A2(n3871), .ZN(n3882) );
  OR2_X1 U3595 ( .A1(n3710), .A2(n3709), .ZN(n3797) );
  AND2_X1 U3596 ( .A1(n4680), .A2(n4566), .ZN(n3456) );
  INV_X1 U3597 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3992) );
  OR2_X1 U3598 ( .A1(n6222), .A2(n3483), .ZN(n3482) );
  INV_X1 U3599 ( .A(n3484), .ZN(n3483) );
  INV_X1 U3600 ( .A(n4443), .ZN(n5869) );
  AND2_X1 U3601 ( .A1(n4196), .A2(n5621), .ZN(n3481) );
  INV_X1 U3602 ( .A(n5631), .ZN(n4196) );
  NAND2_X1 U3603 ( .A1(n3435), .A2(n4156), .ZN(n4165) );
  AND2_X1 U3604 ( .A1(n5433), .A2(n4157), .ZN(n4156) );
  AND2_X1 U3605 ( .A1(n4956), .A2(n4126), .ZN(n4127) );
  AND2_X1 U3606 ( .A1(n3905), .A2(n3878), .ZN(n4049) );
  INV_X1 U3607 ( .A(n3904), .ZN(n3902) );
  NOR2_X1 U3608 ( .A1(n3463), .A2(n3462), .ZN(n3461) );
  INV_X1 U3609 ( .A(n5767), .ZN(n3462) );
  INV_X1 U3610 ( .A(n5695), .ZN(n3463) );
  NAND2_X1 U3611 ( .A1(n5555), .A2(n5450), .ZN(n5580) );
  INV_X1 U3612 ( .A(n5616), .ZN(n5450) );
  AND2_X1 U3613 ( .A1(n6119), .A2(n3450), .ZN(n5555) );
  NOR2_X1 U3614 ( .A1(n3451), .A2(n5554), .ZN(n3450) );
  INV_X1 U3615 ( .A(n3452), .ZN(n3451) );
  NAND2_X1 U3616 ( .A1(n5805), .A2(n5816), .ZN(n5795) );
  AND2_X1 U3617 ( .A1(n5805), .A2(n4965), .ZN(n5796) );
  INV_X1 U3618 ( .A(n4675), .ZN(n3659) );
  NAND2_X1 U3619 ( .A1(n3778), .A2(n3777), .ZN(n3808) );
  OR2_X1 U3620 ( .A1(n3774), .A2(n3449), .ZN(n3778) );
  OAI21_X1 U3621 ( .B1(n5934), .B2(STATE2_REG_0__SCAN_IN), .A(n3760), .ZN(
        n3759) );
  NAND2_X1 U3622 ( .A1(n4636), .A2(n7159), .ZN(n3828) );
  AND2_X1 U3623 ( .A1(n5127), .A2(n5126), .ZN(n7127) );
  NAND2_X1 U3624 ( .A1(n3659), .A2(n3671), .ZN(n3752) );
  NOR2_X2 U3626 ( .A1(n6831), .A2(n5186), .ZN(n6979) );
  AND2_X1 U3627 ( .A1(n5182), .A2(n7176), .ZN(n4615) );
  AND2_X1 U3628 ( .A1(n3487), .A2(n5940), .ZN(n3486) );
  NOR2_X1 U3629 ( .A1(n4424), .A2(n6196), .ZN(n4425) );
  OR2_X1 U3630 ( .A1(n4399), .A2(n6039), .ZN(n4424) );
  NAND2_X1 U3631 ( .A1(n4376), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4397)
         );
  INV_X1 U3632 ( .A(n4375), .ZN(n4376) );
  NAND2_X1 U3633 ( .A1(n6078), .A2(n3477), .ZN(n3476) );
  INV_X1 U3634 ( .A(n3478), .ZN(n3477) );
  NAND2_X1 U3635 ( .A1(n4112), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4109)
         );
  INV_X1 U3636 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U3637 ( .A1(n6002), .A2(n5819), .ZN(n5950) );
  NAND2_X1 U3638 ( .A1(n6009), .A2(n6000), .ZN(n6002) );
  AND2_X1 U3639 ( .A1(n6006), .A2(n6007), .ZN(n6009) );
  AND2_X1 U3640 ( .A1(n5897), .A2(n5896), .ZN(n6182) );
  NAND2_X1 U3641 ( .A1(n6211), .A2(n3445), .ZN(n6183) );
  AOI21_X1 U3642 ( .B1(n3497), .B2(n3499), .A(n3496), .ZN(n3495) );
  OR2_X1 U3643 ( .A1(n4810), .A2(n6442), .ZN(n5653) );
  INV_X1 U3644 ( .A(n5796), .ZN(n5949) );
  NAND2_X1 U3645 ( .A1(n4487), .A2(n4486), .ZN(n4512) );
  INV_X1 U3646 ( .A(n4738), .ZN(n5148) );
  NAND2_X1 U3647 ( .A1(n5148), .A2(n5357), .ZN(n5475) );
  AND4_X1 U3648 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3621)
         );
  INV_X2 U3649 ( .A(n3688), .ZN(n4652) );
  AND4_X1 U3650 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  OR2_X1 U3651 ( .A1(n5222), .A2(n4012), .ZN(n4934) );
  AOI21_X1 U3652 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5927), .A(n4738), .ZN(
        n5266) );
  INV_X1 U3653 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7128) );
  INV_X1 U3654 ( .A(n7164), .ZN(n5993) );
  XNOR2_X1 U3655 ( .A(n5994), .B(n5880), .ZN(n6130) );
  NAND2_X1 U3656 ( .A1(n7108), .A2(n4450), .ZN(n6287) );
  CLKBUF_X1 U3657 ( .A(n3433), .Z(n4431) );
  BUF_X1 U3658 ( .A(n4363), .Z(n5857) );
  AND2_X1 U3659 ( .A1(n3901), .A2(n3900), .ZN(n3904) );
  NAND2_X1 U3660 ( .A1(n3764), .A2(n3763), .ZN(n3802) );
  NOR2_X1 U3661 ( .A1(n4491), .A2(n3752), .ZN(n4465) );
  AND2_X1 U3662 ( .A1(n3730), .A2(n3729), .ZN(n3766) );
  NAND2_X1 U3663 ( .A1(n3427), .A2(n4652), .ZN(n3779) );
  OR2_X1 U3664 ( .A1(n3779), .A2(n7159), .ZN(n3979) );
  INV_X1 U3665 ( .A(n3979), .ZN(n3986) );
  NAND2_X1 U3666 ( .A1(n3985), .A2(n4034), .ZN(n4474) );
  INV_X1 U3667 ( .A(n3991), .ZN(n3985) );
  INV_X1 U3668 ( .A(n4596), .ZN(n3472) );
  AND2_X1 U3669 ( .A1(n4423), .A2(n4449), .ZN(n3489) );
  INV_X1 U3670 ( .A(n6021), .ZN(n4423) );
  NOR2_X1 U3671 ( .A1(n6063), .A2(n6143), .ZN(n3484) );
  INV_X1 U3672 ( .A(n6060), .ZN(n3485) );
  NAND2_X1 U3673 ( .A1(n4243), .A2(n3479), .ZN(n3478) );
  INV_X1 U3674 ( .A(n6089), .ZN(n3479) );
  AND2_X1 U3675 ( .A1(n4127), .A2(n5433), .ZN(n3475) );
  AOI21_X1 U3676 ( .B1(n4863), .B2(n4191), .A(n5941), .ZN(n4597) );
  NOR2_X1 U3677 ( .A1(n4652), .A2(n7159), .ZN(n3923) );
  OR2_X1 U3678 ( .A1(n3726), .A2(n3725), .ZN(n3926) );
  NOR2_X1 U3679 ( .A1(n3441), .A2(n3506), .ZN(n3505) );
  INV_X1 U3680 ( .A(n3936), .ZN(n3506) );
  INV_X1 U3681 ( .A(n5904), .ZN(n3504) );
  INV_X1 U3682 ( .A(n5672), .ZN(n3496) );
  INV_X1 U3683 ( .A(n5795), .ZN(n5809) );
  NOR2_X1 U3684 ( .A1(n3454), .A2(n3453), .ZN(n3452) );
  INV_X1 U3685 ( .A(n4971), .ZN(n3453) );
  INV_X1 U3686 ( .A(n5461), .ZN(n3454) );
  NAND2_X1 U3687 ( .A1(n3885), .A2(n3884), .ZN(n3887) );
  NAND2_X1 U3688 ( .A1(n3457), .A2(n4563), .ZN(n4572) );
  NAND2_X1 U3689 ( .A1(n3456), .A2(n3677), .ZN(n3458) );
  AOI21_X1 U3690 ( .B1(n3670), .B2(n3671), .A(n4680), .ZN(n3693) );
  NAND2_X1 U3691 ( .A1(n3502), .A2(n3671), .ZN(n3691) );
  NOR2_X1 U3692 ( .A1(n3979), .A2(n4488), .ZN(n3999) );
  AND2_X1 U3693 ( .A1(n3779), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3996) );
  NAND2_X1 U3694 ( .A1(n3995), .A2(n3994), .ZN(n4473) );
  INV_X1 U3695 ( .A(n3794), .ZN(n3792) );
  OR2_X1 U3696 ( .A1(n4869), .A2(n4863), .ZN(n4975) );
  AND2_X1 U3697 ( .A1(n4739), .A2(n3776), .ZN(n4646) );
  OAI21_X1 U3698 ( .B1(n5183), .B2(n5925), .A(n7160), .ZN(n4647) );
  INV_X1 U3699 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7124) );
  INV_X1 U3700 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5706) );
  OR2_X1 U3701 ( .A1(n3774), .A2(n5969), .ZN(n3815) );
  NAND2_X1 U3702 ( .A1(n4017), .A2(n4016), .ZN(n4556) );
  NAND2_X1 U3703 ( .A1(n4556), .A2(n4555), .ZN(n4595) );
  OR2_X1 U3704 ( .A1(n6979), .A2(n6823), .ZN(n5195) );
  AND2_X1 U3705 ( .A1(n5693), .A2(n5692), .ZN(n5695) );
  AND2_X1 U3706 ( .A1(n5694), .A2(n5695), .ZN(n5768) );
  NAND2_X1 U3707 ( .A1(n4582), .A2(n4581), .ZN(n4603) );
  INV_X1 U3708 ( .A(n4600), .ZN(n4581) );
  INV_X1 U3709 ( .A(n4064), .ZN(n4065) );
  OAI21_X1 U3710 ( .B1(n4067), .B2(n4063), .A(n4062), .ZN(n4064) );
  AND2_X1 U3711 ( .A1(n4777), .A2(n5990), .ZN(n6672) );
  OR2_X1 U3712 ( .A1(n5162), .A2(n4776), .ZN(n4777) );
  OR2_X1 U3713 ( .A1(n5985), .A2(n7164), .ZN(n4775) );
  INV_X1 U3714 ( .A(n5169), .ZN(n5093) );
  AND2_X1 U3715 ( .A1(n6210), .A2(n3426), .ZN(n4377) );
  OR2_X1 U3716 ( .A1(n4354), .A2(n7090), .ZN(n4375) );
  NOR2_X1 U3717 ( .A1(n4308), .A2(n6244), .ZN(n4309) );
  AND2_X1 U3718 ( .A1(n4293), .A2(n4292), .ZN(n6152) );
  AND2_X1 U3719 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4275), .ZN(n4276)
         );
  NAND2_X1 U3720 ( .A1(n4276), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4308)
         );
  NOR2_X1 U3721 ( .A1(n4239), .A2(n6270), .ZN(n4240) );
  NAND2_X1 U3722 ( .A1(n4240), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4274)
         );
  OR2_X1 U3723 ( .A1(n4211), .A2(n5706), .ZN(n4239) );
  INV_X1 U3724 ( .A(n5681), .ZN(n3480) );
  NOR2_X1 U3725 ( .A1(n4179), .A2(n7042), .ZN(n4197) );
  NAND2_X1 U3726 ( .A1(n5622), .A2(n3481), .ZN(n5682) );
  NOR2_X1 U3727 ( .A1(n4159), .A2(n5547), .ZN(n4160) );
  NAND2_X1 U3728 ( .A1(n4160), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4179)
         );
  NAND2_X1 U3729 ( .A1(n4128), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4159)
         );
  NOR2_X1 U3730 ( .A1(n4109), .A2(n5562), .ZN(n4128) );
  AND2_X1 U3731 ( .A1(n4111), .A2(n4110), .ZN(n5552) );
  OR2_X1 U3732 ( .A1(n5458), .A2(n5459), .ZN(n5551) );
  NAND2_X1 U3733 ( .A1(n4060), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4081)
         );
  AOI21_X1 U3734 ( .B1(n4049), .B2(n4191), .A(n4048), .ZN(n4729) );
  AND2_X1 U3735 ( .A1(n5808), .A2(n5807), .ZN(n6031) );
  OR2_X1 U3736 ( .A1(n6350), .A2(n5804), .ZN(n6050) );
  NAND2_X1 U3737 ( .A1(n6157), .A2(n3468), .ZN(n6350) );
  NOR2_X1 U3738 ( .A1(n6145), .A2(n3469), .ZN(n3468) );
  INV_X1 U3739 ( .A(n6066), .ZN(n3469) );
  NAND2_X1 U3740 ( .A1(n6157), .A2(n6066), .ZN(n6146) );
  AND2_X1 U3741 ( .A1(n6155), .A2(n6154), .ZN(n6157) );
  NOR2_X1 U3742 ( .A1(n6096), .A2(n6082), .ZN(n6155) );
  NAND2_X1 U3743 ( .A1(n5694), .A2(n3459), .ZN(n6096) );
  NOR2_X1 U3744 ( .A1(n6093), .A2(n3460), .ZN(n3459) );
  INV_X1 U3745 ( .A(n3461), .ZN(n3460) );
  NAND2_X1 U3746 ( .A1(n5694), .A2(n3461), .ZN(n6094) );
  AND2_X1 U3747 ( .A1(n5688), .A2(n5687), .ZN(n5690) );
  OR2_X1 U3748 ( .A1(n5636), .A2(n5637), .ZN(n5689) );
  AOI21_X1 U3749 ( .B1(n3442), .B2(n3932), .A(n3498), .ZN(n3497) );
  INV_X1 U3750 ( .A(n5717), .ZN(n3498) );
  INV_X1 U3751 ( .A(n5640), .ZN(n3500) );
  INV_X1 U3752 ( .A(n3932), .ZN(n3499) );
  NOR2_X1 U3753 ( .A1(n5580), .A2(n5579), .ZN(n5629) );
  AND2_X1 U3754 ( .A1(n6248), .A2(n5669), .ZN(n5715) );
  NAND2_X1 U3755 ( .A1(n5641), .A2(n5640), .ZN(n5649) );
  OR2_X1 U3756 ( .A1(n6887), .A2(n5659), .ZN(n5663) );
  NAND2_X1 U3757 ( .A1(n6119), .A2(n3452), .ZN(n5553) );
  NOR2_X1 U3758 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  AND2_X1 U3759 ( .A1(n6119), .A2(n4971), .ZN(n5462) );
  NAND2_X1 U3760 ( .A1(n3910), .A2(n6792), .ZN(n6799) );
  AND2_X1 U3761 ( .A1(n4961), .A2(n4960), .ZN(n5218) );
  NAND2_X1 U3762 ( .A1(n6441), .A2(n7159), .ZN(n4454) );
  NAND2_X1 U3763 ( .A1(n4733), .A2(n4732), .ZN(n5217) );
  INV_X1 U3764 ( .A(n4736), .ZN(n4732) );
  AND2_X1 U3765 ( .A1(n4806), .A2(n5655), .ZN(n6417) );
  XNOR2_X1 U3766 ( .A(n3887), .B(n3886), .ZN(n4802) );
  CLKBUF_X1 U3767 ( .A(n4637), .Z(n4638) );
  OAI211_X1 U3768 ( .C1(n4534), .C2(n4533), .A(n4532), .B(n4531), .ZN(n7119)
         );
  INV_X1 U3769 ( .A(n4834), .ZN(n4828) );
  OR3_X1 U3770 ( .A1(n5222), .A2(n3829), .A3(n5150), .ZN(n5227) );
  NOR2_X1 U3771 ( .A1(n4012), .A2(n4018), .ZN(n5279) );
  AND2_X1 U3772 ( .A1(n4012), .A2(n5931), .ZN(n4981) );
  INV_X1 U3773 ( .A(n4975), .ZN(n4982) );
  AND3_X1 U3774 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7159), .A3(n4647), .ZN(
        n4681) );
  NAND2_X1 U3775 ( .A1(n7159), .A2(n4647), .ZN(n4738) );
  INV_X1 U3776 ( .A(n4644), .ZN(n4740) );
  AND2_X1 U3777 ( .A1(n4005), .A2(n4004), .ZN(n7136) );
  AND2_X1 U3778 ( .A1(n6443), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4002) );
  INV_X1 U3779 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5547) );
  INV_X1 U3780 ( .A(n7097), .ZN(n7071) );
  OR2_X1 U3781 ( .A1(n6979), .A2(n5978), .ZN(n7051) );
  OR2_X1 U3782 ( .A1(n6979), .A2(n5471), .ZN(n7097) );
  INV_X1 U3783 ( .A(n7083), .ZN(n7104) );
  OR2_X1 U3784 ( .A1(n6979), .A2(n5204), .ZN(n7061) );
  OR2_X1 U3785 ( .A1(n6009), .A2(n6008), .ZN(n6136) );
  AND2_X1 U3786 ( .A1(n6785), .A2(n4006), .ZN(n6783) );
  INV_X1 U3787 ( .A(n6776), .ZN(n6782) );
  INV_X1 U3788 ( .A(n6785), .ZN(n6159) );
  AND2_X1 U3789 ( .A1(n4561), .A2(n5993), .ZN(n6785) );
  NAND2_X1 U3790 ( .A1(n6785), .A2(n5974), .ZN(n6776) );
  INV_X1 U3791 ( .A(n6173), .ZN(n7209) );
  INV_X1 U3792 ( .A(n5973), .ZN(n7208) );
  AND2_X1 U3793 ( .A1(n5973), .A2(n5170), .ZN(n7206) );
  OAI21_X1 U3794 ( .B1(n5167), .B2(n5166), .A(n5993), .ZN(n5168) );
  INV_X1 U3795 ( .A(n7206), .ZN(n6180) );
  XNOR2_X1 U3796 ( .A(n5187), .B(n5956), .ZN(n5946) );
  OR2_X1 U3797 ( .A1(n5875), .A2(n5921), .ZN(n5187) );
  XNOR2_X1 U3798 ( .A(n5944), .B(n5943), .ZN(n5975) );
  NAND2_X1 U3799 ( .A1(n6020), .A2(n3486), .ZN(n5944) );
  AND2_X1 U3800 ( .A1(n5824), .A2(n4427), .ZN(n6013) );
  XNOR2_X1 U3801 ( .A(n3948), .B(n3947), .ZN(n6311) );
  NAND2_X1 U3802 ( .A1(n6183), .A2(n5897), .ZN(n3948) );
  INV_X1 U3803 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6244) );
  INV_X1 U3804 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6270) );
  INV_X1 U3805 ( .A(n7108), .ZN(n6810) );
  XNOR2_X1 U3806 ( .A(n5952), .B(n3467), .ZN(n6292) );
  INV_X1 U3807 ( .A(n5953), .ZN(n3467) );
  OAI21_X1 U3808 ( .B1(n6002), .B2(n5951), .A(n5950), .ZN(n5952) );
  AOI22_X1 U3809 ( .A1(n6183), .A2(n6182), .B1(n6277), .B2(n6316), .ZN(n6185)
         );
  INV_X1 U3810 ( .A(n6136), .ZN(n6313) );
  OR2_X1 U3811 ( .A1(n6363), .A2(n5911), .ZN(n6351) );
  OR2_X1 U3812 ( .A1(n4454), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6912) );
  AND2_X1 U3813 ( .A1(n4512), .A2(n4501), .ZN(n6932) );
  INV_X1 U3814 ( .A(n6932), .ZN(n6915) );
  INV_X1 U3815 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5927) );
  INV_X1 U3816 ( .A(n4018), .ZN(n5931) );
  INV_X1 U3817 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5224) );
  INV_X1 U3818 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6443) );
  INV_X1 U3819 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U3820 ( .A1(n5471), .A2(n5985), .ZN(n5965) );
  NOR2_X2 U3821 ( .A1(n5156), .A2(n5046), .ZN(n5342) );
  INV_X1 U3822 ( .A(n5467), .ZN(n5537) );
  NOR2_X2 U3823 ( .A1(n4834), .A2(n4018), .ZN(n4919) );
  INV_X1 U3824 ( .A(n5272), .ZN(n5327) );
  OAI21_X1 U3825 ( .B1(n5426), .B2(n5471), .A(n5402), .ZN(n5425) );
  INV_X1 U3826 ( .A(n5389), .ZN(n5427) );
  CLKBUF_X1 U3827 ( .A(n4640), .Z(n4951) );
  INV_X1 U3828 ( .A(n5278), .ZN(n5496) );
  INV_X1 U3829 ( .A(n5319), .ZN(n5489) );
  INV_X1 U3830 ( .A(n5325), .ZN(n5533) );
  INV_X1 U3831 ( .A(n5332), .ZN(n5482) );
  INV_X1 U3832 ( .A(n5304), .ZN(n5524) );
  INV_X1 U3833 ( .A(n5316), .ZN(n5517) );
  INV_X1 U3834 ( .A(n5322), .ZN(n5510) );
  INV_X1 U3835 ( .A(n5301), .ZN(n5503) );
  INV_X1 U3836 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7159) );
  INV_X1 U3837 ( .A(READY_N), .ZN(n7176) );
  AOI21_X1 U3838 ( .B1(n6130), .B2(n4644), .A(n5922), .ZN(n5923) );
  OAI21_X1 U3839 ( .B1(n6302), .B2(n6892), .A(n3464), .ZN(U2987) );
  INV_X1 U3840 ( .A(n3465), .ZN(n3464) );
  OAI21_X1 U3841 ( .B1(n6292), .B2(n6915), .A(n3466), .ZN(n3465) );
  NOR3_X1 U3842 ( .A1(n6301), .A2(n6300), .A3(n6299), .ZN(n3466) );
  AND3_X1 U3843 ( .A1(n5178), .A2(n5179), .A3(n4127), .ZN(n3435) );
  NAND2_X1 U3844 ( .A1(n3485), .A2(n3484), .ZN(n3436) );
  NAND2_X1 U3845 ( .A1(n6283), .A2(n3443), .ZN(n3437) );
  NAND2_X1 U3846 ( .A1(n6020), .A2(n3489), .ZN(n5842) );
  OR2_X1 U3847 ( .A1(n5697), .A2(n5760), .ZN(n5759) );
  AND2_X1 U3848 ( .A1(n3446), .A2(n3945), .ZN(n3438) );
  INV_X1 U3849 ( .A(n4502), .ZN(n5805) );
  MUX2_X2 U3850 ( .A(n3760), .B(n3759), .S(n3758), .Z(n4018) );
  NOR2_X1 U3851 ( .A1(n5697), .A2(n3478), .ZN(n3439) );
  AND2_X2 U3852 ( .A1(n3529), .A2(n3524), .ZN(n3639) );
  NAND2_X1 U3853 ( .A1(n6211), .A2(n3945), .ZN(n6201) );
  NAND2_X1 U3854 ( .A1(n6283), .A2(n3936), .ZN(n6276) );
  NOR2_X1 U3855 ( .A1(n5697), .A2(n3476), .ZN(n6077) );
  AND2_X1 U3856 ( .A1(n6020), .A2(n4423), .ZN(n4448) );
  AND4_X1 U3857 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3440)
         );
  NAND2_X1 U3858 ( .A1(n3636), .A2(n3655), .ZN(n3670) );
  INV_X1 U3859 ( .A(n3671), .ZN(n4503) );
  AND2_X1 U3860 ( .A1(n6248), .A2(n5684), .ZN(n3441) );
  OR2_X1 U3861 ( .A1(n3500), .A2(n5715), .ZN(n3442) );
  NAND2_X1 U3862 ( .A1(n3485), .A2(n4313), .ZN(n6061) );
  AND2_X1 U3863 ( .A1(n6030), .A2(n6018), .ZN(n6006) );
  AOI21_X1 U3864 ( .B1(n3759), .B2(n3758), .A(n3751), .ZN(n3765) );
  AND2_X1 U3865 ( .A1(n3505), .A2(n3504), .ZN(n3443) );
  INV_X1 U3866 ( .A(n6277), .ZN(n3938) );
  INV_X1 U3867 ( .A(n3829), .ZN(n4933) );
  AND2_X1 U3868 ( .A1(n5178), .A2(n5179), .ZN(n4955) );
  NOR2_X1 U3869 ( .A1(n4623), .A2(n4058), .ZN(n5178) );
  NAND2_X1 U3870 ( .A1(n5622), .A2(n5621), .ZN(n5620) );
  OAI21_X1 U3871 ( .B1(n5641), .B2(n3499), .A(n3497), .ZN(n5671) );
  INV_X1 U3872 ( .A(n4006), .ZN(n5974) );
  NOR2_X1 U3873 ( .A1(n5689), .A2(n5690), .ZN(n5694) );
  INV_X1 U3874 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U3875 ( .A1(n6248), .A2(n6324), .ZN(n3444) );
  INV_X1 U3876 ( .A(n6063), .ZN(n4313) );
  AND2_X1 U3877 ( .A1(n3438), .A2(n3444), .ZN(n3445) );
  AND2_X1 U3878 ( .A1(n4278), .A2(n4277), .ZN(n6078) );
  NAND2_X1 U3879 ( .A1(n6248), .A2(n6337), .ZN(n3446) );
  AND2_X1 U3880 ( .A1(n3481), .A2(n3480), .ZN(n3447) );
  INV_X1 U3881 ( .A(n3455), .ZN(n5816) );
  NAND2_X1 U3882 ( .A1(n3677), .A2(n4680), .ZN(n3455) );
  NOR2_X1 U3883 ( .A1(n4636), .A2(n5934), .ZN(n3448) );
  AND2_X1 U3884 ( .A1(n4599), .A2(n4570), .ZN(n4569) );
  INV_X1 U3885 ( .A(n5895), .ZN(n6193) );
  INV_X2 U3886 ( .A(n6193), .ZN(n6248) );
  INV_X2 U3887 ( .A(n6193), .ZN(n6277) );
  INV_X1 U3888 ( .A(n5760), .ZN(n4243) );
  NAND2_X1 U3889 ( .A1(n4562), .A2(n3458), .ZN(n3457) );
  NAND2_X1 U3890 ( .A1(n4597), .A2(n3470), .ZN(n3471) );
  NAND3_X1 U3891 ( .A1(n4556), .A2(n3472), .A3(n4555), .ZN(n3470) );
  NAND2_X1 U3892 ( .A1(n4165), .A2(n3473), .ZN(n5572) );
  NAND2_X1 U3893 ( .A1(n3474), .A2(n4158), .ZN(n3473) );
  NAND3_X1 U3894 ( .A1(n5178), .A2(n3475), .A3(n5179), .ZN(n3474) );
  NAND2_X1 U3895 ( .A1(n3490), .A2(n3765), .ZN(n3770) );
  XNOR2_X1 U3896 ( .A(n3490), .B(n3765), .ZN(n4011) );
  NAND3_X1 U3897 ( .A1(n3493), .A2(n3491), .A3(n5585), .ZN(n5584) );
  NAND2_X1 U3898 ( .A1(n3492), .A2(n3921), .ZN(n3491) );
  INV_X1 U3899 ( .A(n6798), .ZN(n3492) );
  NAND3_X1 U3900 ( .A1(n3921), .A2(n3910), .A3(n6792), .ZN(n3493) );
  NAND2_X1 U3901 ( .A1(n6797), .A2(n3921), .ZN(n5586) );
  NAND2_X1 U3902 ( .A1(n6799), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U3903 ( .A1(n5641), .A2(n3497), .ZN(n3494) );
  NAND2_X1 U3904 ( .A1(n3494), .A2(n3495), .ZN(n3934) );
  INV_X1 U3905 ( .A(n3676), .ZN(n3503) );
  NAND2_X1 U3906 ( .A1(n6211), .A2(n3438), .ZN(n6191) );
  NAND2_X1 U3907 ( .A1(n6311), .A2(n6810), .ZN(n4460) );
  INV_X1 U3908 ( .A(n6020), .ZN(n6035) );
  INV_X1 U3909 ( .A(n3802), .ZN(n3804) );
  INV_X1 U3910 ( .A(n3959), .ZN(n3672) );
  NAND2_X1 U3911 ( .A1(n3959), .A2(n3561), .ZN(n3669) );
  NAND2_X1 U3912 ( .A1(n5171), .A2(n5973), .ZN(n5639) );
  NAND2_X1 U3913 ( .A1(n3830), .A2(n3796), .ZN(n4639) );
  AND2_X1 U3914 ( .A1(n5649), .A2(n5648), .ZN(n5716) );
  NOR2_X2 U3915 ( .A1(n6243), .A2(n6242), .ZN(n6241) );
  AOI21_X2 U3916 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n3938), .A(n6241), 
        .ZN(n6235) );
  OAI21_X1 U3917 ( .B1(n3430), .B2(n3944), .A(n3943), .ZN(n6213) );
  AOI22_X1 U3918 ( .A1(n3703), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5829), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3553) );
  NAND2_X4 U3919 ( .A1(n3550), .A2(n3549), .ZN(n3655) );
  INV_X1 U3920 ( .A(n3703), .ZN(n3583) );
  OR2_X1 U3921 ( .A1(n3510), .A2(n5899), .ZN(n3509) );
  INV_X1 U3922 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4034) );
  AND2_X1 U3923 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3510) );
  INV_X1 U3924 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5899) );
  NOR2_X1 U3925 ( .A1(n3683), .A2(n7159), .ZN(n3511) );
  INV_X1 U3926 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n7042) );
  INV_X1 U3927 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3803) );
  INV_X1 U3928 ( .A(n4067), .ZN(n5874) );
  NAND2_X1 U3929 ( .A1(n3636), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4030) );
  INV_X1 U3930 ( .A(n4030), .ZN(n4191) );
  INV_X1 U3931 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5471) );
  OR2_X1 U3932 ( .A1(n5390), .A2(n6824), .ZN(n6291) );
  INV_X1 U3933 ( .A(n6291), .ZN(n4644) );
  OR2_X1 U3934 ( .A1(n5614), .A2(n5552), .ZN(n3512) );
  INV_X1 U3935 ( .A(n4181), .ZN(n5941) );
  OR2_X1 U3936 ( .A1(n3899), .A2(n3898), .ZN(n3915) );
  OR2_X1 U3937 ( .A1(n3789), .A2(n3788), .ZN(n3832) );
  INV_X1 U3938 ( .A(n3960), .ZN(n3962) );
  NAND2_X1 U3939 ( .A1(n3952), .A2(n3951), .ZN(n3982) );
  NOR2_X1 U3940 ( .A1(n4006), .A2(n6823), .ZN(n4041) );
  OR2_X1 U3941 ( .A1(n3851), .A2(n3850), .ZN(n3879) );
  OR2_X1 U3942 ( .A1(n3826), .A2(n3825), .ZN(n3853) );
  OR2_X1 U3943 ( .A1(n3993), .A2(n3992), .ZN(n3991) );
  OR2_X1 U3944 ( .A1(n5824), .A2(n5996), .ZN(n5875) );
  INV_X1 U3945 ( .A(n4274), .ZN(n4275) );
  NAND2_X1 U3946 ( .A1(n6436), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4443) );
  INV_X1 U3947 ( .A(n4041), .ZN(n4067) );
  NOR2_X1 U3948 ( .A1(n4081), .A2(n5588), .ZN(n4112) );
  XNOR2_X1 U3949 ( .A(n3861), .B(n3860), .ZN(n4031) );
  OR2_X1 U3950 ( .A1(n3746), .A2(n3745), .ZN(n3798) );
  AND3_X1 U3951 ( .A1(n3923), .A2(n3922), .A3(n3926), .ZN(n3924) );
  AND2_X1 U3952 ( .A1(n5447), .A2(n5446), .ZN(n5554) );
  INV_X1 U3953 ( .A(n4002), .ZN(n3812) );
  NAND2_X1 U3954 ( .A1(n3866), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U3955 ( .A1(n3820), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3704), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U3956 ( .A1(n4576), .A2(n4575), .ZN(n4601) );
  NAND2_X1 U3957 ( .A1(n4662), .A2(n4006), .ZN(n4003) );
  NAND2_X1 U3958 ( .A1(n4425), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5824)
         );
  INV_X1 U3959 ( .A(n3426), .ZN(n5872) );
  AND2_X1 U3960 ( .A1(n4490), .A2(n4489), .ZN(n4540) );
  NAND2_X1 U3961 ( .A1(n3815), .A2(n3814), .ZN(n5141) );
  OR2_X1 U3962 ( .A1(n4508), .A2(n5190), .ZN(n4541) );
  OR4_X1 U3963 ( .A1(n6736), .A2(n6738), .A3(n5882), .A4(n6065), .ZN(n7096) );
  NAND2_X1 U3964 ( .A1(n4197), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4211)
         );
  NAND2_X1 U3965 ( .A1(n5954), .A2(n5192), .ZN(n7041) );
  AND2_X1 U3966 ( .A1(n5786), .A2(n5785), .ZN(n6154) );
  INV_X1 U3967 ( .A(n5555), .ZN(n5617) );
  INV_X1 U3968 ( .A(n5940), .ZN(n5880) );
  OR2_X1 U3969 ( .A1(n4402), .A2(n4401), .ZN(n6037) );
  NAND2_X1 U3970 ( .A1(n4309), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4354)
         );
  NAND2_X1 U3971 ( .A1(n3939), .A2(n3938), .ZN(n3940) );
  AND2_X1 U3972 ( .A1(n4195), .A2(n4194), .ZN(n5631) );
  INV_X1 U3973 ( .A(n5571), .ZN(n4163) );
  INV_X1 U3974 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5588) );
  NOR2_X1 U3975 ( .A1(n4044), .A2(n4043), .ZN(n4050) );
  OR2_X1 U3976 ( .A1(n5936), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U3977 ( .A1(n3934), .A2(n3933), .ZN(n5747) );
  NAND2_X1 U3978 ( .A1(n4512), .A2(n4540), .ZN(n6933) );
  INV_X1 U3979 ( .A(n7115), .ZN(n6438) );
  OR2_X1 U3980 ( .A1(n4934), .A2(n3829), .ZN(n4834) );
  INV_X1 U3981 ( .A(n5383), .ZN(n5013) );
  INV_X2 U3982 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6823) );
  NOR2_X1 U3983 ( .A1(n4775), .A2(n4518), .ZN(n5182) );
  INV_X1 U3984 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6451) );
  INV_X1 U3985 ( .A(n5195), .ZN(n5954) );
  AND2_X1 U3986 ( .A1(n7041), .A2(n6957), .ZN(n6980) );
  INV_X1 U3987 ( .A(n7051), .ZN(n7057) );
  INV_X1 U3988 ( .A(n7073), .ZN(n7105) );
  NAND3_X1 U3989 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A3(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4044) );
  NOR2_X2 U3990 ( .A1(n5195), .A2(n5194), .ZN(n7079) );
  NOR2_X1 U3991 ( .A1(n4615), .A2(n5162), .ZN(n5082) );
  NOR2_X1 U3992 ( .A1(n4775), .A2(n7143), .ZN(n5105) );
  NAND2_X1 U3993 ( .A1(n6823), .A2(n5471), .ZN(n5390) );
  INV_X1 U3994 ( .A(n6815), .ZN(n6805) );
  AND2_X1 U3995 ( .A1(n4050), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4060)
         );
  INV_X1 U3996 ( .A(n6287), .ZN(n6809) );
  AND2_X1 U3997 ( .A1(n6929), .A2(n5906), .ZN(n6835) );
  OAI21_X1 U3998 ( .B1(n6933), .B2(n5658), .A(n6934), .ZN(n6929) );
  AND2_X1 U3999 ( .A1(n6890), .A2(n5661), .ZN(n5662) );
  INV_X1 U4000 ( .A(n6892), .ZN(n6938) );
  OAI21_X1 U4001 ( .B1(n6877), .B2(n6871), .A(n6933), .ZN(n6909) );
  AND2_X1 U4002 ( .A1(n5653), .A2(n5655), .ZN(n6877) );
  NOR2_X1 U4003 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6441) );
  INV_X1 U4004 ( .A(n5289), .ZN(n5341) );
  AND2_X1 U4005 ( .A1(n5280), .A2(n5025), .ZN(n5535) );
  AND2_X1 U4006 ( .A1(n4869), .A2(n5222), .ZN(n5280) );
  NOR2_X2 U4007 ( .A1(n5227), .A2(n5931), .ZN(n5328) );
  NOR2_X2 U4008 ( .A1(n5227), .A2(n4018), .ZN(n5329) );
  INV_X1 U4009 ( .A(n5403), .ZN(n5428) );
  AND2_X1 U4010 ( .A1(n4982), .A2(n4981), .ZN(n5383) );
  INV_X1 U4011 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6820) );
  INV_X1 U4012 ( .A(n6749), .ZN(n6751) );
  OR2_X1 U4013 ( .A1(n5182), .A2(n5181), .ZN(n6831) );
  NAND2_X1 U4014 ( .A1(n5954), .A2(n5199), .ZN(n7083) );
  OR2_X1 U4015 ( .A1(n6979), .A2(n5189), .ZN(n7073) );
  INV_X1 U4016 ( .A(n7079), .ZN(n7094) );
  INV_X2 U4017 ( .A(n6783), .ZN(n6777) );
  NAND2_X1 U4018 ( .A1(n5973), .A2(n5891), .ZN(n6173) );
  NAND2_X1 U4019 ( .A1(n5169), .A2(n5168), .ZN(n5973) );
  INV_X1 U4020 ( .A(n6672), .ZN(n6701) );
  NAND2_X1 U4021 ( .A1(n4615), .A2(n4680), .ZN(n5169) );
  NAND2_X1 U4022 ( .A1(n6287), .A2(n4453), .ZN(n6815) );
  AND2_X1 U4023 ( .A1(n6415), .A2(n5907), .ZN(n6842) );
  NAND2_X1 U4024 ( .A1(n4512), .A2(n4511), .ZN(n6892) );
  NOR2_X1 U4025 ( .A1(n5149), .A2(n5148), .ZN(n6454) );
  INV_X1 U4026 ( .A(n5965), .ZN(n7160) );
  NAND2_X1 U4027 ( .A1(n5280), .A2(n5279), .ZN(n5467) );
  NAND2_X1 U4028 ( .A1(n5280), .A2(n4981), .ZN(n5045) );
  AND2_X1 U4029 ( .A1(n4693), .A2(n4692), .ZN(n4728) );
  NAND2_X1 U4030 ( .A1(n4828), .A2(n4018), .ZN(n4861) );
  INV_X1 U4031 ( .A(n4895), .ZN(n4924) );
  NAND2_X1 U4032 ( .A1(n4982), .A2(n5279), .ZN(n5403) );
  AOI21_X1 U4033 ( .B1(n4978), .B2(n4979), .A(n4977), .ZN(n5018) );
  AND2_X1 U4034 ( .A1(n5355), .A2(n5354), .ZN(n5388) );
  AND2_X1 U4035 ( .A1(n4643), .A2(n4642), .ZN(n4686) );
  AND2_X1 U4036 ( .A1(n5266), .A2(n4743), .ZN(n4774) );
  NAND2_X1 U4037 ( .A1(n4002), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7164) );
  NOR2_X1 U4038 ( .A1(n6820), .A2(STATE_REG_0__SCAN_IN), .ZN(n7183) );
  INV_X1 U4039 ( .A(n6747), .ZN(n6753) );
  NOR2_X4 U4040 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3529) );
  AND2_X4 U4041 ( .A1(n3529), .A2(n3530), .ZN(n4407) );
  NAND2_X1 U4042 ( .A1(n4407), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3517) );
  AND2_X2 U4043 ( .A1(n3513), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3531)
         );
  NAND2_X1 U4044 ( .A1(n3714), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3516)
         );
  AND2_X2 U4045 ( .A1(n3529), .A2(n5124), .ZN(n3704) );
  NAND2_X1 U4046 ( .A1(n3704), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3515)
         );
  AND2_X2 U4047 ( .A1(n3530), .A2(n4535), .ZN(n3866) );
  INV_X1 U4048 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3518) );
  AND2_X2 U4049 ( .A1(n3518), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3532)
         );
  AND2_X2 U4050 ( .A1(n3532), .A2(n3530), .ZN(n4144) );
  NAND2_X1 U4051 ( .A1(n4144), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3523) );
  INV_X1 U4052 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3519) );
  AND2_X2 U4053 ( .A1(n3531), .A2(n3524), .ZN(n3703) );
  NAND2_X1 U4054 ( .A1(n3703), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3522) );
  AND2_X2 U4055 ( .A1(n3524), .A2(n4535), .ZN(n3720) );
  NAND2_X1 U4056 ( .A1(n3720), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3521) );
  NAND2_X1 U4057 ( .A1(n5829), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3520)
         );
  NAND2_X1 U4058 ( .A1(n3702), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3528)
         );
  AND2_X4 U4059 ( .A1(n3532), .A2(n5964), .ZN(n3713) );
  NAND2_X1 U4060 ( .A1(n3713), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3527) );
  AND2_X2 U4061 ( .A1(n3532), .A2(n3524), .ZN(n3640) );
  NAND2_X1 U4062 ( .A1(n3640), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4063 ( .A1(n3639), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3525) );
  AND2_X4 U4064 ( .A1(n4535), .A2(n5964), .ZN(n3820) );
  NAND2_X1 U4065 ( .A1(n3820), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3536)
         );
  AND2_X2 U4066 ( .A1(n5964), .A2(n3529), .ZN(n3645) );
  NAND2_X1 U4067 ( .A1(n3645), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4068 ( .A1(n3719), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U4069 ( .A1(n4096), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3533)
         );
  AOI22_X1 U4070 ( .A1(n3719), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3645), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4071 ( .A1(n4144), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3640), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4072 ( .A1(n3703), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4073 ( .A1(n3820), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3541) );
  AND4_X2 U4074 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3550)
         );
  AOI22_X1 U4075 ( .A1(n3702), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4076 ( .A1(n3714), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4077 ( .A1(n4096), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3704), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4078 ( .A1(n3713), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3720), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3545) );
  AND4_X2 U4079 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3549)
         );
  NAND2_X2 U4080 ( .A1(n3688), .A2(n3655), .ZN(n3959) );
  AOI22_X1 U4081 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n4407), .B1(n3866), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4082 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n3719), .B1(n3640), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4083 ( .A1(n4144), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3720), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4084 ( .A1(n3639), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        INSTQUEUE_REG_13__6__SCAN_IN), .B2(n4096), .ZN(n3557) );
  AOI22_X1 U4085 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n3714), .B1(n3645), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4086 ( .A1(n3713), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3702), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3555) );
  INV_X1 U4087 ( .A(n3657), .ZN(n3636) );
  NAND2_X1 U4088 ( .A1(n3636), .A2(n3688), .ZN(n3561) );
  NAND2_X1 U4089 ( .A1(n3645), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3565) );
  NAND2_X1 U4090 ( .A1(n3719), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3564) );
  NAND2_X1 U4091 ( .A1(n3714), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3563)
         );
  NAND2_X1 U4092 ( .A1(n3820), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3562)
         );
  NAND2_X1 U4093 ( .A1(n4144), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U4094 ( .A1(n3703), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3568) );
  NAND2_X1 U4095 ( .A1(n3640), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4096 ( .A1(n3639), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3566) );
  NAND2_X1 U4097 ( .A1(n3713), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3573) );
  NAND2_X1 U4098 ( .A1(n3702), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3572)
         );
  NAND2_X1 U4099 ( .A1(n3720), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4100 ( .A1(n5829), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3570)
         );
  NAND2_X1 U4101 ( .A1(n4096), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3580)
         );
  NAND2_X1 U4102 ( .A1(n3704), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3579)
         );
  NAND2_X1 U4103 ( .A1(n4407), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4104 ( .A1(n3866), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4105 ( .A1(n3669), .A2(n4006), .ZN(n3624) );
  NAND2_X1 U4106 ( .A1(n3703), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U4107 ( .A1(n4144), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3586) );
  NAND2_X1 U4108 ( .A1(n3713), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3585) );
  NAND2_X1 U4109 ( .A1(n3702), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3584)
         );
  NAND2_X1 U4110 ( .A1(n4096), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3591)
         );
  NAND2_X1 U4111 ( .A1(n3640), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4112 ( .A1(n3719), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4113 ( .A1(n3704), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3588)
         );
  NAND2_X1 U4114 ( .A1(n4363), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3595) );
  NAND2_X1 U4115 ( .A1(n3720), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4116 ( .A1(n3639), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U4117 ( .A1(n3434), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3592)
         );
  AND4_X2 U4118 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3601)
         );
  NAND2_X1 U4119 ( .A1(n3714), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3599)
         );
  NAND2_X1 U4120 ( .A1(n3820), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3598)
         );
  NAND2_X1 U4121 ( .A1(n4407), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3597) );
  NAND2_X1 U4122 ( .A1(n3866), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4123 ( .A1(n3719), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4124 ( .A1(n4096), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3606)
         );
  NAND2_X1 U4125 ( .A1(n3820), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3605)
         );
  NAND2_X1 U4126 ( .A1(n4363), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3604) );
  AND4_X2 U4127 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3623)
         );
  NAND2_X1 U4128 ( .A1(n3713), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4129 ( .A1(n3639), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3609) );
  NAND2_X1 U4130 ( .A1(n3702), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3608)
         );
  NAND3_X1 U4131 ( .A1(n3610), .A2(n3609), .A3(n3608), .ZN(n3611) );
  AOI21_X2 U4132 ( .B1(n3433), .B2(INSTQUEUE_REG_5__0__SCAN_IN), .A(n3611), 
        .ZN(n3622) );
  NAND2_X1 U4133 ( .A1(n4144), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4134 ( .A1(n3703), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U4135 ( .A1(n3720), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3613) );
  NAND2_X1 U4136 ( .A1(n5829), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3612)
         );
  NAND2_X1 U4137 ( .A1(n3714), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3619)
         );
  NAND2_X1 U4138 ( .A1(n4407), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3618) );
  NAND2_X1 U4139 ( .A1(n3704), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3617)
         );
  NAND2_X1 U4140 ( .A1(n3866), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3616) );
  NAND4_X4 U4141 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3677)
         );
  NAND2_X1 U4142 ( .A1(n3624), .A2(n3836), .ZN(n3635) );
  AOI22_X1 U4143 ( .A1(n4144), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3703), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4144 ( .A1(n3713), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4145 ( .A1(n3719), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3704), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4146 ( .A1(n3714), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4147 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3634)
         );
  AOI22_X1 U4148 ( .A1(n3702), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3640), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4149 ( .A1(n4363), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4150 ( .A1(n3720), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5829), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4151 ( .A1(n3820), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3629) );
  NAND4_X1 U4152 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3633)
         );
  AND2_X2 U4153 ( .A1(n3671), .A2(n3661), .ZN(n4502) );
  NAND2_X1 U4154 ( .A1(n3672), .A2(n4502), .ZN(n4536) );
  AND2_X2 U4155 ( .A1(n3635), .A2(n4536), .ZN(n3697) );
  INV_X1 U4156 ( .A(n3670), .ZN(n3637) );
  NAND2_X1 U4157 ( .A1(n3637), .A2(n3688), .ZN(n3638) );
  NAND2_X1 U4158 ( .A1(n3638), .A2(n4006), .ZN(n4491) );
  AOI22_X1 U4159 ( .A1(n4144), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3703), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4160 ( .A1(n3713), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3702), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4161 ( .A1(n3640), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4162 ( .A1(n3720), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5829), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4163 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3651)
         );
  AOI22_X1 U4164 ( .A1(n3719), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4165 ( .A1(n3820), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3645), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4166 ( .A1(n4407), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3704), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4167 ( .A1(n3714), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3646) );
  NAND4_X1 U4168 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3650)
         );
  OR2_X2 U4169 ( .A1(n3651), .A2(n3650), .ZN(n4675) );
  AND2_X1 U4170 ( .A1(n3670), .A2(n3427), .ZN(n4466) );
  INV_X1 U4171 ( .A(n3655), .ZN(n3653) );
  XNOR2_X1 U4172 ( .A(n6451), .B(STATE_REG_1__SCAN_IN), .ZN(n7170) );
  INV_X1 U4173 ( .A(n3678), .ZN(n3652) );
  AOI22_X1 U4174 ( .A1(n4466), .A2(n4652), .B1(n3653), .B2(n3652), .ZN(n3654)
         );
  AND3_X1 U4175 ( .A1(n3697), .A2(n4465), .A3(n3654), .ZN(n3664) );
  NAND2_X1 U4176 ( .A1(n3669), .A2(n4675), .ZN(n3656) );
  NOR2_X1 U4177 ( .A1(n4675), .A2(n3655), .ZN(n3676) );
  NAND2_X1 U4178 ( .A1(n3656), .A2(n3503), .ZN(n3658) );
  NAND2_X1 U4179 ( .A1(n3658), .A2(n5892), .ZN(n3660) );
  NAND2_X1 U4180 ( .A1(n3660), .A2(n4551), .ZN(n3662) );
  NAND2_X1 U4181 ( .A1(n3662), .A2(n3693), .ZN(n3663) );
  NAND2_X1 U4182 ( .A1(n3663), .A2(n4528), .ZN(n3687) );
  NAND2_X1 U4183 ( .A1(n3664), .A2(n3687), .ZN(n3665) );
  NAND2_X2 U4184 ( .A1(n3665), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3774) );
  NAND2_X1 U4185 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5019) );
  OAI21_X1 U4186 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n5019), .ZN(n5232) );
  OR2_X1 U4187 ( .A1(n4454), .A2(n5232), .ZN(n3667) );
  NAND2_X1 U4188 ( .A1(n3812), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3666) );
  OAI21_X1 U4189 ( .B1(n3774), .B2(n3518), .A(n3681), .ZN(n3668) );
  INV_X1 U4190 ( .A(n3668), .ZN(n3680) );
  AND2_X2 U4191 ( .A1(n3670), .A2(n4006), .ZN(n5171) );
  NAND2_X1 U4192 ( .A1(n5171), .A2(n3669), .ZN(n4468) );
  NAND2_X1 U4193 ( .A1(n4462), .A2(n3427), .ZN(n4518) );
  AND2_X1 U4194 ( .A1(n3676), .A2(n4503), .ZN(n4558) );
  NOR2_X1 U4195 ( .A1(n4680), .A2(n3427), .ZN(n4507) );
  NAND2_X1 U4196 ( .A1(n5165), .A2(n5892), .ZN(n4505) );
  OAI211_X2 U4197 ( .C1(n4518), .C2(n3678), .A(n5145), .B(n4505), .ZN(n3684)
         );
  NAND2_X1 U4198 ( .A1(n3684), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3679) );
  INV_X1 U4199 ( .A(n3681), .ZN(n3682) );
  NOR2_X1 U4200 ( .A1(n3682), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3683)
         );
  NAND2_X1 U4201 ( .A1(n3511), .A2(n3684), .ZN(n3685) );
  MUX2_X1 U4202 ( .A(n4454), .B(n4002), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3686) );
  OAI21_X2 U4203 ( .B1(n3774), .B2(n3513), .A(n3686), .ZN(n3731) );
  INV_X1 U4204 ( .A(n3687), .ZN(n3690) );
  INV_X2 U4205 ( .A(n4488), .ZN(n3922) );
  NAND2_X1 U4206 ( .A1(n3922), .A2(n3688), .ZN(n3689) );
  NAND2_X1 U4207 ( .A1(n3690), .A2(n3689), .ZN(n4498) );
  NAND2_X1 U4208 ( .A1(n3691), .A2(n4680), .ZN(n3696) );
  NAND2_X1 U4209 ( .A1(n6441), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7145) );
  INV_X1 U4210 ( .A(n7145), .ZN(n3695) );
  OAI21_X1 U4211 ( .B1(n4551), .B2(n3671), .A(n4528), .ZN(n3692) );
  OAI21_X1 U4212 ( .B1(n3693), .B2(n4675), .A(n3692), .ZN(n3694) );
  NAND2_X1 U4213 ( .A1(n4498), .A2(n3440), .ZN(n3732) );
  NAND2_X1 U4214 ( .A1(n3731), .A2(n3732), .ZN(n3736) );
  NAND2_X1 U4216 ( .A1(n4637), .A2(n7159), .ZN(n3712) );
  AOI22_X1 U4217 ( .A1(n5845), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4218 ( .A1(n4436), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4219 ( .A1(n5855), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4220 ( .A1(n5849), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4221 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3710)
         );
  AOI22_X1 U4222 ( .A1(n5856), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4223 ( .A1(n5860), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4224 ( .A1(n4314), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4225 ( .A1(n5847), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4226 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  NAND2_X1 U4227 ( .A1(n3923), .A2(n3797), .ZN(n3711) );
  NAND2_X1 U4228 ( .A1(n3986), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4229 ( .A1(n5845), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4230 ( .A1(n5856), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4231 ( .A1(n5849), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4232 ( .A1(n3433), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4233 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3726)
         );
  AOI22_X1 U4234 ( .A1(n5855), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4235 ( .A1(n4436), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4236 ( .A1(n4407), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4237 ( .A1(n5966), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5829), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4238 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3725)
         );
  INV_X1 U4239 ( .A(n3926), .ZN(n3728) );
  NOR2_X1 U4240 ( .A1(n3427), .A2(n7159), .ZN(n3727) );
  AOI22_X1 U4241 ( .A1(n3923), .A2(n3728), .B1(n3727), .B2(n3797), .ZN(n3729)
         );
  INV_X1 U4242 ( .A(n3731), .ZN(n3734) );
  INV_X1 U4243 ( .A(n3732), .ZN(n3733) );
  NAND2_X1 U4244 ( .A1(n3734), .A2(n3733), .ZN(n3735) );
  AOI22_X1 U4245 ( .A1(n4144), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4246 ( .A1(n5858), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4247 ( .A1(n3433), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4248 ( .A1(n5847), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4249 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3746)
         );
  AOI22_X1 U4250 ( .A1(n5845), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4251 ( .A1(n4436), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4252 ( .A1(n5966), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4253 ( .A1(n5849), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4254 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3745)
         );
  INV_X1 U4255 ( .A(n3798), .ZN(n3747) );
  XNOR2_X1 U4256 ( .A(n3747), .B(n3926), .ZN(n3748) );
  NAND2_X1 U4257 ( .A1(n3748), .A2(n3923), .ZN(n3760) );
  INV_X1 U4258 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5065) );
  AOI21_X1 U4259 ( .B1(n3688), .B2(n3926), .A(n7159), .ZN(n3750) );
  NAND2_X1 U4260 ( .A1(n4528), .A2(n3798), .ZN(n3749) );
  OAI211_X1 U4261 ( .C1(n3979), .C2(n5065), .A(n3750), .B(n3749), .ZN(n3758)
         );
  AND2_X1 U4262 ( .A1(n3923), .A2(n3926), .ZN(n3751) );
  NAND2_X1 U4263 ( .A1(n4011), .A2(n3922), .ZN(n3757) );
  XNOR2_X1 U4264 ( .A(n3798), .B(n3797), .ZN(n3754) );
  INV_X1 U4265 ( .A(n3836), .ZN(n6827) );
  INV_X1 U4266 ( .A(n3752), .ZN(n3753) );
  OAI211_X1 U4267 ( .C1(n3754), .C2(n6827), .A(n3753), .B(n3655), .ZN(n3755)
         );
  INV_X1 U4268 ( .A(n3755), .ZN(n3756) );
  NAND2_X1 U4269 ( .A1(n4528), .A2(n3671), .ZN(n3799) );
  OAI21_X1 U4270 ( .B1(n6827), .B2(n3798), .A(n3799), .ZN(n3761) );
  INV_X1 U4271 ( .A(n3761), .ZN(n3762) );
  OAI21_X1 U4272 ( .B1(n4018), .B2(n4488), .A(n3762), .ZN(n4514) );
  AND2_X1 U4273 ( .A1(n4514), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4606)
         );
  NAND2_X1 U4274 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3763)
         );
  NAND2_X1 U4275 ( .A1(n3802), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6662)
         );
  INV_X1 U4276 ( .A(n3766), .ZN(n3767) );
  NAND2_X1 U4277 ( .A1(n3770), .A2(n3769), .ZN(n3795) );
  INV_X1 U4278 ( .A(n3795), .ZN(n3793) );
  OAI21_X2 U4279 ( .B1(n3773), .B2(n3432), .A(n3771), .ZN(n3807) );
  INV_X1 U4280 ( .A(n5019), .ZN(n3775) );
  NAND2_X1 U4281 ( .A1(n3775), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U4282 ( .A1(n5019), .A2(n5224), .ZN(n3776) );
  INV_X1 U4283 ( .A(n4454), .ZN(n3813) );
  AOI22_X1 U4284 ( .A1(n4646), .A2(n3813), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3812), .ZN(n3777) );
  INV_X1 U4285 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5059) );
  AOI22_X1 U4286 ( .A1(n4144), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4287 ( .A1(n5860), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4288 ( .A1(n5856), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4289 ( .A1(n5857), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4290 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4291 ( .A1(n5845), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4292 ( .A1(n3820), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4293 ( .A1(n5849), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4294 ( .A1(n5966), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4295 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  NAND2_X1 U4296 ( .A1(n3996), .A2(n3832), .ZN(n3790) );
  OAI21_X1 U4297 ( .B1(n5059), .B2(n3979), .A(n3790), .ZN(n3791) );
  NAND2_X1 U4298 ( .A1(n3795), .A2(n3794), .ZN(n3796) );
  NAND2_X1 U4299 ( .A1(n3798), .A2(n3797), .ZN(n3834) );
  XNOR2_X1 U4300 ( .A(n3834), .B(n3832), .ZN(n3800) );
  OAI21_X1 U4301 ( .B1(n3800), .B2(n6827), .A(n3799), .ZN(n3801) );
  AOI21_X2 U4302 ( .B1(n4863), .B2(n3922), .A(n3801), .ZN(n6664) );
  NAND2_X1 U4303 ( .A1(n6662), .A2(n6664), .ZN(n3805) );
  NAND2_X1 U4304 ( .A1(n3805), .A2(n6663), .ZN(n3840) );
  INV_X1 U4305 ( .A(n3840), .ZN(n3806) );
  INV_X1 U4306 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4307 ( .A1(n3806), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4819)
         );
  INV_X1 U4308 ( .A(n3807), .ZN(n3809) );
  INV_X1 U4309 ( .A(n4739), .ZN(n3810) );
  NAND2_X1 U4310 ( .A1(n3810), .A2(n7128), .ZN(n5333) );
  NAND2_X1 U4311 ( .A1(n4739), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3811) );
  NAND2_X1 U4312 ( .A1(n5333), .A2(n3811), .ZN(n5233) );
  AOI22_X1 U4313 ( .A1(n5233), .A2(n3813), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3812), .ZN(n3814) );
  AOI22_X1 U4314 ( .A1(n5855), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4315 ( .A1(n5845), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4316 ( .A1(n3433), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4317 ( .A1(n5966), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4318 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3826)
         );
  AOI22_X1 U4319 ( .A1(n4436), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4320 ( .A1(n3820), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4321 ( .A1(n5847), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4322 ( .A1(n5849), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4323 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3825)
         );
  AOI22_X1 U4324 ( .A1(n3986), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3996), 
        .B2(n3853), .ZN(n3827) );
  NAND2_X1 U4325 ( .A1(n3830), .A2(n4933), .ZN(n3831) );
  INV_X1 U4326 ( .A(n3832), .ZN(n3833) );
  NAND2_X1 U4327 ( .A1(n3834), .A2(n3833), .ZN(n3854) );
  INV_X1 U4328 ( .A(n3853), .ZN(n3835) );
  XNOR2_X1 U4329 ( .A(n3854), .B(n3835), .ZN(n3837) );
  AND2_X1 U4330 ( .A1(n3837), .A2(n5979), .ZN(n3838) );
  AOI21_X1 U4331 ( .B1(n5156), .B2(n3922), .A(n3838), .ZN(n4821) );
  NAND2_X1 U4332 ( .A1(n4819), .A2(n4821), .ZN(n3841) );
  NAND2_X1 U4333 ( .A1(n3840), .A2(n3839), .ZN(n4820) );
  NAND2_X1 U4334 ( .A1(n3841), .A2(n4820), .ZN(n4797) );
  INV_X1 U4335 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5080) );
  INV_X1 U4336 ( .A(n3583), .ZN(n4430) );
  AOI22_X1 U4337 ( .A1(n5855), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4338 ( .A1(n5845), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4339 ( .A1(n3433), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4340 ( .A1(n5966), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4341 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3851)
         );
  AOI22_X1 U4342 ( .A1(n4436), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4343 ( .A1(n5858), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4344 ( .A1(n5847), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4345 ( .A1(n5849), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4346 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  NAND2_X1 U4347 ( .A1(n3996), .A2(n3879), .ZN(n3852) );
  OAI21_X1 U4348 ( .B1(n3979), .B2(n5080), .A(n3852), .ZN(n3860) );
  NAND2_X1 U4349 ( .A1(n4031), .A2(n3922), .ZN(n3857) );
  NAND2_X1 U4350 ( .A1(n3854), .A2(n3853), .ZN(n3881) );
  XNOR2_X1 U4351 ( .A(n3881), .B(n3879), .ZN(n3855) );
  NAND2_X1 U4352 ( .A1(n3855), .A2(n5979), .ZN(n3856) );
  NAND2_X1 U4353 ( .A1(n3858), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3859)
         );
  INV_X1 U4354 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5074) );
  AOI22_X1 U4355 ( .A1(n3433), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4356 ( .A1(n5855), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4357 ( .A1(n5860), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4358 ( .A1(n5856), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4359 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3872)
         );
  AOI22_X1 U4360 ( .A1(n4436), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4361 ( .A1(n5849), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4362 ( .A1(n5845), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4363 ( .A1(n5848), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4364 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  NAND2_X1 U4365 ( .A1(n3996), .A2(n3882), .ZN(n3873) );
  OAI21_X1 U4366 ( .B1(n3979), .B2(n5074), .A(n3873), .ZN(n3875) );
  NAND2_X1 U4367 ( .A1(n3874), .A2(n3875), .ZN(n3905) );
  INV_X1 U4368 ( .A(n3875), .ZN(n3876) );
  NAND2_X1 U4369 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  NAND2_X1 U4370 ( .A1(n4049), .A2(n3922), .ZN(n3885) );
  INV_X1 U4371 ( .A(n3879), .ZN(n3880) );
  NOR2_X1 U4372 ( .A1(n3881), .A2(n3880), .ZN(n3883) );
  NAND2_X1 U4373 ( .A1(n3883), .A2(n3882), .ZN(n3914) );
  OAI211_X1 U4374 ( .C1(n3883), .C2(n3882), .A(n3914), .B(n5979), .ZN(n3884)
         );
  INV_X1 U4375 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U4376 ( .A1(n4801), .A2(n4802), .ZN(n3889) );
  NAND2_X1 U4377 ( .A1(n3887), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3888)
         );
  NAND2_X1 U4378 ( .A1(n3889), .A2(n3888), .ZN(n6791) );
  INV_X1 U4379 ( .A(n3905), .ZN(n3903) );
  NAND2_X1 U4380 ( .A1(n3986), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4381 ( .A1(n5855), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4382 ( .A1(n5845), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4383 ( .A1(n3433), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4384 ( .A1(n5966), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4385 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3899)
         );
  AOI22_X1 U4386 ( .A1(n4436), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4387 ( .A1(n5858), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4388 ( .A1(n5847), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4389 ( .A1(n5849), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4390 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  NAND2_X1 U4391 ( .A1(n3996), .A2(n3915), .ZN(n3900) );
  NAND2_X1 U4392 ( .A1(n3905), .A2(n3904), .ZN(n4055) );
  NAND3_X1 U4393 ( .A1(n3913), .A2(n4055), .A3(n3922), .ZN(n3908) );
  XNOR2_X1 U4394 ( .A(n3914), .B(n3915), .ZN(n3906) );
  NAND2_X1 U4395 ( .A1(n3906), .A2(n5979), .ZN(n3907) );
  NAND2_X1 U4396 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  NAND2_X1 U4397 ( .A1(n6791), .A2(n6793), .ZN(n3910) );
  NAND2_X1 U4398 ( .A1(n3909), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6792)
         );
  INV_X1 U4399 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U4400 ( .A1(n3996), .A2(n3926), .ZN(n3911) );
  OAI21_X1 U4401 ( .B1(n5068), .B2(n3979), .A(n3911), .ZN(n3912) );
  NAND2_X1 U4402 ( .A1(n4059), .A2(n3922), .ZN(n3919) );
  INV_X1 U4403 ( .A(n3914), .ZN(n3916) );
  NAND2_X1 U4404 ( .A1(n3916), .A2(n3915), .ZN(n3925) );
  XNOR2_X1 U4405 ( .A(n3925), .B(n3926), .ZN(n3917) );
  NAND2_X1 U4406 ( .A1(n3917), .A2(n5979), .ZN(n3918) );
  NAND2_X1 U4407 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  INV_X1 U4408 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6906) );
  XNOR2_X1 U4409 ( .A(n3920), .B(n6906), .ZN(n6798) );
  NAND2_X1 U4410 ( .A1(n3920), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3921)
         );
  INV_X1 U4411 ( .A(n3925), .ZN(n3927) );
  NAND3_X1 U4412 ( .A1(n3927), .A2(n5979), .A3(n3926), .ZN(n3928) );
  NAND2_X1 U4413 ( .A1(n5895), .A2(n3928), .ZN(n3929) );
  INV_X1 U4414 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6900) );
  XNOR2_X1 U4415 ( .A(n3929), .B(n6900), .ZN(n5585) );
  NAND2_X1 U4416 ( .A1(n3929), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3930)
         );
  NAND2_X1 U4417 ( .A1(n5584), .A2(n3930), .ZN(n5607) );
  XNOR2_X1 U4418 ( .A(n6248), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5606)
         );
  INV_X1 U4419 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6927) );
  OR2_X1 U4420 ( .A1(n6248), .A2(n6927), .ZN(n3931) );
  INV_X1 U4421 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U4422 ( .A1(n6277), .A2(n6920), .ZN(n5640) );
  INV_X1 U4423 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5669) );
  OR2_X1 U4424 ( .A1(n6248), .A2(n6920), .ZN(n5648) );
  OR2_X1 U4425 ( .A1(n6248), .A2(n5669), .ZN(n5714) );
  INV_X1 U4426 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5451) );
  OR2_X1 U4427 ( .A1(n6248), .A2(n5451), .ZN(n5718) );
  AND3_X1 U4428 ( .A1(n5648), .A2(n5714), .A3(n5718), .ZN(n3932) );
  NAND2_X1 U4429 ( .A1(n6277), .A2(n5451), .ZN(n5717) );
  XNOR2_X1 U4430 ( .A(n6248), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5672)
         );
  INV_X1 U4431 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U4432 ( .A1(n6277), .A2(n5675), .ZN(n3933) );
  XNOR2_X1 U4433 ( .A(n6277), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5746)
         );
  NAND2_X1 U4434 ( .A1(n5747), .A2(n5746), .ZN(n5745) );
  INV_X1 U4435 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U4436 ( .A1(n6248), .A2(n6419), .ZN(n3935) );
  NAND2_X1 U4437 ( .A1(n5745), .A2(n3935), .ZN(n6285) );
  XNOR2_X1 U4438 ( .A(n6277), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6284)
         );
  INV_X1 U4439 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U4440 ( .A1(n6277), .A2(n6428), .ZN(n3936) );
  INV_X1 U4441 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5684) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6400) );
  INV_X1 U4443 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5762) );
  AND3_X1 U4444 ( .A1(n5684), .A2(n6400), .A3(n5762), .ZN(n3937) );
  NAND2_X1 U4445 ( .A1(n6225), .A2(n3937), .ZN(n3939) );
  NAND2_X1 U4446 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U4447 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6389) );
  NOR2_X1 U4448 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6218) );
  NOR2_X1 U4449 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6353) );
  AND3_X1 U4450 ( .A1(n6389), .A2(n6218), .A3(n6353), .ZN(n3941) );
  NOR2_X1 U4451 ( .A1(n6277), .A2(n3941), .ZN(n3944) );
  AND2_X1 U4452 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6388) );
  AND2_X1 U4453 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4454 ( .A1(n6388), .A2(n3942), .ZN(n5905) );
  NAND2_X1 U4455 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5909) );
  OAI21_X1 U4456 ( .B1(n5905), .B2(n5909), .A(n6277), .ZN(n3943) );
  XNOR2_X1 U4457 ( .A(n6248), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6212)
         );
  NAND2_X1 U4458 ( .A1(n6213), .A2(n6212), .ZN(n6211) );
  INV_X1 U4459 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U4460 ( .A1(n6277), .A2(n6336), .ZN(n3945) );
  INV_X1 U4461 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6337) );
  INV_X1 U4462 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6324) );
  NOR2_X1 U4463 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3946) );
  OR2_X1 U4464 ( .A1(n6248), .A2(n3946), .ZN(n5897) );
  INV_X1 U4465 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6316) );
  XNOR2_X1 U4466 ( .A(n6248), .B(n6316), .ZN(n3947) );
  NAND2_X1 U4467 ( .A1(n5927), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3960) );
  XNOR2_X1 U4468 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3961) );
  NAND2_X1 U4469 ( .A1(n3962), .A2(n3961), .ZN(n3950) );
  NAND2_X1 U4470 ( .A1(n7124), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3949) );
  NAND2_X1 U4471 ( .A1(n3950), .A2(n3949), .ZN(n3954) );
  XNOR2_X1 U4472 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3953) );
  NAND2_X1 U4473 ( .A1(n3954), .A2(n3953), .ZN(n3952) );
  NAND2_X1 U4474 ( .A1(n5224), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3951) );
  XNOR2_X1 U4475 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3981) );
  XNOR2_X1 U4476 ( .A(n3982), .B(n3981), .ZN(n4471) );
  XNOR2_X1 U4477 ( .A(n3954), .B(n3953), .ZN(n4469) );
  AND2_X1 U4478 ( .A1(n3675), .A2(n3655), .ZN(n3955) );
  NOR2_X1 U4479 ( .A1(n4507), .A2(n3955), .ZN(n3969) );
  INV_X1 U4480 ( .A(n3969), .ZN(n3958) );
  INV_X1 U4481 ( .A(n4469), .ZN(n3956) );
  NAND2_X1 U4482 ( .A1(n3996), .A2(n3956), .ZN(n3970) );
  INV_X1 U4483 ( .A(n3970), .ZN(n3957) );
  AOI211_X1 U4484 ( .C1(n3986), .C2(n4469), .A(n3958), .B(n3957), .ZN(n3978)
         );
  OAI21_X1 U4485 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5927), .A(n3960), 
        .ZN(n3966) );
  INV_X1 U4486 ( .A(n3966), .ZN(n3968) );
  XNOR2_X1 U4487 ( .A(n3962), .B(n3961), .ZN(n4470) );
  INV_X1 U4488 ( .A(n3996), .ZN(n3965) );
  OAI21_X1 U4489 ( .B1(n3965), .B2(n3675), .A(n3655), .ZN(n3963) );
  AOI21_X1 U4490 ( .B1(n3986), .B2(n4470), .A(n3963), .ZN(n3972) );
  INV_X1 U4491 ( .A(n4470), .ZN(n3964) );
  NAND2_X1 U4492 ( .A1(n3964), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3973) );
  AOI211_X1 U4493 ( .C1(n3972), .C2(n3973), .A(n3966), .B(n3965), .ZN(n3967)
         );
  NOR2_X1 U4494 ( .A1(n3967), .A2(n3999), .ZN(n3971) );
  AOI211_X1 U4495 ( .C1(n3959), .C2(n3968), .A(n4528), .B(n3971), .ZN(n3976)
         );
  AOI21_X1 U4496 ( .B1(n3971), .B2(n3970), .A(n3969), .ZN(n3975) );
  INV_X1 U4497 ( .A(n3999), .ZN(n3987) );
  AOI21_X1 U4498 ( .B1(n3987), .B2(n3973), .A(n3972), .ZN(n3974) );
  NOR3_X1 U4499 ( .A1(n3976), .A2(n3975), .A3(n3974), .ZN(n3977) );
  AOI211_X1 U4500 ( .C1(n3979), .C2(n4471), .A(n3978), .B(n3977), .ZN(n3980)
         );
  AOI21_X1 U4501 ( .B1(n4471), .B2(n3999), .A(n3980), .ZN(n3989) );
  NAND2_X1 U4502 ( .A1(n3982), .A2(n3981), .ZN(n3984) );
  NAND2_X1 U4503 ( .A1(n7128), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U4504 ( .A1(n3984), .A2(n3983), .ZN(n3993) );
  NOR2_X1 U4505 ( .A1(n3986), .A2(n4474), .ZN(n3988) );
  OAI22_X1 U4506 ( .A1(n3989), .A2(n3988), .B1(n3987), .B2(n4474), .ZN(n3990)
         );
  AOI21_X1 U4507 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7159), .A(n3990), 
        .ZN(n3998) );
  NAND2_X1 U4508 ( .A1(n3991), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U4509 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  NAND2_X1 U4510 ( .A1(n3996), .A2(n4473), .ZN(n3997) );
  NAND2_X1 U4511 ( .A1(n3998), .A2(n3997), .ZN(n4001) );
  NAND2_X1 U4512 ( .A1(n3999), .A2(n4473), .ZN(n4000) );
  NOR2_X1 U4513 ( .A1(n3752), .A2(n4003), .ZN(n4005) );
  NOR2_X1 U4514 ( .A1(n3959), .A2(n4528), .ZN(n4004) );
  OR2_X1 U4515 ( .A1(n4003), .A2(n6823), .ZN(n4035) );
  INV_X1 U4516 ( .A(n4035), .ZN(n4020) );
  NAND2_X1 U4517 ( .A1(n4020), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4010) );
  INV_X1 U4518 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U4519 ( .A1(n6823), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4181) );
  NAND2_X1 U4520 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4024) );
  OAI21_X1 U4521 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4024), .ZN(n6967) );
  NAND2_X1 U4522 ( .A1(n3426), .A2(n6967), .ZN(n4007) );
  OAI21_X1 U4523 ( .B1(n6951), .B2(n4181), .A(n4007), .ZN(n4008) );
  AOI21_X1 U4524 ( .B1(n4041), .B2(EAX_REG_2__SCAN_IN), .A(n4008), .ZN(n4009)
         );
  AND2_X1 U4525 ( .A1(n4010), .A2(n4009), .ZN(n4596) );
  BUF_X1 U4526 ( .A(n4011), .Z(n4012) );
  NAND2_X1 U4527 ( .A1(n4012), .A2(n4191), .ZN(n4017) );
  NAND2_X1 U4528 ( .A1(n4041), .A2(EAX_REG_1__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4529 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4013)
         );
  OAI211_X1 U4530 ( .C1(n4035), .C2(n3518), .A(n4014), .B(n4013), .ZN(n4015)
         );
  INV_X1 U4531 ( .A(n4015), .ZN(n4016) );
  NOR2_X1 U4532 ( .A1(n5974), .A2(n4662), .ZN(n4019) );
  AOI21_X1 U4533 ( .B1(n4018), .B2(n4019), .A(n6823), .ZN(n4568) );
  AOI22_X1 U4534 ( .A1(n4041), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6823), .ZN(n4022) );
  NAND2_X1 U4535 ( .A1(n4020), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4021) );
  OAI211_X1 U4536 ( .C1(n5934), .C2(n4030), .A(n4022), .B(n4021), .ZN(n4567)
         );
  MUX2_X1 U4537 ( .A(n3426), .B(n4568), .S(n4567), .Z(n4555) );
  NAND2_X1 U4538 ( .A1(n4595), .A2(n4596), .ZN(n4023) );
  INV_X1 U4539 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U4540 ( .A1(n6969), .A2(n4024), .ZN(n4025) );
  NAND2_X1 U4541 ( .A1(n4044), .A2(n4025), .ZN(n6968) );
  AOI22_X1 U4542 ( .A1(n3426), .A2(n6968), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4027) );
  NAND2_X1 U4543 ( .A1(n5874), .A2(EAX_REG_3__SCAN_IN), .ZN(n4026) );
  OAI211_X1 U4544 ( .C1(n4035), .C2(n5969), .A(n4027), .B(n4026), .ZN(n4028)
         );
  INV_X1 U4545 ( .A(n4028), .ZN(n4029) );
  OAI21_X1 U4546 ( .B1(n4869), .B2(n4030), .A(n4029), .ZN(n4570) );
  NAND2_X1 U4547 ( .A1(n4031), .A2(n4191), .ZN(n4040) );
  NAND2_X1 U4548 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4033)
         );
  NAND2_X1 U4549 ( .A1(n5874), .A2(EAX_REG_4__SCAN_IN), .ZN(n4032) );
  OAI211_X1 U4550 ( .C1(n4035), .C2(n4034), .A(n4033), .B(n4032), .ZN(n4038)
         );
  INV_X1 U4551 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4036) );
  XNOR2_X1 U4552 ( .A(n4044), .B(n4036), .ZN(n6996) );
  AND2_X1 U4553 ( .A1(n6996), .A2(n3426), .ZN(n4037) );
  AOI21_X1 U4554 ( .B1(n4038), .B2(n5872), .A(n4037), .ZN(n4039) );
  NAND2_X1 U4555 ( .A1(n4040), .A2(n4039), .ZN(n4622) );
  NAND2_X1 U4556 ( .A1(n4569), .A2(n4622), .ZN(n4623) );
  INV_X1 U4557 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4047) );
  INV_X1 U4558 ( .A(n4044), .ZN(n4042) );
  AOI21_X1 U4559 ( .B1(n4042), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U4560 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4043) );
  OR2_X1 U4561 ( .A1(n4045), .A2(n4050), .ZN(n7001) );
  AOI22_X1 U4562 ( .A1(n7001), .A2(n3426), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4046) );
  OAI21_X1 U4563 ( .B1(n4067), .B2(n4047), .A(n4046), .ZN(n4048) );
  INV_X1 U4564 ( .A(n4729), .ZN(n4057) );
  INV_X1 U4565 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4053) );
  NOR2_X1 U4566 ( .A1(n4050), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4051)
         );
  OR2_X1 U4567 ( .A1(n4060), .A2(n4051), .ZN(n7019) );
  AOI22_X1 U4568 ( .A1(n7019), .A2(n3426), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4052) );
  OAI21_X1 U4569 ( .B1(n4067), .B2(n4053), .A(n4052), .ZN(n4054) );
  AOI21_X1 U4570 ( .B1(n4055), .B2(n4191), .A(n4054), .ZN(n5215) );
  INV_X1 U4571 ( .A(n5215), .ZN(n4056) );
  NAND2_X1 U4572 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  NAND2_X1 U4573 ( .A1(n4059), .A2(n4191), .ZN(n4066) );
  INV_X1 U4574 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4063) );
  OR2_X1 U4575 ( .A1(n4060), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U4576 ( .A1(n4061), .A2(n4081), .ZN(n6804) );
  AOI22_X1 U4577 ( .A1(n6804), .A2(n3426), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U4578 ( .A1(n4066), .A2(n4065), .ZN(n5179) );
  XNOR2_X1 U4579 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4081), .ZN(n5592) );
  OAI22_X1 U4580 ( .A1(n5872), .A2(n5592), .B1(n4181), .B2(n5588), .ZN(n4068)
         );
  AOI21_X1 U4581 ( .B1(n5874), .B2(EAX_REG_8__SCAN_IN), .A(n4068), .ZN(n4080)
         );
  AOI22_X1 U4582 ( .A1(n5860), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4583 ( .A1(n5858), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4584 ( .A1(n5845), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4585 ( .A1(n5846), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4069) );
  NAND4_X1 U4586 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4078)
         );
  AOI22_X1 U4587 ( .A1(n5855), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4588 ( .A1(n5856), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U4589 ( .A1(n5849), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U4590 ( .A1(n4430), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U4591 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4077)
         );
  OAI21_X1 U4592 ( .B1(n4078), .B2(n4077), .A(n4191), .ZN(n4079) );
  NAND2_X1 U4593 ( .A1(n4080), .A2(n4079), .ZN(n4956) );
  XOR2_X1 U4594 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4128), .Z(n7023) );
  AOI22_X1 U4595 ( .A1(n5874), .A2(EAX_REG_11__SCAN_IN), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U4596 ( .A1(n5860), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U4597 ( .A1(n4436), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4598 ( .A1(n5966), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4599 ( .A1(n5846), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U4600 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4091)
         );
  AOI22_X1 U4601 ( .A1(n5855), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4602 ( .A1(n5845), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4603 ( .A1(n5858), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4604 ( .A1(n5849), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U4605 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  OAI21_X1 U4606 ( .B1(n4091), .B2(n4090), .A(n4191), .ZN(n4092) );
  OAI211_X1 U4607 ( .C1(n7023), .C2(n5872), .A(n4093), .B(n4092), .ZN(n4094)
         );
  INV_X1 U4608 ( .A(n4094), .ZN(n5614) );
  NOR2_X1 U4609 ( .A1(n4181), .A2(n5562), .ZN(n4095) );
  AOI21_X1 U4610 ( .B1(n5874), .B2(EAX_REG_10__SCAN_IN), .A(n4095), .ZN(n4108)
         );
  AOI22_X1 U4611 ( .A1(n4430), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U4612 ( .A1(n5855), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U4613 ( .A1(n5856), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U4614 ( .A1(n5847), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U4615 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4106)
         );
  AOI22_X1 U4616 ( .A1(n4431), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U4617 ( .A1(n5858), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U4618 ( .A1(n5845), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U4619 ( .A1(n5849), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U4620 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  OAI21_X1 U4621 ( .B1(n4106), .B2(n4105), .A(n4191), .ZN(n4107) );
  AND2_X1 U4622 ( .A1(n4108), .A2(n4107), .ZN(n4111) );
  XNOR2_X1 U4623 ( .A(n4109), .B(n5562), .ZN(n5644) );
  NAND2_X1 U4624 ( .A1(n5644), .A2(n3426), .ZN(n4110) );
  XOR2_X1 U4625 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4112), .Z(n5608) );
  AOI22_X1 U4626 ( .A1(n5874), .A2(EAX_REG_9__SCAN_IN), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U4627 ( .A1(n5845), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U4628 ( .A1(n4436), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U4629 ( .A1(n5849), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U4630 ( .A1(n5855), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4113) );
  NAND4_X1 U4631 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4122)
         );
  AOI22_X1 U4632 ( .A1(n4430), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U4633 ( .A1(n5860), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U4634 ( .A1(n5856), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U4635 ( .A1(n5847), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U4636 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4121)
         );
  OAI21_X1 U4637 ( .B1(n4122), .B2(n4121), .A(n4191), .ZN(n4123) );
  OAI211_X1 U4638 ( .C1(n5608), .C2(n5872), .A(n4124), .B(n4123), .ZN(n4125)
         );
  INV_X1 U4639 ( .A(n4125), .ZN(n5459) );
  NOR2_X1 U4640 ( .A1(n3512), .A2(n5459), .ZN(n4126) );
  XNOR2_X1 U4641 ( .A(n4159), .B(n5547), .ZN(n5722) );
  NAND2_X1 U4642 ( .A1(n5722), .A2(n3426), .ZN(n4143) );
  INV_X1 U4643 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4129) );
  OAI22_X1 U4644 ( .A1(n4067), .A2(n4129), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5547), .ZN(n4141) );
  AOI22_X1 U4645 ( .A1(n5845), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U4646 ( .A1(n5858), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U4647 ( .A1(n5855), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U4648 ( .A1(n5846), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U4649 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4139)
         );
  AOI22_X1 U4650 ( .A1(n5860), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U4651 ( .A1(n5856), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U4652 ( .A1(n5849), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4653 ( .A1(n4430), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4134) );
  NAND4_X1 U4654 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  OR2_X1 U4655 ( .A1(n4139), .A2(n4138), .ZN(n4140) );
  AOI22_X1 U4656 ( .A1(n4141), .A2(n5872), .B1(n4191), .B2(n4140), .ZN(n4142)
         );
  NAND2_X1 U4657 ( .A1(n4143), .A2(n4142), .ZN(n5433) );
  AOI22_X1 U4658 ( .A1(n5845), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U4659 ( .A1(n5860), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U4660 ( .A1(n4436), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U4661 ( .A1(n4430), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4145) );
  NAND4_X1 U4662 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4154)
         );
  AOI22_X1 U4663 ( .A1(n5858), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U4664 ( .A1(n5966), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U4665 ( .A1(n5847), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U4666 ( .A1(n5849), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4149) );
  NAND4_X1 U4667 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4153)
         );
  OR2_X1 U4668 ( .A1(n4154), .A2(n4153), .ZN(n4155) );
  AND2_X1 U4669 ( .A1(n4191), .A2(n4155), .ZN(n4157) );
  INV_X1 U4670 ( .A(n4157), .ZN(n4158) );
  INV_X1 U4671 ( .A(n5572), .ZN(n4164) );
  INV_X1 U4672 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5740) );
  OAI21_X1 U4673 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4160), .A(n4179), 
        .ZN(n7032) );
  NAND2_X1 U4674 ( .A1(n3426), .A2(n7032), .ZN(n4161) );
  OAI21_X1 U4675 ( .B1(n4181), .B2(n5740), .A(n4161), .ZN(n4162) );
  AOI21_X1 U4676 ( .B1(n5874), .B2(EAX_REG_13__SCAN_IN), .A(n4162), .ZN(n5571)
         );
  NAND2_X1 U4677 ( .A1(n4164), .A2(n4163), .ZN(n5574) );
  XOR2_X1 U4678 ( .A(n7042), .B(n4179), .Z(n7047) );
  OAI22_X1 U4679 ( .A1(n7047), .A2(n5872), .B1(n4181), .B2(n7042), .ZN(n4166)
         );
  AOI21_X1 U4680 ( .B1(n5874), .B2(EAX_REG_14__SCAN_IN), .A(n4166), .ZN(n4178)
         );
  AOI22_X1 U4681 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n4430), .B1(n5966), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4682 ( .A1(n5845), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4683 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n4431), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4684 ( .A1(n5858), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U4685 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4176)
         );
  AOI22_X1 U4686 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n5856), .B1(n4436), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4687 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n5857), .B1(n5846), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U4688 ( .A1(n5849), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U4689 ( .A1(n5855), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4171) );
  NAND4_X1 U4690 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4175)
         );
  OAI21_X1 U4691 ( .B1(n4176), .B2(n4175), .A(n4191), .ZN(n4177) );
  NAND2_X1 U4692 ( .A1(n4178), .A2(n4177), .ZN(n5621) );
  INV_X1 U4693 ( .A(n4197), .ZN(n4180) );
  XNOR2_X1 U4694 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4180), .ZN(n7060)
         );
  INV_X1 U4695 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6286) );
  OAI22_X1 U4696 ( .A1(n7060), .A2(n5872), .B1(n4181), .B2(n6286), .ZN(n4182)
         );
  AOI21_X1 U4697 ( .B1(n5874), .B2(EAX_REG_15__SCAN_IN), .A(n4182), .ZN(n4195)
         );
  AOI22_X1 U4698 ( .A1(n5860), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4699 ( .A1(n5856), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U4700 ( .A1(n4430), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U4701 ( .A1(n5847), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4183) );
  NAND4_X1 U4702 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4193)
         );
  AOI22_X1 U4703 ( .A1(n4436), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U4704 ( .A1(n5845), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4705 ( .A1(n5855), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U4706 ( .A1(n5849), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4187) );
  NAND4_X1 U4707 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(n4192)
         );
  OAI21_X1 U4708 ( .B1(n4193), .B2(n4192), .A(n4191), .ZN(n4194) );
  XOR2_X1 U4709 ( .A(n5706), .B(n4211), .Z(n5704) );
  INV_X1 U4710 ( .A(n5704), .ZN(n6280) );
  INV_X1 U4711 ( .A(n4551), .ZN(n6436) );
  AOI22_X1 U4712 ( .A1(n4431), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U4713 ( .A1(n4436), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U4714 ( .A1(n5860), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4715 ( .A1(n5847), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4198) );
  NAND4_X1 U4716 ( .A1(n4201), .A2(n4200), .A3(n4199), .A4(n4198), .ZN(n4207)
         );
  INV_X1 U4717 ( .A(n3583), .ZN(n4314) );
  AOI22_X1 U4718 ( .A1(n4314), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U4719 ( .A1(n5845), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5855), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U4720 ( .A1(n5858), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4721 ( .A1(n5849), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U4722 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4206)
         );
  NOR2_X1 U4723 ( .A1(n4207), .A2(n4206), .ZN(n4209) );
  AOI22_X1 U4724 ( .A1(n5874), .A2(EAX_REG_16__SCAN_IN), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4208) );
  OAI21_X1 U4725 ( .B1(n4443), .B2(n4209), .A(n4208), .ZN(n4210) );
  AOI21_X1 U4726 ( .B1(n6280), .B2(n3426), .A(n4210), .ZN(n5681) );
  XNOR2_X1 U4727 ( .A(n4239), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6272)
         );
  AOI21_X1 U4728 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6270), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4212) );
  AOI21_X1 U4729 ( .B1(n5874), .B2(EAX_REG_17__SCAN_IN), .A(n4212), .ZN(n4224)
         );
  AOI22_X1 U4730 ( .A1(n4314), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U4731 ( .A1(n5856), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U4732 ( .A1(n5849), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U4733 ( .A1(n5857), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U4734 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4222)
         );
  AOI22_X1 U4735 ( .A1(n5845), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U4736 ( .A1(n3433), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U4737 ( .A1(n5855), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U4738 ( .A1(n5858), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U4739 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4221)
         );
  OAI21_X1 U4740 ( .B1(n4222), .B2(n4221), .A(n5869), .ZN(n4223) );
  AOI22_X1 U4741 ( .A1(n6272), .A2(n3426), .B1(n4224), .B2(n4223), .ZN(n5698)
         );
  NAND2_X1 U4742 ( .A1(n5680), .A2(n5698), .ZN(n5697) );
  AOI22_X1 U4743 ( .A1(n5845), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5855), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U4744 ( .A1(n4436), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U4745 ( .A1(n4314), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U4746 ( .A1(n5857), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4225) );
  NAND4_X1 U4747 ( .A1(n4228), .A2(n4227), .A3(n4226), .A4(n4225), .ZN(n4234)
         );
  AOI22_X1 U4748 ( .A1(n4431), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U4749 ( .A1(n5860), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U4750 ( .A1(n5858), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5847), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U4751 ( .A1(n5849), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4229) );
  NAND4_X1 U4752 ( .A1(n4232), .A2(n4231), .A3(n4230), .A4(n4229), .ZN(n4233)
         );
  NOR2_X1 U4753 ( .A1(n4234), .A2(n4233), .ZN(n4238) );
  NAND2_X1 U4754 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4235)
         );
  NAND2_X1 U4755 ( .A1(n5872), .A2(n4235), .ZN(n4236) );
  AOI21_X1 U4756 ( .B1(n5874), .B2(EAX_REG_18__SCAN_IN), .A(n4236), .ZN(n4237)
         );
  OAI21_X1 U4757 ( .B1(n4443), .B2(n4238), .A(n4237), .ZN(n4242) );
  OAI21_X1 U4758 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4240), .A(n4274), 
        .ZN(n6814) );
  OR2_X1 U4759 ( .A1(n5872), .A2(n6814), .ZN(n4241) );
  NAND2_X1 U4760 ( .A1(n4242), .A2(n4241), .ZN(n5760) );
  AOI22_X1 U4761 ( .A1(n4436), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U4762 ( .A1(n5845), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U4763 ( .A1(n4430), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4245) );
  AOI22_X1 U4764 ( .A1(n5858), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4244) );
  NAND4_X1 U4765 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(n4253)
         );
  AOI22_X1 U4766 ( .A1(n5860), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4767 ( .A1(n5855), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4768 ( .A1(n5857), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U4769 ( .A1(n5849), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4248) );
  NAND4_X1 U4770 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4252)
         );
  NOR2_X1 U4771 ( .A1(n4253), .A2(n4252), .ZN(n4257) );
  NAND2_X1 U4772 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4254)
         );
  NAND2_X1 U4773 ( .A1(n5872), .A2(n4254), .ZN(n4255) );
  AOI21_X1 U4774 ( .B1(n5874), .B2(EAX_REG_19__SCAN_IN), .A(n4255), .ZN(n4256)
         );
  OAI21_X1 U4775 ( .B1(n4443), .B2(n4257), .A(n4256), .ZN(n4259) );
  XNOR2_X1 U4776 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4274), .ZN(n6092)
         );
  NAND2_X1 U4777 ( .A1(n3426), .A2(n6092), .ZN(n4258) );
  NAND2_X1 U4778 ( .A1(n4259), .A2(n4258), .ZN(n6089) );
  AOI22_X1 U4779 ( .A1(n5860), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U4780 ( .A1(n4436), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U4781 ( .A1(n5857), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U4782 ( .A1(n5855), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4260) );
  NAND4_X1 U4783 ( .A1(n4263), .A2(n4262), .A3(n4261), .A4(n4260), .ZN(n4269)
         );
  AOI22_X1 U4784 ( .A1(n5845), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4785 ( .A1(n4430), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U4786 ( .A1(n5858), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4265) );
  AOI22_X1 U4787 ( .A1(n5849), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4264) );
  NAND4_X1 U4788 ( .A1(n4267), .A2(n4266), .A3(n4265), .A4(n4264), .ZN(n4268)
         );
  NOR2_X1 U4789 ( .A1(n4269), .A2(n4268), .ZN(n4273) );
  NAND2_X1 U4790 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4270)
         );
  NAND2_X1 U4791 ( .A1(n5872), .A2(n4270), .ZN(n4271) );
  AOI21_X1 U4792 ( .B1(n5874), .B2(EAX_REG_20__SCAN_IN), .A(n4271), .ZN(n4272)
         );
  OAI21_X1 U4793 ( .B1(n4443), .B2(n4273), .A(n4272), .ZN(n4278) );
  OAI21_X1 U4794 ( .B1(n4276), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4308), 
        .ZN(n6251) );
  OR2_X1 U4795 ( .A1(n6251), .A2(n5872), .ZN(n4277) );
  AOI22_X1 U4796 ( .A1(n5860), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U4797 ( .A1(n5849), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U4798 ( .A1(n5856), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U4799 ( .A1(n5966), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4279) );
  NAND4_X1 U4800 ( .A1(n4282), .A2(n4281), .A3(n4280), .A4(n4279), .ZN(n4288)
         );
  AOI22_X1 U4801 ( .A1(n5855), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U4802 ( .A1(n5845), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U4803 ( .A1(n5858), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U4804 ( .A1(n5847), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4283) );
  NAND4_X1 U4805 ( .A1(n4286), .A2(n4285), .A3(n4284), .A4(n4283), .ZN(n4287)
         );
  NOR2_X1 U4806 ( .A1(n4288), .A2(n4287), .ZN(n4291) );
  OAI21_X1 U4807 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6244), .A(n5872), .ZN(
        n4289) );
  AOI21_X1 U4808 ( .B1(n5874), .B2(EAX_REG_21__SCAN_IN), .A(n4289), .ZN(n4290)
         );
  OAI21_X1 U4809 ( .B1(n4443), .B2(n4291), .A(n4290), .ZN(n4293) );
  XNOR2_X1 U4810 ( .A(n4308), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n7070)
         );
  NAND2_X1 U4811 ( .A1(n7070), .A2(n3426), .ZN(n4292) );
  NAND2_X1 U4812 ( .A1(n6077), .A2(n6152), .ZN(n6060) );
  AOI22_X1 U4813 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n4431), .B1(n5860), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U4814 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n5858), .B1(n5857), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U4815 ( .A1(n5845), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4816 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5856), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4294) );
  NAND4_X1 U4817 ( .A1(n4297), .A2(n4296), .A3(n4295), .A4(n4294), .ZN(n4303)
         );
  AOI22_X1 U4818 ( .A1(n5855), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4436), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U4819 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5847), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U4820 ( .A1(n5849), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U4821 ( .A1(n4430), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4298) );
  NAND4_X1 U4822 ( .A1(n4301), .A2(n4300), .A3(n4299), .A4(n4298), .ZN(n4302)
         );
  NOR2_X1 U4823 ( .A1(n4303), .A2(n4302), .ZN(n4307) );
  NAND2_X1 U4824 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4304)
         );
  NAND2_X1 U4825 ( .A1(n5872), .A2(n4304), .ZN(n4305) );
  AOI21_X1 U4826 ( .B1(n5874), .B2(EAX_REG_22__SCAN_IN), .A(n4305), .ZN(n4306)
         );
  OAI21_X1 U4827 ( .B1(n4443), .B2(n4307), .A(n4306), .ZN(n4312) );
  OR2_X1 U4828 ( .A1(n4309), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4310)
         );
  AND2_X1 U4829 ( .A1(n4354), .A2(n4310), .ZN(n6238) );
  NAND2_X1 U4830 ( .A1(n6238), .A2(n3426), .ZN(n4311) );
  NAND2_X1 U4831 ( .A1(n4312), .A2(n4311), .ZN(n6063) );
  AOI22_X1 U4832 ( .A1(n5845), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U4833 ( .A1(n5856), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U4834 ( .A1(n4314), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U4835 ( .A1(n5847), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4315) );
  NAND4_X1 U4836 ( .A1(n4318), .A2(n4317), .A3(n4316), .A4(n4315), .ZN(n4324)
         );
  AOI22_X1 U4837 ( .A1(n5855), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4838 ( .A1(n4436), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4839 ( .A1(n4431), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U4840 ( .A1(n5849), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4319) );
  NAND4_X1 U4841 ( .A1(n4322), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(n4323)
         );
  NOR2_X1 U4842 ( .A1(n4324), .A2(n4323), .ZN(n4341) );
  AOI22_X1 U4843 ( .A1(n5856), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U4844 ( .A1(n3433), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U4845 ( .A1(n5855), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4846 ( .A1(n4407), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4325) );
  NAND4_X1 U4847 ( .A1(n4328), .A2(n4327), .A3(n4326), .A4(n4325), .ZN(n4334)
         );
  AOI22_X1 U4848 ( .A1(n5845), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U4849 ( .A1(n4436), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4850 ( .A1(n4430), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4851 ( .A1(n5849), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4329) );
  NAND4_X1 U4852 ( .A1(n4332), .A2(n4331), .A3(n4330), .A4(n4329), .ZN(n4333)
         );
  NOR2_X1 U4853 ( .A1(n4334), .A2(n4333), .ZN(n4342) );
  XOR2_X1 U4854 ( .A(n4341), .B(n4342), .Z(n4335) );
  NAND2_X1 U4855 ( .A1(n4335), .A2(n5869), .ZN(n4338) );
  INV_X1 U4856 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n7090) );
  OAI21_X1 U4857 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7090), .A(n5872), .ZN(
        n4336) );
  AOI21_X1 U4858 ( .B1(n5874), .B2(EAX_REG_23__SCAN_IN), .A(n4336), .ZN(n4337)
         );
  NAND2_X1 U4859 ( .A1(n4338), .A2(n4337), .ZN(n4340) );
  XNOR2_X1 U4860 ( .A(n4354), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n7080)
         );
  NAND2_X1 U4861 ( .A1(n7080), .A2(n3426), .ZN(n4339) );
  NAND2_X1 U4862 ( .A1(n4340), .A2(n4339), .ZN(n6143) );
  OR2_X1 U4863 ( .A1(n4342), .A2(n4341), .ZN(n4371) );
  AOI22_X1 U4864 ( .A1(n4431), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4865 ( .A1(n5845), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5855), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U4866 ( .A1(n4430), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U4867 ( .A1(n5860), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4343) );
  NAND4_X1 U4868 ( .A1(n4346), .A2(n4345), .A3(n4344), .A4(n4343), .ZN(n4352)
         );
  AOI22_X1 U4869 ( .A1(n5856), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4870 ( .A1(n5849), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4871 ( .A1(n4436), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4872 ( .A1(n5847), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4347) );
  NAND4_X1 U4873 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4351)
         );
  NOR2_X1 U4874 ( .A1(n4352), .A2(n4351), .ZN(n4370) );
  INV_X1 U4875 ( .A(n4370), .ZN(n4353) );
  XNOR2_X1 U4876 ( .A(n4371), .B(n4353), .ZN(n4358) );
  XNOR2_X1 U4877 ( .A(n4375), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n7102)
         );
  NAND2_X1 U4878 ( .A1(n5874), .A2(EAX_REG_24__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U4879 ( .A1(n5941), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4355)
         );
  OAI211_X1 U4880 ( .C1(n7102), .C2(n5872), .A(n4356), .B(n4355), .ZN(n4357)
         );
  AOI21_X1 U4881 ( .B1(n4358), .B2(n5869), .A(n4357), .ZN(n6222) );
  AOI22_X1 U4882 ( .A1(n5855), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U4883 ( .A1(n4436), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U4884 ( .A1(n5966), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U4885 ( .A1(n5846), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4359) );
  NAND4_X1 U4886 ( .A1(n4362), .A2(n4361), .A3(n4360), .A4(n4359), .ZN(n4369)
         );
  AOI22_X1 U4887 ( .A1(n5845), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U4888 ( .A1(n5858), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4363), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U4889 ( .A1(n5860), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4890 ( .A1(n5849), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4364) );
  NAND4_X1 U4891 ( .A1(n4367), .A2(n4366), .A3(n4365), .A4(n4364), .ZN(n4368)
         );
  NOR2_X1 U4892 ( .A1(n4369), .A2(n4368), .ZN(n4381) );
  OR2_X1 U4893 ( .A1(n4371), .A2(n4370), .ZN(n4380) );
  XOR2_X1 U4894 ( .A(n4381), .B(n4380), .Z(n4372) );
  NAND2_X1 U4895 ( .A1(n4372), .A2(n5869), .ZN(n4379) );
  NAND2_X1 U4896 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4373)
         );
  NAND2_X1 U4897 ( .A1(n5872), .A2(n4373), .ZN(n4374) );
  AOI21_X1 U4898 ( .B1(n5874), .B2(EAX_REG_25__SCAN_IN), .A(n4374), .ZN(n4378)
         );
  XNOR2_X1 U4899 ( .A(n4397), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6210)
         );
  AOI21_X1 U4900 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(n6047) );
  NAND2_X1 U4901 ( .A1(n6046), .A2(n6047), .ZN(n6034) );
  NOR2_X1 U4902 ( .A1(n4381), .A2(n4380), .ZN(n4415) );
  AOI22_X1 U4903 ( .A1(n5855), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U4904 ( .A1(n5845), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4905 ( .A1(n4431), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4906 ( .A1(n5966), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4382) );
  NAND4_X1 U4907 ( .A1(n4385), .A2(n4384), .A3(n4383), .A4(n4382), .ZN(n4391)
         );
  AOI22_X1 U4908 ( .A1(n4436), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U4909 ( .A1(n5858), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U4910 ( .A1(n5847), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U4911 ( .A1(n5849), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4386) );
  NAND4_X1 U4912 ( .A1(n4389), .A2(n4388), .A3(n4387), .A4(n4386), .ZN(n4390)
         );
  OR2_X1 U4913 ( .A1(n4391), .A2(n4390), .ZN(n4414) );
  INV_X1 U4914 ( .A(n4414), .ZN(n4392) );
  XNOR2_X1 U4915 ( .A(n4415), .B(n4392), .ZN(n4396) );
  INV_X1 U4916 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U4917 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4393)
         );
  OAI211_X1 U4918 ( .C1(n4067), .C2(n4394), .A(n5872), .B(n4393), .ZN(n4395)
         );
  AOI21_X1 U4919 ( .B1(n4396), .B2(n5869), .A(n4395), .ZN(n4402) );
  INV_X1 U4920 ( .A(n4397), .ZN(n4398) );
  NAND2_X1 U4921 ( .A1(n4398), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4399)
         );
  INV_X1 U4922 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U4923 ( .A1(n4399), .A2(n6039), .ZN(n4400) );
  NAND2_X1 U4924 ( .A1(n4424), .A2(n4400), .ZN(n6204) );
  NOR2_X1 U4925 ( .A1(n6204), .A2(n5872), .ZN(n4401) );
  NOR2_X2 U4926 ( .A1(n6034), .A2(n6037), .ZN(n6020) );
  AOI22_X1 U4927 ( .A1(n5845), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5855), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U4928 ( .A1(n5856), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4929 ( .A1(n4430), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U4930 ( .A1(n5846), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4403) );
  NAND4_X1 U4931 ( .A1(n4406), .A2(n4405), .A3(n4404), .A4(n4403), .ZN(n4413)
         );
  AOI22_X1 U4932 ( .A1(n5860), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4933 ( .A1(n4436), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5858), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4934 ( .A1(n4431), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4935 ( .A1(n5849), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U4936 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4412)
         );
  NOR2_X1 U4937 ( .A1(n4413), .A2(n4412), .ZN(n4429) );
  NAND2_X1 U4938 ( .A1(n4415), .A2(n4414), .ZN(n4428) );
  XOR2_X1 U4939 ( .A(n4429), .B(n4428), .Z(n4419) );
  INV_X1 U4940 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U4941 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4416)
         );
  OAI211_X1 U4942 ( .C1(n4067), .C2(n4417), .A(n5872), .B(n4416), .ZN(n4418)
         );
  AOI21_X1 U4943 ( .B1(n4419), .B2(n5869), .A(n4418), .ZN(n4420) );
  INV_X1 U4944 ( .A(n4420), .ZN(n4422) );
  XNOR2_X1 U4945 ( .A(n4424), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6198)
         );
  NAND2_X1 U4946 ( .A1(n6198), .A2(n3426), .ZN(n4421) );
  NAND2_X1 U4947 ( .A1(n4422), .A2(n4421), .ZN(n6021) );
  INV_X1 U4948 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6196) );
  INV_X1 U4949 ( .A(n4425), .ZN(n4426) );
  INV_X1 U4950 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U4951 ( .A1(n4426), .A2(n4455), .ZN(n4427) );
  OAI21_X1 U4952 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4455), .A(n5872), .ZN(
        n4446) );
  NOR2_X1 U4953 ( .A1(n4429), .A2(n4428), .ZN(n5837) );
  AOI22_X1 U4954 ( .A1(n5855), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U4955 ( .A1(n5845), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5860), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U4956 ( .A1(n4431), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U4957 ( .A1(n5966), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4432) );
  NAND4_X1 U4958 ( .A1(n4435), .A2(n4434), .A3(n4433), .A4(n4432), .ZN(n4442)
         );
  AOI22_X1 U4959 ( .A1(n4436), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U4960 ( .A1(n5858), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U4961 ( .A1(n5847), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U4962 ( .A1(n5849), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4437) );
  NAND4_X1 U4963 ( .A1(n4440), .A2(n4439), .A3(n4438), .A4(n4437), .ZN(n4441)
         );
  OR2_X1 U4964 ( .A1(n4442), .A2(n4441), .ZN(n5836) );
  XNOR2_X1 U4965 ( .A(n5837), .B(n5836), .ZN(n4444) );
  NOR2_X1 U4966 ( .A1(n4444), .A2(n4443), .ZN(n4445) );
  AOI211_X1 U4967 ( .C1(n5874), .C2(EAX_REG_28__SCAN_IN), .A(n4446), .B(n4445), 
        .ZN(n4447) );
  AOI21_X1 U4968 ( .B1(n3426), .B2(n6013), .A(n4447), .ZN(n4449) );
  NOR2_X1 U4969 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6443), .ZN(n5184) );
  NAND2_X1 U4970 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5184), .ZN(n6824) );
  NAND2_X1 U4971 ( .A1(n4454), .A2(n5390), .ZN(n6832) );
  NAND2_X1 U4972 ( .A1(n6832), .A2(n7159), .ZN(n4450) );
  NAND2_X1 U4973 ( .A1(n7159), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4452) );
  INV_X1 U4974 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6463) );
  NAND2_X1 U4975 ( .A1(n6463), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4451) );
  AND2_X1 U4976 ( .A1(n4452), .A2(n4451), .ZN(n4588) );
  INV_X1 U4977 ( .A(n4588), .ZN(n4453) );
  INV_X1 U4978 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U4979 ( .A1(n6912), .A2(n6537), .ZN(n6312) );
  NOR2_X1 U4980 ( .A1(n6287), .A2(n4455), .ZN(n4456) );
  AOI211_X1 U4981 ( .C1(n6805), .C2(n6013), .A(n6312), .B(n4456), .ZN(n4457)
         );
  NAND2_X1 U4982 ( .A1(n4460), .A2(n4459), .ZN(U2958) );
  INV_X1 U4983 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U4984 ( .A1(n7170), .A2(n7177), .ZN(n6821) );
  NAND2_X1 U4985 ( .A1(n3675), .A2(n6821), .ZN(n5191) );
  NAND2_X1 U4986 ( .A1(n5191), .A2(n7176), .ZN(n4461) );
  OR2_X1 U4987 ( .A1(n5985), .A2(n4461), .ZN(n4534) );
  INV_X1 U4988 ( .A(n4462), .ZN(n4482) );
  NOR2_X1 U4989 ( .A1(n4551), .A2(n4488), .ZN(n4480) );
  NAND2_X1 U4990 ( .A1(n4463), .A2(n4528), .ZN(n4464) );
  NAND2_X1 U4991 ( .A1(n4465), .A2(n4464), .ZN(n4508) );
  OR2_X1 U4992 ( .A1(n4466), .A2(n5979), .ZN(n4467) );
  AND2_X1 U4993 ( .A1(n4468), .A2(n4467), .ZN(n4496) );
  INV_X1 U4994 ( .A(n4519), .ZN(n5988) );
  OAI21_X1 U4995 ( .B1(n4508), .B2(n4496), .A(n5988), .ZN(n4529) );
  NAND2_X1 U4996 ( .A1(n4680), .A2(n6821), .ZN(n4477) );
  NOR3_X1 U4997 ( .A1(n4471), .A2(n4470), .A3(n4469), .ZN(n4472) );
  OR2_X1 U4998 ( .A1(n4473), .A2(n4472), .ZN(n4475) );
  NAND2_X1 U4999 ( .A1(n4475), .A2(n4474), .ZN(n5989) );
  NAND2_X1 U5000 ( .A1(n7176), .A2(n5989), .ZN(n4527) );
  INV_X1 U5001 ( .A(n4527), .ZN(n4476) );
  NAND3_X1 U5002 ( .A1(n4477), .A2(n4675), .A3(n4476), .ZN(n4478) );
  NAND2_X1 U5003 ( .A1(n4529), .A2(n4478), .ZN(n4479) );
  AOI21_X1 U5004 ( .B1(n5985), .B2(n4480), .A(n4479), .ZN(n4481) );
  OAI21_X1 U5005 ( .B1(n4534), .B2(n4482), .A(n4481), .ZN(n4483) );
  NAND2_X1 U5006 ( .A1(n4483), .A2(n5993), .ZN(n4487) );
  AOI21_X1 U5007 ( .B1(n4003), .B2(n3677), .A(n4675), .ZN(n4484) );
  NAND2_X1 U5008 ( .A1(n4485), .A2(n4484), .ZN(n4486) );
  INV_X2 U5009 ( .A(n6912), .ZN(n6924) );
  OR2_X1 U5010 ( .A1(n4512), .A2(n6924), .ZN(n4808) );
  AND2_X1 U5011 ( .A1(n4519), .A2(n4680), .ZN(n7115) );
  NAND2_X1 U5012 ( .A1(n4512), .A2(n7115), .ZN(n5655) );
  INV_X1 U5013 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6442) );
  AOI21_X1 U5014 ( .B1(n4808), .B2(n5655), .A(n6442), .ZN(n4517) );
  NOR2_X1 U5015 ( .A1(n4551), .A2(n3752), .ZN(n4490) );
  NOR2_X1 U5016 ( .A1(n4488), .A2(n4528), .ZN(n4489) );
  INV_X1 U5017 ( .A(n4491), .ZN(n4494) );
  OAI211_X1 U5018 ( .C1(n3675), .C2(n4675), .A(n5892), .B(n4528), .ZN(n4492)
         );
  NAND2_X1 U5019 ( .A1(n4492), .A2(n3752), .ZN(n4493) );
  NAND2_X1 U5020 ( .A1(n4494), .A2(n4493), .ZN(n4495) );
  NOR2_X1 U5021 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  NAND2_X1 U5022 ( .A1(n4498), .A2(n4497), .ZN(n4539) );
  NOR2_X1 U5023 ( .A1(n4536), .A2(n3677), .ZN(n4499) );
  OR2_X1 U5024 ( .A1(n4539), .A2(n4499), .ZN(n4500) );
  NAND2_X1 U5025 ( .A1(n4512), .A2(n4500), .ZN(n4810) );
  AND2_X1 U5026 ( .A1(n6933), .A2(n4810), .ZN(n4806) );
  NOR2_X1 U5027 ( .A1(n4806), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4609)
         );
  NAND2_X1 U5028 ( .A1(n4462), .A2(n5979), .ZN(n7143) );
  OAI21_X1 U5029 ( .B1(n4505), .B2(n4652), .A(n7143), .ZN(n4501) );
  NAND2_X1 U5030 ( .A1(n4965), .A2(EBX_REG_0__SCAN_IN), .ZN(n4504) );
  OAI21_X1 U5031 ( .B1(n4502), .B2(EBX_REG_0__SCAN_IN), .A(n4504), .ZN(n4573)
         );
  OAI21_X1 U5032 ( .B1(n5949), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4573), 
        .ZN(n5200) );
  NAND2_X1 U5033 ( .A1(n6924), .A2(REIP_REG_0__SCAN_IN), .ZN(n4589) );
  OAI21_X1 U5034 ( .B1(n6915), .B2(n5200), .A(n4589), .ZN(n4516) );
  OAI21_X1 U5035 ( .B1(n4505), .B2(n3688), .A(n5145), .ZN(n4506) );
  AOI21_X1 U5036 ( .B1(n4462), .B2(n5816), .A(n4506), .ZN(n4510) );
  INV_X1 U5037 ( .A(n4507), .ZN(n5190) );
  INV_X1 U5038 ( .A(n7136), .ZN(n4509) );
  AND2_X1 U5039 ( .A1(n4541), .A2(n4509), .ZN(n5983) );
  NAND2_X1 U5040 ( .A1(n4510), .A2(n5983), .ZN(n4511) );
  INV_X1 U5041 ( .A(n4606), .ZN(n4513) );
  OAI21_X1 U5042 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4514), .A(n4513), 
        .ZN(n4594) );
  NOR2_X1 U5043 ( .A1(n6892), .A2(n4594), .ZN(n4515) );
  OR4_X1 U5044 ( .A1(n4517), .A2(n4609), .A3(n4516), .A4(n4515), .ZN(U3018) );
  NAND2_X1 U5045 ( .A1(n5989), .A2(n4519), .ZN(n4522) );
  AOI22_X1 U5046 ( .A1(n5985), .A2(n5190), .B1(n4518), .B2(n4522), .ZN(n5992)
         );
  AND2_X1 U5047 ( .A1(n5992), .A2(n5993), .ZN(n4521) );
  INV_X1 U5048 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6625) );
  NOR2_X1 U5049 ( .A1(n5390), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5050 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4523), .ZN(n4520) );
  OAI21_X1 U5051 ( .B1(n4521), .B2(n6625), .A(n4520), .ZN(U2790) );
  NOR2_X1 U5052 ( .A1(n4522), .A2(n7164), .ZN(n5181) );
  INV_X1 U5053 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4525) );
  INV_X1 U5054 ( .A(n5182), .ZN(n4524) );
  INV_X1 U5055 ( .A(n4523), .ZN(n5978) );
  OAI211_X1 U5056 ( .C1(n5181), .C2(n4525), .A(n4524), .B(n5978), .ZN(U2788)
         );
  NAND2_X1 U5057 ( .A1(n4518), .A2(n6821), .ZN(n4526) );
  OAI21_X1 U5058 ( .B1(n4462), .B2(n7115), .A(n4526), .ZN(n4533) );
  OAI22_X1 U5059 ( .A1(n5985), .A2(n4541), .B1(n4527), .B2(n5145), .ZN(n5167)
         );
  INV_X1 U5060 ( .A(n5167), .ZN(n4532) );
  NAND2_X1 U5061 ( .A1(n4528), .A2(n4680), .ZN(n5203) );
  NAND2_X1 U5062 ( .A1(n5985), .A2(n4540), .ZN(n4560) );
  OAI211_X1 U5063 ( .C1(n4675), .C2(n5203), .A(n4560), .B(n4529), .ZN(n4530)
         );
  INV_X1 U5064 ( .A(n4530), .ZN(n4531) );
  NOR2_X1 U5065 ( .A1(n6823), .A2(n6443), .ZN(n5925) );
  NAND2_X1 U5066 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5925), .ZN(n7151) );
  INV_X1 U5067 ( .A(n7151), .ZN(n7156) );
  AOI22_X1 U5068 ( .A1(n7119), .A2(n5993), .B1(n7156), .B2(FLUSH_REG_SCAN_IN), 
        .ZN(n7110) );
  OAI21_X1 U5069 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n5471), .A(n7110), .ZN(
        n7114) );
  INV_X1 U5070 ( .A(n7114), .ZN(n5971) );
  NOR2_X1 U5071 ( .A1(n4535), .A2(n7160), .ZN(n6447) );
  NOR2_X1 U5072 ( .A1(n5971), .A2(n6447), .ZN(n5968) );
  INV_X1 U5073 ( .A(n5165), .ZN(n4537) );
  NAND3_X1 U5074 ( .A1(n4537), .A2(n4536), .A3(n5145), .ZN(n4538) );
  OR3_X1 U5075 ( .A1(n4539), .A2(n4462), .A3(n4538), .ZN(n6440) );
  NAND2_X1 U5076 ( .A1(n3429), .A2(n6440), .ZN(n4547) );
  INV_X1 U5077 ( .A(n4540), .ZN(n5982) );
  AND2_X1 U5078 ( .A1(n4541), .A2(n5982), .ZN(n5132) );
  NOR2_X1 U5079 ( .A1(n4535), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5131)
         );
  AND2_X1 U5080 ( .A1(n4535), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4542)
         );
  NOR2_X1 U5081 ( .A1(n5131), .A2(n4542), .ZN(n4544) );
  XNOR2_X1 U5082 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4543) );
  OAI22_X1 U5083 ( .A1(n5132), .A2(n4544), .B1(n6438), .B2(n4543), .ZN(n4545)
         );
  INV_X1 U5084 ( .A(n4545), .ZN(n4546) );
  NAND2_X1 U5085 ( .A1(n4547), .A2(n4546), .ZN(n5125) );
  INV_X1 U5086 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6295) );
  INV_X1 U5087 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U5088 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6295), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6876), .ZN(n6445) );
  NOR3_X1 U5089 ( .A1(n6443), .A2(n6442), .A3(n6445), .ZN(n4549) );
  INV_X1 U5090 ( .A(n4535), .ZN(n6435) );
  NOR3_X1 U5091 ( .A1(n6435), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n7160), 
        .ZN(n4548) );
  AOI211_X1 U5092 ( .C1(n5125), .C2(n6441), .A(n4549), .B(n4548), .ZN(n4550)
         );
  OAI22_X1 U5093 ( .A1(n5968), .A2(n3449), .B1(n5971), .B2(n4550), .ZN(U3459)
         );
  AOI21_X1 U5094 ( .B1(n7115), .B2(n6441), .A(n5971), .ZN(n4554) );
  INV_X1 U5095 ( .A(n6440), .ZN(n5134) );
  OAI22_X1 U5096 ( .A1(n5934), .A2(n5134), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4551), .ZN(n7118) );
  OAI22_X1 U5097 ( .A1(n6443), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7160), .ZN(n4552) );
  AOI21_X1 U5098 ( .B1(n7118), .B2(n6441), .A(n4552), .ZN(n4553) );
  OAI22_X1 U5099 ( .A1(n4554), .A2(n3513), .B1(n5971), .B2(n4553), .ZN(U3461)
         );
  OR2_X1 U5100 ( .A1(n4556), .A2(n4555), .ZN(n4557) );
  AND2_X1 U5101 ( .A1(n4595), .A2(n4557), .ZN(n6948) );
  INV_X1 U5102 ( .A(n6948), .ZN(n5173) );
  AND3_X1 U5103 ( .A1(n3688), .A2(n5974), .A3(n4662), .ZN(n5164) );
  NAND3_X1 U5104 ( .A1(n4558), .A2(n5816), .A3(n5164), .ZN(n4559) );
  NAND2_X1 U5105 ( .A1(n4560), .A2(n4559), .ZN(n4561) );
  INV_X1 U5106 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4566) );
  OAI21_X1 U5107 ( .B1(n4502), .B2(n6876), .A(n4965), .ZN(n4562) );
  NAND2_X1 U5108 ( .A1(n4502), .A2(n4566), .ZN(n4563) );
  XNOR2_X1 U5109 ( .A(n4572), .B(n4573), .ZN(n4564) );
  NAND2_X1 U5110 ( .A1(n4564), .A2(n5816), .ZN(n4576) );
  OR2_X1 U5111 ( .A1(n4564), .A2(n5816), .ZN(n4565) );
  NAND2_X1 U5112 ( .A1(n4576), .A2(n4565), .ZN(n4610) );
  INV_X1 U5113 ( .A(n4610), .ZN(n6943) );
  OAI222_X1 U5114 ( .A1(n5173), .A2(n6777), .B1(n4566), .B2(n6785), .C1(n6776), 
        .C2(n6943), .ZN(U2858) );
  INV_X1 U5115 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5201) );
  XNOR2_X1 U5116 ( .A(n4568), .B(n4567), .ZN(n5211) );
  OAI222_X1 U5117 ( .A1(n5200), .A2(n6776), .B1(n5201), .B2(n6785), .C1(n6777), 
        .C2(n5211), .ZN(U2859) );
  NOR2_X1 U5118 ( .A1(n4599), .A2(n4570), .ZN(n4571) );
  OR2_X1 U5119 ( .A1(n4569), .A2(n4571), .ZN(n5172) );
  INV_X1 U5120 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4587) );
  INV_X1 U5121 ( .A(n4572), .ZN(n4574) );
  NAND2_X1 U5122 ( .A1(n4574), .A2(n4573), .ZN(n4575) );
  INV_X1 U5123 ( .A(n4601), .ZN(n4582) );
  NAND2_X1 U5124 ( .A1(n4965), .A2(n3803), .ZN(n4578) );
  INV_X1 U5125 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U5126 ( .A1(n5816), .A2(n6963), .ZN(n4577) );
  NAND3_X1 U5127 ( .A1(n4578), .A2(n5805), .A3(n4577), .ZN(n4580) );
  NAND2_X1 U5128 ( .A1(n4502), .A2(n6963), .ZN(n4579) );
  AND2_X1 U5129 ( .A1(n4580), .A2(n4579), .ZN(n4600) );
  MUX2_X1 U5130 ( .A(n5795), .B(n5805), .S(EBX_REG_3__SCAN_IN), .Z(n4584) );
  NAND2_X1 U5131 ( .A1(n5796), .A2(n3839), .ZN(n4583) );
  NAND2_X1 U5132 ( .A1(n4584), .A2(n4583), .ZN(n4585) );
  AND2_X1 U5133 ( .A1(n4603), .A2(n4585), .ZN(n4586) );
  OR2_X1 U5134 ( .A1(n4631), .A2(n4586), .ZN(n6973) );
  OAI222_X1 U5135 ( .A1(n5172), .A2(n6777), .B1(n4587), .B2(n6785), .C1(n6776), 
        .C2(n6973), .ZN(U2856) );
  NAND2_X1 U5136 ( .A1(n4588), .A2(n6287), .ZN(n4592) );
  INV_X1 U5137 ( .A(n4589), .ZN(n4591) );
  NOR2_X1 U5138 ( .A1(n5211), .A2(n6291), .ZN(n4590) );
  AOI211_X1 U5139 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4592), .A(n4591), 
        .B(n4590), .ZN(n4593) );
  OAI21_X1 U5140 ( .B1(n7108), .B2(n4594), .A(n4593), .ZN(U2986) );
  AND3_X1 U5141 ( .A1(n4597), .A2(n4596), .A3(n4595), .ZN(n4598) );
  NOR2_X1 U5142 ( .A1(n4599), .A2(n4598), .ZN(n6960) );
  INV_X1 U5143 ( .A(n6960), .ZN(n5176) );
  NAND2_X1 U5144 ( .A1(n4601), .A2(n4600), .ZN(n4602) );
  AND2_X1 U5145 ( .A1(n4603), .A2(n4602), .ZN(n6956) );
  AOI22_X1 U5146 ( .A1(n6782), .A2(n6956), .B1(EBX_REG_2__SCAN_IN), .B2(n6159), 
        .ZN(n4604) );
  OAI21_X1 U5147 ( .B1(n5176), .B2(n6777), .A(n4604), .ZN(U2857) );
  INV_X1 U5148 ( .A(n6933), .ZN(n6886) );
  NAND2_X1 U5149 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6886), .ZN(n6872)
         );
  AOI21_X1 U5150 ( .B1(n6877), .B2(n6872), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4614) );
  XNOR2_X1 U5151 ( .A(n4606), .B(n6876), .ZN(n4607) );
  XNOR2_X1 U5152 ( .A(n3431), .B(n4607), .ZN(n6787) );
  INV_X1 U5153 ( .A(n4808), .ZN(n4608) );
  OAI21_X1 U5154 ( .B1(n4609), .B2(n4608), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4612) );
  AOI22_X1 U5155 ( .A1(n6932), .A2(n4610), .B1(n6924), .B2(REIP_REG_1__SCAN_IN), .ZN(n4611) );
  OAI211_X1 U5156 ( .C1(n6787), .C2(n6892), .A(n4612), .B(n4611), .ZN(n4613)
         );
  OR2_X1 U5157 ( .A1(n4614), .A2(n4613), .ZN(U3017) );
  NAND2_X1 U5158 ( .A1(n5093), .A2(DATAI_5_), .ZN(n5117) );
  AOI22_X1 U5159 ( .A1(n5162), .A2(EAX_REG_21__SCAN_IN), .B1(n5082), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5160 ( .A1(n5117), .A2(n4616), .ZN(U2929) );
  NAND2_X1 U5161 ( .A1(n5093), .A2(DATAI_4_), .ZN(n5119) );
  AOI22_X1 U5162 ( .A1(n5162), .A2(EAX_REG_20__SCAN_IN), .B1(n5082), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U5163 ( .A1(n5119), .A2(n4617), .ZN(U2928) );
  NAND2_X1 U5164 ( .A1(n5093), .A2(DATAI_7_), .ZN(n5113) );
  AOI22_X1 U5165 ( .A1(n5105), .A2(EAX_REG_23__SCAN_IN), .B1(n5082), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5166 ( .A1(n5113), .A2(n4618), .ZN(U2931) );
  NAND2_X1 U5167 ( .A1(n5093), .A2(DATAI_8_), .ZN(n5111) );
  AOI22_X1 U5168 ( .A1(n5162), .A2(EAX_REG_24__SCAN_IN), .B1(n5082), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5169 ( .A1(n5111), .A2(n4619), .ZN(U2932) );
  NAND2_X1 U5170 ( .A1(n5093), .A2(DATAI_6_), .ZN(n5098) );
  AOI22_X1 U5171 ( .A1(n5162), .A2(EAX_REG_22__SCAN_IN), .B1(n5082), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5172 ( .A1(n5098), .A2(n4620), .ZN(U2930) );
  INV_X1 U5173 ( .A(DATAI_9_), .ZN(n5460) );
  OR2_X1 U5174 ( .A1(n5169), .A2(n5460), .ZN(n5109) );
  AOI22_X1 U5175 ( .A1(n5162), .A2(EAX_REG_25__SCAN_IN), .B1(n5082), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5176 ( .A1(n5109), .A2(n4621), .ZN(U2933) );
  OR2_X1 U5177 ( .A1(n4569), .A2(n4622), .ZN(n4624) );
  AND2_X1 U5178 ( .A1(n4624), .A2(n4623), .ZN(n6993) );
  INV_X1 U5179 ( .A(n6993), .ZN(n5177) );
  INV_X1 U5180 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U5181 ( .A1(n4965), .A2(n4807), .ZN(n4626) );
  INV_X1 U5182 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5183 ( .A1(n5816), .A2(n4627), .ZN(n4625) );
  NAND3_X1 U5184 ( .A1(n4626), .A2(n5805), .A3(n4625), .ZN(n4629) );
  NAND2_X1 U5185 ( .A1(n5819), .A2(n4627), .ZN(n4628) );
  NAND2_X1 U5186 ( .A1(n4629), .A2(n4628), .ZN(n4630) );
  NAND2_X1 U5187 ( .A1(n4631), .A2(n4630), .ZN(n4735) );
  OR2_X1 U5188 ( .A1(n4631), .A2(n4630), .ZN(n4632) );
  AND2_X1 U5189 ( .A1(n4735), .A2(n4632), .ZN(n6986) );
  AOI22_X1 U5190 ( .A1(n6782), .A2(n6986), .B1(EBX_REG_4__SCAN_IN), .B2(n6159), 
        .ZN(n4633) );
  OAI21_X1 U5191 ( .B1(n5177), .B2(n6777), .A(n4633), .ZN(U2855) );
  NAND3_X1 U5192 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4745) );
  NOR2_X1 U5193 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4745), .ZN(n4682)
         );
  INV_X1 U5194 ( .A(n4682), .ZN(n4635) );
  OR2_X1 U5195 ( .A1(n5232), .A2(n7128), .ZN(n5392) );
  AND2_X1 U5196 ( .A1(n5392), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5396) );
  NOR2_X1 U5197 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5183) );
  INV_X1 U5198 ( .A(n4646), .ZN(n4634) );
  NAND2_X1 U5199 ( .A1(n4634), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U5200 ( .A1(n5148), .A2(n5477), .ZN(n5348) );
  AOI211_X1 U5201 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4635), .A(n5396), .B(
        n5348), .ZN(n4643) );
  OR2_X1 U5202 ( .A1(n4636), .A2(n5390), .ZN(n5480) );
  INV_X1 U5203 ( .A(n5480), .ZN(n5353) );
  NAND2_X1 U5204 ( .A1(n3429), .A2(n4638), .ZN(n4896) );
  INV_X1 U5205 ( .A(n4896), .ZN(n5269) );
  NOR2_X1 U5206 ( .A1(n5269), .A2(n5390), .ZN(n4889) );
  NOR3_X1 U5207 ( .A1(n4934), .A2(n4933), .A3(n4018), .ZN(n4640) );
  NAND3_X1 U5208 ( .A1(n4863), .A2(n3829), .A3(n4012), .ZN(n4744) );
  NOR2_X2 U5209 ( .A1(n4744), .A2(n5931), .ZN(n4769) );
  OAI21_X1 U5210 ( .B1(n4951), .B2(n4769), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4641) );
  OAI21_X1 U5211 ( .B1(n5353), .B2(n4889), .A(n4641), .ZN(n4642) );
  INV_X1 U5212 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4650) );
  INV_X1 U5213 ( .A(DATAI_27_), .ZN(n4645) );
  NOR2_X2 U5214 ( .A1(n4740), .A2(n4645), .ZN(n5484) );
  INV_X1 U5215 ( .A(DATAI_3_), .ZN(n6606) );
  NOR2_X2 U5216 ( .A1(n6606), .A2(n4738), .ZN(n5481) );
  INV_X1 U5217 ( .A(n5390), .ZN(n5282) );
  AND2_X1 U5218 ( .A1(n4636), .A2(n5282), .ZN(n4890) );
  INV_X1 U5219 ( .A(n4890), .ZN(n5359) );
  NAND2_X1 U5220 ( .A1(n4646), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5357) );
  OAI22_X1 U5221 ( .A1(n5359), .A2(n4896), .B1(n5357), .B2(n5392), .ZN(n4679)
         );
  AOI22_X1 U5222 ( .A1(n4951), .A2(n5484), .B1(n5481), .B2(n4679), .ZN(n4649)
         );
  NAND2_X1 U5223 ( .A1(n4681), .A2(n3671), .ZN(n5332) );
  INV_X1 U5224 ( .A(DATAI_19_), .ZN(n6555) );
  NOR2_X1 U5225 ( .A1(n4740), .A2(n6555), .ZN(n5483) );
  AOI22_X1 U5226 ( .A1(n5482), .A2(n4682), .B1(n5483), .B2(n4769), .ZN(n4648)
         );
  OAI211_X1 U5227 ( .C1(n4686), .C2(n4650), .A(n4649), .B(n4648), .ZN(U3135)
         );
  INV_X1 U5228 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4655) );
  INV_X1 U5229 ( .A(DATAI_28_), .ZN(n4651) );
  NOR2_X2 U5230 ( .A1(n4740), .A2(n4651), .ZN(n5526) );
  INV_X1 U5231 ( .A(DATAI_4_), .ZN(n6503) );
  NOR2_X2 U5232 ( .A1(n6503), .A2(n4738), .ZN(n5523) );
  AOI22_X1 U5233 ( .A1(n4951), .A2(n5526), .B1(n5523), .B2(n4679), .ZN(n4654)
         );
  NAND2_X1 U5234 ( .A1(n4681), .A2(n4652), .ZN(n5304) );
  INV_X1 U5235 ( .A(DATAI_20_), .ZN(n6573) );
  NOR2_X1 U5236 ( .A1(n4740), .A2(n6573), .ZN(n5525) );
  AOI22_X1 U5237 ( .A1(n5524), .A2(n4682), .B1(n5525), .B2(n4769), .ZN(n4653)
         );
  OAI211_X1 U5238 ( .C1(n4686), .C2(n4655), .A(n4654), .B(n4653), .ZN(U3136)
         );
  INV_X1 U5239 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4660) );
  INV_X1 U5240 ( .A(DATAI_29_), .ZN(n4656) );
  NOR2_X2 U5241 ( .A1(n4740), .A2(n4656), .ZN(n5519) );
  INV_X1 U5242 ( .A(DATAI_5_), .ZN(n5174) );
  NOR2_X2 U5243 ( .A1(n5174), .A2(n4738), .ZN(n5516) );
  AOI22_X1 U5244 ( .A1(n4951), .A2(n5519), .B1(n5516), .B2(n4679), .ZN(n4659)
         );
  NAND2_X1 U5245 ( .A1(n4681), .A2(n3655), .ZN(n5316) );
  INV_X1 U5246 ( .A(DATAI_21_), .ZN(n4657) );
  NOR2_X1 U5247 ( .A1(n4740), .A2(n4657), .ZN(n5518) );
  AOI22_X1 U5248 ( .A1(n5517), .A2(n4682), .B1(n5518), .B2(n4769), .ZN(n4658)
         );
  OAI211_X1 U5249 ( .C1(n4686), .C2(n4660), .A(n4659), .B(n4658), .ZN(U3137)
         );
  INV_X1 U5250 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4665) );
  INV_X1 U5251 ( .A(DATAI_30_), .ZN(n4661) );
  NOR2_X2 U5252 ( .A1(n4740), .A2(n4661), .ZN(n5512) );
  INV_X1 U5253 ( .A(DATAI_6_), .ZN(n6500) );
  NOR2_X2 U5254 ( .A1(n6500), .A2(n4738), .ZN(n5509) );
  AOI22_X1 U5255 ( .A1(n4951), .A2(n5512), .B1(n5509), .B2(n4679), .ZN(n4664)
         );
  NAND2_X1 U5256 ( .A1(n4681), .A2(n4662), .ZN(n5322) );
  INV_X1 U5257 ( .A(DATAI_22_), .ZN(n6565) );
  NOR2_X1 U5258 ( .A1(n6291), .A2(n6565), .ZN(n5511) );
  AOI22_X1 U5259 ( .A1(n5510), .A2(n4682), .B1(n5511), .B2(n4769), .ZN(n4663)
         );
  OAI211_X1 U5260 ( .C1(n4686), .C2(n4665), .A(n4664), .B(n4663), .ZN(U3138)
         );
  INV_X1 U5261 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4669) );
  INV_X1 U5262 ( .A(DATAI_24_), .ZN(n4666) );
  NOR2_X2 U5263 ( .A1(n6291), .A2(n4666), .ZN(n5498) );
  INV_X1 U5264 ( .A(DATAI_0_), .ZN(n6511) );
  NOR2_X2 U5265 ( .A1(n6511), .A2(n4738), .ZN(n5495) );
  AOI22_X1 U5266 ( .A1(n4951), .A2(n5498), .B1(n5495), .B2(n4679), .ZN(n4668)
         );
  NAND2_X1 U5267 ( .A1(n4681), .A2(n3427), .ZN(n5278) );
  NOR2_X1 U5268 ( .A1(n4740), .A2(n6582), .ZN(n5497) );
  AOI22_X1 U5269 ( .A1(n5496), .A2(n4682), .B1(n5497), .B2(n4769), .ZN(n4667)
         );
  OAI211_X1 U5270 ( .C1(n4686), .C2(n4669), .A(n4668), .B(n4667), .ZN(U3132)
         );
  INV_X1 U5271 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4673) );
  INV_X1 U5272 ( .A(DATAI_31_), .ZN(n4670) );
  NOR2_X2 U5273 ( .A1(n4740), .A2(n4670), .ZN(n5505) );
  INV_X1 U5274 ( .A(DATAI_7_), .ZN(n6596) );
  NOR2_X2 U5275 ( .A1(n6596), .A2(n4738), .ZN(n5502) );
  AOI22_X1 U5276 ( .A1(n4951), .A2(n5505), .B1(n5502), .B2(n4679), .ZN(n4672)
         );
  NAND2_X1 U5277 ( .A1(n4681), .A2(n4006), .ZN(n5301) );
  INV_X1 U5278 ( .A(DATAI_23_), .ZN(n6566) );
  NOR2_X1 U5279 ( .A1(n4740), .A2(n6566), .ZN(n5504) );
  AOI22_X1 U5280 ( .A1(n5503), .A2(n4682), .B1(n5504), .B2(n4769), .ZN(n4671)
         );
  OAI211_X1 U5281 ( .C1(n4686), .C2(n4673), .A(n4672), .B(n4671), .ZN(U3139)
         );
  INV_X1 U5282 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4678) );
  INV_X1 U5283 ( .A(DATAI_26_), .ZN(n4674) );
  NOR2_X2 U5284 ( .A1(n4740), .A2(n4674), .ZN(n5536) );
  INV_X1 U5285 ( .A(DATAI_2_), .ZN(n6605) );
  NOR2_X2 U5286 ( .A1(n6605), .A2(n4738), .ZN(n5531) );
  AOI22_X1 U5287 ( .A1(n4951), .A2(n5536), .B1(n5531), .B2(n4679), .ZN(n4677)
         );
  NAND2_X1 U5288 ( .A1(n4681), .A2(n4675), .ZN(n5325) );
  NOR2_X1 U5289 ( .A1(n4740), .A2(n6575), .ZN(n5534) );
  AOI22_X1 U5290 ( .A1(n5533), .A2(n4682), .B1(n5534), .B2(n4769), .ZN(n4676)
         );
  OAI211_X1 U5291 ( .C1(n4686), .C2(n4678), .A(n4677), .B(n4676), .ZN(U3134)
         );
  INV_X1 U5292 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4685) );
  INV_X1 U5293 ( .A(DATAI_25_), .ZN(n6563) );
  NOR2_X2 U5294 ( .A1(n4740), .A2(n6563), .ZN(n5491) );
  INV_X1 U5295 ( .A(DATAI_1_), .ZN(n6614) );
  NOR2_X2 U5296 ( .A1(n6614), .A2(n4738), .ZN(n5488) );
  AOI22_X1 U5297 ( .A1(n4951), .A2(n5491), .B1(n5488), .B2(n4679), .ZN(n4684)
         );
  NAND2_X1 U5298 ( .A1(n4681), .A2(n4680), .ZN(n5319) );
  NOR2_X1 U5299 ( .A1(n6291), .A2(n6579), .ZN(n5490) );
  AOI22_X1 U5300 ( .A1(n5489), .A2(n4682), .B1(n5490), .B2(n4769), .ZN(n4683)
         );
  OAI211_X1 U5301 ( .C1(n4686), .C2(n4685), .A(n4684), .B(n4683), .ZN(U3133)
         );
  NAND3_X1 U5302 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7128), .A3(n7124), .ZN(n4831) );
  NOR2_X1 U5303 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4831), .ZN(n4723)
         );
  INV_X1 U5304 ( .A(n4723), .ZN(n4688) );
  INV_X1 U5305 ( .A(n5233), .ZN(n4687) );
  NAND2_X1 U5306 ( .A1(n4687), .A2(n5232), .ZN(n5053) );
  AND2_X1 U5307 ( .A1(n5053), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5051) );
  AOI211_X1 U5308 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4688), .A(n5051), .B(
        n5348), .ZN(n4693) );
  INV_X1 U5309 ( .A(n4638), .ZN(n6944) );
  AND2_X1 U5310 ( .A1(n3429), .A2(n6944), .ZN(n4927) );
  NOR2_X1 U5311 ( .A1(n4927), .A2(n5390), .ZN(n5352) );
  INV_X1 U5312 ( .A(n4861), .ZN(n4690) );
  INV_X1 U5313 ( .A(n5045), .ZN(n4689) );
  OAI21_X1 U5314 ( .B1(n4690), .B2(n4689), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4691) );
  OAI21_X1 U5315 ( .B1(n4890), .B2(n5352), .A(n4691), .ZN(n4692) );
  INV_X1 U5316 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4697) );
  INV_X1 U5317 ( .A(n4927), .ZN(n5358) );
  OAI22_X1 U5318 ( .A1(n5480), .A2(n5358), .B1(n5357), .B2(n5053), .ZN(n4722)
         );
  AOI22_X1 U5319 ( .A1(n5510), .A2(n4723), .B1(n5509), .B2(n4722), .ZN(n4696)
         );
  INV_X1 U5320 ( .A(n5511), .ZN(n5336) );
  INV_X1 U5321 ( .A(n5512), .ZN(n4855) );
  OAI22_X1 U5322 ( .A1(n4861), .A2(n5336), .B1(n5045), .B2(n4855), .ZN(n4694)
         );
  INV_X1 U5323 ( .A(n4694), .ZN(n4695) );
  OAI211_X1 U5324 ( .C1(n4728), .C2(n4697), .A(n4696), .B(n4695), .ZN(U3058)
         );
  INV_X1 U5325 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5326 ( .A1(n5517), .A2(n4723), .B1(n5516), .B2(n4722), .ZN(n4700)
         );
  INV_X1 U5327 ( .A(n5518), .ZN(n5298) );
  INV_X1 U5328 ( .A(n5519), .ZN(n4852) );
  OAI22_X1 U5329 ( .A1(n4861), .A2(n5298), .B1(n5045), .B2(n4852), .ZN(n4698)
         );
  INV_X1 U5330 ( .A(n4698), .ZN(n4699) );
  OAI211_X1 U5331 ( .C1(n4728), .C2(n4701), .A(n4700), .B(n4699), .ZN(U3057)
         );
  INV_X1 U5332 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5333 ( .A1(n5524), .A2(n4723), .B1(n5523), .B2(n4722), .ZN(n4704)
         );
  INV_X1 U5334 ( .A(n5525), .ZN(n5295) );
  INV_X1 U5335 ( .A(n5526), .ZN(n4849) );
  OAI22_X1 U5336 ( .A1(n4861), .A2(n5295), .B1(n5045), .B2(n4849), .ZN(n4702)
         );
  INV_X1 U5337 ( .A(n4702), .ZN(n4703) );
  OAI211_X1 U5338 ( .C1(n4728), .C2(n4705), .A(n4704), .B(n4703), .ZN(U3056)
         );
  INV_X1 U5339 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5340 ( .A1(n5489), .A2(n4723), .B1(n5488), .B2(n4722), .ZN(n4708)
         );
  INV_X1 U5341 ( .A(n5490), .ZN(n5346) );
  INV_X1 U5342 ( .A(n5491), .ZN(n4837) );
  OAI22_X1 U5343 ( .A1(n4861), .A2(n5346), .B1(n5045), .B2(n4837), .ZN(n4706)
         );
  INV_X1 U5344 ( .A(n4706), .ZN(n4707) );
  OAI211_X1 U5345 ( .C1(n4728), .C2(n4709), .A(n4708), .B(n4707), .ZN(U3053)
         );
  INV_X1 U5346 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5347 ( .A1(n5496), .A2(n4723), .B1(n5495), .B2(n4722), .ZN(n4712)
         );
  INV_X1 U5348 ( .A(n5497), .ZN(n5313) );
  INV_X1 U5349 ( .A(n5498), .ZN(n4843) );
  OAI22_X1 U5350 ( .A1(n4861), .A2(n5313), .B1(n5045), .B2(n4843), .ZN(n4710)
         );
  INV_X1 U5351 ( .A(n4710), .ZN(n4711) );
  OAI211_X1 U5352 ( .C1(n4728), .C2(n4713), .A(n4712), .B(n4711), .ZN(U3052)
         );
  INV_X1 U5353 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5354 ( .A1(n5482), .A2(n4723), .B1(n5481), .B2(n4722), .ZN(n4716)
         );
  INV_X1 U5355 ( .A(n5483), .ZN(n5307) );
  INV_X1 U5356 ( .A(n5484), .ZN(n4846) );
  OAI22_X1 U5357 ( .A1(n4861), .A2(n5307), .B1(n5045), .B2(n4846), .ZN(n4714)
         );
  INV_X1 U5358 ( .A(n4714), .ZN(n4715) );
  OAI211_X1 U5359 ( .C1(n4728), .C2(n4717), .A(n4716), .B(n4715), .ZN(U3055)
         );
  INV_X1 U5360 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4721) );
  AOI22_X1 U5361 ( .A1(n5503), .A2(n4723), .B1(n5502), .B2(n4722), .ZN(n4720)
         );
  INV_X1 U5362 ( .A(n5504), .ZN(n5310) );
  INV_X1 U5363 ( .A(n5505), .ZN(n4862) );
  OAI22_X1 U5364 ( .A1(n4861), .A2(n5310), .B1(n5045), .B2(n4862), .ZN(n4718)
         );
  INV_X1 U5365 ( .A(n4718), .ZN(n4719) );
  OAI211_X1 U5366 ( .C1(n4728), .C2(n4721), .A(n4720), .B(n4719), .ZN(U3059)
         );
  INV_X1 U5367 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5368 ( .A1(n5533), .A2(n4723), .B1(n5531), .B2(n4722), .ZN(n4726)
         );
  INV_X1 U5369 ( .A(n5534), .ZN(n5339) );
  INV_X1 U5370 ( .A(n5536), .ZN(n4840) );
  OAI22_X1 U5371 ( .A1(n4861), .A2(n5339), .B1(n5045), .B2(n4840), .ZN(n4724)
         );
  INV_X1 U5372 ( .A(n4724), .ZN(n4725) );
  OAI211_X1 U5373 ( .C1(n4728), .C2(n4727), .A(n4726), .B(n4725), .ZN(U3054)
         );
  NOR2_X1 U5374 ( .A1(n4623), .A2(n4729), .ZN(n5213) );
  AOI21_X1 U5375 ( .B1(n4729), .B2(n4623), .A(n5213), .ZN(n7004) );
  INV_X1 U5376 ( .A(n7004), .ZN(n5175) );
  MUX2_X1 U5377 ( .A(n5795), .B(n5805), .S(EBX_REG_5__SCAN_IN), .Z(n4731) );
  NAND2_X1 U5378 ( .A1(n5796), .A2(n3886), .ZN(n4730) );
  NAND2_X1 U5379 ( .A1(n4731), .A2(n4730), .ZN(n4736) );
  INV_X1 U5380 ( .A(n4735), .ZN(n4733) );
  INV_X1 U5381 ( .A(n5217), .ZN(n4734) );
  AOI21_X1 U5382 ( .B1(n4736), .B2(n4735), .A(n4734), .ZN(n7000) );
  AOI22_X1 U5383 ( .A1(n6782), .A2(n7000), .B1(EBX_REG_5__SCAN_IN), .B2(n6159), 
        .ZN(n4737) );
  OAI21_X1 U5384 ( .B1(n5175), .B2(n6777), .A(n4737), .ZN(U2854) );
  INV_X1 U5385 ( .A(n4636), .ZN(n6972) );
  NOR2_X1 U5386 ( .A1(n6972), .A2(n5934), .ZN(n4928) );
  NOR2_X1 U5387 ( .A1(n4739), .A2(n7128), .ZN(n4770) );
  AOI21_X1 U5388 ( .B1(n4928), .B2(n5269), .A(n4770), .ZN(n4746) );
  INV_X1 U5389 ( .A(n4744), .ZN(n4741) );
  NAND2_X1 U5390 ( .A1(n5282), .A2(n6463), .ZN(n5468) );
  OAI21_X1 U5391 ( .B1(n4741), .B2(n4740), .A(n5468), .ZN(n4742) );
  AOI22_X1 U5392 ( .A1(n4746), .A2(n4742), .B1(n5390), .B2(n4745), .ZN(n4743)
         );
  INV_X1 U5393 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4749) );
  NOR2_X2 U5394 ( .A1(n4744), .A2(n4018), .ZN(n5076) );
  OAI22_X1 U5395 ( .A1(n4746), .A2(n5390), .B1(n4745), .B2(n6823), .ZN(n4768)
         );
  AOI22_X1 U5396 ( .A1(n5076), .A2(n5490), .B1(n5488), .B2(n4768), .ZN(n4748)
         );
  AOI22_X1 U5397 ( .A1(n5489), .A2(n4770), .B1(n5491), .B2(n4769), .ZN(n4747)
         );
  OAI211_X1 U5398 ( .C1(n4774), .C2(n4749), .A(n4748), .B(n4747), .ZN(U3141)
         );
  INV_X1 U5399 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4752) );
  AOI22_X1 U5400 ( .A1(n5076), .A2(n5483), .B1(n5481), .B2(n4768), .ZN(n4751)
         );
  AOI22_X1 U5401 ( .A1(n5482), .A2(n4770), .B1(n5484), .B2(n4769), .ZN(n4750)
         );
  OAI211_X1 U5402 ( .C1(n4774), .C2(n4752), .A(n4751), .B(n4750), .ZN(U3143)
         );
  INV_X1 U5403 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4755) );
  AOI22_X1 U5404 ( .A1(n5076), .A2(n5525), .B1(n5523), .B2(n4768), .ZN(n4754)
         );
  AOI22_X1 U5405 ( .A1(n5524), .A2(n4770), .B1(n5526), .B2(n4769), .ZN(n4753)
         );
  OAI211_X1 U5406 ( .C1(n4774), .C2(n4755), .A(n4754), .B(n4753), .ZN(U3144)
         );
  INV_X1 U5407 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4758) );
  AOI22_X1 U5408 ( .A1(n5076), .A2(n5504), .B1(n5502), .B2(n4768), .ZN(n4757)
         );
  AOI22_X1 U5409 ( .A1(n5503), .A2(n4770), .B1(n5505), .B2(n4769), .ZN(n4756)
         );
  OAI211_X1 U5410 ( .C1(n4774), .C2(n4758), .A(n4757), .B(n4756), .ZN(U3147)
         );
  INV_X1 U5411 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5412 ( .A1(n5076), .A2(n5497), .B1(n5495), .B2(n4768), .ZN(n4760)
         );
  AOI22_X1 U5413 ( .A1(n5496), .A2(n4770), .B1(n5498), .B2(n4769), .ZN(n4759)
         );
  OAI211_X1 U5414 ( .C1(n4774), .C2(n4761), .A(n4760), .B(n4759), .ZN(U3140)
         );
  INV_X1 U5415 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5416 ( .A1(n5076), .A2(n5534), .B1(n5531), .B2(n4768), .ZN(n4763)
         );
  AOI22_X1 U5417 ( .A1(n5533), .A2(n4770), .B1(n5536), .B2(n4769), .ZN(n4762)
         );
  OAI211_X1 U5418 ( .C1(n4774), .C2(n4764), .A(n4763), .B(n4762), .ZN(U3142)
         );
  INV_X1 U5419 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U5420 ( .A1(n5076), .A2(n5511), .B1(n5509), .B2(n4768), .ZN(n4766)
         );
  AOI22_X1 U5421 ( .A1(n5510), .A2(n4770), .B1(n5512), .B2(n4769), .ZN(n4765)
         );
  OAI211_X1 U5422 ( .C1(n4774), .C2(n4767), .A(n4766), .B(n4765), .ZN(U3146)
         );
  INV_X1 U5423 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4773) );
  AOI22_X1 U5424 ( .A1(n5076), .A2(n5518), .B1(n5516), .B2(n4768), .ZN(n4772)
         );
  AOI22_X1 U5425 ( .A1(n5517), .A2(n4770), .B1(n5519), .B2(n4769), .ZN(n4771)
         );
  OAI211_X1 U5426 ( .C1(n4774), .C2(n4773), .A(n4772), .B(n4771), .ZN(U3145)
         );
  INV_X1 U5427 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5428 ( .A1(n4775), .A2(n6438), .ZN(n4776) );
  INV_X1 U5429 ( .A(n6821), .ZN(n5990) );
  NAND2_X1 U5430 ( .A1(n6672), .A2(n3677), .ZN(n5603) );
  NAND2_X1 U5431 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5184), .ZN(n7141) );
  INV_X2 U5432 ( .A(n7141), .ZN(n6699) );
  NOR2_X4 U5433 ( .A1(n6699), .A2(n6672), .ZN(n6455) );
  AOI22_X1 U5434 ( .A1(n6699), .A2(UWORD_REG_4__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4778) );
  OAI21_X1 U5435 ( .B1(n4779), .B2(n5603), .A(n4778), .ZN(U2903) );
  INV_X1 U5436 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5437 ( .A1(n6699), .A2(UWORD_REG_12__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4780) );
  OAI21_X1 U5438 ( .B1(n4781), .B2(n5603), .A(n4780), .ZN(U2895) );
  INV_X1 U5439 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5440 ( .A1(n6699), .A2(UWORD_REG_5__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4782) );
  OAI21_X1 U5441 ( .B1(n4783), .B2(n5603), .A(n4782), .ZN(U2902) );
  INV_X1 U5442 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5443 ( .A1(n6699), .A2(UWORD_REG_6__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4784) );
  OAI21_X1 U5444 ( .B1(n4785), .B2(n5603), .A(n4784), .ZN(U2901) );
  INV_X1 U5445 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4787) );
  AOI22_X1 U5446 ( .A1(n6699), .A2(UWORD_REG_13__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4786) );
  OAI21_X1 U5447 ( .B1(n4787), .B2(n5603), .A(n4786), .ZN(U2894) );
  INV_X1 U5448 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5449 ( .A1(n6699), .A2(UWORD_REG_8__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4788) );
  OAI21_X1 U5450 ( .B1(n4789), .B2(n5603), .A(n4788), .ZN(U2899) );
  INV_X1 U5451 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5452 ( .A1(n6699), .A2(UWORD_REG_7__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4790) );
  OAI21_X1 U5453 ( .B1(n4791), .B2(n5603), .A(n4790), .ZN(U2900) );
  AOI22_X1 U5454 ( .A1(n6699), .A2(UWORD_REG_11__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4792) );
  OAI21_X1 U5455 ( .B1(n4417), .B2(n5603), .A(n4792), .ZN(U2896) );
  AOI22_X1 U5456 ( .A1(n6699), .A2(UWORD_REG_10__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4793) );
  OAI21_X1 U5457 ( .B1(n4394), .B2(n5603), .A(n4793), .ZN(U2897) );
  INV_X1 U5458 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5459 ( .A1(n6699), .A2(UWORD_REG_9__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4794) );
  OAI21_X1 U5460 ( .B1(n4795), .B2(n5603), .A(n4794), .ZN(U2898) );
  XNOR2_X1 U5461 ( .A(n4797), .B(n4796), .ZN(n6847) );
  INV_X1 U5462 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U5463 ( .A1(n6912), .A2(n6707), .ZN(n6844) );
  AOI21_X1 U5464 ( .B1(n6809), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6844), 
        .ZN(n4798) );
  OAI21_X1 U5465 ( .B1(n6996), .B2(n6815), .A(n4798), .ZN(n4799) );
  AOI21_X1 U5466 ( .B1(n4644), .B2(n6993), .A(n4799), .ZN(n4800) );
  OAI21_X1 U5467 ( .B1(n6847), .B2(n7108), .A(n4800), .ZN(U2982) );
  XNOR2_X1 U5468 ( .A(n4801), .B(n4802), .ZN(n4818) );
  AOI22_X1 U5469 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6924), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4803) );
  OAI21_X1 U5470 ( .B1(n7001), .B2(n6815), .A(n4803), .ZN(n4804) );
  AOI21_X1 U5471 ( .B1(n7004), .B2(n4644), .A(n4804), .ZN(n4805) );
  OAI21_X1 U5472 ( .B1(n7108), .B2(n4818), .A(n4805), .ZN(U2981) );
  NOR2_X1 U5473 ( .A1(n4807), .A2(n3839), .ZN(n6851) );
  OAI21_X1 U5474 ( .B1(n6876), .B2(n6442), .A(n3803), .ZN(n6852) );
  NOR2_X1 U5475 ( .A1(n6933), .A2(n6852), .ZN(n6873) );
  OR2_X1 U5476 ( .A1(n4810), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4809)
         );
  NAND2_X1 U5477 ( .A1(n4809), .A2(n4808), .ZN(n6887) );
  NAND2_X1 U5478 ( .A1(n5655), .A2(n4810), .ZN(n6890) );
  NOR2_X1 U5479 ( .A1(n3803), .A2(n6876), .ZN(n6875) );
  INV_X1 U5480 ( .A(n6875), .ZN(n6871) );
  AND2_X1 U5481 ( .A1(n6890), .A2(n6871), .ZN(n4811) );
  OR2_X1 U5482 ( .A1(n6887), .A2(n4811), .ZN(n4812) );
  OR2_X1 U5483 ( .A1(n6873), .A2(n4812), .ZN(n6843) );
  INV_X1 U5484 ( .A(n6843), .ZN(n6862) );
  OAI21_X1 U5485 ( .B1(n6417), .B2(n6851), .A(n6862), .ZN(n6864) );
  NAND2_X1 U5486 ( .A1(n6851), .A2(n6875), .ZN(n5652) );
  NOR3_X1 U5487 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6877), .A3(n5652), 
        .ZN(n6865) );
  INV_X1 U5488 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6997) );
  AND2_X1 U5489 ( .A1(n6852), .A2(n6851), .ZN(n6863) );
  INV_X1 U5490 ( .A(n6863), .ZN(n4813) );
  NOR3_X1 U5491 ( .A1(n6933), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4813), 
        .ZN(n4814) );
  AOI21_X1 U5492 ( .B1(n7000), .B2(n6932), .A(n4814), .ZN(n4815) );
  OAI21_X1 U5493 ( .B1(n6912), .B2(n6997), .A(n4815), .ZN(n4816) );
  AOI211_X1 U5494 ( .C1(INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n6864), .A(n6865), 
        .B(n4816), .ZN(n4817) );
  OAI21_X1 U5495 ( .B1(n6892), .B2(n4818), .A(n4817), .ZN(U3013) );
  NAND2_X1 U5496 ( .A1(n4819), .A2(n4820), .ZN(n4823) );
  INV_X1 U5497 ( .A(n4821), .ZN(n4822) );
  XNOR2_X1 U5498 ( .A(n4823), .B(n4822), .ZN(n6856) );
  INV_X1 U5499 ( .A(n6856), .ZN(n4827) );
  INV_X1 U5500 ( .A(n5172), .ZN(n6971) );
  AOI22_X1 U5501 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6924), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4824) );
  OAI21_X1 U5502 ( .B1(n6968), .B2(n6815), .A(n4824), .ZN(n4825) );
  AOI21_X1 U5503 ( .B1(n4644), .B2(n6971), .A(n4825), .ZN(n4826) );
  OAI21_X1 U5504 ( .B1(n4827), .B2(n7108), .A(n4826), .ZN(U2983) );
  NOR2_X1 U5505 ( .A1(n5927), .A2(n4831), .ZN(n4858) );
  AOI21_X1 U5506 ( .B1(n3448), .B2(n4927), .A(n4858), .ZN(n4833) );
  AOI21_X1 U5507 ( .B1(n4828), .B2(STATEBS16_REG_SCAN_IN), .A(n5390), .ZN(
        n4830) );
  AOI22_X1 U5508 ( .A1(n4833), .A2(n4830), .B1(n5390), .B2(n4831), .ZN(n4829)
         );
  NAND2_X1 U5509 ( .A1(n5266), .A2(n4829), .ZN(n4857) );
  INV_X1 U5510 ( .A(n4830), .ZN(n4832) );
  OAI22_X1 U5511 ( .A1(n4833), .A2(n4832), .B1(n6823), .B2(n4831), .ZN(n4856)
         );
  AOI22_X1 U5512 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4857), .B1(n5488), 
        .B2(n4856), .ZN(n4836) );
  AOI22_X1 U5513 ( .A1(n5489), .A2(n4858), .B1(n5490), .B2(n4919), .ZN(n4835)
         );
  OAI211_X1 U5514 ( .C1(n4837), .C2(n4861), .A(n4836), .B(n4835), .ZN(U3061)
         );
  AOI22_X1 U5515 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n4857), .B1(n5531), 
        .B2(n4856), .ZN(n4839) );
  AOI22_X1 U5516 ( .A1(n5533), .A2(n4858), .B1(n5534), .B2(n4919), .ZN(n4838)
         );
  OAI211_X1 U5517 ( .C1(n4840), .C2(n4861), .A(n4839), .B(n4838), .ZN(U3062)
         );
  AOI22_X1 U5518 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4857), .B1(n5495), 
        .B2(n4856), .ZN(n4842) );
  AOI22_X1 U5519 ( .A1(n5496), .A2(n4858), .B1(n5497), .B2(n4919), .ZN(n4841)
         );
  OAI211_X1 U5520 ( .C1(n4843), .C2(n4861), .A(n4842), .B(n4841), .ZN(U3060)
         );
  AOI22_X1 U5521 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n4857), .B1(n5481), 
        .B2(n4856), .ZN(n4845) );
  AOI22_X1 U5522 ( .A1(n5482), .A2(n4858), .B1(n5483), .B2(n4919), .ZN(n4844)
         );
  OAI211_X1 U5523 ( .C1(n4846), .C2(n4861), .A(n4845), .B(n4844), .ZN(U3063)
         );
  AOI22_X1 U5524 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4857), .B1(n5523), 
        .B2(n4856), .ZN(n4848) );
  AOI22_X1 U5525 ( .A1(n5524), .A2(n4858), .B1(n5525), .B2(n4919), .ZN(n4847)
         );
  OAI211_X1 U5526 ( .C1(n4849), .C2(n4861), .A(n4848), .B(n4847), .ZN(U3064)
         );
  AOI22_X1 U5527 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n4857), .B1(n5516), 
        .B2(n4856), .ZN(n4851) );
  AOI22_X1 U5528 ( .A1(n5517), .A2(n4858), .B1(n5518), .B2(n4919), .ZN(n4850)
         );
  OAI211_X1 U5529 ( .C1(n4852), .C2(n4861), .A(n4851), .B(n4850), .ZN(U3065)
         );
  AOI22_X1 U5530 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n4857), .B1(n5509), 
        .B2(n4856), .ZN(n4854) );
  AOI22_X1 U5531 ( .A1(n5510), .A2(n4858), .B1(n5511), .B2(n4919), .ZN(n4853)
         );
  OAI211_X1 U5532 ( .C1(n4855), .C2(n4861), .A(n4854), .B(n4853), .ZN(U3066)
         );
  AOI22_X1 U5533 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n4857), .B1(n5502), 
        .B2(n4856), .ZN(n4860) );
  AOI22_X1 U5534 ( .A1(n5503), .A2(n4858), .B1(n5504), .B2(n4919), .ZN(n4859)
         );
  OAI211_X1 U5535 ( .C1(n4862), .C2(n4861), .A(n4860), .B(n4859), .ZN(U3067)
         );
  OR2_X1 U5536 ( .A1(n3429), .A2(n4638), .ZN(n5237) );
  INV_X1 U5537 ( .A(n5237), .ZN(n5285) );
  NAND3_X1 U5538 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5224), .A3(n7124), .ZN(n5234) );
  NOR2_X1 U5539 ( .A1(n5927), .A2(n5234), .ZN(n4886) );
  AOI21_X1 U5540 ( .B1(n4928), .B2(n5285), .A(n4886), .ZN(n4867) );
  OR2_X1 U5541 ( .A1(n4012), .A2(n6463), .ZN(n5283) );
  INV_X1 U5542 ( .A(n5283), .ZN(n4864) );
  AOI21_X1 U5543 ( .B1(n4982), .B2(n4864), .A(n5390), .ZN(n4866) );
  AOI22_X1 U5544 ( .A1(n4867), .A2(n4866), .B1(n5390), .B2(n5234), .ZN(n4865)
         );
  NAND2_X1 U5545 ( .A1(n5266), .A2(n4865), .ZN(n4885) );
  INV_X1 U5546 ( .A(n4866), .ZN(n4868) );
  OAI22_X1 U5547 ( .A1(n4868), .A2(n4867), .B1(n6823), .B2(n5234), .ZN(n4884)
         );
  AOI22_X1 U5548 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4885), .B1(n5488), 
        .B2(n4884), .ZN(n4871) );
  INV_X1 U5549 ( .A(n4012), .ZN(n5150) );
  NAND3_X1 U5550 ( .A1(n5222), .A2(n5150), .A3(n4018), .ZN(n5046) );
  NOR2_X2 U5551 ( .A1(n5046), .A2(n4869), .ZN(n5260) );
  AOI22_X1 U5552 ( .A1(n5489), .A2(n4886), .B1(n5491), .B2(n5260), .ZN(n4870)
         );
  OAI211_X1 U5553 ( .C1(n5346), .C2(n5403), .A(n4871), .B(n4870), .ZN(U3093)
         );
  AOI22_X1 U5554 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4885), .B1(n5531), 
        .B2(n4884), .ZN(n4873) );
  AOI22_X1 U5555 ( .A1(n5533), .A2(n4886), .B1(n5536), .B2(n5260), .ZN(n4872)
         );
  OAI211_X1 U5556 ( .C1(n5339), .C2(n5403), .A(n4873), .B(n4872), .ZN(U3094)
         );
  AOI22_X1 U5557 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4885), .B1(n5481), 
        .B2(n4884), .ZN(n4875) );
  AOI22_X1 U5558 ( .A1(n5482), .A2(n4886), .B1(n5484), .B2(n5260), .ZN(n4874)
         );
  OAI211_X1 U5559 ( .C1(n5307), .C2(n5403), .A(n4875), .B(n4874), .ZN(U3095)
         );
  AOI22_X1 U5560 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4885), .B1(n5523), 
        .B2(n4884), .ZN(n4877) );
  AOI22_X1 U5561 ( .A1(n5524), .A2(n4886), .B1(n5526), .B2(n5260), .ZN(n4876)
         );
  OAI211_X1 U5562 ( .C1(n5295), .C2(n5403), .A(n4877), .B(n4876), .ZN(U3096)
         );
  AOI22_X1 U5563 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4885), .B1(n5516), 
        .B2(n4884), .ZN(n4879) );
  AOI22_X1 U5564 ( .A1(n5517), .A2(n4886), .B1(n5519), .B2(n5260), .ZN(n4878)
         );
  OAI211_X1 U5565 ( .C1(n5298), .C2(n5403), .A(n4879), .B(n4878), .ZN(U3097)
         );
  AOI22_X1 U5566 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4885), .B1(n5495), 
        .B2(n4884), .ZN(n4881) );
  AOI22_X1 U5567 ( .A1(n5496), .A2(n4886), .B1(n5498), .B2(n5260), .ZN(n4880)
         );
  OAI211_X1 U5568 ( .C1(n5313), .C2(n5403), .A(n4881), .B(n4880), .ZN(U3092)
         );
  AOI22_X1 U5569 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4885), .B1(n5509), 
        .B2(n4884), .ZN(n4883) );
  AOI22_X1 U5570 ( .A1(n5510), .A2(n4886), .B1(n5512), .B2(n5260), .ZN(n4882)
         );
  OAI211_X1 U5571 ( .C1(n5336), .C2(n5403), .A(n4883), .B(n4882), .ZN(U3098)
         );
  AOI22_X1 U5572 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4885), .B1(n5502), 
        .B2(n4884), .ZN(n4888) );
  AOI22_X1 U5573 ( .A1(n5503), .A2(n4886), .B1(n5505), .B2(n5260), .ZN(n4887)
         );
  OAI211_X1 U5574 ( .C1(n5310), .C2(n5403), .A(n4888), .B(n4887), .ZN(U3099)
         );
  NAND3_X1 U5575 ( .A1(n7128), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5273) );
  NOR2_X1 U5576 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5273), .ZN(n4920)
         );
  OAI21_X1 U5577 ( .B1(n4919), .B2(n5328), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4892) );
  OR2_X1 U5578 ( .A1(n4890), .A2(n4889), .ZN(n4891) );
  AOI21_X1 U5579 ( .B1(n4892), .B2(n4891), .A(n5348), .ZN(n4894) );
  INV_X1 U5580 ( .A(n5232), .ZN(n4893) );
  NAND2_X1 U5581 ( .A1(n4893), .A2(n7128), .ZN(n5478) );
  NAND2_X1 U5582 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5478), .ZN(n5473) );
  OAI211_X1 U5583 ( .C1(n4920), .C2(n5471), .A(n4894), .B(n5473), .ZN(n4895)
         );
  INV_X1 U5584 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4899) );
  OAI22_X1 U5585 ( .A1(n5480), .A2(n4896), .B1(n5478), .B2(n5357), .ZN(n4918)
         );
  AOI22_X1 U5586 ( .A1(n5328), .A2(n5518), .B1(n5516), .B2(n4918), .ZN(n4898)
         );
  AOI22_X1 U5587 ( .A1(n5517), .A2(n4920), .B1(n5519), .B2(n4919), .ZN(n4897)
         );
  OAI211_X1 U5588 ( .C1(n4924), .C2(n4899), .A(n4898), .B(n4897), .ZN(U3073)
         );
  INV_X1 U5589 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4902) );
  AOI22_X1 U5590 ( .A1(n5328), .A2(n5525), .B1(n5523), .B2(n4918), .ZN(n4901)
         );
  AOI22_X1 U5591 ( .A1(n5524), .A2(n4920), .B1(n5526), .B2(n4919), .ZN(n4900)
         );
  OAI211_X1 U5592 ( .C1(n4924), .C2(n4902), .A(n4901), .B(n4900), .ZN(U3072)
         );
  INV_X1 U5593 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4905) );
  AOI22_X1 U5594 ( .A1(n5328), .A2(n5483), .B1(n5481), .B2(n4918), .ZN(n4904)
         );
  AOI22_X1 U5595 ( .A1(n5482), .A2(n4920), .B1(n5484), .B2(n4919), .ZN(n4903)
         );
  OAI211_X1 U5596 ( .C1(n4924), .C2(n4905), .A(n4904), .B(n4903), .ZN(U3071)
         );
  INV_X1 U5597 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4908) );
  AOI22_X1 U5598 ( .A1(n5328), .A2(n5511), .B1(n5509), .B2(n4918), .ZN(n4907)
         );
  AOI22_X1 U5599 ( .A1(n5510), .A2(n4920), .B1(n5512), .B2(n4919), .ZN(n4906)
         );
  OAI211_X1 U5600 ( .C1(n4924), .C2(n4908), .A(n4907), .B(n4906), .ZN(U3074)
         );
  INV_X1 U5601 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U5602 ( .A1(n5328), .A2(n5504), .B1(n5502), .B2(n4918), .ZN(n4910)
         );
  AOI22_X1 U5603 ( .A1(n5503), .A2(n4920), .B1(n5505), .B2(n4919), .ZN(n4909)
         );
  OAI211_X1 U5604 ( .C1(n4924), .C2(n4911), .A(n4910), .B(n4909), .ZN(U3075)
         );
  INV_X1 U5605 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4914) );
  AOI22_X1 U5606 ( .A1(n5328), .A2(n5534), .B1(n5531), .B2(n4918), .ZN(n4913)
         );
  AOI22_X1 U5607 ( .A1(n5533), .A2(n4920), .B1(n5536), .B2(n4919), .ZN(n4912)
         );
  OAI211_X1 U5608 ( .C1(n4924), .C2(n4914), .A(n4913), .B(n4912), .ZN(U3070)
         );
  INV_X1 U5609 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4917) );
  AOI22_X1 U5610 ( .A1(n5328), .A2(n5490), .B1(n5488), .B2(n4918), .ZN(n4916)
         );
  AOI22_X1 U5611 ( .A1(n5489), .A2(n4920), .B1(n5491), .B2(n4919), .ZN(n4915)
         );
  OAI211_X1 U5612 ( .C1(n4924), .C2(n4917), .A(n4916), .B(n4915), .ZN(U3069)
         );
  INV_X1 U5613 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4923) );
  AOI22_X1 U5614 ( .A1(n5328), .A2(n5497), .B1(n5495), .B2(n4918), .ZN(n4922)
         );
  AOI22_X1 U5615 ( .A1(n5496), .A2(n4920), .B1(n5498), .B2(n4919), .ZN(n4921)
         );
  OAI211_X1 U5616 ( .C1(n4924), .C2(n4923), .A(n4922), .B(n4921), .ZN(U3068)
         );
  NAND3_X1 U5617 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n7124), .ZN(n5347) );
  NOR2_X1 U5618 ( .A1(n5927), .A2(n5347), .ZN(n4926) );
  INV_X1 U5619 ( .A(n4926), .ZN(n4954) );
  OR2_X1 U5620 ( .A1(n5222), .A2(n6463), .ZN(n5155) );
  OR2_X1 U5621 ( .A1(n4012), .A2(n4933), .ZN(n4925) );
  NOR2_X1 U5622 ( .A1(n5155), .A2(n4925), .ZN(n5153) );
  NOR2_X1 U5623 ( .A1(n5153), .A2(n5390), .ZN(n4930) );
  AOI21_X1 U5624 ( .B1(n4928), .B2(n4927), .A(n4926), .ZN(n4932) );
  AOI22_X1 U5625 ( .A1(n4930), .A2(n4932), .B1(n5390), .B2(n5347), .ZN(n4929)
         );
  NAND2_X1 U5626 ( .A1(n5266), .A2(n4929), .ZN(n4950) );
  INV_X1 U5627 ( .A(n4930), .ZN(n4931) );
  OAI22_X1 U5628 ( .A1(n4932), .A2(n4931), .B1(n6823), .B2(n5347), .ZN(n4949)
         );
  AOI22_X1 U5629 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4950), .B1(n5509), 
        .B2(n4949), .ZN(n4936) );
  NOR3_X4 U5630 ( .A1(n4934), .A2(n4933), .A3(n5931), .ZN(n5382) );
  AOI22_X1 U5631 ( .A1(n5511), .A2(n4951), .B1(n5382), .B2(n5512), .ZN(n4935)
         );
  OAI211_X1 U5632 ( .C1(n5322), .C2(n4954), .A(n4936), .B(n4935), .ZN(U3130)
         );
  AOI22_X1 U5633 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4950), .B1(n5502), 
        .B2(n4949), .ZN(n4938) );
  AOI22_X1 U5634 ( .A1(n5504), .A2(n4951), .B1(n5382), .B2(n5505), .ZN(n4937)
         );
  OAI211_X1 U5635 ( .C1(n5301), .C2(n4954), .A(n4938), .B(n4937), .ZN(U3131)
         );
  AOI22_X1 U5636 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4950), .B1(n5481), 
        .B2(n4949), .ZN(n4940) );
  AOI22_X1 U5637 ( .A1(n5483), .A2(n4951), .B1(n5382), .B2(n5484), .ZN(n4939)
         );
  OAI211_X1 U5638 ( .C1(n5332), .C2(n4954), .A(n4940), .B(n4939), .ZN(U3127)
         );
  AOI22_X1 U5639 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4950), .B1(n5495), 
        .B2(n4949), .ZN(n4942) );
  AOI22_X1 U5640 ( .A1(n5497), .A2(n4951), .B1(n5382), .B2(n5498), .ZN(n4941)
         );
  OAI211_X1 U5641 ( .C1(n5278), .C2(n4954), .A(n4942), .B(n4941), .ZN(U3124)
         );
  AOI22_X1 U5642 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4950), .B1(n5488), 
        .B2(n4949), .ZN(n4944) );
  AOI22_X1 U5643 ( .A1(n5490), .A2(n4951), .B1(n5382), .B2(n5491), .ZN(n4943)
         );
  OAI211_X1 U5644 ( .C1(n5319), .C2(n4954), .A(n4944), .B(n4943), .ZN(U3125)
         );
  AOI22_X1 U5645 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4950), .B1(n5523), 
        .B2(n4949), .ZN(n4946) );
  AOI22_X1 U5646 ( .A1(n5525), .A2(n4951), .B1(n5382), .B2(n5526), .ZN(n4945)
         );
  OAI211_X1 U5647 ( .C1(n5304), .C2(n4954), .A(n4946), .B(n4945), .ZN(U3128)
         );
  AOI22_X1 U5648 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4950), .B1(n5516), 
        .B2(n4949), .ZN(n4948) );
  AOI22_X1 U5649 ( .A1(n5518), .A2(n4951), .B1(n5382), .B2(n5519), .ZN(n4947)
         );
  OAI211_X1 U5650 ( .C1(n5316), .C2(n4954), .A(n4948), .B(n4947), .ZN(U3129)
         );
  AOI22_X1 U5651 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4950), .B1(n5531), 
        .B2(n4949), .ZN(n4953) );
  AOI22_X1 U5652 ( .A1(n5534), .A2(n4951), .B1(n5382), .B2(n5536), .ZN(n4952)
         );
  OAI211_X1 U5653 ( .C1(n5325), .C2(n4954), .A(n4953), .B(n4952), .ZN(U3126)
         );
  NAND2_X1 U5654 ( .A1(n4955), .A2(n4956), .ZN(n5458) );
  OR2_X1 U5655 ( .A1(n4955), .A2(n4956), .ZN(n4957) );
  NAND2_X1 U5656 ( .A1(n5458), .A2(n4957), .ZN(n5589) );
  INV_X1 U5657 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U5658 ( .A1(n4965), .A2(n6869), .ZN(n4959) );
  INV_X1 U5659 ( .A(EBX_REG_6__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U5660 ( .A1(n5816), .A2(n7015), .ZN(n4958) );
  NAND3_X1 U5661 ( .A1(n4959), .A2(n5805), .A3(n4958), .ZN(n4961) );
  NAND2_X1 U5662 ( .A1(n5819), .A2(n7015), .ZN(n4960) );
  OR2_X2 U5663 ( .A1(n5217), .A2(n5218), .ZN(n6118) );
  INV_X1 U5664 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6781) );
  NAND2_X1 U5665 ( .A1(n5809), .A2(n6781), .ZN(n4964) );
  NAND2_X1 U5666 ( .A1(n5816), .A2(n6781), .ZN(n4962) );
  OAI211_X1 U5667 ( .C1(n5819), .C2(n6906), .A(n4962), .B(n4965), .ZN(n4963)
         );
  NAND2_X1 U5668 ( .A1(n4964), .A2(n4963), .ZN(n6117) );
  NAND2_X1 U5669 ( .A1(n4965), .A2(n6900), .ZN(n4967) );
  INV_X1 U5670 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U5671 ( .A1(n5816), .A2(n4968), .ZN(n4966) );
  NAND3_X1 U5672 ( .A1(n4967), .A2(n5805), .A3(n4966), .ZN(n4970) );
  NAND2_X1 U5673 ( .A1(n5819), .A2(n4968), .ZN(n4969) );
  NAND2_X1 U5674 ( .A1(n4970), .A2(n4969), .ZN(n4971) );
  NOR2_X1 U5675 ( .A1(n6119), .A2(n4971), .ZN(n4972) );
  OR2_X1 U5676 ( .A1(n5462), .A2(n4972), .ZN(n6893) );
  INV_X1 U5677 ( .A(n6893), .ZN(n4973) );
  AOI22_X1 U5678 ( .A1(n6782), .A2(n4973), .B1(EBX_REG_8__SCAN_IN), .B2(n6159), 
        .ZN(n4974) );
  OAI21_X1 U5679 ( .B1(n5589), .B2(n6777), .A(n4974), .ZN(U2851) );
  NAND2_X1 U5680 ( .A1(n4012), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5221) );
  OAI21_X1 U5681 ( .B1(n4975), .B2(n5221), .A(n5282), .ZN(n4980) );
  INV_X1 U5682 ( .A(n4980), .ZN(n4978) );
  OR2_X1 U5683 ( .A1(n3429), .A2(n6944), .ZN(n5479) );
  INV_X1 U5684 ( .A(n5479), .ZN(n5020) );
  AND2_X1 U5685 ( .A1(n5020), .A2(n4636), .ZN(n5397) );
  INV_X1 U5686 ( .A(n5934), .ZN(n5207) );
  NAND3_X1 U5687 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5224), .ZN(n5395) );
  NOR2_X1 U5688 ( .A1(n5927), .A2(n5395), .ZN(n5011) );
  AOI21_X1 U5689 ( .B1(n5397), .B2(n5207), .A(n5011), .ZN(n4979) );
  INV_X1 U5690 ( .A(n5395), .ZN(n4976) );
  OAI21_X1 U5691 ( .B1(n5282), .B2(n4976), .A(n5266), .ZN(n4977) );
  INV_X1 U5692 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4986) );
  OAI22_X1 U5693 ( .A1(n4980), .A2(n4979), .B1(n5395), .B2(n6823), .ZN(n5015)
         );
  AND2_X1 U5694 ( .A1(n4012), .A2(n4018), .ZN(n5025) );
  NAND2_X1 U5695 ( .A1(n4982), .A2(n5025), .ZN(n5389) );
  AOI22_X1 U5696 ( .A1(n5510), .A2(n5011), .B1(n5512), .B2(n5427), .ZN(n4983)
         );
  OAI21_X1 U5697 ( .B1(n5336), .B2(n5013), .A(n4983), .ZN(n4984) );
  AOI21_X1 U5698 ( .B1(n5509), .B2(n5015), .A(n4984), .ZN(n4985) );
  OAI21_X1 U5699 ( .B1(n5018), .B2(n4986), .A(n4985), .ZN(U3114) );
  INV_X1 U5700 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4990) );
  AOI22_X1 U5701 ( .A1(n5503), .A2(n5011), .B1(n5505), .B2(n5427), .ZN(n4987)
         );
  OAI21_X1 U5702 ( .B1(n5310), .B2(n5013), .A(n4987), .ZN(n4988) );
  AOI21_X1 U5703 ( .B1(n5502), .B2(n5015), .A(n4988), .ZN(n4989) );
  OAI21_X1 U5704 ( .B1(n5018), .B2(n4990), .A(n4989), .ZN(U3115) );
  INV_X1 U5705 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4994) );
  AOI22_X1 U5706 ( .A1(n5524), .A2(n5011), .B1(n5526), .B2(n5427), .ZN(n4991)
         );
  OAI21_X1 U5707 ( .B1(n5295), .B2(n5013), .A(n4991), .ZN(n4992) );
  AOI21_X1 U5708 ( .B1(n5523), .B2(n5015), .A(n4992), .ZN(n4993) );
  OAI21_X1 U5709 ( .B1(n5018), .B2(n4994), .A(n4993), .ZN(U3112) );
  INV_X1 U5710 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4998) );
  AOI22_X1 U5711 ( .A1(n5517), .A2(n5011), .B1(n5519), .B2(n5427), .ZN(n4995)
         );
  OAI21_X1 U5712 ( .B1(n5298), .B2(n5013), .A(n4995), .ZN(n4996) );
  AOI21_X1 U5713 ( .B1(n5516), .B2(n5015), .A(n4996), .ZN(n4997) );
  OAI21_X1 U5714 ( .B1(n5018), .B2(n4998), .A(n4997), .ZN(U3113) );
  INV_X1 U5715 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5002) );
  AOI22_X1 U5716 ( .A1(n5496), .A2(n5011), .B1(n5498), .B2(n5427), .ZN(n4999)
         );
  OAI21_X1 U5717 ( .B1(n5313), .B2(n5013), .A(n4999), .ZN(n5000) );
  AOI21_X1 U5718 ( .B1(n5495), .B2(n5015), .A(n5000), .ZN(n5001) );
  OAI21_X1 U5719 ( .B1(n5018), .B2(n5002), .A(n5001), .ZN(U3108) );
  INV_X1 U5720 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n5006) );
  AOI22_X1 U5721 ( .A1(n5489), .A2(n5011), .B1(n5491), .B2(n5427), .ZN(n5003)
         );
  OAI21_X1 U5722 ( .B1(n5346), .B2(n5013), .A(n5003), .ZN(n5004) );
  AOI21_X1 U5723 ( .B1(n5488), .B2(n5015), .A(n5004), .ZN(n5005) );
  OAI21_X1 U5724 ( .B1(n5018), .B2(n5006), .A(n5005), .ZN(U3109) );
  INV_X1 U5725 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U5726 ( .A1(n5533), .A2(n5011), .B1(n5536), .B2(n5427), .ZN(n5007)
         );
  OAI21_X1 U5727 ( .B1(n5339), .B2(n5013), .A(n5007), .ZN(n5008) );
  AOI21_X1 U5728 ( .B1(n5531), .B2(n5015), .A(n5008), .ZN(n5009) );
  OAI21_X1 U5729 ( .B1(n5018), .B2(n5010), .A(n5009), .ZN(U3110) );
  INV_X1 U5730 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5017) );
  AOI22_X1 U5731 ( .A1(n5482), .A2(n5011), .B1(n5484), .B2(n5427), .ZN(n5012)
         );
  OAI21_X1 U5732 ( .B1(n5307), .B2(n5013), .A(n5012), .ZN(n5014) );
  AOI21_X1 U5733 ( .B1(n5481), .B2(n5015), .A(n5014), .ZN(n5016) );
  OAI21_X1 U5734 ( .B1(n5018), .B2(n5017), .A(n5016), .ZN(U3111) );
  INV_X1 U5735 ( .A(n5280), .ZN(n5284) );
  OAI21_X1 U5736 ( .B1(n5284), .B2(n5221), .A(n5282), .ZN(n5023) );
  NAND2_X1 U5737 ( .A1(n7128), .A2(n5224), .ZN(n5281) );
  NOR2_X1 U5738 ( .A1(n5019), .A2(n5281), .ZN(n5042) );
  AOI21_X1 U5739 ( .B1(n3448), .B2(n5020), .A(n5042), .ZN(n5024) );
  INV_X1 U5740 ( .A(n5024), .ZN(n5022) );
  OR2_X1 U5741 ( .A1(n7124), .A2(n5281), .ZN(n5470) );
  NAND2_X1 U5742 ( .A1(n5390), .A2(n5470), .ZN(n5021) );
  OAI211_X1 U5743 ( .C1(n5023), .C2(n5022), .A(n5266), .B(n5021), .ZN(n5041)
         );
  OAI22_X1 U5744 ( .A1(n5024), .A2(n5023), .B1(n6823), .B2(n5470), .ZN(n5040)
         );
  AOI22_X1 U5745 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5041), .B1(n5516), 
        .B2(n5040), .ZN(n5027) );
  AOI22_X1 U5746 ( .A1(n5517), .A2(n5042), .B1(n5519), .B2(n5535), .ZN(n5026)
         );
  OAI211_X1 U5747 ( .C1(n5298), .C2(n5045), .A(n5027), .B(n5026), .ZN(U3049)
         );
  AOI22_X1 U5748 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5041), .B1(n5523), 
        .B2(n5040), .ZN(n5029) );
  AOI22_X1 U5749 ( .A1(n5524), .A2(n5042), .B1(n5526), .B2(n5535), .ZN(n5028)
         );
  OAI211_X1 U5750 ( .C1(n5295), .C2(n5045), .A(n5029), .B(n5028), .ZN(U3048)
         );
  AOI22_X1 U5751 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5041), .B1(n5502), 
        .B2(n5040), .ZN(n5031) );
  AOI22_X1 U5752 ( .A1(n5503), .A2(n5042), .B1(n5505), .B2(n5535), .ZN(n5030)
         );
  OAI211_X1 U5753 ( .C1(n5310), .C2(n5045), .A(n5031), .B(n5030), .ZN(U3051)
         );
  AOI22_X1 U5754 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5041), .B1(n5509), 
        .B2(n5040), .ZN(n5033) );
  AOI22_X1 U5755 ( .A1(n5510), .A2(n5042), .B1(n5512), .B2(n5535), .ZN(n5032)
         );
  OAI211_X1 U5756 ( .C1(n5336), .C2(n5045), .A(n5033), .B(n5032), .ZN(U3050)
         );
  AOI22_X1 U5757 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5041), .B1(n5481), 
        .B2(n5040), .ZN(n5035) );
  AOI22_X1 U5758 ( .A1(n5482), .A2(n5042), .B1(n5484), .B2(n5535), .ZN(n5034)
         );
  OAI211_X1 U5759 ( .C1(n5307), .C2(n5045), .A(n5035), .B(n5034), .ZN(U3047)
         );
  AOI22_X1 U5760 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5041), .B1(n5531), 
        .B2(n5040), .ZN(n5037) );
  AOI22_X1 U5761 ( .A1(n5533), .A2(n5042), .B1(n5536), .B2(n5535), .ZN(n5036)
         );
  OAI211_X1 U5762 ( .C1(n5339), .C2(n5045), .A(n5037), .B(n5036), .ZN(U3046)
         );
  AOI22_X1 U5763 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5041), .B1(n5488), 
        .B2(n5040), .ZN(n5039) );
  AOI22_X1 U5764 ( .A1(n5489), .A2(n5042), .B1(n5491), .B2(n5535), .ZN(n5038)
         );
  OAI211_X1 U5765 ( .C1(n5346), .C2(n5045), .A(n5039), .B(n5038), .ZN(U3045)
         );
  AOI22_X1 U5766 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5041), .B1(n5495), 
        .B2(n5040), .ZN(n5044) );
  AOI22_X1 U5767 ( .A1(n5496), .A2(n5042), .B1(n5498), .B2(n5535), .ZN(n5043)
         );
  OAI211_X1 U5768 ( .C1(n5313), .C2(n5045), .A(n5044), .B(n5043), .ZN(U3044)
         );
  NAND2_X1 U5769 ( .A1(n5237), .A2(n5282), .ZN(n5231) );
  INV_X1 U5770 ( .A(n5076), .ZN(n5048) );
  INV_X1 U5771 ( .A(n5342), .ZN(n5047) );
  AOI21_X1 U5772 ( .B1(n5048), .B2(n5047), .A(n6463), .ZN(n5049) );
  AOI21_X1 U5773 ( .B1(n5359), .B2(n5231), .A(n5049), .ZN(n5052) );
  NOR3_X2 U5774 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n5281), .ZN(n5077) );
  NOR2_X1 U5775 ( .A1(n5471), .A2(n5077), .ZN(n5050) );
  NOR4_X2 U5776 ( .A1(n5052), .A2(n5475), .A3(n5051), .A4(n5050), .ZN(n5081)
         );
  INV_X1 U5777 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5056) );
  OAI22_X1 U5778 ( .A1(n5480), .A2(n5237), .B1(n5053), .B2(n5477), .ZN(n5075)
         );
  AOI22_X1 U5779 ( .A1(n5342), .A2(n5483), .B1(n5481), .B2(n5075), .ZN(n5055)
         );
  AOI22_X1 U5780 ( .A1(n5482), .A2(n5077), .B1(n5484), .B2(n5076), .ZN(n5054)
         );
  OAI211_X1 U5781 ( .C1(n5081), .C2(n5056), .A(n5055), .B(n5054), .ZN(U3023)
         );
  AOI22_X1 U5782 ( .A1(n5342), .A2(n5534), .B1(n5531), .B2(n5075), .ZN(n5058)
         );
  AOI22_X1 U5783 ( .A1(n5533), .A2(n5077), .B1(n5536), .B2(n5076), .ZN(n5057)
         );
  OAI211_X1 U5784 ( .C1(n5081), .C2(n5059), .A(n5058), .B(n5057), .ZN(U3022)
         );
  INV_X1 U5785 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U5786 ( .A1(n5342), .A2(n5490), .B1(n5488), .B2(n5075), .ZN(n5061)
         );
  AOI22_X1 U5787 ( .A1(n5489), .A2(n5077), .B1(n5491), .B2(n5076), .ZN(n5060)
         );
  OAI211_X1 U5788 ( .C1(n5081), .C2(n5062), .A(n5061), .B(n5060), .ZN(U3021)
         );
  AOI22_X1 U5789 ( .A1(n5342), .A2(n5497), .B1(n5495), .B2(n5075), .ZN(n5064)
         );
  AOI22_X1 U5790 ( .A1(n5496), .A2(n5077), .B1(n5498), .B2(n5076), .ZN(n5063)
         );
  OAI211_X1 U5791 ( .C1(n5081), .C2(n5065), .A(n5064), .B(n5063), .ZN(U3020)
         );
  AOI22_X1 U5792 ( .A1(n5342), .A2(n5504), .B1(n5502), .B2(n5075), .ZN(n5067)
         );
  AOI22_X1 U5793 ( .A1(n5503), .A2(n5077), .B1(n5505), .B2(n5076), .ZN(n5066)
         );
  OAI211_X1 U5794 ( .C1(n5081), .C2(n5068), .A(n5067), .B(n5066), .ZN(U3027)
         );
  INV_X1 U5795 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5071) );
  AOI22_X1 U5796 ( .A1(n5342), .A2(n5511), .B1(n5509), .B2(n5075), .ZN(n5070)
         );
  AOI22_X1 U5797 ( .A1(n5510), .A2(n5077), .B1(n5512), .B2(n5076), .ZN(n5069)
         );
  OAI211_X1 U5798 ( .C1(n5081), .C2(n5071), .A(n5070), .B(n5069), .ZN(U3026)
         );
  AOI22_X1 U5799 ( .A1(n5342), .A2(n5518), .B1(n5516), .B2(n5075), .ZN(n5073)
         );
  AOI22_X1 U5800 ( .A1(n5517), .A2(n5077), .B1(n5519), .B2(n5076), .ZN(n5072)
         );
  OAI211_X1 U5801 ( .C1(n5081), .C2(n5074), .A(n5073), .B(n5072), .ZN(U3025)
         );
  AOI22_X1 U5802 ( .A1(n5342), .A2(n5525), .B1(n5523), .B2(n5075), .ZN(n5079)
         );
  AOI22_X1 U5803 ( .A1(n5524), .A2(n5077), .B1(n5526), .B2(n5076), .ZN(n5078)
         );
  OAI211_X1 U5804 ( .C1(n5081), .C2(n5080), .A(n5079), .B(n5078), .ZN(U3024)
         );
  NAND2_X1 U5805 ( .A1(n5093), .A2(DATAI_10_), .ZN(n5090) );
  AOI22_X1 U5806 ( .A1(n5162), .A2(EAX_REG_10__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U5807 ( .A1(n5090), .A2(n5083), .ZN(U2949) );
  NAND2_X1 U5808 ( .A1(n5093), .A2(DATAI_0_), .ZN(n5096) );
  AOI22_X1 U5809 ( .A1(n5162), .A2(EAX_REG_0__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U5810 ( .A1(n5096), .A2(n5084), .ZN(U2939) );
  NAND2_X1 U5811 ( .A1(n5093), .A2(DATAI_14_), .ZN(n5100) );
  AOI22_X1 U5812 ( .A1(n5162), .A2(EAX_REG_30__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U5813 ( .A1(n5100), .A2(n5085), .ZN(U2938) );
  NAND2_X1 U5814 ( .A1(n5093), .A2(DATAI_13_), .ZN(n5102) );
  AOI22_X1 U5815 ( .A1(n5162), .A2(EAX_REG_29__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U5816 ( .A1(n5102), .A2(n5086), .ZN(U2937) );
  NAND2_X1 U5817 ( .A1(n5093), .A2(DATAI_12_), .ZN(n5104) );
  AOI22_X1 U5818 ( .A1(n5162), .A2(EAX_REG_28__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U5819 ( .A1(n5104), .A2(n5087), .ZN(U2936) );
  NAND2_X1 U5820 ( .A1(n5093), .A2(DATAI_11_), .ZN(n5107) );
  AOI22_X1 U5821 ( .A1(n5162), .A2(EAX_REG_27__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5822 ( .A1(n5107), .A2(n5088), .ZN(U2935) );
  AOI22_X1 U5823 ( .A1(n5162), .A2(EAX_REG_26__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5824 ( .A1(n5090), .A2(n5089), .ZN(U2934) );
  NAND2_X1 U5825 ( .A1(n5093), .A2(DATAI_3_), .ZN(n5115) );
  AOI22_X1 U5826 ( .A1(n5162), .A2(EAX_REG_19__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U5827 ( .A1(n5115), .A2(n5091), .ZN(U2927) );
  NAND2_X1 U5828 ( .A1(n5093), .A2(DATAI_2_), .ZN(n5121) );
  AOI22_X1 U5829 ( .A1(n5162), .A2(EAX_REG_18__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U5830 ( .A1(n5121), .A2(n5092), .ZN(U2926) );
  NAND2_X1 U5831 ( .A1(n5093), .A2(DATAI_1_), .ZN(n5123) );
  AOI22_X1 U5832 ( .A1(n5162), .A2(EAX_REG_17__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U5833 ( .A1(n5123), .A2(n5094), .ZN(U2925) );
  AOI22_X1 U5834 ( .A1(n5162), .A2(EAX_REG_16__SCAN_IN), .B1(n5161), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5835 ( .A1(n5096), .A2(n5095), .ZN(U2924) );
  AOI22_X1 U5836 ( .A1(n5162), .A2(EAX_REG_6__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5837 ( .A1(n5098), .A2(n5097), .ZN(U2945) );
  AOI22_X1 U5838 ( .A1(n5105), .A2(EAX_REG_14__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U5839 ( .A1(n5100), .A2(n5099), .ZN(U2953) );
  AOI22_X1 U5840 ( .A1(n5105), .A2(EAX_REG_13__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U5841 ( .A1(n5102), .A2(n5101), .ZN(U2952) );
  AOI22_X1 U5842 ( .A1(n5105), .A2(EAX_REG_12__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5843 ( .A1(n5104), .A2(n5103), .ZN(U2951) );
  AOI22_X1 U5844 ( .A1(n5105), .A2(EAX_REG_11__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U5845 ( .A1(n5107), .A2(n5106), .ZN(U2950) );
  AOI22_X1 U5846 ( .A1(n5162), .A2(EAX_REG_9__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U5847 ( .A1(n5109), .A2(n5108), .ZN(U2948) );
  AOI22_X1 U5848 ( .A1(n5162), .A2(EAX_REG_8__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U5849 ( .A1(n5111), .A2(n5110), .ZN(U2947) );
  AOI22_X1 U5850 ( .A1(n5162), .A2(EAX_REG_7__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U5851 ( .A1(n5113), .A2(n5112), .ZN(U2946) );
  AOI22_X1 U5852 ( .A1(n5162), .A2(EAX_REG_3__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U5853 ( .A1(n5115), .A2(n5114), .ZN(U2942) );
  AOI22_X1 U5854 ( .A1(n5162), .A2(EAX_REG_5__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U5855 ( .A1(n5117), .A2(n5116), .ZN(U2944) );
  AOI22_X1 U5856 ( .A1(n5162), .A2(EAX_REG_4__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U5857 ( .A1(n5119), .A2(n5118), .ZN(U2943) );
  AOI22_X1 U5858 ( .A1(n5162), .A2(EAX_REG_2__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U5859 ( .A1(n5121), .A2(n5120), .ZN(U2941) );
  AOI22_X1 U5860 ( .A1(n5162), .A2(EAX_REG_1__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U5861 ( .A1(n5123), .A2(n5122), .ZN(U2940) );
  INV_X1 U5862 ( .A(n3529), .ZN(n6446) );
  INV_X1 U5863 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7133) );
  NAND2_X1 U5864 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7133), .ZN(n5139) );
  INV_X1 U5865 ( .A(n5124), .ZN(n5138) );
  OR2_X1 U5866 ( .A1(n7119), .A2(n3449), .ZN(n5127) );
  NAND2_X1 U5867 ( .A1(n7119), .A2(n5125), .ZN(n5126) );
  INV_X1 U5868 ( .A(n7127), .ZN(n5136) );
  NAND2_X1 U5869 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5130) );
  INV_X1 U5870 ( .A(n5130), .ZN(n5129) );
  MUX2_X1 U5871 ( .A(n5130), .B(n5129), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n5135) );
  XNOR2_X1 U5872 ( .A(n5131), .B(n5969), .ZN(n5133) );
  OAI222_X1 U5873 ( .A1(n6438), .A2(n5135), .B1(n6972), .B2(n5134), .C1(n5133), 
        .C2(n5132), .ZN(n5967) );
  MUX2_X1 U5874 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5967), .S(n7119), 
        .Z(n7129) );
  NAND3_X1 U5875 ( .A1(n5136), .A2(n7129), .A3(n6443), .ZN(n5137) );
  OAI21_X1 U5876 ( .B1(n5139), .B2(n5138), .A(n5137), .ZN(n7137) );
  MUX2_X1 U5877 ( .A(FLUSH_REG_SCAN_IN), .B(n7119), .S(n6443), .Z(n5140) );
  NOR2_X1 U5878 ( .A1(n5140), .A2(n4034), .ZN(n5146) );
  INV_X1 U5879 ( .A(n5141), .ZN(n5142) );
  NOR2_X1 U5880 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  XNOR2_X1 U5881 ( .A(n5144), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6991)
         );
  NOR3_X1 U5882 ( .A1(n6991), .A2(STATE2_REG_1__SCAN_IN), .A3(n5145), .ZN(
        n7111) );
  NOR2_X1 U5883 ( .A1(n5146), .A2(n7111), .ZN(n7139) );
  INV_X1 U5884 ( .A(n7139), .ZN(n5147) );
  AOI21_X1 U5885 ( .B1(n6446), .B2(n7137), .A(n5147), .ZN(n7157) );
  AOI21_X1 U5886 ( .B1(n7157), .B2(n7133), .A(n7151), .ZN(n5149) );
  INV_X1 U5887 ( .A(n6454), .ZN(n5928) );
  OAI21_X1 U5888 ( .B1(n6443), .B2(STATE2_REG_3__SCAN_IN), .A(n5928), .ZN(
        n5933) );
  NOR2_X1 U5889 ( .A1(n6454), .A2(n5390), .ZN(n5930) );
  OAI21_X1 U5890 ( .B1(n5150), .B2(STATEBS16_REG_SCAN_IN), .A(n5283), .ZN(
        n5151) );
  AOI22_X1 U5891 ( .A1(n5930), .A2(n5151), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6454), .ZN(n5152) );
  OAI21_X1 U5892 ( .B1(n6944), .B2(n5933), .A(n5152), .ZN(U3464) );
  INV_X1 U5893 ( .A(n5153), .ZN(n5158) );
  INV_X1 U5894 ( .A(n5227), .ZN(n5154) );
  NAND2_X1 U5895 ( .A1(n5154), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5267) );
  NAND2_X1 U5896 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND3_X1 U5897 ( .A1(n5158), .A2(n5267), .A3(n5157), .ZN(n5159) );
  AOI22_X1 U5898 ( .A1(n5930), .A2(n5159), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6454), .ZN(n5160) );
  OAI21_X1 U5899 ( .B1(n6972), .B2(n5933), .A(n5160), .ZN(U3462) );
  INV_X1 U5900 ( .A(DATAI_15_), .ZN(n6584) );
  AOI22_X1 U5901 ( .A1(n5162), .A2(EAX_REG_15__SCAN_IN), .B1(n5161), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5163) );
  OAI21_X1 U5902 ( .B1(n5169), .B2(n6584), .A(n5163), .ZN(U2954) );
  AND2_X1 U5903 ( .A1(n5165), .A2(n5164), .ZN(n5166) );
  INV_X1 U5904 ( .A(n5171), .ZN(n5170) );
  INV_X1 U5905 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6680) );
  OAI222_X1 U5906 ( .A1(n5172), .A2(n6180), .B1(n5639), .B2(n6606), .C1(n5973), 
        .C2(n6680), .ZN(U2888) );
  INV_X1 U5907 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6676) );
  OAI222_X1 U5908 ( .A1(n5173), .A2(n6180), .B1(n5639), .B2(n6614), .C1(n5973), 
        .C2(n6676), .ZN(U2890) );
  INV_X1 U5909 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6674) );
  OAI222_X1 U5910 ( .A1(n6180), .A2(n5211), .B1(n5639), .B2(n6511), .C1(n5973), 
        .C2(n6674), .ZN(U2891) );
  OAI222_X1 U5911 ( .A1(n5175), .A2(n6180), .B1(n5639), .B2(n5174), .C1(n5973), 
        .C2(n4047), .ZN(U2886) );
  INV_X1 U5912 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U5913 ( .A1(n5176), .A2(n6180), .B1(n5639), .B2(n6605), .C1(n5973), 
        .C2(n6678), .ZN(U2889) );
  INV_X1 U5914 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6682) );
  OAI222_X1 U5915 ( .A1(n5177), .A2(n6180), .B1(n5639), .B2(n6503), .C1(n5973), 
        .C2(n6682), .ZN(U2887) );
  NOR2_X1 U5916 ( .A1(n5178), .A2(n5179), .ZN(n5180) );
  OR2_X1 U5917 ( .A1(n4955), .A2(n5180), .ZN(n6778) );
  OAI222_X1 U5918 ( .A1(n6778), .A2(n6180), .B1(n5639), .B2(n6596), .C1(n5973), 
        .C2(n4063), .ZN(U2884) );
  INV_X1 U5919 ( .A(DATAI_8_), .ZN(n6594) );
  INV_X1 U5920 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U5921 ( .A1(n5589), .A2(n6180), .B1(n5639), .B2(n6594), .C1(n5973), 
        .C2(n6687), .ZN(U2883) );
  INV_X1 U5922 ( .A(n5183), .ZN(n7161) );
  NOR3_X1 U5923 ( .A1(n7159), .A2(n5471), .A3(n7161), .ZN(n7155) );
  INV_X1 U5924 ( .A(n7155), .ZN(n5185) );
  NAND2_X1 U5925 ( .A1(n3426), .A2(n5184), .ZN(n7149) );
  NAND3_X1 U5926 ( .A1(n6912), .A2(n5185), .A3(n7149), .ZN(n5186) );
  INV_X1 U5927 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5996) );
  INV_X1 U5928 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5921) );
  INV_X1 U5929 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5956) );
  INV_X1 U5930 ( .A(n5946), .ZN(n5188) );
  NAND2_X1 U5931 ( .A1(n5188), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5189) );
  OAI21_X1 U5932 ( .B1(n5195), .B2(n5190), .A(n7073), .ZN(n7003) );
  INV_X1 U5933 ( .A(n7003), .ZN(n5212) );
  NOR2_X1 U5934 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5196) );
  AND3_X1 U5935 ( .A1(n5191), .A2(n5196), .A3(n3427), .ZN(n5192) );
  INV_X1 U5936 ( .A(n6979), .ZN(n6957) );
  INV_X1 U5937 ( .A(n6980), .ZN(n6055) );
  NAND3_X1 U5938 ( .A1(n6463), .A2(n7176), .A3(n5990), .ZN(n7144) );
  NOR2_X1 U5939 ( .A1(n5196), .A2(EBX_REG_31__SCAN_IN), .ZN(n5193) );
  AOI22_X1 U5940 ( .A1(n5979), .A2(n7144), .B1(n5193), .B2(n3677), .ZN(n5194)
         );
  INV_X1 U5941 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U5942 ( .A1(n5197), .A2(EBX_REG_31__SCAN_IN), .ZN(n5198) );
  NOR2_X1 U5943 ( .A1(n3455), .A2(n5198), .ZN(n5199) );
  OAI22_X1 U5944 ( .A1(n7094), .A2(n5201), .B1(n5200), .B2(n7083), .ZN(n5202)
         );
  AOI21_X1 U5945 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6055), .A(n5202), .ZN(n5210)
         );
  INV_X1 U5946 ( .A(n5203), .ZN(n5980) );
  NAND2_X1 U5947 ( .A1(n5954), .A2(n5980), .ZN(n6990) );
  INV_X1 U5948 ( .A(n6990), .ZN(n5208) );
  NAND2_X1 U5949 ( .A1(n5946), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5204) );
  INV_X1 U5950 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5205) );
  AOI21_X1 U5951 ( .B1(n7097), .B2(n7061), .A(n5205), .ZN(n5206) );
  AOI21_X1 U5952 ( .B1(n5208), .B2(n5207), .A(n5206), .ZN(n5209) );
  OAI211_X1 U5953 ( .C1(n5212), .C2(n5211), .A(n5210), .B(n5209), .ZN(U2827)
         );
  INV_X1 U5954 ( .A(n5213), .ZN(n5214) );
  AOI21_X1 U5955 ( .B1(n5215), .B2(n5214), .A(n5178), .ZN(n7017) );
  INV_X1 U5956 ( .A(n7017), .ZN(n5220) );
  INV_X1 U5957 ( .A(n6118), .ZN(n5216) );
  AOI21_X1 U5958 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n7013) );
  AOI22_X1 U5959 ( .A1(n6782), .A2(n7013), .B1(EBX_REG_6__SCAN_IN), .B2(n6159), 
        .ZN(n5219) );
  OAI21_X1 U5960 ( .B1(n5220), .B2(n6777), .A(n5219), .ZN(U2853) );
  OAI222_X1 U5961 ( .A1(n5220), .A2(n6180), .B1(n5639), .B2(n6500), .C1(n5973), 
        .C2(n4053), .ZN(U2885) );
  XNOR2_X1 U5962 ( .A(n5222), .B(n5221), .ZN(n5226) );
  INV_X1 U5963 ( .A(n5930), .ZN(n5225) );
  INV_X1 U5964 ( .A(n3429), .ZN(n6952) );
  OAI222_X1 U5965 ( .A1(n5226), .A2(n5225), .B1(n5933), .B2(n6952), .C1(n5224), 
        .C2(n5928), .ZN(U3463) );
  INV_X1 U5966 ( .A(n5260), .ZN(n5229) );
  INV_X1 U5967 ( .A(n5329), .ZN(n5228) );
  AOI21_X1 U5968 ( .B1(n5229), .B2(n5228), .A(n6463), .ZN(n5230) );
  AOI21_X1 U5969 ( .B1(n5480), .B2(n5231), .A(n5230), .ZN(n5236) );
  NAND2_X1 U5970 ( .A1(n5233), .A2(n5232), .ZN(n5356) );
  AND2_X1 U5971 ( .A1(n5356), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5349) );
  NOR2_X1 U5972 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5234), .ZN(n5261)
         );
  NOR2_X1 U5973 ( .A1(n5261), .A2(n5471), .ZN(n5235) );
  NOR4_X2 U5974 ( .A1(n5236), .A2(n5475), .A3(n5349), .A4(n5235), .ZN(n5265)
         );
  INV_X1 U5975 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5240) );
  OAI22_X1 U5976 ( .A1(n5359), .A2(n5237), .B1(n5356), .B2(n5477), .ZN(n5259)
         );
  AOI22_X1 U5977 ( .A1(n5260), .A2(n5518), .B1(n5516), .B2(n5259), .ZN(n5239)
         );
  AOI22_X1 U5978 ( .A1(n5517), .A2(n5261), .B1(n5519), .B2(n5329), .ZN(n5238)
         );
  OAI211_X1 U5979 ( .C1(n5265), .C2(n5240), .A(n5239), .B(n5238), .ZN(U3089)
         );
  INV_X1 U5980 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5243) );
  AOI22_X1 U5981 ( .A1(n5260), .A2(n5525), .B1(n5523), .B2(n5259), .ZN(n5242)
         );
  AOI22_X1 U5982 ( .A1(n5524), .A2(n5261), .B1(n5526), .B2(n5329), .ZN(n5241)
         );
  OAI211_X1 U5983 ( .C1(n5265), .C2(n5243), .A(n5242), .B(n5241), .ZN(U3088)
         );
  INV_X1 U5984 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U5985 ( .A1(n5260), .A2(n5534), .B1(n5531), .B2(n5259), .ZN(n5245)
         );
  AOI22_X1 U5986 ( .A1(n5533), .A2(n5261), .B1(n5536), .B2(n5329), .ZN(n5244)
         );
  OAI211_X1 U5987 ( .C1(n5265), .C2(n5246), .A(n5245), .B(n5244), .ZN(U3086)
         );
  INV_X1 U5988 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U5989 ( .A1(n5260), .A2(n5504), .B1(n5502), .B2(n5259), .ZN(n5248)
         );
  AOI22_X1 U5990 ( .A1(n5503), .A2(n5261), .B1(n5505), .B2(n5329), .ZN(n5247)
         );
  OAI211_X1 U5991 ( .C1(n5265), .C2(n5249), .A(n5248), .B(n5247), .ZN(U3091)
         );
  INV_X1 U5992 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5252) );
  AOI22_X1 U5993 ( .A1(n5260), .A2(n5497), .B1(n5495), .B2(n5259), .ZN(n5251)
         );
  AOI22_X1 U5994 ( .A1(n5496), .A2(n5261), .B1(n5498), .B2(n5329), .ZN(n5250)
         );
  OAI211_X1 U5995 ( .C1(n5265), .C2(n5252), .A(n5251), .B(n5250), .ZN(U3084)
         );
  INV_X1 U5996 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5255) );
  AOI22_X1 U5997 ( .A1(n5260), .A2(n5511), .B1(n5509), .B2(n5259), .ZN(n5254)
         );
  AOI22_X1 U5998 ( .A1(n5510), .A2(n5261), .B1(n5512), .B2(n5329), .ZN(n5253)
         );
  OAI211_X1 U5999 ( .C1(n5265), .C2(n5255), .A(n5254), .B(n5253), .ZN(U3090)
         );
  INV_X1 U6000 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5258) );
  AOI22_X1 U6001 ( .A1(n5260), .A2(n5490), .B1(n5488), .B2(n5259), .ZN(n5257)
         );
  AOI22_X1 U6002 ( .A1(n5489), .A2(n5261), .B1(n5491), .B2(n5329), .ZN(n5256)
         );
  OAI211_X1 U6003 ( .C1(n5265), .C2(n5258), .A(n5257), .B(n5256), .ZN(U3085)
         );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5264) );
  AOI22_X1 U6005 ( .A1(n5260), .A2(n5483), .B1(n5481), .B2(n5259), .ZN(n5263)
         );
  AOI22_X1 U6006 ( .A1(n5482), .A2(n5261), .B1(n5484), .B2(n5329), .ZN(n5262)
         );
  OAI211_X1 U6007 ( .C1(n5265), .C2(n5264), .A(n5263), .B(n5262), .ZN(U3087)
         );
  INV_X1 U6008 ( .A(n5266), .ZN(n5288) );
  NAND2_X1 U6009 ( .A1(n5267), .A2(n5282), .ZN(n5274) );
  INV_X1 U6010 ( .A(n5333), .ZN(n5268) );
  AOI21_X1 U6011 ( .B1(n3448), .B2(n5269), .A(n5268), .ZN(n5275) );
  INV_X1 U6012 ( .A(n5275), .ZN(n5270) );
  NOR2_X1 U6013 ( .A1(n5274), .A2(n5270), .ZN(n5271) );
  AOI211_X1 U6014 ( .C1(n5390), .C2(n5273), .A(n5288), .B(n5271), .ZN(n5272)
         );
  OAI22_X1 U6015 ( .A1(n5275), .A2(n5274), .B1(n6823), .B2(n5273), .ZN(n5326)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5327), .B1(n5495), 
        .B2(n5326), .ZN(n5277) );
  AOI22_X1 U6017 ( .A1(n5497), .A2(n5329), .B1(n5328), .B2(n5498), .ZN(n5276)
         );
  OAI211_X1 U6018 ( .C1(n5333), .C2(n5278), .A(n5277), .B(n5276), .ZN(U3076)
         );
  OR2_X1 U6019 ( .A1(n5281), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5290)
         );
  OAI21_X1 U6020 ( .B1(n5284), .B2(n5283), .A(n5282), .ZN(n5291) );
  NOR2_X1 U6021 ( .A1(n5927), .A2(n5290), .ZN(n5343) );
  AOI21_X1 U6022 ( .B1(n3448), .B2(n5285), .A(n5343), .ZN(n5292) );
  INV_X1 U6023 ( .A(n5292), .ZN(n5286) );
  NOR2_X1 U6024 ( .A1(n5291), .A2(n5286), .ZN(n5287) );
  AOI211_X1 U6025 ( .C1(n5390), .C2(n5290), .A(n5288), .B(n5287), .ZN(n5289)
         );
  OAI22_X1 U6026 ( .A1(n5292), .A2(n5291), .B1(n6823), .B2(n5290), .ZN(n5340)
         );
  AOI22_X1 U6027 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5341), .B1(n5523), 
        .B2(n5340), .ZN(n5294) );
  AOI22_X1 U6028 ( .A1(n5524), .A2(n5343), .B1(n5342), .B2(n5526), .ZN(n5293)
         );
  OAI211_X1 U6029 ( .C1(n5467), .C2(n5295), .A(n5294), .B(n5293), .ZN(U3032)
         );
  AOI22_X1 U6030 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5341), .B1(n5516), 
        .B2(n5340), .ZN(n5297) );
  AOI22_X1 U6031 ( .A1(n5517), .A2(n5343), .B1(n5342), .B2(n5519), .ZN(n5296)
         );
  OAI211_X1 U6032 ( .C1(n5467), .C2(n5298), .A(n5297), .B(n5296), .ZN(U3033)
         );
  AOI22_X1 U6033 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5327), .B1(n5502), 
        .B2(n5326), .ZN(n5300) );
  AOI22_X1 U6034 ( .A1(n5504), .A2(n5329), .B1(n5328), .B2(n5505), .ZN(n5299)
         );
  OAI211_X1 U6035 ( .C1(n5333), .C2(n5301), .A(n5300), .B(n5299), .ZN(U3083)
         );
  AOI22_X1 U6036 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5327), .B1(n5523), 
        .B2(n5326), .ZN(n5303) );
  AOI22_X1 U6037 ( .A1(n5525), .A2(n5329), .B1(n5328), .B2(n5526), .ZN(n5302)
         );
  OAI211_X1 U6038 ( .C1(n5333), .C2(n5304), .A(n5303), .B(n5302), .ZN(U3080)
         );
  AOI22_X1 U6039 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5341), .B1(n5481), 
        .B2(n5340), .ZN(n5306) );
  AOI22_X1 U6040 ( .A1(n5482), .A2(n5343), .B1(n5342), .B2(n5484), .ZN(n5305)
         );
  OAI211_X1 U6041 ( .C1(n5467), .C2(n5307), .A(n5306), .B(n5305), .ZN(U3031)
         );
  AOI22_X1 U6042 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5341), .B1(n5502), 
        .B2(n5340), .ZN(n5309) );
  AOI22_X1 U6043 ( .A1(n5503), .A2(n5343), .B1(n5342), .B2(n5505), .ZN(n5308)
         );
  OAI211_X1 U6044 ( .C1(n5467), .C2(n5310), .A(n5309), .B(n5308), .ZN(U3035)
         );
  AOI22_X1 U6045 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5341), .B1(n5495), 
        .B2(n5340), .ZN(n5312) );
  AOI22_X1 U6046 ( .A1(n5496), .A2(n5343), .B1(n5498), .B2(n5342), .ZN(n5311)
         );
  OAI211_X1 U6047 ( .C1(n5467), .C2(n5313), .A(n5312), .B(n5311), .ZN(U3028)
         );
  AOI22_X1 U6048 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5327), .B1(n5516), 
        .B2(n5326), .ZN(n5315) );
  AOI22_X1 U6049 ( .A1(n5518), .A2(n5329), .B1(n5328), .B2(n5519), .ZN(n5314)
         );
  OAI211_X1 U6050 ( .C1(n5333), .C2(n5316), .A(n5315), .B(n5314), .ZN(U3081)
         );
  AOI22_X1 U6051 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5327), .B1(n5488), 
        .B2(n5326), .ZN(n5318) );
  AOI22_X1 U6052 ( .A1(n5490), .A2(n5329), .B1(n5328), .B2(n5491), .ZN(n5317)
         );
  OAI211_X1 U6053 ( .C1(n5333), .C2(n5319), .A(n5318), .B(n5317), .ZN(U3077)
         );
  AOI22_X1 U6054 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5327), .B1(n5509), 
        .B2(n5326), .ZN(n5321) );
  AOI22_X1 U6055 ( .A1(n5511), .A2(n5329), .B1(n5328), .B2(n5512), .ZN(n5320)
         );
  OAI211_X1 U6056 ( .C1(n5333), .C2(n5322), .A(n5321), .B(n5320), .ZN(U3082)
         );
  AOI22_X1 U6057 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5327), .B1(n5531), 
        .B2(n5326), .ZN(n5324) );
  AOI22_X1 U6058 ( .A1(n5534), .A2(n5329), .B1(n5328), .B2(n5536), .ZN(n5323)
         );
  OAI211_X1 U6059 ( .C1(n5333), .C2(n5325), .A(n5324), .B(n5323), .ZN(U3078)
         );
  AOI22_X1 U6060 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5327), .B1(n5481), 
        .B2(n5326), .ZN(n5331) );
  AOI22_X1 U6061 ( .A1(n5483), .A2(n5329), .B1(n5328), .B2(n5484), .ZN(n5330)
         );
  OAI211_X1 U6062 ( .C1(n5333), .C2(n5332), .A(n5331), .B(n5330), .ZN(U3079)
         );
  AOI22_X1 U6063 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5341), .B1(n5509), 
        .B2(n5340), .ZN(n5335) );
  AOI22_X1 U6064 ( .A1(n5510), .A2(n5343), .B1(n5342), .B2(n5512), .ZN(n5334)
         );
  OAI211_X1 U6065 ( .C1(n5467), .C2(n5336), .A(n5335), .B(n5334), .ZN(U3034)
         );
  AOI22_X1 U6066 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5341), .B1(n5531), 
        .B2(n5340), .ZN(n5338) );
  AOI22_X1 U6067 ( .A1(n5533), .A2(n5343), .B1(n5342), .B2(n5536), .ZN(n5337)
         );
  OAI211_X1 U6068 ( .C1(n5467), .C2(n5339), .A(n5338), .B(n5337), .ZN(U3030)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5341), .B1(n5488), 
        .B2(n5340), .ZN(n5345) );
  AOI22_X1 U6070 ( .A1(n5489), .A2(n5343), .B1(n5342), .B2(n5491), .ZN(n5344)
         );
  OAI211_X1 U6071 ( .C1(n5467), .C2(n5346), .A(n5345), .B(n5344), .ZN(U3029)
         );
  NOR2_X1 U6072 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5347), .ZN(n5384)
         );
  INV_X1 U6073 ( .A(n5384), .ZN(n5350) );
  AOI211_X1 U6074 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5350), .A(n5349), .B(
        n5348), .ZN(n5355) );
  OAI21_X1 U6075 ( .B1(n5383), .B2(n5382), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5351) );
  OAI21_X1 U6076 ( .B1(n5353), .B2(n5352), .A(n5351), .ZN(n5354) );
  INV_X1 U6077 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5362) );
  OAI22_X1 U6078 ( .A1(n5359), .A2(n5358), .B1(n5357), .B2(n5356), .ZN(n5381)
         );
  AOI22_X1 U6079 ( .A1(n5382), .A2(n5511), .B1(n5509), .B2(n5381), .ZN(n5361)
         );
  AOI22_X1 U6080 ( .A1(n5510), .A2(n5384), .B1(n5512), .B2(n5383), .ZN(n5360)
         );
  OAI211_X1 U6081 ( .C1(n5388), .C2(n5362), .A(n5361), .B(n5360), .ZN(U3122)
         );
  INV_X1 U6082 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5365) );
  AOI22_X1 U6083 ( .A1(n5382), .A2(n5534), .B1(n5531), .B2(n5381), .ZN(n5364)
         );
  AOI22_X1 U6084 ( .A1(n5533), .A2(n5384), .B1(n5536), .B2(n5383), .ZN(n5363)
         );
  OAI211_X1 U6085 ( .C1(n5388), .C2(n5365), .A(n5364), .B(n5363), .ZN(U3118)
         );
  INV_X1 U6086 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5368) );
  AOI22_X1 U6087 ( .A1(n5382), .A2(n5518), .B1(n5516), .B2(n5381), .ZN(n5367)
         );
  AOI22_X1 U6088 ( .A1(n5517), .A2(n5384), .B1(n5519), .B2(n5383), .ZN(n5366)
         );
  OAI211_X1 U6089 ( .C1(n5388), .C2(n5368), .A(n5367), .B(n5366), .ZN(U3121)
         );
  INV_X1 U6090 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5371) );
  AOI22_X1 U6091 ( .A1(n5382), .A2(n5497), .B1(n5495), .B2(n5381), .ZN(n5370)
         );
  AOI22_X1 U6092 ( .A1(n5496), .A2(n5384), .B1(n5498), .B2(n5383), .ZN(n5369)
         );
  OAI211_X1 U6093 ( .C1(n5388), .C2(n5371), .A(n5370), .B(n5369), .ZN(U3116)
         );
  INV_X1 U6094 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5374) );
  AOI22_X1 U6095 ( .A1(n5382), .A2(n5525), .B1(n5523), .B2(n5381), .ZN(n5373)
         );
  AOI22_X1 U6096 ( .A1(n5524), .A2(n5384), .B1(n5526), .B2(n5383), .ZN(n5372)
         );
  OAI211_X1 U6097 ( .C1(n5388), .C2(n5374), .A(n5373), .B(n5372), .ZN(U3120)
         );
  INV_X1 U6098 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5377) );
  AOI22_X1 U6099 ( .A1(n5382), .A2(n5504), .B1(n5502), .B2(n5381), .ZN(n5376)
         );
  AOI22_X1 U6100 ( .A1(n5503), .A2(n5384), .B1(n5505), .B2(n5383), .ZN(n5375)
         );
  OAI211_X1 U6101 ( .C1(n5388), .C2(n5377), .A(n5376), .B(n5375), .ZN(U3123)
         );
  INV_X1 U6102 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5380) );
  AOI22_X1 U6103 ( .A1(n5382), .A2(n5490), .B1(n5488), .B2(n5381), .ZN(n5379)
         );
  AOI22_X1 U6104 ( .A1(n5489), .A2(n5384), .B1(n5491), .B2(n5383), .ZN(n5378)
         );
  OAI211_X1 U6105 ( .C1(n5388), .C2(n5380), .A(n5379), .B(n5378), .ZN(U3117)
         );
  INV_X1 U6106 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5387) );
  AOI22_X1 U6107 ( .A1(n5382), .A2(n5483), .B1(n5481), .B2(n5381), .ZN(n5386)
         );
  AOI22_X1 U6108 ( .A1(n5482), .A2(n5384), .B1(n5484), .B2(n5383), .ZN(n5385)
         );
  OAI211_X1 U6109 ( .C1(n5388), .C2(n5387), .A(n5386), .B(n5385), .ZN(U3119)
         );
  NAND2_X1 U6110 ( .A1(n5403), .A2(n5389), .ZN(n5391) );
  AOI21_X1 U6111 ( .B1(n5391), .B2(STATEBS16_REG_SCAN_IN), .A(n5390), .ZN(
        n5399) );
  INV_X1 U6112 ( .A(n5392), .ZN(n5394) );
  INV_X1 U6113 ( .A(n5477), .ZN(n5393) );
  AOI22_X1 U6114 ( .A1(n5399), .A2(n5397), .B1(n5394), .B2(n5393), .ZN(n5432)
         );
  INV_X1 U6115 ( .A(n5531), .ZN(n5406) );
  NOR2_X1 U6116 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5395), .ZN(n5426)
         );
  NOR2_X1 U6117 ( .A1(n5475), .A2(n5396), .ZN(n5401) );
  INV_X1 U6118 ( .A(n5397), .ZN(n5398) );
  NAND2_X1 U6119 ( .A1(n5399), .A2(n5398), .ZN(n5400) );
  AND2_X1 U6120 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  AOI22_X1 U6121 ( .A1(n5533), .A2(n5426), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5425), .ZN(n5405) );
  AOI22_X1 U6122 ( .A1(n5534), .A2(n5427), .B1(n5428), .B2(n5536), .ZN(n5404)
         );
  OAI211_X1 U6123 ( .C1(n5432), .C2(n5406), .A(n5405), .B(n5404), .ZN(U3102)
         );
  INV_X1 U6124 ( .A(n5481), .ZN(n5409) );
  AOI22_X1 U6125 ( .A1(n5482), .A2(n5426), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5425), .ZN(n5408) );
  AOI22_X1 U6126 ( .A1(n5483), .A2(n5427), .B1(n5428), .B2(n5484), .ZN(n5407)
         );
  OAI211_X1 U6127 ( .C1(n5432), .C2(n5409), .A(n5408), .B(n5407), .ZN(U3103)
         );
  INV_X1 U6128 ( .A(n5502), .ZN(n5412) );
  AOI22_X1 U6129 ( .A1(n5503), .A2(n5426), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5425), .ZN(n5411) );
  AOI22_X1 U6130 ( .A1(n5504), .A2(n5427), .B1(n5428), .B2(n5505), .ZN(n5410)
         );
  OAI211_X1 U6131 ( .C1(n5432), .C2(n5412), .A(n5411), .B(n5410), .ZN(U3107)
         );
  INV_X1 U6132 ( .A(n5516), .ZN(n5415) );
  AOI22_X1 U6133 ( .A1(n5517), .A2(n5426), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5425), .ZN(n5414) );
  AOI22_X1 U6134 ( .A1(n5518), .A2(n5427), .B1(n5428), .B2(n5519), .ZN(n5413)
         );
  OAI211_X1 U6135 ( .C1(n5432), .C2(n5415), .A(n5414), .B(n5413), .ZN(U3105)
         );
  INV_X1 U6136 ( .A(n5523), .ZN(n5418) );
  AOI22_X1 U6137 ( .A1(n5524), .A2(n5426), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5425), .ZN(n5417) );
  AOI22_X1 U6138 ( .A1(n5525), .A2(n5427), .B1(n5428), .B2(n5526), .ZN(n5416)
         );
  OAI211_X1 U6139 ( .C1(n5432), .C2(n5418), .A(n5417), .B(n5416), .ZN(U3104)
         );
  INV_X1 U6140 ( .A(n5509), .ZN(n5421) );
  AOI22_X1 U6141 ( .A1(n5510), .A2(n5426), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5425), .ZN(n5420) );
  AOI22_X1 U6142 ( .A1(n5511), .A2(n5427), .B1(n5428), .B2(n5512), .ZN(n5419)
         );
  OAI211_X1 U6143 ( .C1(n5432), .C2(n5421), .A(n5420), .B(n5419), .ZN(U3106)
         );
  INV_X1 U6144 ( .A(n5488), .ZN(n5424) );
  AOI22_X1 U6145 ( .A1(n5489), .A2(n5426), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5425), .ZN(n5423) );
  AOI22_X1 U6146 ( .A1(n5490), .A2(n5427), .B1(n5428), .B2(n5491), .ZN(n5422)
         );
  OAI211_X1 U6147 ( .C1(n5432), .C2(n5424), .A(n5423), .B(n5422), .ZN(U3101)
         );
  INV_X1 U6148 ( .A(n5495), .ZN(n5431) );
  AOI22_X1 U6149 ( .A1(n5496), .A2(n5426), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5425), .ZN(n5430) );
  AOI22_X1 U6150 ( .A1(n5428), .A2(n5498), .B1(n5427), .B2(n5497), .ZN(n5429)
         );
  OAI211_X1 U6151 ( .C1(n5432), .C2(n5431), .A(n5430), .B(n5429), .ZN(U3100)
         );
  XNOR2_X1 U6152 ( .A(n3435), .B(n5433), .ZN(n5726) );
  INV_X1 U6153 ( .A(DATAI_12_), .ZN(n6593) );
  OAI222_X1 U6154 ( .A1(n6180), .A2(n5726), .B1(n5639), .B2(n6593), .C1(n5973), 
        .C2(n4129), .ZN(U2879) );
  NAND3_X1 U6155 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6987) );
  OR2_X1 U6156 ( .A1(n6987), .A2(n6707), .ZN(n6998) );
  NOR2_X1 U6157 ( .A1(n6998), .A2(n6997), .ZN(n6115) );
  INV_X1 U6158 ( .A(n6115), .ZN(n6114) );
  INV_X1 U6159 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6710) );
  INV_X1 U6160 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6712) );
  NOR3_X1 U6161 ( .A1(n6114), .A2(n6710), .A3(n6712), .ZN(n5436) );
  NAND2_X1 U6162 ( .A1(n5436), .A2(REIP_REG_8__SCAN_IN), .ZN(n5542) );
  INV_X1 U6163 ( .A(n5542), .ZN(n5567) );
  NOR2_X1 U6164 ( .A1(n7041), .A2(n5567), .ZN(n5435) );
  OR2_X1 U6165 ( .A1(n5435), .A2(n6979), .ZN(n6109) );
  INV_X1 U6166 ( .A(n5592), .ZN(n5434) );
  OAI22_X1 U6167 ( .A1(n7083), .A2(n6893), .B1(n5434), .B2(n7061), .ZN(n5439)
         );
  AOI22_X1 U6168 ( .A1(EBX_REG_8__SCAN_IN), .A2(n7079), .B1(n5436), .B2(n5435), 
        .ZN(n5437) );
  OAI211_X1 U6169 ( .C1(n7097), .C2(n5588), .A(n5437), .B(n7051), .ZN(n5438)
         );
  AOI211_X1 U6170 ( .C1(REIP_REG_8__SCAN_IN), .C2(n6109), .A(n5439), .B(n5438), 
        .ZN(n5440) );
  OAI21_X1 U6171 ( .B1(n7073), .B2(n5589), .A(n5440), .ZN(U2819) );
  MUX2_X1 U6172 ( .A(n5809), .B(n5819), .S(EBX_REG_9__SCAN_IN), .Z(n5442) );
  NOR2_X1 U6173 ( .A1(n5949), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5441)
         );
  NOR2_X1 U6174 ( .A1(n5442), .A2(n5441), .ZN(n5461) );
  NAND2_X1 U6175 ( .A1(n4965), .A2(n6920), .ZN(n5444) );
  INV_X1 U6176 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6177 ( .A1(n5816), .A2(n5445), .ZN(n5443) );
  NAND3_X1 U6178 ( .A1(n5444), .A2(n5805), .A3(n5443), .ZN(n5447) );
  NAND2_X1 U6179 ( .A1(n5819), .A2(n5445), .ZN(n5446) );
  MUX2_X1 U6180 ( .A(n5795), .B(n5805), .S(EBX_REG_11__SCAN_IN), .Z(n5449) );
  NAND2_X1 U6181 ( .A1(n5796), .A2(n5669), .ZN(n5448) );
  NAND2_X1 U6182 ( .A1(n5449), .A2(n5448), .ZN(n5616) );
  INV_X1 U6183 ( .A(n5580), .ZN(n5615) );
  OAI21_X1 U6184 ( .B1(n5819), .B2(n5451), .A(n4965), .ZN(n5453) );
  INV_X1 U6185 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6186 ( .A1(n5816), .A2(n5456), .ZN(n5452) );
  NAND2_X1 U6187 ( .A1(n5453), .A2(n5452), .ZN(n5455) );
  NAND2_X1 U6188 ( .A1(n5819), .A2(n5456), .ZN(n5454) );
  NAND2_X1 U6189 ( .A1(n5455), .A2(n5454), .ZN(n5577) );
  XNOR2_X1 U6190 ( .A(n5615), .B(n5577), .ZN(n5543) );
  OAI222_X1 U6191 ( .A1(n6776), .A2(n5543), .B1(n6777), .B2(n5726), .C1(n5456), 
        .C2(n6785), .ZN(U2847) );
  INV_X1 U6192 ( .A(n5551), .ZN(n5457) );
  AOI21_X1 U6193 ( .B1(n5459), .B2(n5458), .A(n5457), .ZN(n6104) );
  INV_X1 U6194 ( .A(n6104), .ZN(n5466) );
  INV_X1 U6195 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6689) );
  OAI222_X1 U6196 ( .A1(n5466), .A2(n6180), .B1(n5639), .B2(n5460), .C1(n5973), 
        .C2(n6689), .ZN(U2882) );
  INV_X1 U6197 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5465) );
  OR2_X1 U6198 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  AND2_X1 U6199 ( .A1(n5553), .A2(n5463), .ZN(n6923) );
  INV_X1 U6200 ( .A(n6923), .ZN(n5464) );
  OAI222_X1 U6201 ( .A1(n5466), .A2(n6777), .B1(n6785), .B2(n5465), .C1(n5464), 
        .C2(n6776), .ZN(U2850) );
  OAI21_X1 U6202 ( .B1(n5537), .B2(n5535), .A(n5468), .ZN(n5469) );
  OAI21_X1 U6203 ( .B1(n4636), .B2(n5479), .A(n5469), .ZN(n5472) );
  NOR2_X1 U6204 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5470), .ZN(n5532)
         );
  AOI21_X1 U6205 ( .B1(n5472), .B2(n5471), .A(n5532), .ZN(n5476) );
  INV_X1 U6206 ( .A(n5473), .ZN(n5474) );
  NOR3_X2 U6207 ( .A1(n5476), .A2(n5475), .A3(n5474), .ZN(n5541) );
  INV_X1 U6208 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5487) );
  OAI22_X1 U6209 ( .A1(n5480), .A2(n5479), .B1(n5478), .B2(n5477), .ZN(n5530)
         );
  AOI22_X1 U6210 ( .A1(n5482), .A2(n5532), .B1(n5481), .B2(n5530), .ZN(n5486)
         );
  AOI22_X1 U6211 ( .A1(n5537), .A2(n5484), .B1(n5535), .B2(n5483), .ZN(n5485)
         );
  OAI211_X1 U6212 ( .C1(n5541), .C2(n5487), .A(n5486), .B(n5485), .ZN(U3039)
         );
  INV_X1 U6213 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5494) );
  AOI22_X1 U6214 ( .A1(n5489), .A2(n5532), .B1(n5488), .B2(n5530), .ZN(n5493)
         );
  AOI22_X1 U6215 ( .A1(n5537), .A2(n5491), .B1(n5535), .B2(n5490), .ZN(n5492)
         );
  OAI211_X1 U6216 ( .C1(n5541), .C2(n5494), .A(n5493), .B(n5492), .ZN(U3037)
         );
  INV_X1 U6217 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5501) );
  AOI22_X1 U6218 ( .A1(n5496), .A2(n5532), .B1(n5495), .B2(n5530), .ZN(n5500)
         );
  AOI22_X1 U6219 ( .A1(n5537), .A2(n5498), .B1(n5535), .B2(n5497), .ZN(n5499)
         );
  OAI211_X1 U6220 ( .C1(n5541), .C2(n5501), .A(n5500), .B(n5499), .ZN(U3036)
         );
  INV_X1 U6221 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5508) );
  AOI22_X1 U6222 ( .A1(n5503), .A2(n5532), .B1(n5502), .B2(n5530), .ZN(n5507)
         );
  AOI22_X1 U6223 ( .A1(n5537), .A2(n5505), .B1(n5535), .B2(n5504), .ZN(n5506)
         );
  OAI211_X1 U6224 ( .C1(n5541), .C2(n5508), .A(n5507), .B(n5506), .ZN(U3043)
         );
  INV_X1 U6225 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5515) );
  AOI22_X1 U6226 ( .A1(n5510), .A2(n5532), .B1(n5509), .B2(n5530), .ZN(n5514)
         );
  AOI22_X1 U6227 ( .A1(n5537), .A2(n5512), .B1(n5535), .B2(n5511), .ZN(n5513)
         );
  OAI211_X1 U6228 ( .C1(n5541), .C2(n5515), .A(n5514), .B(n5513), .ZN(U3042)
         );
  INV_X1 U6229 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5522) );
  AOI22_X1 U6230 ( .A1(n5517), .A2(n5532), .B1(n5516), .B2(n5530), .ZN(n5521)
         );
  AOI22_X1 U6231 ( .A1(n5537), .A2(n5519), .B1(n5535), .B2(n5518), .ZN(n5520)
         );
  OAI211_X1 U6232 ( .C1(n5541), .C2(n5522), .A(n5521), .B(n5520), .ZN(U3041)
         );
  INV_X1 U6233 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5529) );
  AOI22_X1 U6234 ( .A1(n5524), .A2(n5532), .B1(n5523), .B2(n5530), .ZN(n5528)
         );
  AOI22_X1 U6235 ( .A1(n5537), .A2(n5526), .B1(n5535), .B2(n5525), .ZN(n5527)
         );
  OAI211_X1 U6236 ( .C1(n5541), .C2(n5529), .A(n5528), .B(n5527), .ZN(U3040)
         );
  INV_X1 U6237 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5540) );
  AOI22_X1 U6238 ( .A1(n5533), .A2(n5532), .B1(n5531), .B2(n5530), .ZN(n5539)
         );
  AOI22_X1 U6239 ( .A1(n5537), .A2(n5536), .B1(n5535), .B2(n5534), .ZN(n5538)
         );
  OAI211_X1 U6240 ( .C1(n5541), .C2(n5540), .A(n5539), .B(n5538), .ZN(U3038)
         );
  INV_X1 U6241 ( .A(n5722), .ZN(n5549) );
  INV_X1 U6242 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6715) );
  NOR2_X1 U6243 ( .A1(n5542), .A2(n6715), .ZN(n5560) );
  AND2_X1 U6244 ( .A1(n5560), .A2(REIP_REG_10__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U6245 ( .A1(n7021), .A2(REIP_REG_11__SCAN_IN), .ZN(n5544) );
  INV_X1 U6246 ( .A(n5544), .ZN(n5701) );
  NOR2_X1 U6247 ( .A1(n7041), .A2(n5701), .ZN(n7020) );
  OR2_X1 U6248 ( .A1(n7020), .A2(n6979), .ZN(n7035) );
  AOI22_X1 U6249 ( .A1(EBX_REG_12__SCAN_IN), .A2(n7079), .B1(
        REIP_REG_12__SCAN_IN), .B2(n7035), .ZN(n5546) );
  INV_X1 U6250 ( .A(n5543), .ZN(n6931) );
  NOR3_X1 U6251 ( .A1(n7041), .A2(REIP_REG_12__SCAN_IN), .A3(n5544), .ZN(n7036) );
  AOI211_X1 U6252 ( .C1(n7104), .C2(n6931), .A(n7057), .B(n7036), .ZN(n5545)
         );
  OAI211_X1 U6253 ( .C1(n5547), .C2(n7097), .A(n5546), .B(n5545), .ZN(n5548)
         );
  AOI21_X1 U6254 ( .B1(n7101), .B2(n5549), .A(n5548), .ZN(n5550) );
  OAI21_X1 U6255 ( .B1(n5726), .B2(n7073), .A(n5550), .ZN(U2815) );
  NOR2_X1 U6256 ( .A1(n5551), .A2(n5552), .ZN(n5612) );
  AOI21_X1 U6257 ( .B1(n5552), .B2(n5551), .A(n5612), .ZN(n5646) );
  INV_X1 U6258 ( .A(n5646), .ZN(n5583) );
  INV_X1 U6259 ( .A(n5553), .ZN(n5557) );
  INV_X1 U6260 ( .A(n5554), .ZN(n5556) );
  OAI21_X1 U6261 ( .B1(n5557), .B2(n5556), .A(n5617), .ZN(n6914) );
  INV_X1 U6262 ( .A(n6914), .ZN(n5558) );
  AOI22_X1 U6263 ( .A1(n6782), .A2(n5558), .B1(EBX_REG_10__SCAN_IN), .B2(n6159), .ZN(n5559) );
  OAI21_X1 U6264 ( .B1(n5583), .B2(n6777), .A(n5559), .ZN(U2849) );
  INV_X1 U6265 ( .A(n5644), .ZN(n5564) );
  INV_X1 U6266 ( .A(n7041), .ZN(n6124) );
  INV_X1 U6267 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6913) );
  NAND3_X1 U6268 ( .A1(n6124), .A2(n6913), .A3(n5560), .ZN(n5561) );
  OAI211_X1 U6269 ( .C1(n7097), .C2(n5562), .A(n7051), .B(n5561), .ZN(n5563)
         );
  AOI21_X1 U6270 ( .B1(n7101), .B2(n5564), .A(n5563), .ZN(n5565) );
  OAI21_X1 U6271 ( .B1(n7083), .B2(n6914), .A(n5565), .ZN(n5566) );
  AOI21_X1 U6272 ( .B1(n7079), .B2(EBX_REG_10__SCAN_IN), .A(n5566), .ZN(n5570)
         );
  NAND2_X1 U6273 ( .A1(n5567), .A2(n6715), .ZN(n5568) );
  NOR2_X1 U6274 ( .A1(n7041), .A2(n5568), .ZN(n6108) );
  OAI21_X1 U6275 ( .B1(n6109), .B2(n6108), .A(REIP_REG_10__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U6276 ( .C1(n5583), .C2(n7073), .A(n5570), .B(n5569), .ZN(U2817)
         );
  NAND2_X1 U6277 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  NAND2_X1 U6278 ( .A1(n5574), .A2(n5573), .ZN(n7033) );
  MUX2_X1 U6279 ( .A(n5795), .B(n5805), .S(EBX_REG_13__SCAN_IN), .Z(n5576) );
  NAND2_X1 U6280 ( .A1(n5796), .A2(n5675), .ZN(n5575) );
  AND2_X1 U6281 ( .A1(n5576), .A2(n5575), .ZN(n5578) );
  AOI21_X1 U6282 ( .B1(n5615), .B2(n5577), .A(n5578), .ZN(n5581) );
  NAND2_X1 U6283 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  NOR2_X1 U6284 ( .A1(n5581), .A2(n5629), .ZN(n7029) );
  AOI22_X1 U6285 ( .A1(n6782), .A2(n7029), .B1(EBX_REG_13__SCAN_IN), .B2(n6159), .ZN(n5582) );
  OAI21_X1 U6286 ( .B1(n7033), .B2(n6777), .A(n5582), .ZN(U2846) );
  INV_X1 U6287 ( .A(DATAI_10_), .ZN(n6599) );
  INV_X1 U6288 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6691) );
  OAI222_X1 U6289 ( .A1(n5583), .A2(n6180), .B1(n5639), .B2(n6599), .C1(n5973), 
        .C2(n6691), .ZN(U2881) );
  OAI21_X1 U6290 ( .B1(n5586), .B2(n5585), .A(n5584), .ZN(n6891) );
  INV_X1 U6291 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5587) );
  OAI22_X1 U6292 ( .A1(n6287), .A2(n5588), .B1(n6912), .B2(n5587), .ZN(n5591)
         );
  NOR2_X1 U6293 ( .A1(n5589), .A2(n6291), .ZN(n5590) );
  AOI211_X1 U6294 ( .C1(n6805), .C2(n5592), .A(n5591), .B(n5590), .ZN(n5593)
         );
  OAI21_X1 U6295 ( .B1(n7108), .B2(n6891), .A(n5593), .ZN(U2978) );
  INV_X1 U6296 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5595) );
  AOI22_X1 U6297 ( .A1(n6699), .A2(UWORD_REG_2__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5594) );
  OAI21_X1 U6298 ( .B1(n5595), .B2(n5603), .A(n5594), .ZN(U2905) );
  INV_X1 U6299 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5597) );
  AOI22_X1 U6300 ( .A1(n6699), .A2(UWORD_REG_1__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5596) );
  OAI21_X1 U6301 ( .B1(n5597), .B2(n5603), .A(n5596), .ZN(U2906) );
  INV_X1 U6302 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5599) );
  AOI22_X1 U6303 ( .A1(n6699), .A2(UWORD_REG_3__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5598) );
  OAI21_X1 U6304 ( .B1(n5599), .B2(n5603), .A(n5598), .ZN(U2904) );
  INV_X1 U6305 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5601) );
  AOI22_X1 U6306 ( .A1(n6699), .A2(UWORD_REG_0__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5600) );
  OAI21_X1 U6307 ( .B1(n5601), .B2(n5603), .A(n5600), .ZN(U2907) );
  INV_X1 U6308 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5604) );
  AOI22_X1 U6309 ( .A1(n6699), .A2(UWORD_REG_14__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5602) );
  OAI21_X1 U6310 ( .B1(n5604), .B2(n5603), .A(n5602), .ZN(U2893) );
  INV_X1 U6311 ( .A(DATAI_13_), .ZN(n6590) );
  INV_X1 U6312 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6696) );
  OAI222_X1 U6313 ( .A1(n7033), .A2(n6180), .B1(n5639), .B2(n6590), .C1(n5973), 
        .C2(n6696), .ZN(U2878) );
  OAI21_X1 U6314 ( .B1(n5607), .B2(n5606), .A(n5605), .ZN(n6921) );
  INV_X1 U6315 ( .A(n5608), .ZN(n6106) );
  AOI22_X1 U6316 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6924), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5609) );
  OAI21_X1 U6317 ( .B1(n6815), .B2(n6106), .A(n5609), .ZN(n5610) );
  AOI21_X1 U6318 ( .B1(n6104), .B2(n4644), .A(n5610), .ZN(n5611) );
  OAI21_X1 U6319 ( .B1(n6921), .B2(n7108), .A(n5611), .ZN(U2977) );
  INV_X1 U6320 ( .A(n5612), .ZN(n5613) );
  AOI21_X1 U6321 ( .B1(n5614), .B2(n5613), .A(n3435), .ZN(n7024) );
  INV_X1 U6322 ( .A(n7024), .ZN(n5619) );
  AOI21_X1 U6323 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n7022) );
  AOI22_X1 U6324 ( .A1(n6782), .A2(n7022), .B1(EBX_REG_11__SCAN_IN), .B2(n6159), .ZN(n5618) );
  OAI21_X1 U6325 ( .B1(n5619), .B2(n6777), .A(n5618), .ZN(U2848) );
  INV_X1 U6326 ( .A(DATAI_11_), .ZN(n6598) );
  INV_X1 U6327 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6693) );
  OAI222_X1 U6328 ( .A1(n5619), .A2(n6180), .B1(n5639), .B2(n6598), .C1(n5973), 
        .C2(n6693), .ZN(U2880) );
  OR2_X1 U6329 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  NAND2_X1 U6330 ( .A1(n5620), .A2(n5623), .ZN(n7049) );
  INV_X1 U6331 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5630) );
  OAI21_X1 U6332 ( .B1(n5819), .B2(n6419), .A(n4965), .ZN(n5625) );
  NAND2_X1 U6333 ( .A1(n5816), .A2(n5630), .ZN(n5624) );
  NAND2_X1 U6334 ( .A1(n5625), .A2(n5624), .ZN(n5627) );
  NAND2_X1 U6335 ( .A1(n5819), .A2(n5630), .ZN(n5626) );
  NAND2_X1 U6336 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  NAND2_X1 U6337 ( .A1(n5629), .A2(n5628), .ZN(n5636) );
  OAI21_X1 U6338 ( .B1(n5629), .B2(n5628), .A(n5636), .ZN(n7043) );
  OAI222_X1 U6339 ( .A1(n7049), .A2(n6777), .B1(n5630), .B2(n6785), .C1(n6776), 
        .C2(n7043), .ZN(U2845) );
  INV_X1 U6340 ( .A(DATAI_14_), .ZN(n6587) );
  INV_X1 U6341 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6698) );
  OAI222_X1 U6342 ( .A1(n7049), .A2(n6180), .B1(n5639), .B2(n6587), .C1(n5973), 
        .C2(n6698), .ZN(U2877) );
  NAND2_X1 U6343 ( .A1(n5620), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U6344 ( .A1(n5682), .A2(n5632), .ZN(n7063) );
  MUX2_X1 U6345 ( .A(n5795), .B(n5805), .S(EBX_REG_15__SCAN_IN), .Z(n5634) );
  NAND2_X1 U6346 ( .A1(n5796), .A2(n6428), .ZN(n5633) );
  NAND2_X1 U6347 ( .A1(n5634), .A2(n5633), .ZN(n5637) );
  INV_X1 U6348 ( .A(n5689), .ZN(n5635) );
  AOI21_X1 U6349 ( .B1(n5637), .B2(n5636), .A(n5635), .ZN(n7056) );
  AOI22_X1 U6350 ( .A1(n6782), .A2(n7056), .B1(EBX_REG_15__SCAN_IN), .B2(n6159), .ZN(n5638) );
  OAI21_X1 U6351 ( .B1(n7063), .B2(n6777), .A(n5638), .ZN(U2844) );
  INV_X1 U6352 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6702) );
  OAI222_X1 U6353 ( .A1(n7063), .A2(n6180), .B1(n5639), .B2(n6584), .C1(n5973), 
        .C2(n6702), .ZN(U2876) );
  NAND2_X1 U6354 ( .A1(n5648), .A2(n5640), .ZN(n5642) );
  XOR2_X1 U6355 ( .A(n5642), .B(n5641), .Z(n6908) );
  AOI22_X1 U6356 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6924), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5643) );
  OAI21_X1 U6357 ( .B1(n5644), .B2(n6815), .A(n5643), .ZN(n5645) );
  AOI21_X1 U6358 ( .B1(n5646), .B2(n4644), .A(n5645), .ZN(n5647) );
  OAI21_X1 U6359 ( .B1(n6908), .B2(n7108), .A(n5647), .ZN(U2976) );
  INV_X1 U6360 ( .A(n5715), .ZN(n5650) );
  NAND2_X1 U6361 ( .A1(n5650), .A2(n5714), .ZN(n5651) );
  XNOR2_X1 U6362 ( .A(n5716), .B(n5651), .ZN(n6808) );
  NAND2_X1 U6363 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6897) );
  NAND3_X1 U6364 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6863), .ZN(n6896) );
  NOR2_X1 U6365 ( .A1(n6897), .A2(n6896), .ZN(n6910) );
  NOR2_X1 U6366 ( .A1(n6920), .A2(n6927), .ZN(n6911) );
  NAND2_X1 U6367 ( .A1(n6910), .A2(n6911), .ZN(n5658) );
  OR3_X1 U6368 ( .A1(n6869), .A2(n3886), .A3(n5652), .ZN(n6889) );
  NOR2_X1 U6369 ( .A1(n6897), .A2(n6889), .ZN(n5660) );
  NAND2_X1 U6370 ( .A1(n5660), .A2(n6911), .ZN(n5654) );
  NOR2_X1 U6371 ( .A1(n5653), .A2(n5654), .ZN(n5657) );
  NOR2_X1 U6372 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  NOR2_X1 U6373 ( .A1(n5657), .A2(n5656), .ZN(n6934) );
  NOR2_X1 U6374 ( .A1(n6933), .A2(n6910), .ZN(n5659) );
  INV_X1 U6375 ( .A(n5660), .ZN(n5661) );
  NOR2_X1 U6376 ( .A1(n5663), .A2(n5662), .ZN(n6926) );
  NAND2_X1 U6377 ( .A1(n6926), .A2(n6911), .ZN(n5666) );
  INV_X1 U6378 ( .A(n5663), .ZN(n5664) );
  NAND2_X1 U6379 ( .A1(n5664), .A2(n6417), .ZN(n5665) );
  NAND2_X1 U6380 ( .A1(n5666), .A2(n5665), .ZN(n6415) );
  AOI22_X1 U6381 ( .A1(n6932), .A2(n7022), .B1(n6924), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U6382 ( .B1(n6415), .B2(n5669), .A(n5667), .ZN(n5668) );
  AOI21_X1 U6383 ( .B1(n6929), .B2(n5669), .A(n5668), .ZN(n5670) );
  OAI21_X1 U6384 ( .B1(n6808), .B2(n6892), .A(n5670), .ZN(U3007) );
  XOR2_X1 U6385 ( .A(n5671), .B(n5672), .Z(n5739) );
  INV_X1 U6386 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6722) );
  NOR2_X1 U6387 ( .A1(n6912), .A2(n6722), .ZN(n5678) );
  NAND3_X1 U6389 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6420) );
  INV_X1 U6390 ( .A(n6417), .ZN(n5673) );
  INV_X1 U6391 ( .A(n6415), .ZN(n6935) );
  AOI21_X1 U6392 ( .B1(n6420), .B2(n5673), .A(n6935), .ZN(n5753) );
  INV_X1 U6393 ( .A(n6929), .ZN(n6421) );
  NAND2_X1 U6394 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5674) );
  OAI33_X1 U6395 ( .A1(1'b0), .A2(n5753), .A3(n5675), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6421), .B3(n5674), .ZN(n5677)
         );
  AOI211_X1 U6396 ( .C1(n6932), .C2(n7029), .A(n5678), .B(n5677), .ZN(n5679)
         );
  OAI21_X1 U6397 ( .B1(n5739), .B2(n6892), .A(n5679), .ZN(U3005) );
  AND2_X1 U6398 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  NOR2_X1 U6399 ( .A1(n5680), .A2(n5683), .ZN(n7185) );
  INV_X1 U6400 ( .A(n7185), .ZN(n5713) );
  NAND2_X1 U6401 ( .A1(n4965), .A2(n5684), .ZN(n5686) );
  INV_X1 U6402 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6403 ( .A1(n5816), .A2(n5709), .ZN(n5685) );
  NAND3_X1 U6404 ( .A1(n5686), .A2(n5805), .A3(n5685), .ZN(n5688) );
  NAND2_X1 U6405 ( .A1(n5819), .A2(n5709), .ZN(n5687) );
  AOI21_X1 U6406 ( .B1(n5690), .B2(n5689), .A(n5694), .ZN(n6418) );
  AOI22_X1 U6407 ( .A1(n6418), .A2(n6782), .B1(EBX_REG_16__SCAN_IN), .B2(n6159), .ZN(n5691) );
  OAI21_X1 U6408 ( .B1(n5713), .B2(n6777), .A(n5691), .ZN(U2843) );
  MUX2_X1 U6409 ( .A(n5795), .B(n5805), .S(EBX_REG_17__SCAN_IN), .Z(n5693) );
  NAND2_X1 U6410 ( .A1(n5796), .A2(n6400), .ZN(n5692) );
  NOR2_X1 U6411 ( .A1(n5694), .A2(n5695), .ZN(n5696) );
  OR2_X1 U6412 ( .A1(n5768), .A2(n5696), .ZN(n6406) );
  INV_X1 U6413 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5700) );
  OR2_X1 U6414 ( .A1(n5680), .A2(n5698), .ZN(n5699) );
  NAND2_X1 U6415 ( .A1(n5697), .A2(n5699), .ZN(n6275) );
  OAI222_X1 U6416 ( .A1(n6406), .A2(n6776), .B1(n6785), .B2(n5700), .C1(n6275), 
        .C2(n6777), .ZN(U2842) );
  INV_X1 U6417 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6726) );
  INV_X1 U6418 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U6419 ( .A1(n5701), .A2(REIP_REG_12__SCAN_IN), .ZN(n7030) );
  NOR2_X1 U6420 ( .A1(n7030), .A2(n6722), .ZN(n7045) );
  NAND2_X1 U6421 ( .A1(n7045), .A2(REIP_REG_14__SCAN_IN), .ZN(n5727) );
  NOR2_X1 U6422 ( .A1(n7041), .A2(n5727), .ZN(n7059) );
  INV_X1 U6423 ( .A(n7059), .ZN(n5702) );
  AOI21_X1 U6424 ( .B1(n6726), .B2(n7058), .A(n5702), .ZN(n5703) );
  NAND2_X1 U6425 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5728) );
  AOI22_X1 U6426 ( .A1(n5704), .A2(n7101), .B1(n5703), .B2(n5728), .ZN(n5712)
         );
  INV_X1 U6427 ( .A(n5727), .ZN(n5705) );
  OAI21_X1 U6428 ( .B1(n7041), .B2(n5705), .A(n6957), .ZN(n7055) );
  OAI21_X1 U6429 ( .B1(n7097), .B2(n5706), .A(n7051), .ZN(n5707) );
  AOI21_X1 U6430 ( .B1(n7104), .B2(n6418), .A(n5707), .ZN(n5708) );
  OAI21_X1 U6431 ( .B1(n5709), .B2(n7094), .A(n5708), .ZN(n5710) );
  AOI21_X1 U6432 ( .B1(REIP_REG_16__SCAN_IN), .B2(n7055), .A(n5710), .ZN(n5711) );
  OAI211_X1 U6433 ( .C1(n5713), .C2(n7073), .A(n5712), .B(n5711), .ZN(U2811)
         );
  OAI21_X1 U6434 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5720) );
  NAND2_X1 U6435 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  XNOR2_X1 U6436 ( .A(n5720), .B(n5719), .ZN(n6939) );
  NAND2_X1 U6437 ( .A1(n6939), .A2(n6810), .ZN(n5725) );
  INV_X1 U6438 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5721) );
  NOR2_X1 U6439 ( .A1(n6912), .A2(n5721), .ZN(n6930) );
  NOR2_X1 U6440 ( .A1(n6815), .A2(n5722), .ZN(n5723) );
  AOI211_X1 U6441 ( .C1(n6809), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6930), 
        .B(n5723), .ZN(n5724) );
  OAI211_X1 U6442 ( .C1(n5726), .C2(n6291), .A(n5725), .B(n5724), .ZN(U2974)
         );
  NOR2_X1 U6443 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  NAND2_X1 U6444 ( .A1(n5729), .A2(REIP_REG_17__SCAN_IN), .ZN(n5882) );
  NOR2_X1 U6445 ( .A1(n5882), .A2(n6979), .ZN(n6070) );
  OR2_X1 U6446 ( .A1(n6980), .A2(n6070), .ZN(n6090) );
  AOI21_X1 U6447 ( .B1(n6124), .B2(n5729), .A(REIP_REG_17__SCAN_IN), .ZN(n5738) );
  INV_X1 U6448 ( .A(n6275), .ZN(n7188) );
  NAND2_X1 U6449 ( .A1(n7188), .A2(n7105), .ZN(n5737) );
  OAI21_X1 U6450 ( .B1(n7097), .B2(n6270), .A(n7051), .ZN(n5732) );
  INV_X1 U6451 ( .A(n6272), .ZN(n5730) );
  NOR2_X1 U6452 ( .A1(n7061), .A2(n5730), .ZN(n5731) );
  NOR2_X1 U6453 ( .A1(n5732), .A2(n5731), .ZN(n5734) );
  NAND2_X1 U6454 ( .A1(n7079), .A2(EBX_REG_17__SCAN_IN), .ZN(n5733) );
  OAI211_X1 U6455 ( .C1(n6406), .C2(n7083), .A(n5734), .B(n5733), .ZN(n5735)
         );
  INV_X1 U6456 ( .A(n5735), .ZN(n5736) );
  OAI211_X1 U6457 ( .C1(n6090), .C2(n5738), .A(n5737), .B(n5736), .ZN(U2810)
         );
  OR2_X1 U6458 ( .A1(n5739), .A2(n7108), .ZN(n5744) );
  INV_X1 U6459 ( .A(n7032), .ZN(n5742) );
  OAI22_X1 U6460 ( .A1(n6287), .A2(n5740), .B1(n6912), .B2(n6722), .ZN(n5741)
         );
  AOI21_X1 U6461 ( .B1(n6805), .B2(n5742), .A(n5741), .ZN(n5743) );
  OAI211_X1 U6462 ( .C1(n6291), .C2(n7033), .A(n5744), .B(n5743), .ZN(U2973)
         );
  OAI21_X1 U6463 ( .B1(n5747), .B2(n5746), .A(n5745), .ZN(n5754) );
  NAND2_X1 U6464 ( .A1(n5754), .A2(n6938), .ZN(n5752) );
  NOR2_X1 U6465 ( .A1(n6421), .A2(n6420), .ZN(n5750) );
  INV_X1 U6466 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5748) );
  NOR2_X1 U6467 ( .A1(n6912), .A2(n5748), .ZN(n5756) );
  NOR2_X1 U6468 ( .A1(n6915), .A2(n7043), .ZN(n5749) );
  AOI211_X1 U6469 ( .C1(n5750), .C2(n6419), .A(n5756), .B(n5749), .ZN(n5751)
         );
  OAI211_X1 U6470 ( .C1(n5753), .C2(n6419), .A(n5752), .B(n5751), .ZN(U3004)
         );
  NAND2_X1 U6471 ( .A1(n5754), .A2(n6810), .ZN(n5758) );
  NOR2_X1 U6472 ( .A1(n6287), .A2(n7042), .ZN(n5755) );
  AOI211_X1 U6473 ( .C1(n6805), .C2(n7047), .A(n5756), .B(n5755), .ZN(n5757)
         );
  OAI211_X1 U6474 ( .C1(n6291), .C2(n7049), .A(n5758), .B(n5757), .ZN(U2972)
         );
  NAND2_X1 U6475 ( .A1(n5697), .A2(n5760), .ZN(n5761) );
  AND2_X1 U6476 ( .A1(n5759), .A2(n5761), .ZN(n7191) );
  INV_X1 U6477 ( .A(n7191), .ZN(n5775) );
  INV_X1 U6478 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5776) );
  INV_X1 U6479 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6728) );
  OAI22_X1 U6480 ( .A1(n7094), .A2(n5776), .B1(n6728), .B2(n6090), .ZN(n5773)
         );
  NOR2_X1 U6481 ( .A1(n7041), .A2(n5882), .ZN(n6080) );
  NAND2_X1 U6482 ( .A1(n6080), .A2(n6728), .ZN(n6091) );
  OAI211_X1 U6483 ( .C1(n7061), .C2(n6814), .A(n6091), .B(n7051), .ZN(n5772)
         );
  NAND2_X1 U6484 ( .A1(n4965), .A2(n5762), .ZN(n5764) );
  NAND2_X1 U6485 ( .A1(n5816), .A2(n5776), .ZN(n5763) );
  NAND3_X1 U6486 ( .A1(n5764), .A2(n5805), .A3(n5763), .ZN(n5766) );
  NAND2_X1 U6487 ( .A1(n5819), .A2(n5776), .ZN(n5765) );
  NAND2_X1 U6488 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  OR2_X1 U6489 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  NAND2_X1 U6490 ( .A1(n6094), .A2(n5769), .ZN(n6398) );
  INV_X1 U6491 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5770) );
  OAI22_X1 U6492 ( .A1(n7083), .A2(n6398), .B1(n5770), .B2(n7097), .ZN(n5771)
         );
  NOR3_X1 U6493 ( .A1(n5773), .A2(n5772), .A3(n5771), .ZN(n5774) );
  OAI21_X1 U6494 ( .B1(n5775), .B2(n7073), .A(n5774), .ZN(U2809) );
  OAI22_X1 U6495 ( .A1(n6398), .A2(n6776), .B1(n5776), .B2(n6785), .ZN(n5777)
         );
  AOI21_X1 U6496 ( .B1(n7191), .B2(n6783), .A(n5777), .ZN(n5778) );
  INV_X1 U6497 ( .A(n5778), .ZN(U2841) );
  OAI22_X1 U6498 ( .A1(n5949), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n3455), .ZN(n5951) );
  INV_X1 U6499 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U6500 ( .A1(n5809), .A2(n6161), .ZN(n5781) );
  INV_X1 U6501 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U6502 ( .A1(n5816), .A2(n6161), .ZN(n5779) );
  OAI211_X1 U6503 ( .C1(n5819), .C2(n6841), .A(n5779), .B(n4965), .ZN(n5780)
         );
  NAND2_X1 U6504 ( .A1(n5781), .A2(n5780), .ZN(n6093) );
  INV_X1 U6505 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6384) );
  OAI21_X1 U6506 ( .B1(n5819), .B2(n6384), .A(n4965), .ZN(n5783) );
  INV_X1 U6507 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U6508 ( .A1(n5816), .A2(n6083), .ZN(n5782) );
  AOI22_X1 U6509 ( .A1(n5783), .A2(n5782), .B1(n5819), .B2(n6083), .ZN(n6082)
         );
  INV_X1 U6510 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U6511 ( .A1(n5809), .A2(n6158), .ZN(n5786) );
  INV_X1 U6512 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U6513 ( .A1(n5816), .A2(n6158), .ZN(n5784) );
  OAI211_X1 U6514 ( .C1(n5819), .C2(n6366), .A(n5784), .B(n4965), .ZN(n5785)
         );
  INV_X1 U6515 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U6516 ( .A1(n4965), .A2(n6233), .ZN(n5788) );
  INV_X1 U6517 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6518 ( .A1(n5816), .A2(n5789), .ZN(n5787) );
  NAND3_X1 U6519 ( .A1(n5788), .A2(n5805), .A3(n5787), .ZN(n5791) );
  NAND2_X1 U6520 ( .A1(n5819), .A2(n5789), .ZN(n5790) );
  NAND2_X1 U6521 ( .A1(n5791), .A2(n5790), .ZN(n6066) );
  MUX2_X1 U6522 ( .A(n5795), .B(n5805), .S(EBX_REG_23__SCAN_IN), .Z(n5794) );
  INV_X1 U6523 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6524 ( .A1(n5796), .A2(n5792), .ZN(n5793) );
  NAND2_X1 U6525 ( .A1(n5794), .A2(n5793), .ZN(n6145) );
  MUX2_X1 U6526 ( .A(n5795), .B(n5805), .S(EBX_REG_25__SCAN_IN), .Z(n5798) );
  NAND2_X1 U6527 ( .A1(n5796), .A2(n6336), .ZN(n5797) );
  NAND2_X1 U6528 ( .A1(n5798), .A2(n5797), .ZN(n6048) );
  INV_X1 U6529 ( .A(n6048), .ZN(n5803) );
  INV_X1 U6530 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U6531 ( .A1(n4965), .A2(n6354), .ZN(n5800) );
  INV_X1 U6532 ( .A(EBX_REG_24__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U6533 ( .A1(n5816), .A2(n7093), .ZN(n5799) );
  NAND3_X1 U6534 ( .A1(n5800), .A2(n5805), .A3(n5799), .ZN(n5802) );
  NAND2_X1 U6535 ( .A1(n5819), .A2(n7093), .ZN(n5801) );
  NAND2_X1 U6536 ( .A1(n5802), .A2(n5801), .ZN(n6349) );
  NAND2_X1 U6537 ( .A1(n5803), .A2(n6349), .ZN(n5804) );
  NAND2_X1 U6538 ( .A1(n4965), .A2(n6337), .ZN(n5806) );
  OAI211_X1 U6539 ( .C1(EBX_REG_26__SCAN_IN), .C2(n3455), .A(n5806), .B(n5805), 
        .ZN(n5808) );
  INV_X1 U6540 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U6541 ( .A1(n5819), .A2(n6140), .ZN(n5807) );
  INV_X1 U6542 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U6543 ( .A1(n5809), .A2(n6138), .ZN(n5812) );
  NAND2_X1 U6544 ( .A1(n5816), .A2(n6138), .ZN(n5810) );
  OAI211_X1 U6545 ( .C1(n5819), .C2(n6324), .A(n5810), .B(n4965), .ZN(n5811)
         );
  AND2_X1 U6546 ( .A1(n5812), .A2(n5811), .ZN(n6018) );
  NAND2_X1 U6547 ( .A1(n4965), .A2(n6316), .ZN(n5813) );
  OAI211_X1 U6548 ( .C1(EBX_REG_28__SCAN_IN), .C2(n3455), .A(n5813), .B(n5805), 
        .ZN(n5815) );
  INV_X1 U6549 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U6550 ( .A1(n5819), .A2(n6137), .ZN(n5814) );
  NAND2_X1 U6551 ( .A1(n5815), .A2(n5814), .ZN(n6007) );
  INV_X1 U6552 ( .A(n6009), .ZN(n5822) );
  OR2_X1 U6553 ( .A1(n5949), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5818)
         );
  INV_X1 U6554 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U6555 ( .A1(n5816), .A2(n6134), .ZN(n5817) );
  NAND2_X1 U6556 ( .A1(n5818), .A2(n5817), .ZN(n5821) );
  NAND2_X1 U6557 ( .A1(n5819), .A2(n6134), .ZN(n5820) );
  OAI21_X1 U6558 ( .B1(n5821), .B2(n5819), .A(n5820), .ZN(n6000) );
  OAI21_X1 U6559 ( .B1(n5822), .B2(n5821), .A(n5950), .ZN(n5823) );
  XOR2_X1 U6560 ( .A(n5951), .B(n5823), .Z(n6131) );
  XOR2_X1 U6561 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n5824), .Z(n6187) );
  AOI22_X1 U6562 ( .A1(n4430), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5966), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5828) );
  AOI22_X1 U6563 ( .A1(n5855), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5827) );
  AOI22_X1 U6564 ( .A1(n5856), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5826) );
  AOI22_X1 U6565 ( .A1(n5847), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5825) );
  NAND4_X1 U6566 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n5835)
         );
  AOI22_X1 U6567 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n5860), .B1(n4436), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5833) );
  AOI22_X1 U6568 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n5858), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5832) );
  AOI22_X1 U6569 ( .A1(n5845), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5831) );
  AOI22_X1 U6570 ( .A1(n5849), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5830) );
  NAND4_X1 U6571 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n5834)
         );
  NOR2_X1 U6572 ( .A1(n5835), .A2(n5834), .ZN(n5844) );
  NAND2_X1 U6573 ( .A1(n5837), .A2(n5836), .ZN(n5843) );
  XOR2_X1 U6574 ( .A(n5844), .B(n5843), .Z(n5838) );
  NAND2_X1 U6575 ( .A1(n5838), .A2(n5869), .ZN(n5840) );
  AOI21_X1 U6576 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6823), .A(n3426), 
        .ZN(n5839) );
  OAI211_X1 U6577 ( .C1(n4067), .C2(n4787), .A(n5840), .B(n5839), .ZN(n5841)
         );
  OAI21_X1 U6578 ( .B1(n5872), .B2(n6187), .A(n5841), .ZN(n5995) );
  NOR2_X1 U6579 ( .A1(n5844), .A2(n5843), .ZN(n5868) );
  AOI22_X1 U6580 ( .A1(n5845), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5854) );
  AOI22_X1 U6581 ( .A1(n5847), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5846), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5853) );
  AOI22_X1 U6582 ( .A1(n5849), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5848), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5852) );
  AOI22_X1 U6583 ( .A1(n5966), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5850), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5851) );
  NAND4_X1 U6584 ( .A1(n5854), .A2(n5853), .A3(n5852), .A4(n5851), .ZN(n5866)
         );
  AOI22_X1 U6585 ( .A1(n5855), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5864) );
  AOI22_X1 U6586 ( .A1(n4436), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5856), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5863) );
  AOI22_X1 U6587 ( .A1(n5858), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5857), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5862) );
  AOI22_X1 U6588 ( .A1(n5860), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5859), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5861) );
  NAND4_X1 U6589 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(n5865)
         );
  NOR2_X1 U6590 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  XNOR2_X1 U6591 ( .A(n5868), .B(n5867), .ZN(n5870) );
  NAND2_X1 U6592 ( .A1(n5870), .A2(n5869), .ZN(n5879) );
  NAND2_X1 U6593 ( .A1(n6823), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5871)
         );
  NAND2_X1 U6594 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  AOI21_X1 U6595 ( .B1(n5874), .B2(EAX_REG_30__SCAN_IN), .A(n5873), .ZN(n5878)
         );
  XNOR2_X1 U6596 ( .A(n5875), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5918)
         );
  AND2_X1 U6597 ( .A1(n5918), .A2(n3426), .ZN(n5877) );
  AOI21_X1 U6598 ( .B1(n5879), .B2(n5878), .A(n5877), .ZN(n5940) );
  NAND2_X1 U6599 ( .A1(n6130), .A2(n7105), .ZN(n5890) );
  INV_X1 U6600 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6551) );
  INV_X1 U6601 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U6602 ( .A1(n6551), .A2(n6750), .ZN(n5886) );
  NAND2_X1 U6603 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6025) );
  NAND2_X1 U6604 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n5881) );
  NOR2_X1 U6605 ( .A1(n6025), .A2(n5881), .ZN(n5958) );
  INV_X1 U6606 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7092) );
  INV_X1 U6607 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6736) );
  INV_X1 U6608 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6738) );
  INV_X1 U6609 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6733) );
  INV_X1 U6610 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6730) );
  NOR3_X1 U6611 ( .A1(n6733), .A2(n6728), .A3(n6730), .ZN(n6071) );
  NAND2_X1 U6612 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6071), .ZN(n6065) );
  NOR2_X1 U6613 ( .A1(n7092), .A2(n7096), .ZN(n5957) );
  NAND2_X1 U6614 ( .A1(n5958), .A2(n5957), .ZN(n5883) );
  OAI21_X1 U6615 ( .B1(n6979), .B2(n5883), .A(n6055), .ZN(n5885) );
  OAI21_X1 U6616 ( .B1(n5886), .B2(n7041), .A(n5885), .ZN(n5961) );
  INV_X1 U6617 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6132) );
  AOI22_X1 U6618 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7071), .B1(n7101), 
        .B2(n5918), .ZN(n5884) );
  OAI21_X1 U6619 ( .B1(n7094), .B2(n6132), .A(n5884), .ZN(n5888) );
  INV_X1 U6620 ( .A(n5885), .ZN(n6011) );
  NOR4_X1 U6621 ( .A1(n6011), .A2(n5886), .A3(n7041), .A4(n6750), .ZN(n5887)
         );
  AOI211_X1 U6622 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5961), .A(n5888), .B(n5887), .ZN(n5889) );
  OAI211_X1 U6623 ( .C1(n6131), .C2(n7083), .A(n5890), .B(n5889), .ZN(U2797)
         );
  NOR2_X1 U6624 ( .A1(n5974), .A2(n3655), .ZN(n5891) );
  NAND2_X1 U6625 ( .A1(n6130), .A2(n7206), .ZN(n5894) );
  AND2_X1 U6626 ( .A1(n5973), .A2(n5892), .ZN(n7205) );
  AOI22_X1 U6627 ( .A1(n7205), .A2(DATAI_30_), .B1(n7208), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5893) );
  OAI211_X1 U6628 ( .C1(n6173), .C2(n6587), .A(n5894), .B(n5893), .ZN(U2861)
         );
  AND2_X1 U6629 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U6630 ( .A1(n6303), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6298) );
  AND2_X1 U6631 ( .A1(n6248), .A2(n6298), .ZN(n5898) );
  NAND2_X1 U6632 ( .A1(n3938), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6633 ( .A1(n6193), .A2(n5899), .ZN(n5900) );
  NAND2_X1 U6634 ( .A1(n5936), .A2(n5895), .ZN(n5901) );
  NAND2_X1 U6635 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  XNOR2_X1 U6636 ( .A(n5903), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5924)
         );
  INV_X1 U6637 ( .A(n6131), .ZN(n5916) );
  NOR2_X1 U6638 ( .A1(n6419), .A2(n6420), .ZN(n6416) );
  NAND3_X1 U6639 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6416), .ZN(n6410) );
  NOR2_X1 U6640 ( .A1(n6410), .A2(n5904), .ZN(n5906) );
  INV_X1 U6641 ( .A(n5905), .ZN(n6226) );
  NAND2_X1 U6642 ( .A1(n6835), .A2(n6226), .ZN(n6360) );
  NOR2_X1 U6643 ( .A1(n6360), .A2(n5909), .ZN(n6334) );
  AND2_X1 U6644 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U6645 ( .A1(n6334), .A2(n6335), .ZN(n6328) );
  OR3_X1 U6646 ( .A1(n6328), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6298), 
        .ZN(n5914) );
  OR2_X1 U6647 ( .A1(n6417), .A2(n5906), .ZN(n5907) );
  OR2_X1 U6648 ( .A1(n6417), .A2(n6226), .ZN(n5908) );
  NAND2_X1 U6649 ( .A1(n6842), .A2(n5908), .ZN(n6363) );
  INV_X1 U6650 ( .A(n5909), .ZN(n5910) );
  AOI21_X1 U6651 ( .B1(n6877), .B2(n6933), .A(n5910), .ZN(n5911) );
  NOR2_X1 U6652 ( .A1(n6417), .A2(n6335), .ZN(n5912) );
  NOR2_X1 U6653 ( .A1(n6351), .A2(n5912), .ZN(n6325) );
  OAI211_X1 U6654 ( .C1(n6303), .C2(n6417), .A(n6325), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U6655 ( .A1(n6325), .A2(n6417), .ZN(n6293) );
  NAND3_X1 U6656 ( .A1(n6308), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6293), .ZN(n5913) );
  NAND2_X1 U6657 ( .A1(n6924), .A2(REIP_REG_30__SCAN_IN), .ZN(n5919) );
  NAND3_X1 U6658 ( .A1(n5914), .A2(n5913), .A3(n5919), .ZN(n5915) );
  AOI21_X1 U6659 ( .B1(n5916), .B2(n6932), .A(n5915), .ZN(n5917) );
  OAI21_X1 U6660 ( .B1(n5924), .B2(n6892), .A(n5917), .ZN(U2988) );
  NAND2_X1 U6661 ( .A1(n6805), .A2(n5918), .ZN(n5920) );
  OAI211_X1 U6662 ( .C1(n5921), .C2(n6287), .A(n5920), .B(n5919), .ZN(n5922)
         );
  OAI21_X1 U6663 ( .B1(n5924), .B2(n7108), .A(n5923), .ZN(U2956) );
  NAND3_X1 U6664 ( .A1(n5928), .A2(n7157), .A3(n5925), .ZN(n5926) );
  OAI21_X1 U6665 ( .B1(n5928), .B2(n5927), .A(n5926), .ZN(n5929) );
  AOI21_X1 U6666 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(n5932) );
  OAI21_X1 U6667 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(U3465) );
  NAND2_X1 U6668 ( .A1(n6183), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U6669 ( .A(n6277), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6184)
         );
  NAND2_X1 U6670 ( .A1(n6184), .A2(n3509), .ZN(n5935) );
  AOI21_X1 U6671 ( .B1(n5936), .B2(n5899), .A(n5935), .ZN(n5937) );
  NAND2_X1 U6672 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  XNOR2_X1 U6673 ( .A(n5939), .B(n6295), .ZN(n6302) );
  AOI22_X1 U6674 ( .A1(n4041), .A2(EAX_REG_31__SCAN_IN), .B1(n5941), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5942) );
  INV_X1 U6675 ( .A(n5942), .ZN(n5943) );
  INV_X1 U6676 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U6677 ( .A1(n6912), .A2(n6754), .ZN(n6300) );
  AOI21_X1 U6678 ( .B1(n6809), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6300), 
        .ZN(n5945) );
  OAI21_X1 U6679 ( .B1(n6815), .B2(n5946), .A(n5945), .ZN(n5947) );
  AOI21_X1 U6680 ( .B1(n5975), .B2(n4644), .A(n5947), .ZN(n5948) );
  OAI21_X1 U6681 ( .B1(n6302), .B2(n7108), .A(n5948), .ZN(U2955) );
  OAI22_X1 U6682 ( .A1(n5949), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3455), .ZN(n5953) );
  NAND2_X1 U6683 ( .A1(n5975), .A2(n7105), .ZN(n5963) );
  NAND4_X1 U6684 ( .A1(n5954), .A2(n5979), .A3(EBX_REG_31__SCAN_IN), .A4(n7144), .ZN(n5955) );
  OAI21_X1 U6685 ( .B1(n7097), .B2(n5956), .A(n5955), .ZN(n5960) );
  INV_X1 U6686 ( .A(n5957), .ZN(n6022) );
  NOR2_X1 U6687 ( .A1(n7041), .A2(n6022), .ZN(n6010) );
  NAND2_X1 U6688 ( .A1(n6010), .A2(n5958), .ZN(n5999) );
  NOR4_X1 U6689 ( .A1(n5999), .A2(REIP_REG_31__SCAN_IN), .A3(n6551), .A4(n6750), .ZN(n5959) );
  AOI211_X1 U6690 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5961), .A(n5960), .B(n5959), .ZN(n5962) );
  OAI211_X1 U6691 ( .C1(n6292), .C2(n7083), .A(n5963), .B(n5962), .ZN(U2796)
         );
  INV_X1 U6692 ( .A(n5964), .ZN(n5972) );
  AOI22_X1 U6693 ( .A1(n5967), .A2(n6441), .B1(n5966), .B2(n5965), .ZN(n5970)
         );
  OAI222_X1 U6694 ( .A1(n7160), .A2(n5972), .B1(n5971), .B2(n5970), .C1(n5969), 
        .C2(n5968), .ZN(U3456) );
  NAND3_X1 U6695 ( .A1(n5975), .A2(n5974), .A3(n5973), .ZN(n5977) );
  AOI22_X1 U6696 ( .A1(n7205), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7208), .ZN(n5976) );
  NAND2_X1 U6697 ( .A1(n5977), .A2(n5976), .ZN(U2860) );
  INV_X1 U6698 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6623) );
  NAND2_X1 U6699 ( .A1(n5978), .A2(n6623), .ZN(n5981) );
  NOR2_X1 U6700 ( .A1(n5980), .A2(n5979), .ZN(n5991) );
  MUX2_X1 U6701 ( .A(n5981), .B(n5991), .S(n6831), .Z(U3474) );
  OR2_X1 U6702 ( .A1(n5985), .A2(n5982), .ZN(n5987) );
  NAND2_X1 U6703 ( .A1(n5983), .A2(n4518), .ZN(n5984) );
  NAND2_X1 U6704 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  OAI211_X1 U6705 ( .C1(n5989), .C2(n5988), .A(n5987), .B(n5986), .ZN(n7134)
         );
  NOR2_X1 U6706 ( .A1(n5991), .A2(n5990), .ZN(n6829) );
  OAI21_X1 U6707 ( .B1(READY_N), .B2(n6829), .A(n5992), .ZN(n7131) );
  AND2_X1 U6708 ( .A1(n7131), .A2(n5993), .ZN(n7109) );
  MUX2_X1 U6709 ( .A(MORE_REG_SCAN_IN), .B(n7134), .S(n7109), .Z(U3471) );
  AOI21_X1 U6710 ( .B1(n5995), .B2(n5842), .A(n5994), .ZN(n6189) );
  INV_X1 U6711 ( .A(n6189), .ZN(n6135) );
  OAI22_X1 U6712 ( .A1(n5996), .A2(n7097), .B1(n7061), .B2(n6187), .ZN(n5997)
         );
  AOI21_X1 U6713 ( .B1(n7079), .B2(EBX_REG_29__SCAN_IN), .A(n5997), .ZN(n5998)
         );
  OAI21_X1 U6714 ( .B1(n5999), .B2(REIP_REG_29__SCAN_IN), .A(n5998), .ZN(n6004) );
  OR2_X1 U6715 ( .A1(n6009), .A2(n6000), .ZN(n6001) );
  NAND2_X1 U6716 ( .A1(n6002), .A2(n6001), .ZN(n6304) );
  NOR2_X1 U6717 ( .A1(n6304), .A2(n7083), .ZN(n6003) );
  AOI211_X1 U6718 ( .C1(n6011), .C2(REIP_REG_29__SCAN_IN), .A(n6004), .B(n6003), .ZN(n6005) );
  OAI21_X1 U6719 ( .B1(n6135), .B2(n7073), .A(n6005), .ZN(U2798) );
  NOR2_X1 U6720 ( .A1(n6006), .A2(n6007), .ZN(n6008) );
  INV_X1 U6721 ( .A(n6010), .ZN(n6054) );
  INV_X1 U6722 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6745) );
  NOR3_X1 U6723 ( .A1(n6054), .A2(n6745), .A3(n6025), .ZN(n6012) );
  OAI21_X1 U6724 ( .B1(n6012), .B2(REIP_REG_28__SCAN_IN), .A(n6011), .ZN(n6015) );
  AOI22_X1 U6725 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n7071), .B1(n7101), 
        .B2(n6013), .ZN(n6014) );
  OAI211_X1 U6726 ( .C1(n6137), .C2(n7094), .A(n6015), .B(n6014), .ZN(n6016)
         );
  AOI21_X1 U6727 ( .B1(n6313), .B2(n7104), .A(n6016), .ZN(n6017) );
  OAI21_X1 U6728 ( .B1(n6168), .B2(n7073), .A(n6017), .ZN(U2799) );
  NOR2_X1 U6729 ( .A1(n6030), .A2(n6018), .ZN(n6019) );
  OR2_X1 U6730 ( .A1(n6006), .A2(n6019), .ZN(n6321) );
  AOI21_X1 U6731 ( .B1(n6021), .B2(n6035), .A(n4448), .ZN(n6195) );
  NAND2_X1 U6732 ( .A1(n6195), .A2(n7105), .ZN(n6029) );
  NOR3_X1 U6733 ( .A1(n6979), .A2(n6022), .A3(n6025), .ZN(n6023) );
  NOR2_X1 U6734 ( .A1(n6980), .A2(n6023), .ZN(n6042) );
  AOI22_X1 U6735 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n7071), .B1(n7101), 
        .B2(n6198), .ZN(n6024) );
  OAI21_X1 U6736 ( .B1(n7094), .B2(n6138), .A(n6024), .ZN(n6027) );
  NOR3_X1 U6737 ( .A1(n6054), .A2(REIP_REG_27__SCAN_IN), .A3(n6025), .ZN(n6026) );
  AOI211_X1 U6738 ( .C1(n6042), .C2(REIP_REG_27__SCAN_IN), .A(n6027), .B(n6026), .ZN(n6028) );
  OAI211_X1 U6739 ( .C1(n7083), .C2(n6321), .A(n6029), .B(n6028), .ZN(U2800)
         );
  INV_X1 U6740 ( .A(n6030), .ZN(n6033) );
  NAND2_X1 U6741 ( .A1(n6050), .A2(n6031), .ZN(n6032) );
  NAND2_X1 U6742 ( .A1(n6033), .A2(n6032), .ZN(n6333) );
  INV_X1 U6743 ( .A(n6035), .ZN(n6036) );
  AOI21_X1 U6744 ( .B1(n6037), .B2(n6034), .A(n6036), .ZN(n6206) );
  NAND2_X1 U6745 ( .A1(n6206), .A2(n7105), .ZN(n6045) );
  INV_X1 U6746 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6742) );
  INV_X1 U6747 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U6748 ( .B1(n6054), .B2(n6742), .A(n6038), .ZN(n6043) );
  OAI22_X1 U6749 ( .A1(n6039), .A2(n7097), .B1(n7061), .B2(n6204), .ZN(n6041)
         );
  NOR2_X1 U6750 ( .A1(n7094), .A2(n6140), .ZN(n6040) );
  AOI211_X1 U6751 ( .C1(n6043), .C2(n6042), .A(n6041), .B(n6040), .ZN(n6044)
         );
  OAI211_X1 U6752 ( .C1(n7083), .C2(n6333), .A(n6045), .B(n6044), .ZN(U2801)
         );
  OAI21_X1 U6753 ( .B1(n6046), .B2(n6047), .A(n6034), .ZN(n6216) );
  INV_X1 U6754 ( .A(n6349), .ZN(n6049) );
  OAI21_X1 U6755 ( .B1(n6350), .B2(n6049), .A(n6048), .ZN(n6051) );
  NAND2_X1 U6756 ( .A1(n6051), .A2(n6050), .ZN(n6344) );
  INV_X1 U6757 ( .A(n6344), .ZN(n6058) );
  AOI22_X1 U6758 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n7071), .B1(n7101), 
        .B2(n6210), .ZN(n6053) );
  NAND2_X1 U6759 ( .A1(n7079), .A2(EBX_REG_25__SCAN_IN), .ZN(n6052) );
  OAI211_X1 U6760 ( .C1(n6054), .C2(REIP_REG_25__SCAN_IN), .A(n6053), .B(n6052), .ZN(n6057) );
  OAI21_X1 U6761 ( .B1(n6979), .B2(n7096), .A(n6055), .ZN(n7091) );
  NAND2_X1 U6762 ( .A1(n6124), .A2(n7092), .ZN(n7095) );
  AOI21_X1 U6763 ( .B1(n7091), .B2(n7095), .A(n6742), .ZN(n6056) );
  AOI211_X1 U6764 ( .C1(n6058), .C2(n7104), .A(n6057), .B(n6056), .ZN(n6059)
         );
  OAI21_X1 U6765 ( .B1(n6216), .B2(n7073), .A(n6059), .ZN(U2802) );
  INV_X1 U6766 ( .A(n6061), .ZN(n6062) );
  AOI21_X1 U6767 ( .B1(n6063), .B2(n6060), .A(n6062), .ZN(n7202) );
  INV_X1 U6768 ( .A(n7202), .ZN(n6151) );
  INV_X1 U6769 ( .A(n6080), .ZN(n6064) );
  NOR2_X1 U6770 ( .A1(n6065), .A2(n6064), .ZN(n7082) );
  OAI21_X1 U6771 ( .B1(n6157), .B2(n6066), .A(n6146), .ZN(n6149) );
  AOI22_X1 U6772 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n7071), .B1(n7101), 
        .B2(n6238), .ZN(n6068) );
  NAND2_X1 U6773 ( .A1(n7079), .A2(EBX_REG_22__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U6774 ( .C1(n6149), .C2(n7083), .A(n6068), .B(n6067), .ZN(n6075)
         );
  INV_X1 U6775 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6069) );
  NAND3_X1 U6776 ( .A1(n6071), .A2(n6080), .A3(n6069), .ZN(n7075) );
  AND2_X1 U6777 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  NOR2_X1 U6778 ( .A1(n6980), .A2(n6072), .ZN(n7069) );
  INV_X1 U6779 ( .A(n7069), .ZN(n6073) );
  AOI21_X1 U6780 ( .B1(n7075), .B2(n6073), .A(n6736), .ZN(n6074) );
  AOI211_X1 U6781 ( .C1(n6736), .C2(n7082), .A(n6075), .B(n6074), .ZN(n6076)
         );
  OAI21_X1 U6782 ( .B1(n6151), .B2(n7073), .A(n6076), .ZN(U2805) );
  NOR2_X1 U6783 ( .A1(n3439), .A2(n6078), .ZN(n6079) );
  OR2_X1 U6784 ( .A1(n6077), .A2(n6079), .ZN(n7194) );
  NAND2_X1 U6785 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6080), .ZN(n6097) );
  OAI21_X1 U6786 ( .B1(n6730), .B2(n6097), .A(n6733), .ZN(n6087) );
  INV_X1 U6787 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6081) );
  OAI22_X1 U6788 ( .A1(n6081), .A2(n7097), .B1(n6251), .B2(n7061), .ZN(n6086)
         );
  AOI21_X1 U6789 ( .B1(n6082), .B2(n6096), .A(n6155), .ZN(n6387) );
  INV_X1 U6790 ( .A(n6387), .ZN(n6084) );
  OAI22_X1 U6791 ( .A1(n6084), .A2(n7083), .B1(n7094), .B2(n6083), .ZN(n6085)
         );
  AOI211_X1 U6792 ( .C1(n6087), .C2(n7069), .A(n6086), .B(n6085), .ZN(n6088)
         );
  OAI21_X1 U6793 ( .B1(n7194), .B2(n7073), .A(n6088), .ZN(U2807) );
  AOI21_X1 U6794 ( .B1(n6089), .B2(n5759), .A(n3439), .ZN(n6261) );
  OAI221_X1 U6795 ( .B1(n6730), .B2(n6091), .C1(n6730), .C2(n6090), .A(n7051), 
        .ZN(n6102) );
  INV_X1 U6796 ( .A(n6092), .ZN(n6259) );
  NAND2_X1 U6797 ( .A1(n6094), .A2(n6093), .ZN(n6095) );
  AND2_X1 U6798 ( .A1(n6096), .A2(n6095), .ZN(n6837) );
  AOI22_X1 U6799 ( .A1(n7104), .A2(n6837), .B1(n7079), .B2(EBX_REG_19__SCAN_IN), .ZN(n6100) );
  INV_X1 U6800 ( .A(n6097), .ZN(n6098) );
  AOI22_X1 U6801 ( .A1(n7071), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6730), 
        .B2(n6098), .ZN(n6099) );
  OAI211_X1 U6802 ( .C1(n6259), .C2(n7061), .A(n6100), .B(n6099), .ZN(n6101)
         );
  AOI211_X1 U6803 ( .C1(n6261), .C2(n7105), .A(n6102), .B(n6101), .ZN(n6103)
         );
  INV_X1 U6804 ( .A(n6103), .ZN(U2808) );
  NAND2_X1 U6805 ( .A1(n6104), .A2(n7105), .ZN(n6113) );
  AOI22_X1 U6806 ( .A1(n7104), .A2(n6923), .B1(n7079), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n6112) );
  NAND2_X1 U6807 ( .A1(n7071), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6105)
         );
  OAI211_X1 U6808 ( .C1(n7061), .C2(n6106), .A(n6105), .B(n7051), .ZN(n6107)
         );
  NOR2_X1 U6809 ( .A1(n6108), .A2(n6107), .ZN(n6111) );
  NAND2_X1 U6810 ( .A1(n6109), .A2(REIP_REG_9__SCAN_IN), .ZN(n6110) );
  NAND4_X1 U6811 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(U2818)
         );
  NOR3_X1 U6812 ( .A1(n7041), .A2(REIP_REG_6__SCAN_IN), .A3(n6114), .ZN(n7008)
         );
  OAI21_X1 U6813 ( .B1(n7041), .B2(n6115), .A(n6957), .ZN(n7009) );
  OAI21_X1 U6814 ( .B1(n7008), .B2(n7009), .A(REIP_REG_7__SCAN_IN), .ZN(n6128)
         );
  NAND2_X1 U6815 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6115), .ZN(n6116) );
  NOR2_X1 U6816 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6116), .ZN(n6123) );
  AND2_X1 U6817 ( .A1(n6118), .A2(n6117), .ZN(n6120) );
  OR2_X1 U6818 ( .A1(n6120), .A2(n6119), .ZN(n6775) );
  INV_X1 U6819 ( .A(n6775), .ZN(n6901) );
  AOI22_X1 U6820 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n7071), .B1(n7104), 
        .B2(n6901), .ZN(n6121) );
  OAI211_X1 U6821 ( .C1(n7061), .C2(n6804), .A(n6121), .B(n7051), .ZN(n6122)
         );
  AOI21_X1 U6822 ( .B1(n6124), .B2(n6123), .A(n6122), .ZN(n6127) );
  INV_X1 U6823 ( .A(n6778), .ZN(n6801) );
  NAND2_X1 U6824 ( .A1(n6801), .A2(n7105), .ZN(n6126) );
  NAND2_X1 U6825 ( .A1(n7079), .A2(EBX_REG_7__SCAN_IN), .ZN(n6125) );
  NAND4_X1 U6826 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(U2820)
         );
  INV_X1 U6827 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6129) );
  OAI22_X1 U6828 ( .A1(n6292), .A2(n6776), .B1(n6785), .B2(n6129), .ZN(U2828)
         );
  INV_X1 U6829 ( .A(n6130), .ZN(n6133) );
  OAI222_X1 U6830 ( .A1(n6133), .A2(n6777), .B1(n6132), .B2(n6785), .C1(n6776), 
        .C2(n6131), .ZN(U2829) );
  OAI222_X1 U6831 ( .A1(n6777), .A2(n6135), .B1(n6134), .B2(n6785), .C1(n6304), 
        .C2(n6776), .ZN(U2830) );
  OAI222_X1 U6832 ( .A1(n6777), .A2(n6168), .B1(n6137), .B2(n6785), .C1(n6136), 
        .C2(n6776), .ZN(U2831) );
  INV_X1 U6833 ( .A(n6195), .ZN(n6139) );
  OAI222_X1 U6834 ( .A1(n6777), .A2(n6139), .B1(n6138), .B2(n6785), .C1(n6321), 
        .C2(n6776), .ZN(U2832) );
  INV_X1 U6835 ( .A(n6206), .ZN(n6141) );
  OAI222_X1 U6836 ( .A1(n6777), .A2(n6141), .B1(n6140), .B2(n6785), .C1(n6333), 
        .C2(n6776), .ZN(U2833) );
  INV_X1 U6837 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6142) );
  OAI222_X1 U6838 ( .A1(n6216), .A2(n6777), .B1(n6142), .B2(n6785), .C1(n6344), 
        .C2(n6776), .ZN(U2834) );
  NAND2_X1 U6839 ( .A1(n6061), .A2(n6143), .ZN(n6144) );
  NAND2_X1 U6840 ( .A1(n3436), .A2(n6144), .ZN(n7081) );
  INV_X1 U6841 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U6842 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  NAND2_X1 U6843 ( .A1(n6350), .A2(n6147), .ZN(n7084) );
  OAI222_X1 U6844 ( .A1(n6777), .A2(n7081), .B1(n6148), .B2(n6785), .C1(n7084), 
        .C2(n6776), .ZN(U2836) );
  INV_X1 U6845 ( .A(n6149), .ZN(n6369) );
  AOI22_X1 U6846 ( .A1(n6369), .A2(n6782), .B1(EBX_REG_22__SCAN_IN), .B2(n6159), .ZN(n6150) );
  OAI21_X1 U6847 ( .B1(n6151), .B2(n6777), .A(n6150), .ZN(U2837) );
  OR2_X1 U6848 ( .A1(n6077), .A2(n6152), .ZN(n6153) );
  NAND2_X1 U6849 ( .A1(n6060), .A2(n6153), .ZN(n7198) );
  NOR2_X1 U6850 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  OR2_X1 U6851 ( .A1(n6157), .A2(n6156), .ZN(n7072) );
  OAI222_X1 U6852 ( .A1(n7198), .A2(n6777), .B1(n6158), .B2(n6785), .C1(n6776), 
        .C2(n7072), .ZN(U2838) );
  AOI22_X1 U6853 ( .A1(n6387), .A2(n6782), .B1(EBX_REG_20__SCAN_IN), .B2(n6159), .ZN(n6160) );
  OAI21_X1 U6854 ( .B1(n7194), .B2(n6777), .A(n6160), .ZN(U2839) );
  INV_X1 U6855 ( .A(n6261), .ZN(n6181) );
  NOR2_X1 U6856 ( .A1(n6785), .A2(n6161), .ZN(n6162) );
  AOI21_X1 U6857 ( .B1(n6837), .B2(n6782), .A(n6162), .ZN(n6163) );
  OAI21_X1 U6858 ( .B1(n6181), .B2(n6777), .A(n6163), .ZN(U2840) );
  NAND2_X1 U6859 ( .A1(n6189), .A2(n7206), .ZN(n6165) );
  AOI22_X1 U6860 ( .A1(n7205), .A2(DATAI_29_), .B1(n7208), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6164) );
  OAI211_X1 U6861 ( .C1(n6173), .C2(n6590), .A(n6165), .B(n6164), .ZN(U2862)
         );
  AOI22_X1 U6862 ( .A1(n7205), .A2(DATAI_28_), .B1(n7208), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U6863 ( .A1(n7209), .A2(DATAI_12_), .ZN(n6166) );
  OAI211_X1 U6864 ( .C1(n6168), .C2(n6180), .A(n6167), .B(n6166), .ZN(U2863)
         );
  NAND2_X1 U6865 ( .A1(n6195), .A2(n7206), .ZN(n6170) );
  AOI22_X1 U6866 ( .A1(n7205), .A2(DATAI_27_), .B1(n7208), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6169) );
  OAI211_X1 U6867 ( .C1(n6173), .C2(n6598), .A(n6170), .B(n6169), .ZN(U2864)
         );
  NAND2_X1 U6868 ( .A1(n6206), .A2(n7206), .ZN(n6172) );
  AOI22_X1 U6869 ( .A1(n7205), .A2(DATAI_26_), .B1(n7208), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6171) );
  OAI211_X1 U6870 ( .C1(n6173), .C2(n6599), .A(n6172), .B(n6171), .ZN(U2865)
         );
  AOI22_X1 U6871 ( .A1(n7205), .A2(DATAI_25_), .B1(n7208), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U6872 ( .A1(n7209), .A2(DATAI_9_), .ZN(n6174) );
  OAI211_X1 U6873 ( .C1(n6216), .C2(n6180), .A(n6175), .B(n6174), .ZN(U2866)
         );
  AOI22_X1 U6874 ( .A1(n7205), .A2(DATAI_23_), .B1(n7208), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U6875 ( .A1(n7209), .A2(DATAI_7_), .ZN(n6176) );
  OAI211_X1 U6876 ( .C1(n7081), .C2(n6180), .A(n6177), .B(n6176), .ZN(U2868)
         );
  AOI22_X1 U6877 ( .A1(n7205), .A2(DATAI_19_), .B1(n7208), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U6878 ( .A1(n7209), .A2(DATAI_3_), .ZN(n6178) );
  OAI211_X1 U6879 ( .C1(n6181), .C2(n6180), .A(n6179), .B(n6178), .ZN(U2872)
         );
  XNOR2_X1 U6880 ( .A(n6185), .B(n6184), .ZN(n6310) );
  NOR2_X1 U6881 ( .A1(n6912), .A2(n6750), .ZN(n6306) );
  AOI21_X1 U6882 ( .B1(n6809), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6306), 
        .ZN(n6186) );
  OAI21_X1 U6883 ( .B1(n6187), .B2(n6815), .A(n6186), .ZN(n6188) );
  AOI21_X1 U6884 ( .B1(n6189), .B2(n4644), .A(n6188), .ZN(n6190) );
  OAI21_X1 U6885 ( .B1(n7108), .B2(n6310), .A(n6190), .ZN(U2957) );
  NAND2_X1 U6886 ( .A1(n3938), .A2(n6337), .ZN(n6192) );
  MUX2_X1 U6887 ( .A(n6193), .B(n6192), .S(n6191), .Z(n6194) );
  XNOR2_X1 U6888 ( .A(n6194), .B(n6324), .ZN(n6331) );
  NAND2_X1 U6889 ( .A1(n6195), .A2(n4644), .ZN(n6200) );
  NOR2_X1 U6890 ( .A1(n6912), .A2(n6745), .ZN(n6322) );
  NOR2_X1 U6891 ( .A1(n6287), .A2(n6196), .ZN(n6197) );
  AOI211_X1 U6892 ( .C1(n6805), .C2(n6198), .A(n6322), .B(n6197), .ZN(n6199)
         );
  OAI211_X1 U6893 ( .C1(n6331), .C2(n7108), .A(n6200), .B(n6199), .ZN(U2959)
         );
  XNOR2_X1 U6894 ( .A(n5895), .B(n6337), .ZN(n6202) );
  XNOR2_X1 U6895 ( .A(n6201), .B(n6202), .ZN(n6341) );
  NAND2_X1 U6896 ( .A1(n6924), .A2(REIP_REG_26__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U6897 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6203)
         );
  OAI211_X1 U6898 ( .C1(n6815), .C2(n6204), .A(n6332), .B(n6203), .ZN(n6205)
         );
  AOI21_X1 U6899 ( .B1(n6206), .B2(n4644), .A(n6205), .ZN(n6207) );
  OAI21_X1 U6900 ( .B1(n7108), .B2(n6341), .A(n6207), .ZN(U2960) );
  INV_X1 U6901 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U6902 ( .A1(n6924), .A2(REIP_REG_25__SCAN_IN), .ZN(n6343) );
  OAI21_X1 U6903 ( .B1(n6287), .B2(n6208), .A(n6343), .ZN(n6209) );
  AOI21_X1 U6904 ( .B1(n6805), .B2(n6210), .A(n6209), .ZN(n6215) );
  OAI21_X1 U6905 ( .B1(n6213), .B2(n6212), .A(n6211), .ZN(n6342) );
  NAND2_X1 U6906 ( .A1(n6342), .A2(n6810), .ZN(n6214) );
  OAI211_X1 U6907 ( .C1(n6216), .C2(n6291), .A(n6215), .B(n6214), .ZN(U2961)
         );
  XNOR2_X1 U6908 ( .A(n3938), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6256)
         );
  NOR2_X2 U6909 ( .A1(n6257), .A2(n6256), .ZN(n6255) );
  OAI21_X1 U6910 ( .B1(n6277), .B2(n6384), .A(n6255), .ZN(n6217) );
  XNOR2_X1 U6911 ( .A(n3938), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6242)
         );
  NAND3_X1 U6912 ( .A1(n6248), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6219) );
  NAND4_X1 U6913 ( .A1(n6255), .A2(n3938), .A3(n6218), .A4(n6384), .ZN(n6228)
         );
  OAI22_X1 U6914 ( .A1(n6235), .A2(n6219), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6228), .ZN(n6220) );
  XNOR2_X1 U6915 ( .A(n6220), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6358)
         );
  NOR2_X1 U6916 ( .A1(n6912), .A2(n7092), .ZN(n6356) );
  INV_X1 U6917 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n7098) );
  NOR2_X1 U6918 ( .A1(n6287), .A2(n7098), .ZN(n6221) );
  AOI211_X1 U6919 ( .C1(n6805), .C2(n7102), .A(n6356), .B(n6221), .ZN(n6224)
         );
  AOI21_X1 U6920 ( .B1(n6222), .B2(n3436), .A(n6046), .ZN(n7207) );
  NAND2_X1 U6921 ( .A1(n7207), .A2(n4644), .ZN(n6223) );
  OAI211_X1 U6922 ( .C1(n6358), .C2(n7108), .A(n6224), .B(n6223), .ZN(U2962)
         );
  NAND2_X1 U6923 ( .A1(n6277), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6266) );
  NOR2_X1 U6924 ( .A1(n6225), .A2(n6266), .ZN(n6394) );
  NAND3_X1 U6925 ( .A1(n6394), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6226), .ZN(n6227) );
  NAND2_X1 U6926 ( .A1(n6228), .A2(n6227), .ZN(n6229) );
  XNOR2_X1 U6927 ( .A(n6229), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6365)
         );
  NAND2_X1 U6928 ( .A1(n6924), .A2(REIP_REG_23__SCAN_IN), .ZN(n6359) );
  OAI21_X1 U6929 ( .B1(n6287), .B2(n7090), .A(n6359), .ZN(n6231) );
  NOR2_X1 U6930 ( .A1(n7081), .A2(n6291), .ZN(n6230) );
  AOI211_X1 U6931 ( .C1(n6805), .C2(n7080), .A(n6231), .B(n6230), .ZN(n6232)
         );
  OAI21_X1 U6932 ( .B1(n6365), .B2(n7108), .A(n6232), .ZN(U2963) );
  XNOR2_X1 U6933 ( .A(n5895), .B(n6233), .ZN(n6234) );
  XNOR2_X1 U6934 ( .A(n6235), .B(n6234), .ZN(n6374) );
  NOR2_X1 U6935 ( .A1(n6912), .A2(n6736), .ZN(n6368) );
  INV_X1 U6936 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6236) );
  NOR2_X1 U6937 ( .A1(n6287), .A2(n6236), .ZN(n6237) );
  AOI211_X1 U6938 ( .C1(n6805), .C2(n6238), .A(n6368), .B(n6237), .ZN(n6240)
         );
  NAND2_X1 U6939 ( .A1(n7202), .A2(n4644), .ZN(n6239) );
  OAI211_X1 U6940 ( .C1(n6374), .C2(n7108), .A(n6240), .B(n6239), .ZN(U2964)
         );
  INV_X1 U6941 ( .A(n6241), .ZN(n6376) );
  NAND2_X1 U6942 ( .A1(n6243), .A2(n6242), .ZN(n6375) );
  NAND3_X1 U6943 ( .A1(n6376), .A2(n6810), .A3(n6375), .ZN(n6247) );
  NAND2_X1 U6944 ( .A1(n6924), .A2(REIP_REG_21__SCAN_IN), .ZN(n6377) );
  OAI21_X1 U6945 ( .B1(n6287), .B2(n6244), .A(n6377), .ZN(n6245) );
  AOI21_X1 U6946 ( .B1(n6805), .B2(n7070), .A(n6245), .ZN(n6246) );
  OAI211_X1 U6947 ( .C1(n6291), .C2(n7198), .A(n6247), .B(n6246), .ZN(U2965)
         );
  NOR2_X1 U6948 ( .A1(n6255), .A2(n6841), .ZN(n6249) );
  MUX2_X1 U6949 ( .A(n6255), .B(n6249), .S(n6248), .Z(n6250) );
  XNOR2_X1 U6950 ( .A(n6250), .B(n6384), .ZN(n6383) );
  NAND2_X1 U6951 ( .A1(n6383), .A2(n6810), .ZN(n6254) );
  AND2_X1 U6952 ( .A1(n6924), .A2(REIP_REG_20__SCAN_IN), .ZN(n6386) );
  NOR2_X1 U6953 ( .A1(n6815), .A2(n6251), .ZN(n6252) );
  AOI211_X1 U6954 ( .C1(n6809), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n6386), 
        .B(n6252), .ZN(n6253) );
  OAI211_X1 U6955 ( .C1(n6291), .C2(n7194), .A(n6254), .B(n6253), .ZN(U2966)
         );
  AOI21_X1 U6956 ( .B1(n3430), .B2(n6256), .A(n6255), .ZN(n6836) );
  AOI22_X1 U6957 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6924), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U6958 ( .B1(n6259), .B2(n6815), .A(n6258), .ZN(n6260) );
  AOI21_X1 U6959 ( .B1(n6261), .B2(n4644), .A(n6260), .ZN(n6262) );
  OAI21_X1 U6960 ( .B1(n6836), .B2(n7108), .A(n6262), .ZN(U2967) );
  OAI21_X1 U6961 ( .B1(n5684), .B2(n6277), .A(n6225), .ZN(n6264) );
  NAND2_X1 U6962 ( .A1(n3938), .A2(n6400), .ZN(n6263) );
  NOR2_X1 U6963 ( .A1(n6264), .A2(n6263), .ZN(n6395) );
  INV_X1 U6964 ( .A(n6395), .ZN(n6268) );
  NAND2_X1 U6965 ( .A1(n6263), .A2(n6266), .ZN(n6265) );
  MUX2_X1 U6966 ( .A(n6266), .B(n6265), .S(n6264), .Z(n6267) );
  NAND2_X1 U6967 ( .A1(n6268), .A2(n6267), .ZN(n6405) );
  NAND2_X1 U6968 ( .A1(n6405), .A2(n6810), .ZN(n6274) );
  INV_X1 U6969 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6269) );
  NOR2_X1 U6970 ( .A1(n6912), .A2(n6269), .ZN(n6408) );
  NOR2_X1 U6971 ( .A1(n6287), .A2(n6270), .ZN(n6271) );
  AOI211_X1 U6972 ( .C1(n6805), .C2(n6272), .A(n6408), .B(n6271), .ZN(n6273)
         );
  OAI211_X1 U6973 ( .C1(n6291), .C2(n6275), .A(n6274), .B(n6273), .ZN(U2969)
         );
  MUX2_X1 U6974 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n5684), .S(n6277), 
        .Z(n6278) );
  XNOR2_X1 U6975 ( .A(n6276), .B(n6278), .ZN(n6426) );
  AOI22_X1 U6976 ( .A1(n6809), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6924), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n6279) );
  OAI21_X1 U6977 ( .B1(n6280), .B2(n6815), .A(n6279), .ZN(n6281) );
  AOI21_X1 U6978 ( .B1(n7185), .B2(n4644), .A(n6281), .ZN(n6282) );
  OAI21_X1 U6979 ( .B1(n6426), .B2(n7108), .A(n6282), .ZN(U2970) );
  OAI21_X1 U6980 ( .B1(n6285), .B2(n6284), .A(n6283), .ZN(n6427) );
  NAND2_X1 U6981 ( .A1(n6427), .A2(n6810), .ZN(n6290) );
  NOR2_X1 U6982 ( .A1(n6912), .A2(n7058), .ZN(n6431) );
  NOR2_X1 U6983 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  AOI211_X1 U6984 ( .C1(n6805), .C2(n7060), .A(n6431), .B(n6288), .ZN(n6289)
         );
  OAI211_X1 U6985 ( .C1(n6291), .C2(n7063), .A(n6290), .B(n6289), .ZN(U2971)
         );
  INV_X1 U6986 ( .A(n6308), .ZN(n6296) );
  INV_X1 U6987 ( .A(n6293), .ZN(n6294) );
  AOI211_X1 U6988 ( .C1(n6296), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6295), .B(n6294), .ZN(n6301) );
  INV_X1 U6989 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6297) );
  NOR4_X1 U6990 ( .A1(n6328), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6298), 
        .A4(n6297), .ZN(n6299) );
  INV_X1 U6991 ( .A(n6303), .ZN(n6314) );
  OAI21_X1 U6992 ( .B1(n6328), .B2(n6314), .A(n5899), .ZN(n6307) );
  NOR2_X1 U6993 ( .A1(n6304), .A2(n6915), .ZN(n6305) );
  AOI211_X1 U6994 ( .C1(n6308), .C2(n6307), .A(n6306), .B(n6305), .ZN(n6309)
         );
  OAI21_X1 U6995 ( .B1(n6310), .B2(n6892), .A(n6309), .ZN(U2989) );
  NAND2_X1 U6996 ( .A1(n6311), .A2(n6938), .ZN(n6320) );
  AOI21_X1 U6997 ( .B1(n6313), .B2(n6932), .A(n6312), .ZN(n6319) );
  OAI21_X1 U6998 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A(n6314), .ZN(n6315) );
  OR2_X1 U6999 ( .A1(n6328), .A2(n6315), .ZN(n6318) );
  OR2_X1 U7000 ( .A1(n6325), .A2(n6316), .ZN(n6317) );
  NAND4_X1 U7001 ( .A1(n6320), .A2(n6319), .A3(n6318), .A4(n6317), .ZN(U2990)
         );
  INV_X1 U7002 ( .A(n6321), .ZN(n6323) );
  AOI21_X1 U7003 ( .B1(n6323), .B2(n6932), .A(n6322), .ZN(n6327) );
  OR2_X1 U7004 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  OAI211_X1 U7005 ( .C1(n6328), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6327), .B(n6326), .ZN(n6329) );
  INV_X1 U7006 ( .A(n6329), .ZN(n6330) );
  OAI21_X1 U7007 ( .B1(n6331), .B2(n6892), .A(n6330), .ZN(U2991) );
  OAI21_X1 U7008 ( .B1(n6333), .B2(n6915), .A(n6332), .ZN(n6339) );
  INV_X1 U7009 ( .A(n6334), .ZN(n6348) );
  AOI211_X1 U7010 ( .C1(n6337), .C2(n6336), .A(n6335), .B(n6348), .ZN(n6338)
         );
  AOI211_X1 U7011 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n6351), .A(n6339), .B(n6338), .ZN(n6340) );
  OAI21_X1 U7012 ( .B1(n6341), .B2(n6892), .A(n6340), .ZN(U2992) );
  NAND2_X1 U7013 ( .A1(n6342), .A2(n6938), .ZN(n6347) );
  OAI21_X1 U7014 ( .B1(n6344), .B2(n6915), .A(n6343), .ZN(n6345) );
  AOI21_X1 U7015 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n6351), .A(n6345), 
        .ZN(n6346) );
  OAI211_X1 U7016 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n6348), .A(n6347), .B(n6346), .ZN(U2993) );
  XNOR2_X1 U7017 ( .A(n6350), .B(n6349), .ZN(n7103) );
  INV_X1 U7018 ( .A(n6351), .ZN(n6352) );
  AOI211_X1 U7019 ( .C1(n6354), .C2(n6360), .A(n6353), .B(n6352), .ZN(n6355)
         );
  AOI211_X1 U7020 ( .C1(n6932), .C2(n7103), .A(n6356), .B(n6355), .ZN(n6357)
         );
  OAI21_X1 U7021 ( .B1(n6358), .B2(n6892), .A(n6357), .ZN(U2994) );
  OAI21_X1 U7022 ( .B1(n7084), .B2(n6915), .A(n6359), .ZN(n6362) );
  NOR2_X1 U7023 ( .A1(n6360), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6361)
         );
  AOI211_X1 U7024 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n6363), .A(n6362), .B(n6361), .ZN(n6364) );
  OAI21_X1 U7025 ( .B1(n6365), .B2(n6892), .A(n6364), .ZN(U2995) );
  INV_X1 U7026 ( .A(n6835), .ZN(n6390) );
  INV_X1 U7027 ( .A(n6388), .ZN(n6370) );
  NOR4_X1 U7028 ( .A1(n6390), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n6370), 
        .A4(n6366), .ZN(n6367) );
  AOI211_X1 U7029 ( .C1(n6932), .C2(n6369), .A(n6368), .B(n6367), .ZN(n6373)
         );
  NOR3_X1 U7030 ( .A1(n6390), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n6370), 
        .ZN(n6378) );
  OR2_X1 U7031 ( .A1(n6417), .A2(n6388), .ZN(n6371) );
  NAND2_X1 U7032 ( .A1(n6842), .A2(n6371), .ZN(n6380) );
  OAI21_X1 U7033 ( .B1(n6378), .B2(n6380), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n6372) );
  OAI211_X1 U7034 ( .C1(n6374), .C2(n6892), .A(n6373), .B(n6372), .ZN(U2996)
         );
  NAND3_X1 U7035 ( .A1(n6376), .A2(n6938), .A3(n6375), .ZN(n6382) );
  OAI21_X1 U7036 ( .B1(n7072), .B2(n6915), .A(n6377), .ZN(n6379) );
  AOI211_X1 U7037 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n6380), .A(n6379), .B(n6378), .ZN(n6381) );
  NAND2_X1 U7038 ( .A1(n6382), .A2(n6381), .ZN(U2997) );
  INV_X1 U7039 ( .A(n6383), .ZN(n6393) );
  NOR2_X1 U7040 ( .A1(n6842), .A2(n6384), .ZN(n6385) );
  AOI211_X1 U7041 ( .C1(n6932), .C2(n6387), .A(n6386), .B(n6385), .ZN(n6392)
         );
  OR3_X1 U7042 ( .A1(n6390), .A2(n6389), .A3(n6388), .ZN(n6391) );
  OAI211_X1 U7043 ( .C1(n6393), .C2(n6892), .A(n6392), .B(n6391), .ZN(U2998)
         );
  NOR2_X1 U7044 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  XNOR2_X1 U7045 ( .A(n6396), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6811)
         );
  INV_X1 U7046 ( .A(n6811), .ZN(n6404) );
  NOR2_X1 U7047 ( .A1(n6400), .A2(n6410), .ZN(n6397) );
  OAI21_X1 U7048 ( .B1(n6417), .B2(n6397), .A(n6415), .ZN(n6409) );
  OAI22_X1 U7049 ( .A1(n6915), .A2(n6398), .B1(n6912), .B2(n6728), .ZN(n6399)
         );
  AOI21_X1 U7050 ( .B1(n6409), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6399), 
        .ZN(n6403) );
  NOR3_X1 U7051 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6400), .A3(n6410), 
        .ZN(n6401) );
  NAND2_X1 U7052 ( .A1(n6929), .A2(n6401), .ZN(n6402) );
  OAI211_X1 U7053 ( .C1(n6404), .C2(n6892), .A(n6403), .B(n6402), .ZN(U3000)
         );
  INV_X1 U7054 ( .A(n6405), .ZN(n6414) );
  NOR2_X1 U7055 ( .A1(n6915), .A2(n6406), .ZN(n6407) );
  AOI211_X1 U7056 ( .C1(n6409), .C2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6408), .B(n6407), .ZN(n6413) );
  NOR2_X1 U7057 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6410), .ZN(n6411)
         );
  NAND2_X1 U7058 ( .A1(n6929), .A2(n6411), .ZN(n6412) );
  OAI211_X1 U7059 ( .C1(n6414), .C2(n6892), .A(n6413), .B(n6412), .ZN(U3001)
         );
  OAI21_X1 U7060 ( .B1(n6417), .B2(n6416), .A(n6415), .ZN(n6430) );
  NAND2_X1 U7061 ( .A1(n6418), .A2(n6932), .ZN(n6423) );
  NOR3_X1 U7062 ( .A1(n6421), .A2(n6420), .A3(n6419), .ZN(n6429) );
  OAI221_X1 U7063 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n5684), .C2(n6428), .A(n6429), 
        .ZN(n6422) );
  OAI211_X1 U7064 ( .C1(n6726), .C2(n6912), .A(n6423), .B(n6422), .ZN(n6424)
         );
  AOI21_X1 U7065 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6430), .A(n6424), 
        .ZN(n6425) );
  OAI21_X1 U7066 ( .B1(n6426), .B2(n6892), .A(n6425), .ZN(U3002) );
  INV_X1 U7067 ( .A(n6427), .ZN(n6434) );
  AOI22_X1 U7068 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6430), .B1(n6429), .B2(n6428), .ZN(n6433) );
  AOI21_X1 U7069 ( .B1(n6932), .B2(n7056), .A(n6431), .ZN(n6432) );
  OAI211_X1 U7070 ( .C1(n6434), .C2(n6892), .A(n6433), .B(n6432), .ZN(U3003)
         );
  NAND3_X1 U7071 ( .A1(n6436), .A2(n6435), .A3(n6446), .ZN(n6437) );
  OAI21_X1 U7072 ( .B1(n6438), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n6437), 
        .ZN(n6439) );
  AOI21_X1 U7073 ( .B1(n4638), .B2(n6440), .A(n6439), .ZN(n7121) );
  INV_X1 U7074 ( .A(n6441), .ZN(n6449) );
  NOR2_X1 U7075 ( .A1(n6443), .A2(n6442), .ZN(n6444) );
  AOI22_X1 U7076 ( .A1(n6447), .A2(n6446), .B1(n6445), .B2(n6444), .ZN(n6448)
         );
  OAI21_X1 U7077 ( .B1(n7121), .B2(n6449), .A(n6448), .ZN(n6450) );
  MUX2_X1 U7078 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n6450), .S(n7114), 
        .Z(U3460) );
  INV_X1 U7079 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6452) );
  AOI21_X1 U7080 ( .B1(n6451), .B2(STATE_REG_1__SCAN_IN), .A(n7177), .ZN(n6456) );
  INV_X1 U7081 ( .A(BS16_N), .ZN(n6616) );
  NAND2_X1 U7082 ( .A1(n6451), .A2(n7177), .ZN(n6817) );
  AOI21_X1 U7083 ( .B1(n6616), .B2(n6817), .A(n6453), .ZN(n7167) );
  AOI21_X1 U7084 ( .B1(n6452), .B2(n6453), .A(n7167), .ZN(U3451) );
  AND2_X1 U7085 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6453), .ZN(U3180) );
  AND2_X1 U7086 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6453), .ZN(U3179) );
  AND2_X1 U7087 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6453), .ZN(U3178) );
  AND2_X1 U7088 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6453), .ZN(U3177) );
  AND2_X1 U7089 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6453), .ZN(U3176) );
  AND2_X1 U7090 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6453), .ZN(U3175) );
  AND2_X1 U7091 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6453), .ZN(U3174) );
  AND2_X1 U7092 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6453), .ZN(U3173) );
  AND2_X1 U7093 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6453), .ZN(U3172) );
  AND2_X1 U7094 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6453), .ZN(U3171) );
  AND2_X1 U7095 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6453), .ZN(U3170) );
  AND2_X1 U7096 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6453), .ZN(U3169) );
  AND2_X1 U7097 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6453), .ZN(U3168) );
  AND2_X1 U7098 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6453), .ZN(U3167) );
  AND2_X1 U7099 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6453), .ZN(U3166) );
  AND2_X1 U7100 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6453), .ZN(U3165) );
  AND2_X1 U7101 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6453), .ZN(U3164) );
  AND2_X1 U7102 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6453), .ZN(U3163) );
  AND2_X1 U7103 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6453), .ZN(U3162) );
  AND2_X1 U7104 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6453), .ZN(U3161) );
  AND2_X1 U7105 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6453), .ZN(U3160) );
  AND2_X1 U7106 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6453), .ZN(U3159) );
  AND2_X1 U7107 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6453), .ZN(U3158) );
  AND2_X1 U7108 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6453), .ZN(U3157) );
  AND2_X1 U7109 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6453), .ZN(U3156) );
  AND2_X1 U7110 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6453), .ZN(U3155) );
  AND2_X1 U7111 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6453), .ZN(U3154) );
  AND2_X1 U7112 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6453), .ZN(U3153) );
  AND2_X1 U7113 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6453), .ZN(U3152) );
  AND2_X1 U7114 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6453), .ZN(U3151) );
  AND2_X1 U7115 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6454), .ZN(U3019)
         );
  AND2_X1 U7116 ( .A1(n6455), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7117 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6519) );
  AOI21_X1 U7118 ( .B1(n6456), .B2(n6519), .A(n7183), .ZN(U2789) );
  OAI22_X1 U7119 ( .A1(n6733), .A2(keyinput_62), .B1(keyinput_61), .B2(
        REIP_REG_21__SCAN_IN), .ZN(n6457) );
  AOI221_X1 U7120 ( .B1(n6733), .B2(keyinput_62), .C1(REIP_REG_21__SCAN_IN), 
        .C2(keyinput_61), .A(n6457), .ZN(n6661) );
  INV_X1 U7121 ( .A(keyinput_60), .ZN(n6546) );
  OAI22_X1 U7122 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_51), .B1(
        REIP_REG_29__SCAN_IN), .B2(keyinput_53), .ZN(n6458) );
  AOI221_X1 U7123 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_51), .C1(
        keyinput_53), .C2(REIP_REG_29__SCAN_IN), .A(n6458), .ZN(n6535) );
  INV_X1 U7124 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6460) );
  OAI22_X1 U7125 ( .A1(n6460), .A2(keyinput_50), .B1(keyinput_48), .B2(
        BYTEENABLE_REG_1__SCAN_IN), .ZN(n6459) );
  AOI221_X1 U7126 ( .B1(n6460), .B2(keyinput_50), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_48), .A(n6459), .ZN(n6534) );
  OAI22_X1 U7127 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_52), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .ZN(n6461) );
  AOI221_X1 U7128 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_52), .C1(
        keyinput_49), .C2(BYTEENABLE_REG_2__SCAN_IN), .A(n6461), .ZN(n6533) );
  INV_X1 U7129 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7130 ( .A1(n6819), .A2(keyinput_42), .B1(n6463), .B2(keyinput_43), 
        .ZN(n6462) );
  OAI221_X1 U7131 ( .B1(n6819), .B2(keyinput_42), .C1(n6463), .C2(keyinput_43), 
        .A(n6462), .ZN(n6531) );
  OAI22_X1 U7132 ( .A1(n6623), .A2(keyinput_37), .B1(HOLD), .B2(keyinput_36), 
        .ZN(n6464) );
  AOI221_X1 U7133 ( .B1(n6623), .B2(keyinput_37), .C1(keyinput_36), .C2(HOLD), 
        .A(n6464), .ZN(n6522) );
  INV_X1 U7134 ( .A(keyinput_35), .ZN(n6517) );
  INV_X1 U7135 ( .A(keyinput_30), .ZN(n6509) );
  INV_X1 U7136 ( .A(keyinput_25), .ZN(n6501) );
  INV_X1 U7137 ( .A(keyinput_18), .ZN(n6491) );
  INV_X1 U7138 ( .A(keyinput_17), .ZN(n6489) );
  INV_X1 U7139 ( .A(keyinput_16), .ZN(n6487) );
  INV_X1 U7140 ( .A(keyinput_15), .ZN(n6485) );
  INV_X1 U7141 ( .A(DATAI_16_), .ZN(n6582) );
  INV_X1 U7142 ( .A(keyinput_14), .ZN(n6483) );
  INV_X1 U7143 ( .A(DATAI_17_), .ZN(n6579) );
  INV_X1 U7144 ( .A(DATAI_18_), .ZN(n6575) );
  INV_X1 U7145 ( .A(keyinput_13), .ZN(n6481) );
  OAI22_X1 U7146 ( .A1(n6573), .A2(keyinput_11), .B1(keyinput_10), .B2(
        DATAI_21_), .ZN(n6465) );
  AOI221_X1 U7147 ( .B1(n6573), .B2(keyinput_11), .C1(DATAI_21_), .C2(
        keyinput_10), .A(n6465), .ZN(n6478) );
  AOI22_X1 U7148 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n6466) );
  OAI221_X1 U7149 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n6466), .ZN(n6471) );
  AOI22_X1 U7150 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(n4651), .B2(keyinput_3), .ZN(n6467) );
  OAI221_X1 U7151 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(n4651), .C2(
        keyinput_3), .A(n6467), .ZN(n6470) );
  AOI22_X1 U7152 ( .A1(n4656), .A2(keyinput_2), .B1(keyinput_4), .B2(n4645), 
        .ZN(n6468) );
  OAI221_X1 U7153 ( .B1(n4656), .B2(keyinput_2), .C1(n4645), .C2(keyinput_4), 
        .A(n6468), .ZN(n6469) );
  NOR3_X1 U7154 ( .A1(n6471), .A2(n6470), .A3(n6469), .ZN(n6476) );
  AOI22_X1 U7155 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(n6563), .B2(keyinput_6), .ZN(n6472) );
  OAI221_X1 U7156 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(n6563), .C2(
        keyinput_6), .A(n6472), .ZN(n6475) );
  OAI22_X1 U7157 ( .A1(n6566), .A2(keyinput_8), .B1(keyinput_9), .B2(DATAI_22_), .ZN(n6473) );
  AOI221_X1 U7158 ( .B1(n6566), .B2(keyinput_8), .C1(DATAI_22_), .C2(
        keyinput_9), .A(n6473), .ZN(n6474) );
  OAI21_X1 U7159 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(n6477) );
  OAI211_X1 U7160 ( .C1(DATAI_19_), .C2(keyinput_12), .A(n6478), .B(n6477), 
        .ZN(n6479) );
  AOI21_X1 U7161 ( .B1(DATAI_19_), .B2(keyinput_12), .A(n6479), .ZN(n6480) );
  AOI221_X1 U7162 ( .B1(DATAI_18_), .B2(keyinput_13), .C1(n6575), .C2(n6481), 
        .A(n6480), .ZN(n6482) );
  AOI221_X1 U7163 ( .B1(DATAI_17_), .B2(n6483), .C1(n6579), .C2(keyinput_14), 
        .A(n6482), .ZN(n6484) );
  AOI221_X1 U7164 ( .B1(DATAI_16_), .B2(n6485), .C1(n6582), .C2(keyinput_15), 
        .A(n6484), .ZN(n6486) );
  AOI221_X1 U7165 ( .B1(DATAI_15_), .B2(keyinput_16), .C1(n6584), .C2(n6487), 
        .A(n6486), .ZN(n6488) );
  AOI221_X1 U7166 ( .B1(DATAI_14_), .B2(keyinput_17), .C1(n6587), .C2(n6489), 
        .A(n6488), .ZN(n6490) );
  AOI221_X1 U7167 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(n6590), .C2(n6491), 
        .A(n6490), .ZN(n6498) );
  AOI22_X1 U7168 ( .A1(DATAI_10_), .A2(keyinput_21), .B1(DATAI_11_), .B2(
        keyinput_20), .ZN(n6492) );
  OAI221_X1 U7169 ( .B1(DATAI_10_), .B2(keyinput_21), .C1(DATAI_11_), .C2(
        keyinput_20), .A(n6492), .ZN(n6497) );
  AOI22_X1 U7170 ( .A1(DATAI_9_), .A2(keyinput_22), .B1(n6593), .B2(
        keyinput_19), .ZN(n6493) );
  OAI221_X1 U7171 ( .B1(DATAI_9_), .B2(keyinput_22), .C1(n6593), .C2(
        keyinput_19), .A(n6493), .ZN(n6496) );
  AOI22_X1 U7172 ( .A1(n6596), .A2(keyinput_24), .B1(n6594), .B2(keyinput_23), 
        .ZN(n6494) );
  OAI221_X1 U7173 ( .B1(n6596), .B2(keyinput_24), .C1(n6594), .C2(keyinput_23), 
        .A(n6494), .ZN(n6495) );
  NOR4_X1 U7174 ( .A1(n6498), .A2(n6497), .A3(n6496), .A4(n6495), .ZN(n6499)
         );
  AOI221_X1 U7175 ( .B1(DATAI_6_), .B2(n6501), .C1(n6500), .C2(keyinput_25), 
        .A(n6499), .ZN(n6507) );
  AOI22_X1 U7176 ( .A1(n6606), .A2(keyinput_28), .B1(n6503), .B2(keyinput_27), 
        .ZN(n6502) );
  OAI221_X1 U7177 ( .B1(n6606), .B2(keyinput_28), .C1(n6503), .C2(keyinput_27), 
        .A(n6502), .ZN(n6506) );
  AOI22_X1 U7178 ( .A1(DATAI_2_), .A2(keyinput_29), .B1(DATAI_5_), .B2(
        keyinput_26), .ZN(n6504) );
  OAI221_X1 U7179 ( .B1(DATAI_2_), .B2(keyinput_29), .C1(DATAI_5_), .C2(
        keyinput_26), .A(n6504), .ZN(n6505) );
  NOR3_X1 U7180 ( .A1(n6507), .A2(n6506), .A3(n6505), .ZN(n6508) );
  AOI221_X1 U7181 ( .B1(DATAI_1_), .B2(keyinput_30), .C1(n6614), .C2(n6509), 
        .A(n6508), .ZN(n6515) );
  AOI22_X1 U7182 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_32), .B1(n6511), 
        .B2(keyinput_31), .ZN(n6510) );
  OAI221_X1 U7183 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_32), .C1(n6511), 
        .C2(keyinput_31), .A(n6510), .ZN(n6514) );
  INV_X1 U7184 ( .A(NA_N), .ZN(n7174) );
  OAI22_X1 U7185 ( .A1(n6616), .A2(keyinput_34), .B1(n7174), .B2(keyinput_33), 
        .ZN(n6512) );
  AOI221_X1 U7186 ( .B1(n6616), .B2(keyinput_34), .C1(keyinput_33), .C2(n7174), 
        .A(n6512), .ZN(n6513) );
  OAI21_X1 U7187 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6516) );
  OAI221_X1 U7188 ( .B1(READY_N), .B2(keyinput_35), .C1(n7176), .C2(n6517), 
        .A(n6516), .ZN(n6521) );
  AOI22_X1 U7189 ( .A1(n6519), .A2(keyinput_38), .B1(n6625), .B2(keyinput_39), 
        .ZN(n6518) );
  OAI221_X1 U7190 ( .B1(n6519), .B2(keyinput_38), .C1(n6625), .C2(keyinput_39), 
        .A(n6518), .ZN(n6520) );
  AOI21_X1 U7191 ( .B1(n6522), .B2(n6521), .A(n6520), .ZN(n6525) );
  XOR2_X1 U7192 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_40), .Z(n6524) );
  INV_X1 U7193 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6633) );
  XOR2_X1 U7194 ( .A(n6633), .B(keyinput_41), .Z(n6523) );
  OAI21_X1 U7195 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6530) );
  OAI22_X1 U7196 ( .A1(n7133), .A2(keyinput_45), .B1(keyinput_47), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6526) );
  AOI221_X1 U7197 ( .B1(n7133), .B2(keyinput_45), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_47), .A(n6526), .ZN(n6529) );
  OAI22_X1 U7198 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_44), .B1(
        W_R_N_REG_SCAN_IN), .B2(keyinput_46), .ZN(n6527) );
  AOI221_X1 U7199 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_44), .C1(keyinput_46), 
        .C2(W_R_N_REG_SCAN_IN), .A(n6527), .ZN(n6528) );
  OAI211_X1 U7200 ( .C1(n6531), .C2(n6530), .A(n6529), .B(n6528), .ZN(n6532)
         );
  NAND4_X1 U7201 ( .A1(n6535), .A2(n6534), .A3(n6533), .A4(n6532), .ZN(n6540)
         );
  OAI22_X1 U7202 ( .A1(n6537), .A2(keyinput_54), .B1(keyinput_55), .B2(
        REIP_REG_27__SCAN_IN), .ZN(n6536) );
  AOI221_X1 U7203 ( .B1(n6537), .B2(keyinput_54), .C1(REIP_REG_27__SCAN_IN), 
        .C2(keyinput_55), .A(n6536), .ZN(n6539) );
  NOR2_X1 U7204 ( .A1(keyinput_57), .A2(REIP_REG_25__SCAN_IN), .ZN(n6538) );
  AOI221_X1 U7205 ( .B1(n6540), .B2(n6539), .C1(REIP_REG_25__SCAN_IN), .C2(
        keyinput_57), .A(n6538), .ZN(n6543) );
  OAI22_X1 U7206 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_58), .B1(
        keyinput_56), .B2(REIP_REG_26__SCAN_IN), .ZN(n6541) );
  AOI221_X1 U7207 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_58), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_56), .A(n6541), .ZN(n6542) );
  AOI22_X1 U7208 ( .A1(n6543), .A2(n6542), .B1(keyinput_59), .B2(
        REIP_REG_23__SCAN_IN), .ZN(n6544) );
  OAI21_X1 U7209 ( .B1(keyinput_59), .B2(REIP_REG_23__SCAN_IN), .A(n6544), 
        .ZN(n6545) );
  OAI221_X1 U7210 ( .B1(REIP_REG_22__SCAN_IN), .B2(n6546), .C1(n6736), .C2(
        keyinput_60), .A(n6545), .ZN(n6660) );
  XNOR2_X1 U7211 ( .A(n6736), .B(keyinput_124), .ZN(n6653) );
  AOI22_X1 U7212 ( .A1(n7092), .A2(keyinput_122), .B1(keyinput_121), .B2(n6742), .ZN(n6547) );
  OAI221_X1 U7213 ( .B1(n7092), .B2(keyinput_122), .C1(n6742), .C2(
        keyinput_121), .A(n6547), .ZN(n6648) );
  OAI22_X1 U7214 ( .A1(n6745), .A2(keyinput_119), .B1(keyinput_118), .B2(
        REIP_REG_28__SCAN_IN), .ZN(n6548) );
  AOI221_X1 U7215 ( .B1(n6745), .B2(keyinput_119), .C1(REIP_REG_28__SCAN_IN), 
        .C2(keyinput_118), .A(n6548), .ZN(n6645) );
  OAI22_X1 U7216 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_115), .B1(
        keyinput_112), .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6549) );
  AOI221_X1 U7217 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_115), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_112), .A(n6549), .ZN(n6643)
         );
  OAI22_X1 U7218 ( .A1(n6551), .A2(keyinput_116), .B1(keyinput_114), .B2(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6550) );
  AOI221_X1 U7219 ( .B1(n6551), .B2(keyinput_116), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_114), .A(n6550), .ZN(n6642)
         );
  INV_X1 U7220 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6768) );
  OAI22_X1 U7221 ( .A1(n6750), .A2(keyinput_117), .B1(n6768), .B2(keyinput_113), .ZN(n6552) );
  AOI221_X1 U7222 ( .B1(n6750), .B2(keyinput_117), .C1(keyinput_113), .C2(
        n6768), .A(n6552), .ZN(n6641) );
  XOR2_X1 U7223 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_104), .Z(n6630) );
  INV_X1 U7224 ( .A(keyinput_99), .ZN(n6621) );
  OAI22_X1 U7225 ( .A1(DATAI_0_), .A2(keyinput_95), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_96), .ZN(n6553) );
  AOI221_X1 U7226 ( .B1(DATAI_0_), .B2(keyinput_95), .C1(keyinput_96), .C2(
        MEMORYFETCH_REG_SCAN_IN), .A(n6553), .ZN(n6619) );
  INV_X1 U7227 ( .A(keyinput_94), .ZN(n6613) );
  INV_X1 U7228 ( .A(keyinput_82), .ZN(n6591) );
  INV_X1 U7229 ( .A(keyinput_81), .ZN(n6588) );
  INV_X1 U7230 ( .A(keyinput_80), .ZN(n6585) );
  INV_X1 U7231 ( .A(keyinput_79), .ZN(n6581) );
  INV_X1 U7232 ( .A(keyinput_78), .ZN(n6578) );
  INV_X1 U7233 ( .A(keyinput_77), .ZN(n6576) );
  OAI22_X1 U7234 ( .A1(n6555), .A2(keyinput_76), .B1(DATAI_21_), .B2(
        keyinput_74), .ZN(n6554) );
  AOI221_X1 U7235 ( .B1(n6555), .B2(keyinput_76), .C1(keyinput_74), .C2(
        DATAI_21_), .A(n6554), .ZN(n6571) );
  AOI22_X1 U7236 ( .A1(DATAI_28_), .A2(keyinput_67), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n6556) );
  OAI221_X1 U7237 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n6556), .ZN(n6561) );
  AOI22_X1 U7238 ( .A1(DATAI_26_), .A2(keyinput_69), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n6557) );
  OAI221_X1 U7239 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(DATAI_30_), .C2(
        keyinput_65), .A(n6557), .ZN(n6560) );
  AOI22_X1 U7240 ( .A1(DATAI_27_), .A2(keyinput_68), .B1(DATAI_29_), .B2(
        keyinput_66), .ZN(n6558) );
  OAI221_X1 U7241 ( .B1(DATAI_27_), .B2(keyinput_68), .C1(DATAI_29_), .C2(
        keyinput_66), .A(n6558), .ZN(n6559) );
  NOR3_X1 U7242 ( .A1(n6561), .A2(n6560), .A3(n6559), .ZN(n6569) );
  AOI22_X1 U7243 ( .A1(DATAI_24_), .A2(keyinput_71), .B1(n6563), .B2(
        keyinput_70), .ZN(n6562) );
  OAI221_X1 U7244 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(n6563), .C2(
        keyinput_70), .A(n6562), .ZN(n6568) );
  OAI22_X1 U7245 ( .A1(n6566), .A2(keyinput_72), .B1(n6565), .B2(keyinput_73), 
        .ZN(n6564) );
  AOI221_X1 U7246 ( .B1(n6566), .B2(keyinput_72), .C1(keyinput_73), .C2(n6565), 
        .A(n6564), .ZN(n6567) );
  OAI21_X1 U7247 ( .B1(n6569), .B2(n6568), .A(n6567), .ZN(n6570) );
  OAI211_X1 U7248 ( .C1(n6573), .C2(keyinput_75), .A(n6571), .B(n6570), .ZN(
        n6572) );
  AOI21_X1 U7249 ( .B1(n6573), .B2(keyinput_75), .A(n6572), .ZN(n6574) );
  AOI221_X1 U7250 ( .B1(DATAI_18_), .B2(n6576), .C1(n6575), .C2(keyinput_77), 
        .A(n6574), .ZN(n6577) );
  AOI221_X1 U7251 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(n6579), .C2(n6578), 
        .A(n6577), .ZN(n6580) );
  AOI221_X1 U7252 ( .B1(DATAI_16_), .B2(keyinput_79), .C1(n6582), .C2(n6581), 
        .A(n6580), .ZN(n6583) );
  AOI221_X1 U7253 ( .B1(DATAI_15_), .B2(n6585), .C1(n6584), .C2(keyinput_80), 
        .A(n6583), .ZN(n6586) );
  AOI221_X1 U7254 ( .B1(DATAI_14_), .B2(n6588), .C1(n6587), .C2(keyinput_81), 
        .A(n6586), .ZN(n6589) );
  AOI221_X1 U7255 ( .B1(DATAI_13_), .B2(n6591), .C1(n6590), .C2(keyinput_82), 
        .A(n6589), .ZN(n6603) );
  AOI22_X1 U7256 ( .A1(n6594), .A2(keyinput_87), .B1(n6593), .B2(keyinput_83), 
        .ZN(n6592) );
  OAI221_X1 U7257 ( .B1(n6594), .B2(keyinput_87), .C1(n6593), .C2(keyinput_83), 
        .A(n6592), .ZN(n6602) );
  AOI22_X1 U7258 ( .A1(DATAI_9_), .A2(keyinput_86), .B1(n6596), .B2(
        keyinput_88), .ZN(n6595) );
  OAI221_X1 U7259 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(n6596), .C2(
        keyinput_88), .A(n6595), .ZN(n6601) );
  AOI22_X1 U7260 ( .A1(n6599), .A2(keyinput_85), .B1(n6598), .B2(keyinput_84), 
        .ZN(n6597) );
  OAI221_X1 U7261 ( .B1(n6599), .B2(keyinput_85), .C1(n6598), .C2(keyinput_84), 
        .A(n6597), .ZN(n6600) );
  NOR4_X1 U7262 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n6611)
         );
  XOR2_X1 U7263 ( .A(keyinput_89), .B(DATAI_6_), .Z(n6610) );
  OAI22_X1 U7264 ( .A1(n6606), .A2(keyinput_92), .B1(n6605), .B2(keyinput_93), 
        .ZN(n6604) );
  AOI221_X1 U7265 ( .B1(n6606), .B2(keyinput_92), .C1(keyinput_93), .C2(n6605), 
        .A(n6604), .ZN(n6609) );
  OAI22_X1 U7266 ( .A1(DATAI_5_), .A2(keyinput_90), .B1(keyinput_91), .B2(
        DATAI_4_), .ZN(n6607) );
  AOI221_X1 U7267 ( .B1(DATAI_5_), .B2(keyinput_90), .C1(DATAI_4_), .C2(
        keyinput_91), .A(n6607), .ZN(n6608) );
  OAI211_X1 U7268 ( .C1(n6611), .C2(n6610), .A(n6609), .B(n6608), .ZN(n6612)
         );
  OAI221_X1 U7269 ( .B1(DATAI_1_), .B2(keyinput_94), .C1(n6614), .C2(n6613), 
        .A(n6612), .ZN(n6618) );
  AOI22_X1 U7270 ( .A1(NA_N), .A2(keyinput_97), .B1(n6616), .B2(keyinput_98), 
        .ZN(n6615) );
  OAI221_X1 U7271 ( .B1(NA_N), .B2(keyinput_97), .C1(n6616), .C2(keyinput_98), 
        .A(n6615), .ZN(n6617) );
  AOI21_X1 U7272 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(n6620) );
  AOI221_X1 U7273 ( .B1(READY_N), .B2(keyinput_99), .C1(n7176), .C2(n6621), 
        .A(n6620), .ZN(n6628) );
  AOI22_X1 U7274 ( .A1(keyinput_100), .A2(HOLD), .B1(n6623), .B2(keyinput_101), 
        .ZN(n6622) );
  OAI221_X1 U7275 ( .B1(keyinput_100), .B2(HOLD), .C1(n6623), .C2(keyinput_101), .A(n6622), .ZN(n6627) );
  OAI22_X1 U7276 ( .A1(n6625), .A2(keyinput_103), .B1(keyinput_102), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6624) );
  AOI221_X1 U7277 ( .B1(n6625), .B2(keyinput_103), .C1(ADS_N_REG_SCAN_IN), 
        .C2(keyinput_102), .A(n6624), .ZN(n6626) );
  OAI21_X1 U7278 ( .B1(n6628), .B2(n6627), .A(n6626), .ZN(n6629) );
  AOI22_X1 U7279 ( .A1(n6630), .A2(n6629), .B1(STATEBS16_REG_SCAN_IN), .B2(
        keyinput_107), .ZN(n6631) );
  OAI21_X1 U7280 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_107), .A(n6631), 
        .ZN(n6639) );
  AOI22_X1 U7281 ( .A1(keyinput_106), .A2(REQUESTPENDING_REG_SCAN_IN), .B1(
        n6633), .B2(keyinput_105), .ZN(n6632) );
  OAI221_X1 U7282 ( .B1(keyinput_106), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(
        n6633), .C2(keyinput_105), .A(n6632), .ZN(n6638) );
  INV_X1 U7283 ( .A(MORE_REG_SCAN_IN), .ZN(n7132) );
  OAI22_X1 U7284 ( .A1(n7133), .A2(keyinput_109), .B1(n7132), .B2(keyinput_108), .ZN(n6634) );
  AOI221_X1 U7285 ( .B1(n7133), .B2(keyinput_109), .C1(keyinput_108), .C2(
        n7132), .A(n6634), .ZN(n6637) );
  INV_X1 U7286 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6818) );
  OAI22_X1 U7287 ( .A1(n6818), .A2(keyinput_110), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_111), .ZN(n6635) );
  AOI221_X1 U7288 ( .B1(n6818), .B2(keyinput_110), .C1(keyinput_111), .C2(
        BYTEENABLE_REG_0__SCAN_IN), .A(n6635), .ZN(n6636) );
  OAI211_X1 U7289 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n6636), .ZN(n6640)
         );
  NAND4_X1 U7290 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6644)
         );
  AOI22_X1 U7291 ( .A1(n6645), .A2(n6644), .B1(REIP_REG_26__SCAN_IN), .B2(
        keyinput_120), .ZN(n6646) );
  OAI21_X1 U7292 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_120), .A(n6646), 
        .ZN(n6647) );
  OAI22_X1 U7293 ( .A1(n6648), .A2(n6647), .B1(keyinput_123), .B2(
        REIP_REG_23__SCAN_IN), .ZN(n6649) );
  AOI21_X1 U7294 ( .B1(keyinput_123), .B2(REIP_REG_23__SCAN_IN), .A(n6649), 
        .ZN(n6652) );
  OAI22_X1 U7295 ( .A1(n6733), .A2(keyinput_126), .B1(keyinput_125), .B2(
        REIP_REG_21__SCAN_IN), .ZN(n6650) );
  AOI221_X1 U7296 ( .B1(n6733), .B2(keyinput_126), .C1(REIP_REG_21__SCAN_IN), 
        .C2(keyinput_125), .A(n6650), .ZN(n6651) );
  OAI21_X1 U7297 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n6655) );
  INV_X1 U7298 ( .A(keyinput_63), .ZN(n6657) );
  AOI21_X1 U7299 ( .B1(keyinput_127), .B2(n6655), .A(n6657), .ZN(n6658) );
  INV_X1 U7300 ( .A(keyinput_127), .ZN(n6654) );
  AOI21_X1 U7301 ( .B1(n6655), .B2(n6654), .A(REIP_REG_19__SCAN_IN), .ZN(n6656) );
  AOI22_X1 U7302 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6658), .B1(n6657), .B2(
        n6656), .ZN(n6659) );
  AOI21_X1 U7303 ( .B1(n6661), .B2(n6660), .A(n6659), .ZN(n6671) );
  AOI22_X1 U7304 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6809), .B1(n6924), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U7305 ( .A1(n6663), .A2(n6662), .ZN(n6665) );
  XNOR2_X1 U7306 ( .A(n6665), .B(n6664), .ZN(n6881) );
  OR2_X1 U7307 ( .A1(n6881), .A2(n7108), .ZN(n6667) );
  NAND2_X1 U7308 ( .A1(n6960), .A2(n4644), .ZN(n6666) );
  AND2_X1 U7309 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  OAI211_X1 U7310 ( .C1(n6815), .C2(n6967), .A(n6669), .B(n6668), .ZN(n6670)
         );
  XOR2_X1 U7311 ( .A(n6671), .B(n6670), .Z(U2984) );
  AOI22_X1 U7312 ( .A1(n6699), .A2(LWORD_REG_0__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6673) );
  OAI21_X1 U7313 ( .B1(n6674), .B2(n6701), .A(n6673), .ZN(U2923) );
  AOI22_X1 U7314 ( .A1(n6699), .A2(LWORD_REG_1__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6675) );
  OAI21_X1 U7315 ( .B1(n6676), .B2(n6701), .A(n6675), .ZN(U2922) );
  AOI22_X1 U7316 ( .A1(n6699), .A2(LWORD_REG_2__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6677) );
  OAI21_X1 U7317 ( .B1(n6678), .B2(n6701), .A(n6677), .ZN(U2921) );
  AOI22_X1 U7318 ( .A1(n6699), .A2(LWORD_REG_3__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U7319 ( .B1(n6680), .B2(n6701), .A(n6679), .ZN(U2920) );
  AOI22_X1 U7320 ( .A1(n6699), .A2(LWORD_REG_4__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6681) );
  OAI21_X1 U7321 ( .B1(n6682), .B2(n6701), .A(n6681), .ZN(U2919) );
  AOI22_X1 U7322 ( .A1(n6699), .A2(LWORD_REG_5__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6683) );
  OAI21_X1 U7323 ( .B1(n4047), .B2(n6701), .A(n6683), .ZN(U2918) );
  AOI22_X1 U7324 ( .A1(n6699), .A2(LWORD_REG_6__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6684) );
  OAI21_X1 U7325 ( .B1(n4053), .B2(n6701), .A(n6684), .ZN(U2917) );
  AOI22_X1 U7326 ( .A1(n6699), .A2(LWORD_REG_7__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6685) );
  OAI21_X1 U7327 ( .B1(n4063), .B2(n6701), .A(n6685), .ZN(U2916) );
  AOI22_X1 U7328 ( .A1(n6699), .A2(LWORD_REG_8__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6686) );
  OAI21_X1 U7329 ( .B1(n6687), .B2(n6701), .A(n6686), .ZN(U2915) );
  AOI22_X1 U7330 ( .A1(n6699), .A2(LWORD_REG_9__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U7331 ( .B1(n6689), .B2(n6701), .A(n6688), .ZN(U2914) );
  AOI22_X1 U7332 ( .A1(n6699), .A2(LWORD_REG_10__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6690) );
  OAI21_X1 U7333 ( .B1(n6691), .B2(n6701), .A(n6690), .ZN(U2913) );
  AOI22_X1 U7334 ( .A1(n6699), .A2(LWORD_REG_11__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6692) );
  OAI21_X1 U7335 ( .B1(n6693), .B2(n6701), .A(n6692), .ZN(U2912) );
  AOI22_X1 U7336 ( .A1(n6699), .A2(LWORD_REG_12__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6694) );
  OAI21_X1 U7337 ( .B1(n4129), .B2(n6701), .A(n6694), .ZN(U2911) );
  AOI22_X1 U7338 ( .A1(n6699), .A2(LWORD_REG_13__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6695) );
  OAI21_X1 U7339 ( .B1(n6696), .B2(n6701), .A(n6695), .ZN(U2910) );
  AOI22_X1 U7340 ( .A1(n6699), .A2(LWORD_REG_14__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6697) );
  OAI21_X1 U7341 ( .B1(n6698), .B2(n6701), .A(n6697), .ZN(U2909) );
  AOI22_X1 U7342 ( .A1(n6699), .A2(LWORD_REG_15__SCAN_IN), .B1(n6455), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6700) );
  OAI21_X1 U7343 ( .B1(n6702), .B2(n6701), .A(n6700), .ZN(U2908) );
  INV_X1 U7344 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6704) );
  INV_X2 U7345 ( .A(n7183), .ZN(n6740) );
  NOR2_X1 U7346 ( .A1(n6740), .A2(STATE_REG_2__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U7347 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7183), .ZN(n6749) );
  AOI22_X1 U7348 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6740), .ZN(n6703) );
  OAI21_X1 U7349 ( .B1(n6704), .B2(n6753), .A(n6703), .ZN(U3184) );
  INV_X1 U7350 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6853) );
  AOI22_X1 U7351 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6740), .ZN(n6705) );
  OAI21_X1 U7352 ( .B1(n6853), .B2(n6753), .A(n6705), .ZN(U3185) );
  AOI22_X1 U7353 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6740), .ZN(n6706) );
  OAI21_X1 U7354 ( .B1(n6707), .B2(n6753), .A(n6706), .ZN(U3186) );
  AOI22_X1 U7355 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6740), .ZN(n6708) );
  OAI21_X1 U7356 ( .B1(n6997), .B2(n6753), .A(n6708), .ZN(U3187) );
  AOI22_X1 U7357 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6740), .ZN(n6709) );
  OAI21_X1 U7358 ( .B1(n6710), .B2(n6753), .A(n6709), .ZN(U3188) );
  AOI22_X1 U7359 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6740), .ZN(n6711) );
  OAI21_X1 U7360 ( .B1(n6712), .B2(n6753), .A(n6711), .ZN(U3189) );
  AOI22_X1 U7361 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6740), .ZN(n6713) );
  OAI21_X1 U7362 ( .B1(n5587), .B2(n6753), .A(n6713), .ZN(U3190) );
  AOI22_X1 U7363 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6740), .ZN(n6714) );
  OAI21_X1 U7364 ( .B1(n6715), .B2(n6753), .A(n6714), .ZN(U3191) );
  AOI22_X1 U7365 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6740), .ZN(n6716) );
  OAI21_X1 U7366 ( .B1(n6913), .B2(n6753), .A(n6716), .ZN(U3192) );
  INV_X1 U7367 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U7368 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6740), .ZN(n6717) );
  OAI21_X1 U7369 ( .B1(n6719), .B2(n6753), .A(n6717), .ZN(U3193) );
  AOI22_X1 U7370 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6740), .ZN(n6718) );
  OAI21_X1 U7371 ( .B1(n6719), .B2(n6749), .A(n6718), .ZN(U3194) );
  AOI22_X1 U7372 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6740), .ZN(n6720) );
  OAI21_X1 U7373 ( .B1(n6722), .B2(n6753), .A(n6720), .ZN(U3195) );
  AOI22_X1 U7374 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6740), .ZN(n6721) );
  OAI21_X1 U7375 ( .B1(n6722), .B2(n6749), .A(n6721), .ZN(U3196) );
  AOI22_X1 U7376 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6740), .ZN(n6723) );
  OAI21_X1 U7377 ( .B1(n7058), .B2(n6753), .A(n6723), .ZN(U3197) );
  AOI22_X1 U7378 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6740), .ZN(n6724) );
  OAI21_X1 U7379 ( .B1(n6726), .B2(n6753), .A(n6724), .ZN(U3198) );
  AOI22_X1 U7380 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6740), .ZN(n6725) );
  OAI21_X1 U7381 ( .B1(n6726), .B2(n6749), .A(n6725), .ZN(U3199) );
  AOI22_X1 U7382 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6740), .ZN(n6727) );
  OAI21_X1 U7383 ( .B1(n6728), .B2(n6753), .A(n6727), .ZN(U3200) );
  AOI22_X1 U7384 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6740), .ZN(n6729) );
  OAI21_X1 U7385 ( .B1(n6730), .B2(n6753), .A(n6729), .ZN(U3201) );
  AOI22_X1 U7386 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6740), .ZN(n6731) );
  OAI21_X1 U7387 ( .B1(n6733), .B2(n6753), .A(n6731), .ZN(U3202) );
  AOI22_X1 U7388 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6740), .ZN(n6732) );
  OAI21_X1 U7389 ( .B1(n6733), .B2(n6749), .A(n6732), .ZN(U3203) );
  AOI22_X1 U7390 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6740), .ZN(n6734) );
  OAI21_X1 U7391 ( .B1(n6736), .B2(n6753), .A(n6734), .ZN(U3204) );
  AOI22_X1 U7392 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6740), .ZN(n6735) );
  OAI21_X1 U7393 ( .B1(n6736), .B2(n6749), .A(n6735), .ZN(U3205) );
  AOI22_X1 U7394 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6740), .ZN(n6737) );
  OAI21_X1 U7395 ( .B1(n6738), .B2(n6749), .A(n6737), .ZN(U3206) );
  AOI22_X1 U7396 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6740), .ZN(n6739) );
  OAI21_X1 U7397 ( .B1(n6742), .B2(n6753), .A(n6739), .ZN(U3207) );
  AOI22_X1 U7398 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6740), .ZN(n6741) );
  OAI21_X1 U7399 ( .B1(n6742), .B2(n6749), .A(n6741), .ZN(U3208) );
  AOI22_X1 U7400 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6740), .ZN(n6743) );
  OAI21_X1 U7401 ( .B1(n6745), .B2(n6753), .A(n6743), .ZN(U3209) );
  AOI22_X1 U7402 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6740), .ZN(n6744) );
  OAI21_X1 U7403 ( .B1(n6745), .B2(n6749), .A(n6744), .ZN(U3210) );
  AOI22_X1 U7404 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6740), .ZN(n6746) );
  OAI21_X1 U7405 ( .B1(n6750), .B2(n6753), .A(n6746), .ZN(U3211) );
  AOI22_X1 U7406 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6747), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6740), .ZN(n6748) );
  OAI21_X1 U7407 ( .B1(n6750), .B2(n6749), .A(n6748), .ZN(U3212) );
  AOI22_X1 U7408 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6751), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6740), .ZN(n6752) );
  OAI21_X1 U7409 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(U3213) );
  MUX2_X1 U7410 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6740), .Z(U3445) );
  AOI221_X1 U7411 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6765) );
  NOR4_X1 U7412 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6758) );
  NOR4_X1 U7413 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6757) );
  NOR4_X1 U7414 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6756) );
  NOR4_X1 U7415 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6755) );
  NAND4_X1 U7416 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6764)
         );
  NOR4_X1 U7417 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6762) );
  AOI211_X1 U7418 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_31__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6761) );
  NOR4_X1 U7419 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6760) );
  NOR4_X1 U7420 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6759) );
  NAND4_X1 U7421 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6763)
         );
  NOR2_X1 U7422 ( .A1(n6764), .A2(n6763), .ZN(n6774) );
  MUX2_X1 U7423 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n6765), .S(n6774), .Z(
        U2795) );
  MUX2_X1 U7424 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6740), .Z(U3446) );
  AOI21_X1 U7425 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6766) );
  INV_X1 U7426 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6953) );
  OAI221_X1 U7427 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6766), .C1(n6953), .C2(
        REIP_REG_0__SCAN_IN), .A(n6774), .ZN(n6767) );
  OAI21_X1 U7428 ( .B1(n6774), .B2(n6768), .A(n6767), .ZN(U3468) );
  MUX2_X1 U7429 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6740), .Z(U3447) );
  INV_X1 U7430 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6771) );
  NOR3_X1 U7431 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6769) );
  OAI21_X1 U7432 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6769), .A(n6774), .ZN(n6770)
         );
  OAI21_X1 U7433 ( .B1(n6774), .B2(n6771), .A(n6770), .ZN(U2794) );
  MUX2_X1 U7434 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6740), .Z(U3448) );
  INV_X1 U7435 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6773) );
  OAI21_X1 U7436 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6774), .ZN(n6772) );
  OAI21_X1 U7437 ( .B1(n6774), .B2(n6773), .A(n6772), .ZN(U3469) );
  OAI22_X1 U7438 ( .A1(n6778), .A2(n6777), .B1(n6776), .B2(n6775), .ZN(n6779)
         );
  INV_X1 U7439 ( .A(n6779), .ZN(n6780) );
  OAI21_X1 U7440 ( .B1(n6785), .B2(n6781), .A(n6780), .ZN(U2852) );
  AOI22_X1 U7441 ( .A1(n7207), .A2(n6783), .B1(n6782), .B2(n7103), .ZN(n6784)
         );
  OAI21_X1 U7442 ( .B1(n6785), .B2(n7093), .A(n6784), .ZN(U2835) );
  AOI22_X1 U7443 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6809), .B1(n6924), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U7444 ( .A1(n6948), .A2(n4644), .ZN(n6786) );
  OAI21_X1 U7445 ( .B1(n7108), .B2(n6787), .A(n6786), .ZN(n6788) );
  INV_X1 U7446 ( .A(n6788), .ZN(n6789) );
  OAI211_X1 U7447 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6815), .A(n6790), 
        .B(n6789), .ZN(U2985) );
  AOI22_X1 U7448 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6809), .B1(n6924), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U7449 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  XNOR2_X1 U7450 ( .A(n6791), .B(n6794), .ZN(n6866) );
  AOI22_X1 U7451 ( .A1(n6866), .A2(n6810), .B1(n7017), .B2(n4644), .ZN(n6795)
         );
  OAI211_X1 U7452 ( .C1(n6815), .C2(n7019), .A(n6796), .B(n6795), .ZN(U2980)
         );
  AOI22_X1 U7453 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6809), .B1(n6924), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6803) );
  OAI21_X1 U7454 ( .B1(n6799), .B2(n6798), .A(n6797), .ZN(n6800) );
  INV_X1 U7455 ( .A(n6800), .ZN(n6903) );
  AOI22_X1 U7456 ( .A1(n6903), .A2(n6810), .B1(n4644), .B2(n6801), .ZN(n6802)
         );
  OAI211_X1 U7457 ( .C1(n6815), .C2(n6804), .A(n6803), .B(n6802), .ZN(U2979)
         );
  AOI22_X1 U7458 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6809), .B1(n6924), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6807) );
  AOI22_X1 U7459 ( .A1(n7024), .A2(n4644), .B1(n6805), .B2(n7023), .ZN(n6806)
         );
  OAI211_X1 U7460 ( .C1(n7108), .C2(n6808), .A(n6807), .B(n6806), .ZN(U2975)
         );
  AOI22_X1 U7461 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6809), .B1(n6924), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U7462 ( .A1(n6811), .A2(n6810), .B1(n4644), .B2(n7191), .ZN(n6812)
         );
  OAI211_X1 U7463 ( .C1(n6815), .C2(n6814), .A(n6813), .B(n6812), .ZN(U2968)
         );
  NOR2_X1 U7464 ( .A1(n7183), .A2(D_C_N_REG_SCAN_IN), .ZN(n6816) );
  AOI22_X1 U7465 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7183), .B1(n6817), .B2(
        n6816), .ZN(U2791) );
  AOI22_X1 U7466 ( .A1(n7183), .A2(READREQUEST_REG_SCAN_IN), .B1(n6818), .B2(
        n6740), .ZN(U3470) );
  AND2_X1 U7467 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7171) );
  NOR2_X1 U7468 ( .A1(n7177), .A2(n6819), .ZN(n7175) );
  AOI21_X1 U7469 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7175), .ZN(n6822)
         );
  NOR2_X1 U7470 ( .A1(n6820), .A2(n7176), .ZN(n7169) );
  INV_X1 U7471 ( .A(n7169), .ZN(n7181) );
  OAI211_X1 U7472 ( .C1(n7171), .C2(n6822), .A(n6821), .B(n7181), .ZN(U3182)
         );
  NOR2_X1 U7473 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6826) );
  NAND2_X1 U7474 ( .A1(READY_N), .A2(n6823), .ZN(n7153) );
  NAND3_X1 U7475 ( .A1(n7161), .A2(n7153), .A3(n7151), .ZN(n6825) );
  OAI21_X1 U7476 ( .B1(n6826), .B2(n6825), .A(n6824), .ZN(U3150) );
  OAI211_X1 U7477 ( .C1(n6827), .C2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .B(n7176), .ZN(n6828) );
  OAI21_X1 U7478 ( .B1(n6829), .B2(n6828), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6830) );
  NAND2_X1 U7479 ( .A1(n6830), .A2(n7161), .ZN(n6834) );
  AOI211_X1 U7480 ( .C1(n6699), .C2(n7176), .A(n6832), .B(n6831), .ZN(n6833)
         );
  MUX2_X1 U7481 ( .A(n6834), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6833), .Z(
        U3472) );
  AOI22_X1 U7482 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6924), .B1(n6835), .B2(
        n6841), .ZN(n6840) );
  INV_X1 U7483 ( .A(n6836), .ZN(n6838) );
  AOI22_X1 U7484 ( .A1(n6838), .A2(n6938), .B1(n6932), .B2(n6837), .ZN(n6839)
         );
  OAI211_X1 U7485 ( .C1(n6842), .C2(n6841), .A(n6840), .B(n6839), .ZN(U2999)
         );
  OAI211_X1 U7486 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6909), .B(n6852), .ZN(n6850) );
  NAND2_X1 U7487 ( .A1(n6843), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6846)
         );
  AOI21_X1 U7488 ( .B1(n6932), .B2(n6986), .A(n6844), .ZN(n6845) );
  OAI211_X1 U7489 ( .C1(n6847), .C2(n6892), .A(n6846), .B(n6845), .ZN(n6848)
         );
  INV_X1 U7490 ( .A(n6848), .ZN(n6849) );
  OAI21_X1 U7491 ( .B1(n6851), .B2(n6850), .A(n6849), .ZN(U3014) );
  NAND2_X1 U7492 ( .A1(n6909), .A2(n6852), .ZN(n6859) );
  INV_X1 U7493 ( .A(n6973), .ZN(n6855) );
  NOR2_X1 U7494 ( .A1(n6912), .A2(n6853), .ZN(n6854) );
  AOI21_X1 U7495 ( .B1(n6932), .B2(n6855), .A(n6854), .ZN(n6858) );
  NAND2_X1 U7496 ( .A1(n6856), .A2(n6938), .ZN(n6857) );
  OAI211_X1 U7497 ( .C1(n6859), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6858), 
        .B(n6857), .ZN(n6860) );
  INV_X1 U7498 ( .A(n6860), .ZN(n6861) );
  OAI21_X1 U7499 ( .B1(n6862), .B2(n3839), .A(n6861), .ZN(U3015) );
  NAND3_X1 U7500 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6863), .A3(n6909), 
        .ZN(n6870) );
  AOI211_X1 U7501 ( .C1(n6886), .C2(n3886), .A(n6865), .B(n6864), .ZN(n6868)
         );
  AOI222_X1 U7502 ( .A1(n6866), .A2(n6938), .B1(n6932), .B2(n7013), .C1(
        REIP_REG_6__SCAN_IN), .C2(n6924), .ZN(n6867) );
  OAI221_X1 U7503 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6870), .C1(n6869), .C2(n6868), .A(n6867), .ZN(U3012) );
  AOI21_X1 U7504 ( .B1(n6890), .B2(n6871), .A(n6887), .ZN(n6885) );
  INV_X1 U7505 ( .A(n6872), .ZN(n6874) );
  AOI21_X1 U7506 ( .B1(n6875), .B2(n6874), .A(n6873), .ZN(n6884) );
  NOR3_X1 U7507 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6877), .A3(n6876), 
        .ZN(n6878) );
  AOI21_X1 U7508 ( .B1(n6924), .B2(REIP_REG_2__SCAN_IN), .A(n6878), .ZN(n6880)
         );
  NAND2_X1 U7509 ( .A1(n6932), .A2(n6956), .ZN(n6879) );
  OAI211_X1 U7510 ( .C1(n6881), .C2(n6892), .A(n6880), .B(n6879), .ZN(n6882)
         );
  INV_X1 U7511 ( .A(n6882), .ZN(n6883) );
  OAI211_X1 U7512 ( .C1(n6885), .C2(n3803), .A(n6884), .B(n6883), .ZN(U3016)
         );
  AND2_X1 U7513 ( .A1(n6896), .A2(n6886), .ZN(n6888) );
  AOI211_X1 U7514 ( .C1(n6890), .C2(n6889), .A(n6888), .B(n6887), .ZN(n6907)
         );
  OAI222_X1 U7515 ( .A1(n6893), .A2(n6915), .B1(n6912), .B2(n5587), .C1(n6892), 
        .C2(n6891), .ZN(n6894) );
  INV_X1 U7516 ( .A(n6894), .ZN(n6899) );
  INV_X1 U7517 ( .A(n6909), .ZN(n6895) );
  NOR2_X1 U7518 ( .A1(n6896), .A2(n6895), .ZN(n6902) );
  OAI211_X1 U7519 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6902), .B(n6897), .ZN(n6898) );
  OAI211_X1 U7520 ( .C1(n6907), .C2(n6900), .A(n6899), .B(n6898), .ZN(U3010)
         );
  AOI22_X1 U7521 ( .A1(n6932), .A2(n6901), .B1(n6924), .B2(REIP_REG_7__SCAN_IN), .ZN(n6905) );
  AOI22_X1 U7522 ( .A1(n6903), .A2(n6938), .B1(n6902), .B2(n6906), .ZN(n6904)
         );
  OAI211_X1 U7523 ( .C1(n6907), .C2(n6906), .A(n6905), .B(n6904), .ZN(U3011)
         );
  INV_X1 U7524 ( .A(n6908), .ZN(n6918) );
  NAND2_X1 U7525 ( .A1(n6910), .A2(n6909), .ZN(n6928) );
  AOI211_X1 U7526 ( .C1(n6920), .C2(n6927), .A(n6911), .B(n6928), .ZN(n6917)
         );
  OAI22_X1 U7527 ( .A1(n6915), .A2(n6914), .B1(n6913), .B2(n6912), .ZN(n6916)
         );
  AOI211_X1 U7528 ( .C1(n6918), .C2(n6938), .A(n6917), .B(n6916), .ZN(n6919)
         );
  OAI21_X1 U7529 ( .B1(n6926), .B2(n6920), .A(n6919), .ZN(U3008) );
  INV_X1 U7530 ( .A(n6921), .ZN(n6922) );
  AOI222_X1 U7531 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6924), .B1(n6932), .B2(
        n6923), .C1(n6938), .C2(n6922), .ZN(n6925) );
  OAI221_X1 U7532 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6928), .C1(n6927), .C2(n6926), .A(n6925), .ZN(U3009) );
  NAND2_X1 U7533 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6929), .ZN(n6942) );
  AOI21_X1 U7534 ( .B1(n6932), .B2(n6931), .A(n6930), .ZN(n6941) );
  AOI21_X1 U7535 ( .B1(n6934), .B2(n6933), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6936) );
  OR2_X1 U7536 ( .A1(n6936), .A2(n6935), .ZN(n6937) );
  AOI22_X1 U7537 ( .A1(n6939), .A2(n6938), .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6937), .ZN(n6940) );
  OAI211_X1 U7538 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n6942), .A(n6941), .B(n6940), .ZN(U3006) );
  OR2_X1 U7539 ( .A1(n7041), .A2(REIP_REG_1__SCAN_IN), .ZN(n6958) );
  OR2_X1 U7540 ( .A1(n7083), .A2(n6943), .ZN(n6947) );
  OR2_X1 U7541 ( .A1(n6990), .A2(n6944), .ZN(n6946) );
  AOI22_X1 U7542 ( .A1(n7071), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6979), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6945) );
  AND4_X1 U7543 ( .A1(n6958), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n6950)
         );
  AOI22_X1 U7544 ( .A1(n7079), .A2(EBX_REG_1__SCAN_IN), .B1(n7003), .B2(n6948), 
        .ZN(n6949) );
  OAI211_X1 U7545 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n7061), .A(n6950), 
        .B(n6949), .ZN(U2826) );
  OAI22_X1 U7546 ( .A1(n6990), .A2(n6952), .B1(n7097), .B2(n6951), .ZN(n6955)
         );
  NOR3_X1 U7547 ( .A1(n7041), .A2(n6953), .A3(REIP_REG_2__SCAN_IN), .ZN(n6954)
         );
  AOI211_X1 U7548 ( .C1(n6956), .C2(n7104), .A(n6955), .B(n6954), .ZN(n6966)
         );
  NAND2_X1 U7549 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  NAND2_X1 U7550 ( .A1(n6959), .A2(REIP_REG_2__SCAN_IN), .ZN(n6962) );
  NAND2_X1 U7551 ( .A1(n7003), .A2(n6960), .ZN(n6961) );
  OAI211_X1 U7552 ( .C1(n7094), .C2(n6963), .A(n6962), .B(n6961), .ZN(n6964)
         );
  INV_X1 U7553 ( .A(n6964), .ZN(n6965) );
  OAI211_X1 U7554 ( .C1(n6967), .C2(n7061), .A(n6966), .B(n6965), .ZN(U2825)
         );
  OAI22_X1 U7555 ( .A1(n6969), .A2(n7097), .B1(n7061), .B2(n6968), .ZN(n6970)
         );
  INV_X1 U7556 ( .A(n6970), .ZN(n6977) );
  NAND2_X1 U7557 ( .A1(n7003), .A2(n6971), .ZN(n6976) );
  OR2_X1 U7558 ( .A1(n6990), .A2(n6972), .ZN(n6975) );
  OR2_X1 U7559 ( .A1(n7083), .A2(n6973), .ZN(n6974) );
  AND4_X1 U7560 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n6983)
         );
  NAND2_X1 U7561 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .ZN(
        n6978) );
  NOR2_X1 U7562 ( .A1(n6979), .A2(n6978), .ZN(n6981) );
  AOI21_X1 U7563 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6981), .A(n6980), .ZN(n6984)
         );
  OAI21_X1 U7564 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6981), .A(n6984), .ZN(n6982)
         );
  OAI211_X1 U7565 ( .C1(n7094), .C2(n4587), .A(n6983), .B(n6982), .ZN(U2824)
         );
  AOI22_X1 U7566 ( .A1(EBX_REG_4__SCAN_IN), .A2(n7079), .B1(
        REIP_REG_4__SCAN_IN), .B2(n6984), .ZN(n6995) );
  OAI21_X1 U7567 ( .B1(n7097), .B2(n4036), .A(n7051), .ZN(n6985) );
  AOI21_X1 U7568 ( .B1(n7104), .B2(n6986), .A(n6985), .ZN(n6989) );
  OR3_X1 U7569 ( .A1(n7041), .A2(REIP_REG_4__SCAN_IN), .A3(n6987), .ZN(n6988)
         );
  OAI211_X1 U7570 ( .C1(n6991), .C2(n6990), .A(n6989), .B(n6988), .ZN(n6992)
         );
  AOI21_X1 U7571 ( .B1(n6993), .B2(n7003), .A(n6992), .ZN(n6994) );
  OAI211_X1 U7572 ( .C1(n6996), .C2(n7061), .A(n6995), .B(n6994), .ZN(U2823)
         );
  OAI21_X1 U7573 ( .B1(n7041), .B2(n6998), .A(n6997), .ZN(n6999) );
  AOI22_X1 U7574 ( .A1(EBX_REG_5__SCAN_IN), .A2(n7079), .B1(n7009), .B2(n6999), 
        .ZN(n7007) );
  AOI22_X1 U7575 ( .A1(n7104), .A2(n7000), .B1(PHYADDRPOINTER_REG_5__SCAN_IN), 
        .B2(n7071), .ZN(n7006) );
  INV_X1 U7576 ( .A(n7001), .ZN(n7002) );
  AOI22_X1 U7577 ( .A1(n7004), .A2(n7003), .B1(n7002), .B2(n7101), .ZN(n7005)
         );
  NAND4_X1 U7578 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7051), .ZN(U2822)
         );
  INV_X1 U7579 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7011) );
  AOI211_X1 U7580 ( .C1(REIP_REG_6__SCAN_IN), .C2(n7009), .A(n7008), .B(n7057), 
        .ZN(n7010) );
  OAI21_X1 U7581 ( .B1(n7097), .B2(n7011), .A(n7010), .ZN(n7012) );
  AOI21_X1 U7582 ( .B1(n7104), .B2(n7013), .A(n7012), .ZN(n7014) );
  OAI21_X1 U7583 ( .B1(n7015), .B2(n7094), .A(n7014), .ZN(n7016) );
  AOI21_X1 U7584 ( .B1(n7105), .B2(n7017), .A(n7016), .ZN(n7018) );
  OAI21_X1 U7585 ( .B1(n7019), .B2(n7061), .A(n7018), .ZN(U2821) );
  AOI22_X1 U7586 ( .A1(n7021), .A2(n7020), .B1(REIP_REG_11__SCAN_IN), .B2(
        n7035), .ZN(n7028) );
  AOI22_X1 U7587 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7071), .B1(
        EBX_REG_11__SCAN_IN), .B2(n7079), .ZN(n7027) );
  AOI21_X1 U7588 ( .B1(n7104), .B2(n7022), .A(n7057), .ZN(n7026) );
  AOI22_X1 U7589 ( .A1(n7024), .A2(n7105), .B1(n7101), .B2(n7023), .ZN(n7025)
         );
  NAND4_X1 U7590 ( .A1(n7028), .A2(n7027), .A3(n7026), .A4(n7025), .ZN(U2816)
         );
  AOI22_X1 U7591 ( .A1(n7104), .A2(n7029), .B1(n7079), .B2(EBX_REG_13__SCAN_IN), .ZN(n7040) );
  NOR3_X1 U7592 ( .A1(n7041), .A2(REIP_REG_13__SCAN_IN), .A3(n7030), .ZN(n7031) );
  AOI211_X1 U7593 ( .C1(n7071), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n7057), 
        .B(n7031), .ZN(n7039) );
  OAI22_X1 U7594 ( .A1(n7033), .A2(n7073), .B1(n7032), .B2(n7061), .ZN(n7034)
         );
  INV_X1 U7595 ( .A(n7034), .ZN(n7038) );
  OAI21_X1 U7596 ( .B1(n7036), .B2(n7035), .A(REIP_REG_13__SCAN_IN), .ZN(n7037) );
  NAND4_X1 U7597 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), .ZN(U2814)
         );
  AOI22_X1 U7598 ( .A1(EBX_REG_14__SCAN_IN), .A2(n7079), .B1(
        REIP_REG_14__SCAN_IN), .B2(n7055), .ZN(n7054) );
  NOR2_X1 U7599 ( .A1(n7041), .A2(REIP_REG_14__SCAN_IN), .ZN(n7046) );
  OAI22_X1 U7600 ( .A1(n7083), .A2(n7043), .B1(n7042), .B2(n7097), .ZN(n7044)
         );
  AOI21_X1 U7601 ( .B1(n7046), .B2(n7045), .A(n7044), .ZN(n7053) );
  INV_X1 U7602 ( .A(n7047), .ZN(n7048) );
  OAI22_X1 U7603 ( .A1(n7049), .A2(n7073), .B1(n7061), .B2(n7048), .ZN(n7050)
         );
  INV_X1 U7604 ( .A(n7050), .ZN(n7052) );
  NAND4_X1 U7605 ( .A1(n7054), .A2(n7053), .A3(n7052), .A4(n7051), .ZN(U2813)
         );
  AOI22_X1 U7606 ( .A1(EBX_REG_15__SCAN_IN), .A2(n7079), .B1(
        REIP_REG_15__SCAN_IN), .B2(n7055), .ZN(n7068) );
  AOI22_X1 U7607 ( .A1(n7104), .A2(n7056), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .B2(n7071), .ZN(n7067) );
  AOI21_X1 U7608 ( .B1(n7059), .B2(n7058), .A(n7057), .ZN(n7066) );
  INV_X1 U7609 ( .A(n7060), .ZN(n7062) );
  OAI22_X1 U7610 ( .A1(n7063), .A2(n7073), .B1(n7062), .B2(n7061), .ZN(n7064)
         );
  INV_X1 U7611 ( .A(n7064), .ZN(n7065) );
  NAND4_X1 U7612 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), .ZN(U2812)
         );
  AOI22_X1 U7613 ( .A1(EBX_REG_21__SCAN_IN), .A2(n7079), .B1(
        REIP_REG_21__SCAN_IN), .B2(n7069), .ZN(n7078) );
  AOI22_X1 U7614 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n7071), .B1(n7070), 
        .B2(n7101), .ZN(n7077) );
  OAI22_X1 U7615 ( .A1(n7198), .A2(n7073), .B1(n7083), .B2(n7072), .ZN(n7074)
         );
  INV_X1 U7616 ( .A(n7074), .ZN(n7076) );
  NAND4_X1 U7617 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(U2806)
         );
  AOI22_X1 U7618 ( .A1(n7080), .A2(n7101), .B1(EBX_REG_23__SCAN_IN), .B2(n7079), .ZN(n7089) );
  INV_X1 U7619 ( .A(n7081), .ZN(n7087) );
  AOI21_X1 U7620 ( .B1(REIP_REG_22__SCAN_IN), .B2(n7082), .A(
        REIP_REG_23__SCAN_IN), .ZN(n7085) );
  OAI22_X1 U7621 ( .A1(n7091), .A2(n7085), .B1(n7084), .B2(n7083), .ZN(n7086)
         );
  AOI21_X1 U7622 ( .B1(n7087), .B2(n7105), .A(n7086), .ZN(n7088) );
  OAI211_X1 U7623 ( .C1(n7090), .C2(n7097), .A(n7089), .B(n7088), .ZN(U2804)
         );
  OAI22_X1 U7624 ( .A1(n7094), .A2(n7093), .B1(n7092), .B2(n7091), .ZN(n7100)
         );
  OAI22_X1 U7625 ( .A1(n7098), .A2(n7097), .B1(n7096), .B2(n7095), .ZN(n7099)
         );
  AOI211_X1 U7626 ( .C1(n7102), .C2(n7101), .A(n7100), .B(n7099), .ZN(n7107)
         );
  AOI22_X1 U7627 ( .A1(n7207), .A2(n7105), .B1(n7104), .B2(n7103), .ZN(n7106)
         );
  NAND2_X1 U7628 ( .A1(n7107), .A2(n7106), .ZN(U2803) );
  OAI21_X1 U7629 ( .B1(n7109), .B2(n7133), .A(n7108), .ZN(U2793) );
  INV_X1 U7630 ( .A(n7110), .ZN(n7112) );
  NAND3_X1 U7631 ( .A1(n7112), .A2(n5471), .A3(n7111), .ZN(n7113) );
  OAI21_X1 U7632 ( .B1(n7114), .B2(n4034), .A(n7113), .ZN(U3455) );
  NAND2_X1 U7633 ( .A1(n7115), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U7634 ( .A1(n7116), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7117) );
  NOR2_X1 U7635 ( .A1(n7118), .A2(n7117), .ZN(n7120) );
  INV_X1 U7636 ( .A(n7120), .ZN(n7125) );
  INV_X1 U7637 ( .A(n7119), .ZN(n7122) );
  OAI22_X1 U7638 ( .A1(n7122), .A2(n7121), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7120), .ZN(n7123) );
  OAI21_X1 U7639 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n7126) );
  AOI222_X1 U7640 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7127), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7126), .C1(n7127), .C2(n7126), 
        .ZN(n7130) );
  AOI222_X1 U7641 ( .A1(n7130), .A2(n7129), .B1(n7130), .B2(n7128), .C1(n7129), 
        .C2(n7128), .ZN(n7140) );
  AOI21_X1 U7642 ( .B1(n7133), .B2(n7132), .A(n7131), .ZN(n7135) );
  NOR4_X1 U7643 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n7134), .ZN(n7138)
         );
  OAI211_X1 U7644 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7140), .A(n7139), .B(n7138), .ZN(n7152) );
  OAI22_X1 U7645 ( .A1(n7152), .A2(n7164), .B1(n7141), .B2(n7176), .ZN(n7142)
         );
  OAI21_X1 U7646 ( .B1(n7144), .B2(n7143), .A(n7142), .ZN(n7158) );
  OAI21_X1 U7647 ( .B1(READY_N), .B2(n7145), .A(n7164), .ZN(n7148) );
  OAI21_X1 U7648 ( .B1(STATE2_REG_0__SCAN_IN), .B2(STATE2_REG_2__SCAN_IN), .A(
        STATE2_REG_1__SCAN_IN), .ZN(n7146) );
  AOI21_X1 U7649 ( .B1(n7153), .B2(n7158), .A(n7146), .ZN(n7147) );
  AOI21_X1 U7650 ( .B1(n7158), .B2(n7148), .A(n7147), .ZN(n7150) );
  NAND2_X1 U7651 ( .A1(n7150), .A2(n7149), .ZN(U3149) );
  OAI221_X1 U7652 ( .B1(n5471), .B2(STATE2_REG_0__SCAN_IN), .C1(n5471), .C2(
        n7158), .A(n7151), .ZN(U3453) );
  INV_X1 U7653 ( .A(n7152), .ZN(n7165) );
  AOI21_X1 U7654 ( .B1(n7158), .B2(n7153), .A(n7159), .ZN(n7154) );
  AOI211_X1 U7655 ( .C1(n7157), .C2(n7156), .A(n7155), .B(n7154), .ZN(n7163)
         );
  OAI211_X1 U7656 ( .C1(n7161), .C2(n7160), .A(n7159), .B(n7158), .ZN(n7162)
         );
  OAI211_X1 U7657 ( .C1(n7165), .C2(n7164), .A(n7163), .B(n7162), .ZN(U3148)
         );
  AOI21_X1 U7658 ( .B1(n6453), .B2(STATEBS16_REG_SCAN_IN), .A(n7167), .ZN(
        n7166) );
  INV_X1 U7659 ( .A(n7166), .ZN(U2792) );
  AOI21_X1 U7660 ( .B1(n6453), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n7167), .ZN(
        n7168) );
  INV_X1 U7661 ( .A(n7168), .ZN(U3452) );
  NAND2_X1 U7662 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7173) );
  AOI221_X1 U7663 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7174), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7179) );
  AOI221_X1 U7664 ( .B1(n7171), .B2(n7170), .C1(n7169), .C2(n7170), .A(n7179), 
        .ZN(n7172) );
  OAI221_X1 U7665 ( .B1(n7183), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7183), 
        .C2(n7173), .A(n7172), .ZN(U3181) );
  AOI21_X1 U7666 ( .B1(n7175), .B2(n7174), .A(STATE_REG_2__SCAN_IN), .ZN(n7182) );
  AOI221_X1 U7667 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7176), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7178) );
  AOI221_X1 U7668 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7178), .C2(HOLD), .A(n7177), .ZN(n7180) );
  OAI22_X1 U7669 ( .A1(n7182), .A2(n7181), .B1(n7180), .B2(n7179), .ZN(U3183)
         );
  OAI22_X1 U7670 ( .A1(n6740), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n7183), .ZN(n7184) );
  INV_X1 U7671 ( .A(n7184), .ZN(U3473) );
  AOI22_X1 U7672 ( .A1(n7185), .A2(n7206), .B1(n7205), .B2(DATAI_16_), .ZN(
        n7187) );
  AOI22_X1 U7673 ( .A1(n7209), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n7208), .ZN(n7186) );
  NAND2_X1 U7674 ( .A1(n7187), .A2(n7186), .ZN(U2875) );
  AOI22_X1 U7675 ( .A1(n7188), .A2(n7206), .B1(n7205), .B2(DATAI_17_), .ZN(
        n7190) );
  AOI22_X1 U7676 ( .A1(n7209), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7208), .ZN(n7189) );
  NAND2_X1 U7677 ( .A1(n7190), .A2(n7189), .ZN(U2874) );
  AOI22_X1 U7678 ( .A1(n7191), .A2(n7206), .B1(n7205), .B2(DATAI_18_), .ZN(
        n7193) );
  AOI22_X1 U7679 ( .A1(n7209), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n7208), .ZN(n7192) );
  NAND2_X1 U7680 ( .A1(n7193), .A2(n7192), .ZN(U2873) );
  INV_X1 U7681 ( .A(n7194), .ZN(n7195) );
  AOI22_X1 U7682 ( .A1(n7195), .A2(n7206), .B1(n7205), .B2(DATAI_20_), .ZN(
        n7197) );
  AOI22_X1 U7683 ( .A1(n7209), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n7208), .ZN(n7196) );
  NAND2_X1 U7684 ( .A1(n7197), .A2(n7196), .ZN(U2871) );
  INV_X1 U7685 ( .A(n7198), .ZN(n7199) );
  AOI22_X1 U7686 ( .A1(n7199), .A2(n7206), .B1(n7205), .B2(DATAI_21_), .ZN(
        n7201) );
  AOI22_X1 U7687 ( .A1(n7209), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7208), .ZN(n7200) );
  NAND2_X1 U7688 ( .A1(n7201), .A2(n7200), .ZN(U2870) );
  AOI22_X1 U7689 ( .A1(n7202), .A2(n7206), .B1(n7205), .B2(DATAI_22_), .ZN(
        n7204) );
  AOI22_X1 U7690 ( .A1(n7209), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7208), .ZN(n7203) );
  NAND2_X1 U7691 ( .A1(n7204), .A2(n7203), .ZN(U2869) );
  AOI22_X1 U7692 ( .A1(n7207), .A2(n7206), .B1(n7205), .B2(DATAI_24_), .ZN(
        n7211) );
  AOI22_X1 U7693 ( .A1(n7209), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n7208), .ZN(n7210) );
  NAND2_X1 U7694 ( .A1(n7211), .A2(n7210), .ZN(U2867) );
  NAND4_X2 U3493 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3661)
         );
  INV_X1 U4215 ( .A(n3736), .ZN(n3773) );
  CLKBUF_X1 U34730 ( .A(n4407), .Z(n5847) );
  CLKBUF_X1 U3482 ( .A(n3836), .Z(n5979) );
  CLKBUF_X1 U3495 ( .A(n5082), .Z(n5161) );
  CLKBUF_X1 U3496 ( .A(n5223), .Z(n3429) );
endmodule

