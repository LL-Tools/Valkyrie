

module b14_C_gen_AntiSAT_k_128_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702;

  OR2_X1 U2285 ( .A1(n3383), .A2(n3485), .ZN(n3384) );
  OR2_X1 U2286 ( .A1(n3075), .A2(n3074), .ZN(n3174) );
  INV_X2 U2287 ( .A(n2952), .ZN(n2903) );
  NAND2_X1 U2288 ( .A1(n4354), .A2(n2772), .ZN(n2337) );
  INV_X1 U2289 ( .A(n3681), .ZN(n3663) );
  AND2_X1 U2290 ( .A1(n2849), .A2(n2847), .ZN(n3662) );
  CLKBUF_X3 U2291 ( .A(n3682), .Z(n3645) );
  INV_X1 U2292 ( .A(n3662), .ZN(n3682) );
  INV_X1 U2293 ( .A(n3418), .ZN(n2549) );
  OAI21_X1 U2294 ( .B1(n4075), .B2(n2196), .A(n2194), .ZN(n4038) );
  NOR2_X1 U2295 ( .A1(n3293), .A2(n3281), .ZN(n3344) );
  NAND2_X1 U2296 ( .A1(n2776), .A2(IR_REG_31__SCAN_IN), .ZN(n2312) );
  XNOR2_X1 U2297 ( .A(n2312), .B(IR_REG_30__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U2298 ( .A1(n2582), .A2(n2581), .ZN(n4024) );
  NOR2_X2 U2299 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2392)
         );
  OAI21_X2 U2300 ( .B1(n2165), .B2(n2164), .A(n2163), .ZN(n2357) );
  XNOR2_X1 U2301 ( .A(n2634), .B(n3496), .ZN(n3962) );
  AND2_X1 U2302 ( .A1(n4026), .A2(n4016), .ZN(n4011) );
  OAI21_X1 U2303 ( .B1(n3046), .B2(n3045), .A(n3499), .ZN(n3066) );
  OR2_X1 U2304 ( .A1(n3027), .A2(n3022), .ZN(n3051) );
  AND2_X1 U2305 ( .A1(n3515), .A2(n3518), .ZN(n3476) );
  NAND2_X1 U2306 ( .A1(n3511), .A2(n3514), .ZN(n3475) );
  NAND2_X2 U2307 ( .A1(n2755), .A2(n4470), .ZN(n4473) );
  NAND2_X1 U2308 ( .A1(n2365), .A2(n2364), .ZN(n3860) );
  NAND2_X1 U2309 ( .A1(n2045), .A2(n2350), .ZN(n3864) );
  OR2_X1 U2310 ( .A1(n2808), .A2(n2807), .ZN(n2185) );
  INV_X1 U2311 ( .A(n3148), .ZN(n3859) );
  OR2_X2 U2312 ( .A1(n2345), .A2(n2344), .ZN(n3862) );
  NAND2_X1 U2313 ( .A1(n2105), .A2(n2355), .ZN(n3861) );
  NAND2_X1 U2314 ( .A1(n2340), .A2(n2339), .ZN(n2345) );
  AND4_X1 U2315 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n3148)
         );
  NAND2_X1 U2316 ( .A1(n2343), .A2(n2342), .ZN(n2344) );
  AOI21_X1 U2317 ( .B1(n2805), .B2(REG2_REG_4__SCAN_IN), .A(n2059), .ZN(n2808)
         );
  NAND2_X2 U2318 ( .A1(n2847), .A2(n2910), .ZN(n3681) );
  NAND2_X2 U2319 ( .A1(n2772), .A2(n2320), .ZN(n3418) );
  INV_X2 U2320 ( .A(n2341), .ZN(n3415) );
  INV_X1 U2321 ( .A(n2314), .ZN(n2772) );
  AOI21_X1 U2322 ( .B1(n3896), .B2(REG2_REG_3__SCAN_IN), .A(n2052), .ZN(n2803)
         );
  NAND2_X1 U2323 ( .A1(n2545), .A2(IR_REG_31__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U2324 ( .A1(n2229), .A2(n2057), .ZN(n2674) );
  NAND2_X1 U2325 ( .A1(n2801), .A2(n2802), .ZN(n3884) );
  XNOR2_X1 U2326 ( .A(n2088), .B(IR_REG_1__SCAN_IN), .ZN(n4365) );
  INV_X1 U2327 ( .A(IR_REG_7__SCAN_IN), .ZN(n2423) );
  NOR2_X1 U2328 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2230)
         );
  INV_X1 U2329 ( .A(IR_REG_8__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U2330 ( .A1(n2432), .A2(n2423), .ZN(n2287) );
  XNOR2_X1 U2331 ( .A(n2312), .B(n2309), .ZN(n2320) );
  INV_X1 U2332 ( .A(IR_REG_30__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U2333 ( .A1(n2647), .A2(n4356), .ZN(n2910) );
  NAND2_X1 U2334 ( .A1(n2305), .A2(n2269), .ZN(n2268) );
  INV_X1 U2335 ( .A(IR_REG_26__SCAN_IN), .ZN(n2269) );
  NAND2_X1 U2336 ( .A1(n2696), .A2(n2695), .ZN(n2847) );
  INV_X1 U2337 ( .A(n2337), .ZN(n2633) );
  OR2_X1 U2338 ( .A1(n4265), .A2(n4140), .ZN(n2537) );
  NAND2_X1 U2339 ( .A1(n3321), .A2(n2498), .ZN(n3386) );
  OR2_X1 U2340 ( .A1(n2886), .A2(n2647), .ZN(n4274) );
  NOR2_X1 U2341 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2296)
         );
  NOR2_X1 U2342 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2294)
         );
  NOR2_X1 U2343 ( .A1(n4430), .A2(n2176), .ZN(n3915) );
  AND2_X1 U2344 ( .A1(n3920), .A2(REG2_REG_15__SCAN_IN), .ZN(n2176) );
  OR2_X1 U2345 ( .A1(n4224), .A2(n4049), .ZN(n3461) );
  INV_X1 U2346 ( .A(n2268), .ZN(n2267) );
  INV_X1 U2347 ( .A(IR_REG_9__SCAN_IN), .ZN(n2288) );
  AND2_X1 U2348 ( .A1(n2911), .A2(n2910), .ZN(n3666) );
  AOI22_X1 U2349 ( .A1(n3615), .A2(n2072), .B1(n2127), .B2(n2125), .ZN(n2123)
         );
  NAND2_X1 U2350 ( .A1(n3752), .A2(n2068), .ZN(n2124) );
  NAND2_X1 U2351 ( .A1(n2128), .A2(n3729), .ZN(n2125) );
  NAND2_X1 U2352 ( .A1(n2139), .A2(n2251), .ZN(n2258) );
  AOI21_X1 U2353 ( .B1(n2255), .B2(n3093), .A(n2063), .ZN(n2251) );
  NAND2_X1 U2354 ( .A1(n3094), .A2(n2255), .ZN(n2139) );
  INV_X1 U2355 ( .A(n3094), .ZN(n2253) );
  AOI22_X1 U2356 ( .A1(n2979), .A2(IR_REG_0__SCAN_IN), .B1(n3662), .B2(n2952), 
        .ZN(n2850) );
  NAND2_X1 U2357 ( .A1(n2848), .A2(n3864), .ZN(n2851) );
  OR2_X1 U2358 ( .A1(n2882), .A2(n4357), .ZN(n2911) );
  XNOR2_X1 U2359 ( .A(n3910), .B(n4491), .ZN(n4401) );
  NAND2_X1 U2360 ( .A1(n2173), .A2(n2171), .ZN(n2732) );
  AOI21_X1 U2361 ( .B1(n2044), .B2(n3552), .A(n2172), .ZN(n2171) );
  INV_X1 U2362 ( .A(n3423), .ZN(n2172) );
  NOR2_X1 U2363 ( .A1(n2597), .A2(n2219), .ZN(n2218) );
  INV_X1 U2364 ( .A(n2590), .ZN(n2219) );
  NAND2_X1 U2365 ( .A1(n4038), .A2(n2282), .ZN(n2582) );
  NAND2_X1 U2366 ( .A1(n2104), .A2(n4176), .ZN(n2160) );
  INV_X1 U2367 ( .A(n3384), .ZN(n2104) );
  OR2_X1 U2368 ( .A1(n4184), .A2(n4288), .ZN(n2511) );
  NAND2_X1 U2369 ( .A1(n2486), .A2(n2075), .ZN(n2212) );
  NAND2_X1 U2370 ( .A1(n3711), .A2(n3793), .ZN(n2214) );
  AND2_X1 U2371 ( .A1(n3048), .A2(n2399), .ZN(n2400) );
  OR2_X1 U2372 ( .A1(n2779), .A2(D_REG_1__SCAN_IN), .ZN(n2879) );
  NAND2_X1 U2373 ( .A1(n2674), .A2(n2164), .ZN(n2163) );
  OR2_X1 U2374 ( .A1(n2779), .A2(D_REG_0__SCAN_IN), .ZN(n2714) );
  AND2_X1 U2375 ( .A1(n2605), .A2(n2604), .ZN(n4218) );
  NAND2_X1 U2376 ( .A1(n2311), .A2(n2776), .ZN(n2314) );
  MUX2_X1 U2377 ( .A(IR_REG_31__SCAN_IN), .B(n2310), .S(IR_REG_29__SCAN_IN), 
        .Z(n2311) );
  INV_X1 U2378 ( .A(IR_REG_20__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U2379 ( .A1(n2639), .A2(IR_REG_31__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U2380 ( .A1(n2521), .A2(n2535), .ZN(n2544) );
  INV_X1 U2381 ( .A(n3711), .ZN(n3849) );
  NAND2_X1 U2382 ( .A1(n2175), .A2(n2044), .ZN(n3983) );
  NAND2_X1 U2383 ( .A1(n2175), .A2(n3558), .ZN(n3981) );
  AND2_X1 U2384 ( .A1(n2553), .A2(REG3_REG_21__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2385 ( .A1(n2240), .A2(n2243), .ZN(n2238) );
  INV_X1 U2386 ( .A(n2281), .ZN(n2272) );
  NAND2_X1 U2387 ( .A1(n2279), .A2(n2278), .ZN(n2277) );
  INV_X1 U2388 ( .A(n3772), .ZN(n2279) );
  NAND2_X1 U2389 ( .A1(n3884), .A2(n2178), .ZN(n2177) );
  NAND2_X1 U2390 ( .A1(n4364), .A2(REG2_REG_2__SCAN_IN), .ZN(n2178) );
  NAND2_X1 U2391 ( .A1(n2221), .A2(n2217), .ZN(n2216) );
  INV_X1 U2392 ( .A(n2218), .ZN(n2217) );
  AND2_X1 U2393 ( .A1(n2451), .A2(n2064), .ZN(n2209) );
  NAND2_X1 U2394 ( .A1(n3861), .A2(n2931), .ZN(n3518) );
  NAND3_X1 U2395 ( .A1(n2193), .A2(n2192), .A3(n3008), .ZN(n3514) );
  NOR2_X1 U2396 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2297)
         );
  NAND2_X1 U2397 ( .A1(n2521), .A2(n2058), .ZN(n2229) );
  AND4_X1 U2398 ( .A1(n2303), .A2(n2302), .A3(n2301), .A4(n2300), .ZN(n2304)
         );
  NOR2_X1 U2399 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2303)
         );
  NOR2_X1 U2400 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2302)
         );
  NOR2_X1 U2401 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2301)
         );
  NOR2_X1 U2402 ( .A1(n2334), .A2(IR_REG_13__SCAN_IN), .ZN(n2496) );
  NOR2_X1 U2403 ( .A1(n3182), .A2(n3183), .ZN(n2265) );
  AOI21_X1 U2404 ( .B1(n2062), .B2(n3182), .A(n2264), .ZN(n2263) );
  NOR2_X1 U2405 ( .A1(n3132), .A2(n2266), .ZN(n2264) );
  NAND2_X1 U2406 ( .A1(n2563), .A2(REG3_REG_22__SCAN_IN), .ZN(n2573) );
  INV_X1 U2407 ( .A(n2121), .ZN(n2115) );
  INV_X1 U2408 ( .A(n3250), .ZN(n2117) );
  INV_X1 U2409 ( .A(n3853), .ZN(n3259) );
  INV_X1 U2410 ( .A(n3778), .ZN(n2243) );
  NAND2_X1 U2411 ( .A1(n3752), .A2(n3830), .ZN(n3617) );
  INV_X1 U2412 ( .A(n3093), .ZN(n2254) );
  AND2_X1 U2413 ( .A1(n2259), .A2(n2256), .ZN(n2255) );
  INV_X1 U2414 ( .A(n3096), .ZN(n2256) );
  OR2_X1 U2415 ( .A1(n3092), .A2(n3091), .ZN(n2259) );
  NAND2_X1 U2416 ( .A1(n2122), .A2(n3207), .ZN(n2121) );
  INV_X1 U2417 ( .A(n3224), .ZN(n2122) );
  INV_X1 U2418 ( .A(n2120), .ZN(n2119) );
  OAI21_X1 U2419 ( .B1(n2260), .B2(n2121), .A(n3223), .ZN(n2120) );
  INV_X1 U2420 ( .A(n3799), .ZN(n2138) );
  XNOR2_X1 U2421 ( .A(n2234), .B(n2972), .ZN(n2926) );
  NAND2_X1 U2422 ( .A1(n2345), .A2(n3662), .ZN(n2233) );
  NAND2_X1 U2423 ( .A1(n2344), .A2(n3662), .ZN(n2232) );
  NAND2_X1 U2424 ( .A1(n2079), .A2(n3624), .ZN(n2249) );
  NAND2_X1 U2425 ( .A1(n2258), .A2(n2257), .ZN(n3133) );
  INV_X1 U2426 ( .A(n3146), .ZN(n2257) );
  AND2_X1 U2427 ( .A1(n2403), .A2(REG3_REG_6__SCAN_IN), .ZN(n2415) );
  INV_X1 U2428 ( .A(n2847), .ZN(n2979) );
  AOI21_X1 U2429 ( .B1(n2271), .B2(n2137), .A(n2135), .ZN(n2134) );
  INV_X1 U2430 ( .A(n2275), .ZN(n2135) );
  AOI21_X1 U2431 ( .B1(n3660), .B2(n3772), .A(n2276), .ZN(n2275) );
  AND2_X1 U2432 ( .A1(n3657), .A2(n3658), .ZN(n2276) );
  INV_X1 U2433 ( .A(n3744), .ZN(n2132) );
  NOR2_X1 U2434 ( .A1(n2241), .A2(n3644), .ZN(n2239) );
  NAND2_X1 U2435 ( .A1(n2326), .A2(REG3_REG_14__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U2436 ( .A1(n3615), .A2(n3614), .ZN(n3829) );
  NAND2_X1 U2437 ( .A1(n4372), .A2(n3906), .ZN(n3907) );
  NAND2_X1 U2438 ( .A1(n4385), .A2(n3932), .ZN(n4390) );
  NAND2_X1 U2439 ( .A1(n4390), .A2(n4391), .ZN(n4389) );
  NAND2_X1 U2440 ( .A1(n4392), .A2(n3909), .ZN(n3910) );
  NAND2_X1 U2441 ( .A1(n4401), .A2(REG2_REG_12__SCAN_IN), .ZN(n4400) );
  OAI21_X1 U2442 ( .B1(n4413), .B2(n4409), .A(n2180), .ZN(n3912) );
  OR2_X1 U2443 ( .A1(n3921), .A2(REG2_REG_13__SCAN_IN), .ZN(n2180) );
  NAND2_X1 U2444 ( .A1(n4435), .A2(n3941), .ZN(n3943) );
  NAND2_X1 U2445 ( .A1(n4441), .A2(n3916), .ZN(n4449) );
  NAND2_X1 U2446 ( .A1(n4449), .A2(n4451), .ZN(n4450) );
  NOR2_X1 U2447 ( .A1(n2190), .A2(n4461), .ZN(n4460) );
  INV_X1 U2448 ( .A(n4022), .ZN(n2103) );
  NAND2_X1 U2449 ( .A1(n2215), .A2(n2067), .ZN(n2220) );
  AOI21_X1 U2450 ( .B1(n2197), .B2(n2195), .A(n2077), .ZN(n2194) );
  INV_X1 U2451 ( .A(n2197), .ZN(n2196) );
  NAND2_X1 U2452 ( .A1(n4075), .A2(n2562), .ZN(n2198) );
  OAI21_X1 U2453 ( .B1(n4088), .B2(n3457), .A(n3458), .ZN(n4075) );
  AOI21_X1 U2454 ( .B1(n4176), .B2(n2226), .A(n2073), .ZN(n2225) );
  AOI21_X1 U2455 ( .B1(n4176), .B2(n2162), .A(n3435), .ZN(n2161) );
  INV_X1 U2456 ( .A(n3504), .ZN(n2162) );
  NOR2_X1 U2457 ( .A1(n4268), .A2(n4273), .ZN(n2228) );
  NOR2_X1 U2458 ( .A1(n4175), .A2(n4176), .ZN(n4174) );
  NAND2_X1 U2459 ( .A1(n3438), .A2(n2211), .ZN(n2658) );
  NOR2_X1 U2460 ( .A1(n2211), .A2(n2488), .ZN(n2210) );
  OR2_X1 U2461 ( .A1(n3850), .A2(n3281), .ZN(n2485) );
  AOI21_X1 U2462 ( .B1(n2051), .B2(n2209), .A(n2208), .ZN(n2207) );
  NOR2_X1 U2463 ( .A1(n3316), .A2(n3265), .ZN(n2208) );
  NAND2_X1 U2464 ( .A1(n3162), .A2(n2209), .ZN(n2206) );
  INV_X1 U2465 ( .A(n2453), .ZN(n2317) );
  OAI21_X1 U2466 ( .B1(n3070), .B2(n2651), .A(n3531), .ZN(n3166) );
  NAND2_X1 U2467 ( .A1(n2402), .A2(n2202), .ZN(n2201) );
  NOR2_X1 U2468 ( .A1(n2413), .A2(n2203), .ZN(n2202) );
  NAND2_X1 U2469 ( .A1(n2744), .A2(n2360), .ZN(n3013) );
  OR2_X1 U2470 ( .A1(n3418), .A2(n2346), .ZN(n2350) );
  NAND2_X1 U2471 ( .A1(n4011), .A2(n3998), .ZN(n3997) );
  NOR2_X2 U2472 ( .A1(n4048), .A2(n4223), .ZN(n4026) );
  NAND2_X1 U2473 ( .A1(n2109), .A2(n3317), .ZN(n3293) );
  AND4_X1 U2474 ( .A1(n2466), .A2(n2465), .A3(n2464), .A4(n2463), .ZN(n3376)
         );
  NAND2_X1 U2475 ( .A1(n2672), .A2(n3451), .ZN(n4171) );
  NAND2_X1 U2476 ( .A1(n2694), .A2(n2766), .ZN(n2779) );
  NAND2_X1 U2477 ( .A1(n4484), .A2(n2847), .ZN(n2895) );
  NAND2_X1 U2478 ( .A1(n2107), .A2(n2060), .ZN(n2165) );
  AND2_X1 U2479 ( .A1(n2144), .A2(n2142), .ZN(n2141) );
  INV_X1 U2480 ( .A(IR_REG_23__SCAN_IN), .ZN(n2698) );
  NAND2_X1 U2481 ( .A1(n2521), .A2(n2144), .ZN(n2688) );
  NOR2_X1 U2482 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2642)
         );
  INV_X1 U2483 ( .A(n2145), .ZN(n2143) );
  NOR2_X2 U2484 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2112)
         );
  AND2_X1 U2485 ( .A1(n2978), .A2(n2977), .ZN(n3094) );
  NAND2_X1 U2486 ( .A1(n2976), .A2(n2933), .ZN(n2977) );
  NOR2_X1 U2487 ( .A1(n2913), .A2(n2286), .ZN(n2918) );
  AND2_X1 U2488 ( .A1(n2589), .A2(n2588), .ZN(n3747) );
  INV_X1 U2489 ( .A(n3860), .ZN(n3099) );
  AND2_X1 U2490 ( .A1(n2560), .A2(n2559), .ZN(n4096) );
  INV_X1 U2491 ( .A(n3852), .ZN(n3316) );
  INV_X1 U2492 ( .A(n3820), .ZN(n3098) );
  OR2_X1 U2493 ( .A1(n2922), .A2(n2898), .ZN(n3822) );
  NAND2_X1 U2494 ( .A1(n2595), .A2(n2594), .ZN(n4029) );
  INV_X1 U2495 ( .A(n4277), .ZN(n4184) );
  INV_X1 U2496 ( .A(n3792), .ZN(n3850) );
  OAI21_X1 U2497 ( .B1(n4365), .B2(n2799), .A(n2087), .ZN(n3869) );
  NAND2_X1 U2498 ( .A1(n4365), .A2(n2799), .ZN(n2087) );
  NAND2_X1 U2499 ( .A1(n4373), .A2(n4374), .ZN(n4372) );
  NAND2_X1 U2500 ( .A1(n4393), .A2(n4394), .ZN(n4392) );
  NOR2_X1 U2501 ( .A1(n4446), .A2(n3944), .ZN(n4455) );
  OAI21_X1 U2502 ( .B1(n4460), .B2(n2188), .A(n2187), .ZN(n2186) );
  AOI21_X1 U2503 ( .B1(n4463), .B2(ADDR_REG_18__SCAN_IN), .A(n4462), .ZN(n2187) );
  NAND2_X1 U2504 ( .A1(n2189), .A2(n4411), .ZN(n2188) );
  NAND2_X1 U2505 ( .A1(n2190), .A2(n4461), .ZN(n2189) );
  NAND2_X1 U2506 ( .A1(n2152), .A2(n2153), .ZN(n4464) );
  NOR2_X1 U2507 ( .A1(n2155), .A2(n2154), .ZN(n2153) );
  INV_X1 U2508 ( .A(n4466), .ZN(n2154) );
  AND2_X1 U2509 ( .A1(n2809), .A2(n2806), .ZN(n4465) );
  AND4_X1 U2510 ( .A1(n2333), .A2(n2332), .A3(n2331), .A4(n2330), .ZN(n3711)
         );
  MUX2_X1 U2511 ( .A(DATAI_1_), .B(n4365), .S(n2357), .Z(n3008) );
  AND2_X1 U2512 ( .A1(n3965), .A2(n2168), .ZN(n2725) );
  AOI21_X1 U2513 ( .B1(n3962), .B2(n4506), .A(n2169), .ZN(n2168) );
  NAND2_X1 U2514 ( .A1(n2683), .A2(n2084), .ZN(n2169) );
  INV_X1 U2515 ( .A(n2725), .ZN(n2167) );
  NAND2_X1 U2516 ( .A1(n2093), .A2(n2092), .ZN(n2091) );
  AOI21_X1 U2517 ( .B1(n4207), .B2(n4289), .A(n4206), .ZN(n2092) );
  OR2_X1 U2518 ( .A1(n4208), .A2(n4262), .ZN(n2093) );
  NAND2_X1 U2519 ( .A1(n2160), .A2(n2158), .ZN(n4113) );
  NOR2_X1 U2520 ( .A1(n2159), .A2(n3432), .ZN(n2158) );
  INV_X1 U2521 ( .A(n2161), .ZN(n2159) );
  NAND2_X1 U2522 ( .A1(n3862), .A2(n2915), .ZN(n3511) );
  NOR2_X1 U2523 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2300)
         );
  NAND2_X1 U2524 ( .A1(n2246), .A2(n3729), .ZN(n2127) );
  INV_X1 U2525 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2318) );
  NOR2_X1 U2526 ( .A1(n2475), .A2(n2474), .ZN(n2327) );
  AND2_X1 U2527 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2370) );
  NAND2_X1 U2528 ( .A1(n3778), .A2(n3633), .ZN(n2242) );
  AND2_X1 U2529 ( .A1(n2327), .A2(REG3_REG_13__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2530 ( .A1(n2149), .A2(n2148), .ZN(n3925) );
  NAND2_X1 U2531 ( .A1(n4359), .A2(REG1_REG_7__SCAN_IN), .ZN(n2148) );
  OR2_X1 U2532 ( .A1(n2871), .A2(n2870), .ZN(n2149) );
  NOR2_X1 U2533 ( .A1(n2606), .A2(n2222), .ZN(n2221) );
  INV_X1 U2534 ( .A(n2596), .ZN(n2222) );
  INV_X1 U2535 ( .A(n2562), .ZN(n2195) );
  NOR2_X1 U2536 ( .A1(n4113), .A2(n3431), .ZN(n4091) );
  NOR2_X1 U2537 ( .A1(n2514), .A2(n2513), .ZN(n2528) );
  INV_X1 U2538 ( .A(n2228), .ZN(n2226) );
  INV_X1 U2539 ( .A(n3503), .ZN(n2100) );
  NAND2_X1 U2540 ( .A1(n2353), .A2(REG0_REG_0__SCAN_IN), .ZN(n2348) );
  NOR3_X1 U2541 ( .A1(n3997), .A2(n3974), .A3(n2717), .ZN(n2718) );
  AND2_X1 U2542 ( .A1(n4065), .A2(n2070), .ZN(n2197) );
  INV_X1 U2543 ( .A(n4104), .ZN(n4094) );
  NOR2_X1 U2544 ( .A1(n3387), .A2(n4288), .ZN(n2110) );
  NAND3_X1 U2545 ( .A1(n2096), .A2(n3514), .A3(n3511), .ZN(n2947) );
  OR2_X1 U2546 ( .A1(n2779), .A2(n2710), .ZN(n2750) );
  NOR2_X1 U2547 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2295)
         );
  NAND2_X1 U2548 ( .A1(n2521), .A2(n2043), .ZN(n2676) );
  INV_X1 U2549 ( .A(n2229), .ZN(n2306) );
  INV_X1 U2550 ( .A(IR_REG_27__SCAN_IN), .ZN(n2307) );
  NOR2_X1 U2551 ( .A1(n2061), .A2(n2145), .ZN(n2144) );
  NAND2_X1 U2552 ( .A1(n2535), .A2(n2146), .ZN(n2145) );
  INV_X1 U2553 ( .A(IR_REG_18__SCAN_IN), .ZN(n2146) );
  INV_X1 U2554 ( .A(IR_REG_17__SCAN_IN), .ZN(n2535) );
  OR2_X1 U2555 ( .A1(n2467), .A2(n2290), .ZN(n2334) );
  AND2_X1 U2556 ( .A1(n2247), .A2(n3755), .ZN(n2128) );
  NOR2_X1 U2557 ( .A1(n3807), .A2(n2248), .ZN(n2247) );
  INV_X1 U2558 ( .A(n3624), .ZN(n2248) );
  OR2_X1 U2559 ( .A1(n2619), .A2(n3690), .ZN(n2629) );
  INV_X1 U2560 ( .A(n3202), .ZN(n2261) );
  INV_X1 U2561 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2474) );
  OR2_X1 U2562 ( .A1(n2502), .A2(n2318), .ZN(n2514) );
  AND2_X1 U2563 ( .A1(n2854), .A2(n2855), .ZN(n2913) );
  INV_X1 U2564 ( .A(n2237), .ZN(n2236) );
  OAI22_X1 U2565 ( .A1(n3644), .A2(n2238), .B1(n3642), .B2(n3643), .ZN(n2237)
         );
  XNOR2_X1 U2566 ( .A(n2930), .B(n2972), .ZN(n2974) );
  AND2_X1 U2567 ( .A1(n2370), .A2(REG3_REG_5__SCAN_IN), .ZN(n2403) );
  OR2_X1 U2568 ( .A1(n2583), .A2(n4654), .ZN(n2599) );
  AND3_X1 U2569 ( .A1(n2543), .A2(n2542), .A3(n2541), .ZN(n3782) );
  XNOR2_X1 U2570 ( .A(n2177), .B(n2816), .ZN(n3896) );
  INV_X1 U2571 ( .A(IR_REG_5__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U2572 ( .A1(n2185), .A2(n2184), .ZN(n2183) );
  NAND2_X1 U2573 ( .A1(n4361), .A2(REG2_REG_5__SCAN_IN), .ZN(n2184) );
  AOI21_X1 U2574 ( .B1(n2840), .B2(REG2_REG_6__SCAN_IN), .A(n2181), .ZN(n2842)
         );
  AND2_X1 U2575 ( .A1(n2183), .A2(n4360), .ZN(n2181) );
  XNOR2_X1 U2576 ( .A(n3925), .B(n2147), .ZN(n3928) );
  NAND2_X1 U2577 ( .A1(n4389), .A2(n3933), .ZN(n3935) );
  XNOR2_X1 U2578 ( .A(n3915), .B(n3942), .ZN(n4442) );
  NAND2_X1 U2579 ( .A1(n4442), .A2(n2313), .ZN(n4441) );
  INV_X1 U2580 ( .A(n4454), .ZN(n2157) );
  NAND2_X1 U2581 ( .A1(n4450), .A2(n2191), .ZN(n2190) );
  NAND2_X1 U2582 ( .A1(n4487), .A2(n2516), .ZN(n2191) );
  NAND2_X1 U2583 ( .A1(n2718), .A2(n3968), .ZN(n4199) );
  OR2_X1 U2584 ( .A1(n4005), .A2(n3552), .ZN(n2175) );
  NAND2_X1 U2585 ( .A1(n2666), .A2(n3461), .ZN(n4022) );
  CLKBUF_X1 U2586 ( .A(n4088), .Z(n4089) );
  AND3_X1 U2587 ( .A1(n2534), .A2(n2533), .A3(n2532), .ZN(n4119) );
  NAND2_X1 U2588 ( .A1(n2528), .A2(REG3_REG_18__SCAN_IN), .ZN(n2539) );
  OAI21_X1 U2589 ( .B1(n2652), .B2(n2101), .A(n2098), .ZN(n3438) );
  INV_X1 U2590 ( .A(n2654), .ZN(n2101) );
  AND2_X1 U2591 ( .A1(n3542), .A2(n2099), .ZN(n2098) );
  NAND2_X1 U2592 ( .A1(n2654), .A2(n2100), .ZN(n2099) );
  INV_X1 U2593 ( .A(n3486), .ZN(n2205) );
  INV_X1 U2594 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U2595 ( .A1(n2652), .A2(n3503), .ZN(n3298) );
  OAI21_X1 U2596 ( .B1(n3156), .B2(n3155), .A(n3534), .ZN(n3244) );
  AND2_X1 U2597 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2315) );
  INV_X1 U2598 ( .A(n2440), .ZN(n2316) );
  NAND2_X1 U2599 ( .A1(n2170), .A2(n3530), .ZN(n3156) );
  NAND2_X1 U2600 ( .A1(n3166), .A2(n3533), .ZN(n2170) );
  NAND2_X1 U2601 ( .A1(n2649), .A2(n3527), .ZN(n3070) );
  OAI21_X1 U2602 ( .B1(n3021), .B2(n2648), .A(n3525), .ZN(n3046) );
  NAND2_X1 U2603 ( .A1(n2382), .A2(n2381), .ZN(n3048) );
  AND2_X1 U2604 ( .A1(n2750), .A2(n2780), .ZN(n2880) );
  NAND2_X1 U2605 ( .A1(n2991), .A2(n3520), .ZN(n3021) );
  NOR2_X1 U2606 ( .A1(n2095), .A2(n2903), .ZN(n2094) );
  INV_X1 U2607 ( .A(n2350), .ZN(n2095) );
  AOI22_X1 U2608 ( .A1(n2682), .A2(n4171), .B1(n3957), .B2(n3844), .ZN(n3965)
         );
  AOI21_X1 U2609 ( .B1(n2732), .B2(n3421), .A(n2670), .ZN(n2671) );
  AND2_X1 U2610 ( .A1(n2615), .A2(n2614), .ZN(n3993) );
  OR2_X1 U2611 ( .A1(n3975), .A2(n2337), .ZN(n2615) );
  NOR2_X1 U2612 ( .A1(n3419), .A2(n4534), .ZN(n4214) );
  NAND2_X1 U2613 ( .A1(n4102), .A2(n2049), .ZN(n4048) );
  NAND2_X1 U2614 ( .A1(n4102), .A2(n2048), .ZN(n4062) );
  NAND2_X1 U2615 ( .A1(n2198), .A2(n2197), .ZN(n4238) );
  AND2_X1 U2616 ( .A1(n4102), .A2(n4082), .ZN(n4076) );
  NOR2_X1 U2617 ( .A1(n3419), .A2(n2561), .ZN(n4242) );
  NAND2_X1 U2618 ( .A1(n2308), .A2(DATAI_20_), .ZN(n4104) );
  NAND2_X1 U2619 ( .A1(n4159), .A2(n4147), .ZN(n4145) );
  INV_X1 U2620 ( .A(n2716), .ZN(n4125) );
  NAND2_X1 U2621 ( .A1(n2110), .A2(n4273), .ZN(n4181) );
  INV_X1 U2622 ( .A(n2110), .ZN(n4179) );
  INV_X1 U2623 ( .A(n3836), .ZN(n4288) );
  NAND2_X1 U2624 ( .A1(n3346), .A2(n3712), .ZN(n3387) );
  INV_X1 U2625 ( .A(n3324), .ZN(n3712) );
  AND2_X1 U2626 ( .A1(n3344), .A2(n3793), .ZN(n3346) );
  NAND2_X1 U2627 ( .A1(n3217), .A2(n3265), .ZN(n2108) );
  INV_X1 U2628 ( .A(n3252), .ZN(n3265) );
  NOR3_X1 U2629 ( .A1(n3174), .A2(n3226), .A3(n3175), .ZN(n3238) );
  NOR2_X1 U2630 ( .A1(n3174), .A2(n3175), .ZN(n3173) );
  INV_X1 U2631 ( .A(n3110), .ZN(n3138) );
  AND4_X1 U2632 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n3137)
         );
  AND2_X1 U2633 ( .A1(n2904), .A2(n2647), .ZN(n4146) );
  INV_X1 U2634 ( .A(n4243), .ZN(n4293) );
  AND2_X1 U2635 ( .A1(n2510), .A2(n2509), .ZN(n3920) );
  AND2_X1 U2636 ( .A1(n2450), .A2(n2467), .ZN(n3923) );
  AND4_X1 U2637 ( .A1(n2506), .A2(n2505), .A3(n2504), .A4(n2503), .ZN(n4277)
         );
  NOR2_X1 U2638 ( .A1(n2262), .A2(n2114), .ZN(n2113) );
  OAI21_X1 U2639 ( .B1(n2119), .B2(n2117), .A(n2071), .ZN(n2116) );
  NAND2_X1 U2640 ( .A1(n2115), .A2(n3250), .ZN(n2114) );
  AND3_X1 U2641 ( .A1(n2552), .A2(n2551), .A3(n2550), .ZN(n3739) );
  NAND2_X1 U2642 ( .A1(n2118), .A2(n3207), .ZN(n3225) );
  NAND2_X1 U2643 ( .A1(n2262), .A2(n2260), .ZN(n2118) );
  AND2_X1 U2644 ( .A1(n2570), .A2(n2569), .ZN(n4247) );
  OAI21_X1 U2645 ( .B1(n3635), .B2(n2243), .A(n2240), .ZN(n3737) );
  AND2_X1 U2646 ( .A1(n2564), .A2(n2555), .ZN(n4079) );
  NAND2_X1 U2647 ( .A1(n2129), .A2(n2134), .ZN(n3746) );
  OR2_X1 U2648 ( .A1(n2235), .A2(n2270), .ZN(n2129) );
  INV_X1 U2649 ( .A(n3133), .ZN(n3145) );
  OAI21_X1 U2650 ( .B1(n3718), .B2(n3657), .A(n3658), .ZN(n3770) );
  NAND2_X1 U2651 ( .A1(n2274), .A2(n2273), .ZN(n3769) );
  INV_X1 U2652 ( .A(n3660), .ZN(n2273) );
  AND2_X1 U2653 ( .A1(n2252), .A2(n2255), .ZN(n3125) );
  NAND2_X1 U2654 ( .A1(n2254), .A2(n2253), .ZN(n2252) );
  AND4_X1 U2655 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n3231)
         );
  NAND2_X1 U2656 ( .A1(n2308), .A2(DATAI_0_), .ZN(n2111) );
  NAND2_X1 U2657 ( .A1(n3419), .A2(IR_REG_0__SCAN_IN), .ZN(n2351) );
  INV_X1 U2658 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4520) );
  AND4_X1 U2659 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n3792)
         );
  NAND2_X1 U2660 ( .A1(n2235), .A2(n2236), .ZN(n3798) );
  NOR2_X1 U2661 ( .A1(n2929), .A2(n2928), .ZN(n2935) );
  AND4_X1 U2662 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n4276)
         );
  INV_X1 U2663 ( .A(n4140), .ZN(n4147) );
  AND2_X1 U2664 ( .A1(n2244), .A2(n2249), .ZN(n3811) );
  AND4_X1 U2665 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n3216)
         );
  AND2_X1 U2666 ( .A1(n3133), .A2(n3132), .ZN(n3184) );
  NOR2_X1 U2667 ( .A1(n2893), .A2(n4186), .ZN(n3820) );
  NAND2_X1 U2668 ( .A1(n2983), .A2(n2982), .ZN(n3825) );
  INV_X1 U2669 ( .A(n2131), .ZN(n2130) );
  OAI21_X1 U2670 ( .B1(n2134), .B2(n2069), .A(n2132), .ZN(n2131) );
  AND4_X1 U2671 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n4294)
         );
  INV_X1 U2672 ( .A(n3098), .ZN(n3837) );
  INV_X1 U2673 ( .A(n3827), .ZN(n3832) );
  INV_X1 U2674 ( .A(n3825), .ZN(n3843) );
  NOR2_X1 U2675 ( .A1(n3656), .A2(n2884), .ZN(n3574) );
  INV_X1 U2676 ( .A(n4357), .ZN(n3952) );
  INV_X1 U2677 ( .A(n3993), .ZN(n3846) );
  INV_X1 U2678 ( .A(n3747), .ZN(n4215) );
  NAND2_X1 U2679 ( .A1(n2579), .A2(n2578), .ZN(n4224) );
  INV_X1 U2680 ( .A(n3782), .ZN(n4141) );
  INV_X1 U2681 ( .A(n4119), .ZN(n4265) );
  INV_X1 U2682 ( .A(n4276), .ZN(n4182) );
  INV_X1 U2683 ( .A(n3376), .ZN(n3851) );
  INV_X1 U2684 ( .A(n3231), .ZN(n3854) );
  INV_X1 U2685 ( .A(n3216), .ZN(n3855) );
  CLKBUF_X1 U2686 ( .A(U4043), .Z(n3856) );
  NOR2_X1 U2687 ( .A1(n2363), .A2(n2056), .ZN(n2364) );
  NAND2_X1 U2688 ( .A1(n3869), .A2(n2800), .ZN(n3881) );
  INV_X1 U2689 ( .A(n2185), .ZN(n2825) );
  XNOR2_X1 U2690 ( .A(n2183), .B(n2182), .ZN(n2840) );
  INV_X1 U2691 ( .A(n4360), .ZN(n2182) );
  NOR2_X1 U2692 ( .A1(n2836), .A2(n2150), .ZN(n2871) );
  AND2_X1 U2693 ( .A1(n2837), .A2(n4360), .ZN(n2150) );
  INV_X1 U2694 ( .A(n3928), .ZN(n3924) );
  OAI21_X1 U2695 ( .B1(n3905), .B2(n4472), .A(n2085), .ZN(n4373) );
  NAND2_X1 U2696 ( .A1(n2086), .A2(n2147), .ZN(n2085) );
  NAND2_X1 U2697 ( .A1(n4380), .A2(n3908), .ZN(n4393) );
  XNOR2_X1 U2698 ( .A(n3935), .B(n4491), .ZN(n4406) );
  NAND2_X1 U2699 ( .A1(n4400), .A2(n3911), .ZN(n4413) );
  XNOR2_X1 U2700 ( .A(n3912), .B(n2179), .ZN(n4423) );
  NAND2_X1 U2701 ( .A1(n4426), .A2(n3940), .ZN(n4436) );
  NAND2_X1 U2702 ( .A1(n4436), .A2(n4437), .ZN(n4435) );
  XNOR2_X1 U2703 ( .A(n3943), .B(n3942), .ZN(n4445) );
  AOI21_X1 U2704 ( .B1(n2729), .B2(n2731), .A(n2628), .ZN(n2634) );
  NAND2_X1 U2705 ( .A1(n2223), .A2(n2596), .ZN(n3986) );
  NAND2_X1 U2706 ( .A1(n2220), .A2(n2218), .ZN(n2223) );
  INV_X1 U2707 ( .A(n4214), .ZN(n4016) );
  NAND2_X1 U2708 ( .A1(n2220), .A2(n2590), .ZN(n4008) );
  AND2_X1 U2709 ( .A1(n2198), .A2(n2070), .ZN(n4066) );
  INV_X1 U2710 ( .A(n4242), .ZN(n4082) );
  NAND2_X1 U2711 ( .A1(n2160), .A2(n2161), .ZN(n4155) );
  NOR2_X1 U2712 ( .A1(n4174), .A2(n2228), .ZN(n4158) );
  NAND2_X1 U2713 ( .A1(n4173), .A2(n4176), .ZN(n4172) );
  NAND2_X1 U2714 ( .A1(n3384), .A2(n3504), .ZN(n4173) );
  AND2_X1 U2715 ( .A1(n2212), .A2(n2213), .ZN(n3323) );
  NAND2_X1 U2716 ( .A1(n2486), .A2(n2485), .ZN(n3343) );
  NAND4_X1 U2717 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(n3852)
         );
  OAI21_X1 U2718 ( .B1(n3162), .B2(n2051), .A(n2451), .ZN(n3237) );
  NOR2_X1 U2719 ( .A1(n3528), .A2(n2200), .ZN(n2199) );
  INV_X1 U2720 ( .A(n2204), .ZN(n2200) );
  NAND2_X1 U2721 ( .A1(n2201), .A2(n2204), .ZN(n3081) );
  INV_X1 U2722 ( .A(n4127), .ZN(n4476) );
  OR2_X1 U2723 ( .A1(n4148), .A2(n4283), .ZN(n4127) );
  OR2_X1 U2724 ( .A1(n2895), .A2(n2754), .ZN(n4470) );
  NOR2_X1 U2725 ( .A1(n2054), .A2(n2106), .ZN(n2105) );
  AND2_X1 U2726 ( .A1(n4473), .A2(n4243), .ZN(n4185) );
  AND3_X1 U2727 ( .A1(n3357), .A2(n3356), .A3(n3355), .ZN(n3360) );
  OR2_X1 U2728 ( .A1(n2724), .A2(n2881), .ZN(n4511) );
  NAND2_X1 U2729 ( .A1(n2107), .A2(n2693), .ZN(n2783) );
  NAND2_X1 U2730 ( .A1(n2779), .A2(n2778), .ZN(n4483) );
  INV_X1 U2731 ( .A(IR_REG_29__SCAN_IN), .ZN(n2102) );
  INV_X1 U2732 ( .A(IR_REG_31__SCAN_IN), .ZN(n2775) );
  INV_X1 U2733 ( .A(n2165), .ZN(n2673) );
  INV_X1 U2734 ( .A(n2783), .ZN(n2766) );
  NAND2_X1 U2735 ( .A1(n2689), .A2(IR_REG_31__SCAN_IN), .ZN(n2690) );
  INV_X1 U2736 ( .A(n2882), .ZN(n4355) );
  XNOR2_X1 U2737 ( .A(n2645), .B(IR_REG_21__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U2738 ( .A1(n2644), .A2(IR_REG_31__SCAN_IN), .ZN(n2645) );
  XNOR2_X1 U2739 ( .A(n2638), .B(IR_REG_19__SCAN_IN), .ZN(n4357) );
  INV_X1 U2740 ( .A(n3920), .ZN(n4489) );
  INV_X1 U2741 ( .A(n3934), .ZN(n4491) );
  AND2_X1 U2742 ( .A1(n2378), .A2(n2368), .ZN(n4363) );
  NAND2_X1 U2743 ( .A1(n2151), .A2(IR_REG_31__SCAN_IN), .ZN(n2356) );
  INV_X1 U2744 ( .A(n2112), .ZN(n2151) );
  NAND2_X1 U2745 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2088)
         );
  NOR2_X1 U2746 ( .A1(n4455), .A2(n4454), .ZN(n4456) );
  INV_X1 U2747 ( .A(n2186), .ZN(n4468) );
  AOI21_X1 U2748 ( .B1(n4307), .B2(n4518), .A(n2089), .ZN(n4209) );
  INV_X1 U2749 ( .A(n2090), .ZN(n2089) );
  AOI22_X1 U2750 ( .A1(n4309), .A2(n2720), .B1(REG1_REG_27__SCAN_IN), .B2(
        n4516), .ZN(n2090) );
  NAND2_X1 U2751 ( .A1(n2167), .A2(n4513), .ZN(n2166) );
  AND3_X1 U2752 ( .A1(n2047), .A2(n2304), .A3(n2164), .ZN(n2043) );
  AND2_X1 U2753 ( .A1(n2277), .A2(n2272), .ZN(n2271) );
  AND2_X1 U2754 ( .A1(n2174), .A2(n3558), .ZN(n2044) );
  INV_X1 U2755 ( .A(n3183), .ZN(n2266) );
  NAND2_X1 U2756 ( .A1(n2112), .A2(n2231), .ZN(n2366) );
  NOR2_X1 U2757 ( .A1(n2053), .A2(n2097), .ZN(n2045) );
  XNOR2_X1 U2758 ( .A(n2356), .B(IR_REG_2__SCAN_IN), .ZN(n4364) );
  NAND2_X1 U2759 ( .A1(n2216), .A2(n2076), .ZN(n2046) );
  INV_X1 U2760 ( .A(n2271), .ZN(n2270) );
  AND2_X1 U2761 ( .A1(n2267), .A2(n2307), .ZN(n2047) );
  AND2_X1 U2762 ( .A1(n3849), .A2(n2487), .ZN(n2488) );
  INV_X1 U2763 ( .A(n3297), .ZN(n3317) );
  AND2_X1 U2764 ( .A1(n2425), .A2(n2431), .ZN(n4359) );
  AND2_X1 U2765 ( .A1(n4082), .A2(n4060), .ZN(n2048) );
  AND2_X1 U2766 ( .A1(n2048), .A2(n4049), .ZN(n2049) );
  XNOR2_X1 U2767 ( .A(n2641), .B(n2640), .ZN(n2647) );
  BUF_X1 U2768 ( .A(n3682), .Z(n3656) );
  INV_X4 U2769 ( .A(n2347), .ZN(n2353) );
  NOR2_X1 U2770 ( .A1(n3997), .A2(n3974), .ZN(n2050) );
  NAND2_X1 U2771 ( .A1(n2351), .A2(n2111), .ZN(n2952) );
  AND2_X1 U2772 ( .A1(n3853), .A2(n3226), .ZN(n2051) );
  INV_X1 U2773 ( .A(n2975), .ZN(n2933) );
  AND2_X1 U2774 ( .A1(n2177), .A2(n4363), .ZN(n2052) );
  INV_X1 U2775 ( .A(n3861), .ZN(n2932) );
  NAND2_X1 U2776 ( .A1(n2126), .A2(n2245), .ZN(n3728) );
  AND2_X1 U2777 ( .A1(n2133), .A2(n2130), .ZN(n3816) );
  NOR2_X1 U2778 ( .A1(n2337), .A2(n2902), .ZN(n2053) );
  NOR2_X1 U2779 ( .A1(n3719), .A2(n2281), .ZN(n3718) );
  INV_X1 U2780 ( .A(n3718), .ZN(n2274) );
  NAND2_X1 U2781 ( .A1(n2521), .A2(n2304), .ZN(n2684) );
  AND2_X1 U2782 ( .A1(n2353), .A2(REG0_REG_2__SCAN_IN), .ZN(n2054) );
  AND2_X1 U2783 ( .A1(n3777), .A2(n3778), .ZN(n2055) );
  NOR2_X1 U2784 ( .A1(n2347), .A2(n2998), .ZN(n2056) );
  NAND2_X1 U2785 ( .A1(n2307), .A2(n2775), .ZN(n2057) );
  AND2_X1 U2786 ( .A1(n2047), .A2(n2304), .ZN(n2058) );
  AND2_X1 U2787 ( .A1(n2804), .A2(n4362), .ZN(n2059) );
  AND2_X1 U2788 ( .A1(n2650), .A2(n3531), .ZN(n3528) );
  AND2_X1 U2789 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2060)
         );
  OR2_X1 U2790 ( .A1(IR_REG_21__SCAN_IN), .A2(n2635), .ZN(n2061) );
  AND2_X1 U2791 ( .A1(n3284), .A2(n3286), .ZN(n3486) );
  OR2_X1 U2792 ( .A1(n3131), .A2(n3183), .ZN(n2062) );
  AND2_X1 U2793 ( .A1(n3124), .A2(n3123), .ZN(n2063) );
  OR2_X1 U2794 ( .A1(n2684), .A2(n2268), .ZN(n2107) );
  OR2_X1 U2795 ( .A1(n3852), .A2(n3252), .ZN(n2064) );
  AND2_X1 U2796 ( .A1(n2207), .A2(n2205), .ZN(n2065) );
  NAND2_X1 U2797 ( .A1(n2250), .A2(n3622), .ZN(n3761) );
  NAND2_X1 U2798 ( .A1(n3635), .A2(n3634), .ZN(n3777) );
  INV_X1 U2799 ( .A(n2156), .ZN(n2155) );
  AOI21_X1 U2800 ( .B1(n3944), .B2(n2157), .A(n3946), .ZN(n2156) );
  AND2_X1 U2801 ( .A1(n2152), .A2(n2156), .ZN(n2066) );
  INV_X1 U2802 ( .A(IR_REG_28__SCAN_IN), .ZN(n2164) );
  INV_X1 U2803 ( .A(IR_REG_25__SCAN_IN), .ZN(n2305) );
  INV_X1 U2804 ( .A(n3658), .ZN(n2278) );
  INV_X1 U2805 ( .A(n3980), .ZN(n2174) );
  NOR2_X1 U2806 ( .A1(n2421), .A2(n2287), .ZN(n2299) );
  INV_X1 U2807 ( .A(n3226), .ZN(n3232) );
  INV_X1 U2808 ( .A(n4268), .ZN(n4290) );
  OR2_X1 U2809 ( .A1(n3747), .A2(n4033), .ZN(n2067) );
  INV_X1 U2810 ( .A(IR_REG_22__SCAN_IN), .ZN(n2142) );
  INV_X1 U2811 ( .A(n3322), .ZN(n2211) );
  AND2_X1 U2812 ( .A1(n2127), .A2(n3830), .ZN(n2068) );
  AND2_X1 U2813 ( .A1(n3670), .A2(n3669), .ZN(n2069) );
  INV_X1 U2814 ( .A(n3217), .ZN(n3175) );
  NAND2_X1 U2815 ( .A1(n4096), .A2(n4082), .ZN(n2070) );
  OR2_X1 U2816 ( .A1(n3249), .A2(n3248), .ZN(n2071) );
  AND2_X1 U2817 ( .A1(n2127), .A2(n3614), .ZN(n2072) );
  INV_X1 U2818 ( .A(n3633), .ZN(n3634) );
  AND2_X1 U2819 ( .A1(n4276), .A2(n4166), .ZN(n2073) );
  INV_X1 U2820 ( .A(n2137), .ZN(n2136) );
  NAND2_X1 U2821 ( .A1(n2236), .A2(n2138), .ZN(n2137) );
  AND2_X1 U2822 ( .A1(n2221), .A2(n2067), .ZN(n2074) );
  AND2_X1 U2823 ( .A1(n2485), .A2(n2214), .ZN(n2075) );
  NAND2_X1 U2824 ( .A1(n4218), .A2(n3998), .ZN(n2076) );
  INV_X1 U2825 ( .A(n2241), .ZN(n2240) );
  NAND2_X1 U2826 ( .A1(n2242), .A2(n3780), .ZN(n2241) );
  NOR2_X1 U2827 ( .A1(n4247), .A2(n4060), .ZN(n2077) );
  INV_X1 U2828 ( .A(n2524), .ZN(n2227) );
  NAND2_X1 U2829 ( .A1(n2045), .A2(n2094), .ZN(n3510) );
  INV_X1 U2830 ( .A(n2246), .ZN(n2245) );
  OAI21_X1 U2831 ( .B1(n2249), .B2(n3807), .A(n3808), .ZN(n2246) );
  OR2_X1 U2832 ( .A1(n3762), .A2(n3763), .ZN(n2078) );
  NAND2_X1 U2833 ( .A1(n2078), .A2(n3622), .ZN(n2079) );
  AND2_X1 U2834 ( .A1(n3782), .A2(n4125), .ZN(n2080) );
  OR2_X1 U2835 ( .A1(n2225), .A2(n2524), .ZN(n2081) );
  AND2_X1 U2836 ( .A1(n2227), .A2(n2226), .ZN(n2082) );
  XNOR2_X1 U2837 ( .A(n2690), .B(IR_REG_24__SCAN_IN), .ZN(n2696) );
  INV_X2 U2838 ( .A(n4516), .ZN(n4518) );
  OR2_X1 U2839 ( .A1(n2724), .A2(n2752), .ZN(n4516) );
  OAI21_X1 U2840 ( .B1(n2262), .B2(n2121), .A(n2119), .ZN(n3251) );
  OR2_X1 U2841 ( .A1(n4513), .A2(n2726), .ZN(n2083) );
  NAND2_X1 U2842 ( .A1(n2252), .A2(n2259), .ZN(n3095) );
  NAND2_X1 U2843 ( .A1(n2206), .A2(n2207), .ZN(n3294) );
  INV_X1 U2844 ( .A(n2109), .ZN(n3292) );
  NOR3_X1 U2845 ( .A1(n3174), .A2(n2108), .A3(n3226), .ZN(n2109) );
  NAND2_X1 U2846 ( .A1(n2140), .A2(IR_REG_31__SCAN_IN), .ZN(n2697) );
  INV_X1 U2847 ( .A(n3938), .ZN(n2179) );
  INV_X1 U2848 ( .A(n3862), .ZN(n2916) );
  AND2_X1 U2849 ( .A1(n2809), .A2(n3573), .ZN(n4411) );
  NOR2_X1 U2850 ( .A1(n3419), .A2(n2580), .ZN(n3647) );
  OR2_X1 U2851 ( .A1(n3968), .A2(n4274), .ZN(n2084) );
  INV_X1 U2852 ( .A(n2488), .ZN(n2213) );
  INV_X1 U2853 ( .A(n3945), .ZN(n4487) );
  INV_X1 U2854 ( .A(n4358), .ZN(n2147) );
  INV_X1 U2855 ( .A(IR_REG_3__SCAN_IN), .ZN(n4618) );
  INV_X1 U2856 ( .A(n3904), .ZN(n2086) );
  XNOR2_X1 U2857 ( .A(n3904), .B(n4358), .ZN(n3905) );
  OR2_X2 U2858 ( .A1(n4205), .A2(n2091), .ZN(n4307) );
  INV_X1 U2859 ( .A(n3864), .ZN(n2946) );
  INV_X1 U2860 ( .A(n3510), .ZN(n2096) );
  NAND2_X1 U2861 ( .A1(n2349), .A2(n2348), .ZN(n2097) );
  NAND3_X1 U2862 ( .A1(n2521), .A2(n2043), .A3(n2102), .ZN(n2776) );
  NAND2_X2 U2863 ( .A1(n2103), .A2(n3455), .ZN(n4005) );
  OAI21_X1 U2864 ( .B1(n3418), .B2(n2813), .A(n2354), .ZN(n2106) );
  AND2_X2 U2865 ( .A1(n2299), .A2(n2298), .ZN(n2521) );
  NOR2_X2 U2866 ( .A1(n4181), .A2(n4264), .ZN(n4159) );
  INV_X4 U2867 ( .A(n2308), .ZN(n3419) );
  NAND4_X1 U2868 ( .A1(n2112), .A2(n2392), .A3(n2231), .A4(n2230), .ZN(n2421)
         );
  NOR2_X2 U2869 ( .A1(n2741), .A2(n2847), .ZN(U4043) );
  NAND2_X1 U2870 ( .A1(n2935), .A2(n2934), .ZN(n2978) );
  NOR2_X1 U2871 ( .A1(n2917), .A2(n2918), .ZN(n2929) );
  XNOR2_X1 U2872 ( .A(n2927), .B(n2926), .ZN(n2917) );
  NOR2_X1 U2873 ( .A1(n2116), .A2(n2113), .ZN(n3258) );
  NAND2_X1 U2874 ( .A1(n2124), .A2(n2123), .ZN(n3635) );
  NAND3_X1 U2875 ( .A1(n3617), .A2(n3829), .A3(n2128), .ZN(n2126) );
  OR3_X1 U2876 ( .A1(n2235), .A2(n2270), .A3(n2069), .ZN(n2133) );
  AND2_X1 U2877 ( .A1(n2235), .A2(n2136), .ZN(n3719) );
  AND2_X1 U2878 ( .A1(n2521), .A2(n2143), .ZN(n2643) );
  NAND2_X1 U2879 ( .A1(n2521), .A2(n2141), .ZN(n2140) );
  NAND2_X1 U2880 ( .A1(n4446), .A2(n2157), .ZN(n2152) );
  AOI22_X1 U2881 ( .A1(n3663), .A2(n2952), .B1(n3864), .B2(n3662), .ZN(n2912)
         );
  NAND3_X1 U2882 ( .A1(n2166), .A2(n2728), .A3(n2083), .ZN(U3515) );
  NAND2_X1 U2883 ( .A1(n4005), .A2(n2044), .ZN(n2173) );
  NAND2_X1 U2884 ( .A1(n2947), .A2(n3514), .ZN(n2746) );
  NAND2_X1 U2885 ( .A1(n2662), .A2(n3549), .ZN(n4072) );
  OAI21_X1 U2886 ( .B1(n4072), .B2(n2665), .A(n3441), .ZN(n2666) );
  NAND2_X2 U2887 ( .A1(n4354), .A2(n2314), .ZN(n2341) );
  NAND2_X1 U2888 ( .A1(n2746), .A2(n3476), .ZN(n2745) );
  INV_X2 U2889 ( .A(n2357), .ZN(n2308) );
  INV_X1 U2890 ( .A(n2344), .ZN(n2192) );
  INV_X1 U2891 ( .A(n2345), .ZN(n2193) );
  NAND2_X1 U2892 ( .A1(n2201), .A2(n2199), .ZN(n3080) );
  NAND2_X1 U2893 ( .A1(n2402), .A2(n2401), .ZN(n3059) );
  INV_X1 U2894 ( .A(n2401), .ZN(n2203) );
  OR2_X1 U2895 ( .A1(n3857), .A2(n3110), .ZN(n2204) );
  NAND2_X1 U2896 ( .A1(n2206), .A2(n2065), .ZN(n3295) );
  NAND2_X1 U2897 ( .A1(n2212), .A2(n2210), .ZN(n3321) );
  AOI21_X2 U2898 ( .B1(n2215), .B2(n2074), .A(n2046), .ZN(n3973) );
  INV_X1 U2899 ( .A(n4024), .ZN(n2215) );
  NAND2_X1 U2900 ( .A1(n4175), .A2(n2082), .ZN(n2224) );
  NAND2_X1 U2901 ( .A1(n2224), .A2(n2081), .ZN(n4136) );
  OR2_X1 U2902 ( .A1(n2337), .A2(n3004), .ZN(n2340) );
  INV_X1 U2903 ( .A(IR_REG_2__SCAN_IN), .ZN(n2231) );
  NAND3_X1 U2904 ( .A1(n2233), .A2(n2914), .A3(n2232), .ZN(n2234) );
  NAND2_X1 U2905 ( .A1(n3635), .A2(n2239), .ZN(n2235) );
  NAND4_X1 U2906 ( .A1(n3617), .A2(n3829), .A3(n3755), .A4(n3624), .ZN(n2244)
         );
  NAND3_X1 U2907 ( .A1(n3617), .A2(n3829), .A3(n3755), .ZN(n2250) );
  INV_X1 U2908 ( .A(n2258), .ZN(n3144) );
  OAI21_X1 U2909 ( .B1(n3133), .B2(n2265), .A(n2263), .ZN(n3203) );
  AOI21_X1 U2910 ( .B1(n2263), .B2(n2265), .A(n2261), .ZN(n2260) );
  NAND2_X1 U2911 ( .A1(n3133), .A2(n2263), .ZN(n2262) );
  OR2_X1 U2912 ( .A1(n2684), .A2(IR_REG_25__SCAN_IN), .ZN(n2686) );
  OAI22_X1 U2913 ( .A1(n2931), .A2(n3681), .B1(n2932), .B2(n3682), .ZN(n2930)
         );
  OR2_X1 U2914 ( .A1(n3418), .A2(n2338), .ZN(n2339) );
  NAND2_X1 U2915 ( .A1(n2353), .A2(REG0_REG_1__SCAN_IN), .ZN(n2342) );
  INV_X1 U2916 ( .A(n2978), .ZN(n2936) );
  OR2_X1 U2917 ( .A1(n4277), .A2(n3836), .ZN(n2280) );
  OR2_X1 U2918 ( .A1(n3720), .A2(n3721), .ZN(n2281) );
  OR2_X1 U2919 ( .A1(n4224), .A2(n3647), .ZN(n2282) );
  OR2_X1 U2920 ( .A1(n3589), .A2(n4299), .ZN(n2283) );
  INV_X1 U2921 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2513) );
  INV_X1 U2922 ( .A(n4299), .ZN(n2720) );
  OR2_X1 U2923 ( .A1(n3792), .A2(n3377), .ZN(n2284) );
  OR2_X1 U2924 ( .A1(n3589), .A2(n4347), .ZN(n2285) );
  INV_X1 U2925 ( .A(n4347), .ZN(n2727) );
  INV_X1 U2926 ( .A(n3966), .ZN(n2721) );
  NAND2_X1 U2927 ( .A1(n2320), .A2(n2314), .ZN(n2347) );
  AOI22_X1 U2928 ( .A1(n3606), .A2(n3788), .B1(n3605), .B2(n3604), .ZN(n3706)
         );
  AND2_X1 U2929 ( .A1(n2912), .A2(n3666), .ZN(n2286) );
  NAND2_X1 U2930 ( .A1(n3663), .A2(n3008), .ZN(n2914) );
  NOR2_X1 U2931 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  AND4_X1 U2932 ( .A1(n2297), .A2(n2296), .A3(n2295), .A4(n2294), .ZN(n2298)
         );
  NOR2_X1 U2933 ( .A1(n2547), .A2(n4520), .ZN(n2553) );
  INV_X1 U2934 ( .A(n3613), .ZN(n3614) );
  INV_X1 U2935 ( .A(n4356), .ZN(n3466) );
  NOR2_X1 U2936 ( .A1(n2783), .A2(n2765), .ZN(n2695) );
  OR2_X1 U2937 ( .A1(n4215), .A2(n4033), .ZN(n3455) );
  AND2_X1 U2938 ( .A1(n4244), .A2(n4094), .ZN(n3457) );
  AND2_X1 U2939 ( .A1(n4182), .A2(n4264), .ZN(n2524) );
  OR2_X1 U2940 ( .A1(n3848), .A2(n3324), .ZN(n2498) );
  INV_X1 U2941 ( .A(n4166), .ZN(n4264) );
  INV_X1 U2942 ( .A(n3149), .ZN(n3084) );
  AND2_X1 U2943 ( .A1(n2468), .A2(IR_REG_31__SCAN_IN), .ZN(n2469) );
  OR2_X1 U2944 ( .A1(n2573), .A2(n3723), .ZN(n2583) );
  OR2_X1 U2945 ( .A1(n2539), .A2(n2538), .ZN(n2547) );
  OR2_X1 U2946 ( .A1(n3206), .A2(n3205), .ZN(n3207) );
  OR2_X1 U2947 ( .A1(n2599), .A2(n2598), .ZN(n2608) );
  AND2_X1 U2948 ( .A1(n2981), .A2(n3577), .ZN(n2982) );
  NAND2_X1 U2949 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
  INV_X1 U2950 ( .A(n4362), .ZN(n2865) );
  INV_X1 U2951 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3834) );
  INV_X1 U2952 ( .A(n4178), .ZN(n4273) );
  INV_X1 U2953 ( .A(n3857), .ZN(n3187) );
  INV_X1 U2954 ( .A(n4275), .ZN(n4289) );
  INV_X1 U2955 ( .A(n2994), .ZN(n3038) );
  INV_X1 U2956 ( .A(n4204), .ZN(n3974) );
  INV_X1 U2957 ( .A(n2572), .ZN(n4060) );
  INV_X1 U2958 ( .A(n3377), .ZN(n3281) );
  INV_X1 U2959 ( .A(n4171), .ZN(n4122) );
  NAND2_X1 U2960 ( .A1(n2415), .A2(REG3_REG_7__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U2961 ( .A1(n2317), .A2(REG3_REG_10__SCAN_IN), .ZN(n2461) );
  AND2_X1 U2962 ( .A1(n2629), .A2(n2620), .ZN(n3695) );
  AND2_X1 U2963 ( .A1(n2599), .A2(n2584), .ZN(n4030) );
  NAND2_X1 U2964 ( .A1(n2316), .A2(n2315), .ZN(n2453) );
  OR2_X1 U2965 ( .A1(n2461), .A2(n2460), .ZN(n2475) );
  AND2_X1 U2966 ( .A1(n2608), .A2(n2600), .ZN(n3999) );
  OR2_X1 U2967 ( .A1(n2500), .A2(n3834), .ZN(n2502) );
  AND2_X1 U2968 ( .A1(n2626), .A2(n2625), .ZN(n3684) );
  AND4_X1 U2969 ( .A1(n2325), .A2(n2324), .A3(n2323), .A4(n2322), .ZN(n4268)
         );
  NAND2_X1 U2970 ( .A1(n3415), .A2(REG2_REG_0__SCAN_IN), .ZN(n2349) );
  NOR2_X1 U2971 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4445), .ZN(n4446) );
  OR2_X1 U2972 ( .A1(n2678), .A2(n2677), .ZN(n2897) );
  INV_X1 U2973 ( .A(n4274), .ZN(n4287) );
  AND2_X1 U2974 ( .A1(n3439), .A2(n3506), .ZN(n4176) );
  INV_X1 U2975 ( .A(n4154), .ZN(n4177) );
  AND2_X1 U2976 ( .A1(n4473), .A2(n4289), .ZN(n4183) );
  INV_X1 U2977 ( .A(n4470), .ZN(n4186) );
  NAND2_X1 U2978 ( .A1(n2714), .A2(n2713), .ZN(n2752) );
  NAND2_X1 U2979 ( .A1(n4100), .A2(n4497), .ZN(n4506) );
  AND2_X1 U2980 ( .A1(n3020), .A2(n3019), .ZN(n4505) );
  INV_X1 U2981 ( .A(n2752), .ZN(n2881) );
  XNOR2_X1 U2982 ( .A(n2636), .B(n2142), .ZN(n2882) );
  AND2_X1 U2983 ( .A1(n2472), .A2(n2482), .ZN(n3922) );
  AND2_X1 U2984 ( .A1(n2791), .A2(n2789), .ZN(n4463) );
  OR2_X1 U2985 ( .A1(n2922), .A2(n2896), .ZN(n3827) );
  INV_X1 U2986 ( .A(n3684), .ZN(n4207) );
  INV_X1 U2987 ( .A(n3739), .ZN(n4244) );
  INV_X1 U2988 ( .A(n4294), .ZN(n3848) );
  NAND2_X1 U2989 ( .A1(n2809), .A2(n2897), .ZN(n4469) );
  INV_X1 U2990 ( .A(n4411), .ZN(n4459) );
  INV_X1 U2991 ( .A(n4473), .ZN(n4087) );
  INV_X1 U2992 ( .A(n4473), .ZN(n4482) );
  NAND2_X1 U2993 ( .A1(n4473), .A2(n3034), .ZN(n4154) );
  NAND2_X1 U2994 ( .A1(n2721), .A2(n2720), .ZN(n2722) );
  NAND2_X1 U2995 ( .A1(n4518), .A2(n4146), .ZN(n4299) );
  NAND2_X1 U2996 ( .A1(n2721), .A2(n2727), .ZN(n2728) );
  NAND2_X1 U2997 ( .A1(n4513), .A2(n4146), .ZN(n4347) );
  AND3_X1 U2998 ( .A1(n4510), .A2(n4509), .A3(n4508), .ZN(n4517) );
  INV_X2 U2999 ( .A(n4511), .ZN(n4513) );
  INV_X1 U3000 ( .A(n2696), .ZN(n2784) );
  AND2_X1 U3001 ( .A1(n2787), .A2(STATE_REG_SCAN_IN), .ZN(n4484) );
  INV_X1 U3002 ( .A(n3921), .ZN(n4490) );
  INV_X1 U3003 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3004 ( .A1(n2299), .A2(n2288), .ZN(n2467) );
  INV_X1 U3005 ( .A(IR_REG_12__SCAN_IN), .ZN(n2289) );
  NAND2_X1 U3006 ( .A1(n2297), .A2(n2289), .ZN(n2290) );
  INV_X1 U3007 ( .A(IR_REG_14__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U3008 ( .A1(n2496), .A2(n2291), .ZN(n2292) );
  NAND2_X1 U3009 ( .A1(n2292), .A2(IR_REG_31__SCAN_IN), .ZN(n2508) );
  INV_X1 U3010 ( .A(IR_REG_15__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3011 ( .A1(n2508), .A2(n2507), .ZN(n2510) );
  NAND2_X1 U3012 ( .A1(n2510), .A2(IR_REG_31__SCAN_IN), .ZN(n2293) );
  XNOR2_X1 U3013 ( .A(n2293), .B(IR_REG_16__SCAN_IN), .ZN(n3942) );
  MUX2_X1 U3014 ( .A(DATAI_16_), .B(n3942), .S(n3419), .Z(n4178) );
  NAND2_X1 U3015 ( .A1(n2676), .A2(IR_REG_31__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U3016 ( .A1(n2353), .A2(REG0_REG_16__SCAN_IN), .ZN(n2325) );
  INV_X1 U3017 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2313) );
  OR2_X1 U3018 ( .A1(n2341), .A2(n2313), .ZN(n2324) );
  NAND2_X1 U3019 ( .A1(n2502), .A2(n2318), .ZN(n2319) );
  NAND2_X1 U3020 ( .A1(n2514), .A2(n2319), .ZN(n3756) );
  OR2_X1 U3021 ( .A1(n2337), .A2(n3756), .ZN(n2323) );
  INV_X1 U3022 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2321) );
  OR2_X1 U3023 ( .A1(n3418), .A2(n2321), .ZN(n2322) );
  NAND2_X1 U3024 ( .A1(n2353), .A2(REG0_REG_13__SCAN_IN), .ZN(n2333) );
  INV_X1 U3025 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4410) );
  OR2_X1 U3026 ( .A1(n2341), .A2(n4410), .ZN(n2332) );
  INV_X1 U3027 ( .A(n2326), .ZN(n2489) );
  INV_X1 U3028 ( .A(n2327), .ZN(n2477) );
  INV_X1 U3029 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U3030 ( .A1(n2477), .A2(n2328), .ZN(n2329) );
  NAND2_X1 U3031 ( .A1(n2489), .A2(n2329), .ZN(n3797) );
  OR2_X1 U3032 ( .A1(n2337), .A2(n3797), .ZN(n2331) );
  INV_X1 U3033 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3409) );
  OR2_X1 U3034 ( .A1(n3418), .A2(n3409), .ZN(n2330) );
  INV_X1 U3035 ( .A(DATAI_13_), .ZN(n2336) );
  NAND2_X1 U3036 ( .A1(n2334), .A2(IR_REG_31__SCAN_IN), .ZN(n2335) );
  XNOR2_X1 U3037 ( .A(n2335), .B(IR_REG_13__SCAN_IN), .ZN(n3921) );
  MUX2_X1 U3038 ( .A(n2336), .B(n4490), .S(n3419), .Z(n3793) );
  INV_X1 U3039 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3004) );
  INV_X1 U3040 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2338) );
  NAND2_X1 U3041 ( .A1(n3415), .A2(REG2_REG_1__SCAN_IN), .ZN(n2343) );
  INV_X1 U3042 ( .A(n3008), .ZN(n2915) );
  INV_X1 U3043 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2902) );
  INV_X1 U3044 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2346) );
  AND2_X1 U3045 ( .A1(n3864), .A2(n2952), .ZN(n2942) );
  NAND2_X1 U3046 ( .A1(n3475), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U3047 ( .A1(n3862), .A2(n3008), .ZN(n2352) );
  NAND2_X1 U3048 ( .A1(n2944), .A2(n2352), .ZN(n2742) );
  INV_X1 U3049 ( .A(n2742), .ZN(n2359) );
  INV_X1 U3050 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3874) );
  OR2_X1 U3051 ( .A1(n2337), .A2(n3874), .ZN(n2355) );
  INV_X1 U3052 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2813) );
  OR2_X1 U3053 ( .A1(n2341), .A2(n3879), .ZN(n2354) );
  MUX2_X1 U3054 ( .A(DATAI_2_), .B(n4364), .S(n2357), .Z(n2961) );
  NAND2_X1 U3055 ( .A1(n2932), .A2(n2961), .ZN(n3515) );
  INV_X1 U3056 ( .A(n2961), .ZN(n2931) );
  INV_X1 U3057 ( .A(n3476), .ZN(n2358) );
  NAND2_X1 U3058 ( .A1(n2359), .A2(n2358), .ZN(n2744) );
  NAND2_X1 U3059 ( .A1(n2932), .A2(n2931), .ZN(n2360) );
  INV_X1 U3060 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3895) );
  OR2_X1 U3061 ( .A1(n2341), .A2(n3895), .ZN(n2365) );
  NAND2_X1 U3062 ( .A1(n2549), .A2(REG1_REG_3__SCAN_IN), .ZN(n2362) );
  OR2_X1 U3063 ( .A1(n2337), .A2(REG3_REG_3__SCAN_IN), .ZN(n2361) );
  INV_X1 U3064 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3065 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3066 ( .A1(n2367), .A2(n4618), .ZN(n2378) );
  OR2_X1 U3067 ( .A1(n2367), .A2(n4618), .ZN(n2368) );
  MUX2_X1 U3068 ( .A(DATAI_3_), .B(n4363), .S(n3419), .Z(n2994) );
  NAND2_X1 U3069 ( .A1(n3860), .A2(n2994), .ZN(n3012) );
  NAND2_X1 U3070 ( .A1(n3415), .A2(REG2_REG_4__SCAN_IN), .ZN(n2377) );
  INV_X1 U3071 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2369) );
  OR2_X1 U3072 ( .A1(n2347), .A2(n2369), .ZN(n2376) );
  INV_X1 U3073 ( .A(n2370), .ZN(n2384) );
  INV_X1 U3074 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2984) );
  INV_X1 U3075 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3076 ( .A1(n2984), .A2(n2371), .ZN(n2372) );
  NAND2_X1 U3077 ( .A1(n2384), .A2(n2372), .ZN(n3105) );
  OR2_X1 U3078 ( .A1(n2337), .A2(n3105), .ZN(n2375) );
  INV_X1 U3079 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2373) );
  OR2_X1 U3080 ( .A1(n3418), .A2(n2373), .ZN(n2374) );
  NAND2_X1 U3081 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2379) );
  XNOR2_X1 U3082 ( .A(n2379), .B(IR_REG_4__SCAN_IN), .ZN(n4362) );
  MUX2_X1 U3083 ( .A(DATAI_4_), .B(n4362), .S(n3419), .Z(n3022) );
  NAND2_X1 U3084 ( .A1(n3859), .A2(n3022), .ZN(n2381) );
  AND2_X1 U3085 ( .A1(n3012), .A2(n2381), .ZN(n2380) );
  NAND2_X1 U3086 ( .A1(n3013), .A2(n2380), .ZN(n3049) );
  INV_X1 U3087 ( .A(n3022), .ZN(n3100) );
  NAND2_X1 U3088 ( .A1(n3859), .A2(n3100), .ZN(n3525) );
  NAND2_X1 U3089 ( .A1(n3148), .A2(n3022), .ZN(n3521) );
  NAND2_X1 U3090 ( .A1(n3525), .A2(n3521), .ZN(n3017) );
  NAND2_X1 U3091 ( .A1(n3099), .A2(n3038), .ZN(n3015) );
  AND2_X1 U3092 ( .A1(n3017), .A2(n3015), .ZN(n3014) );
  INV_X1 U3093 ( .A(n3014), .ZN(n2382) );
  NAND2_X1 U3094 ( .A1(n2353), .A2(REG0_REG_5__SCAN_IN), .ZN(n2391) );
  INV_X1 U3095 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2828) );
  OR2_X1 U3096 ( .A1(n3418), .A2(n2828), .ZN(n2390) );
  INV_X1 U3097 ( .A(n2403), .ZN(n2386) );
  INV_X1 U3098 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U3099 ( .A1(n2384), .A2(n2383), .ZN(n2385) );
  NAND2_X1 U3100 ( .A1(n2386), .A2(n2385), .ZN(n3154) );
  OR2_X1 U3101 ( .A1(n2337), .A2(n3154), .ZN(n2389) );
  INV_X1 U3102 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2387) );
  OR2_X1 U3103 ( .A1(n2341), .A2(n2387), .ZN(n2388) );
  INV_X1 U3104 ( .A(DATAI_5_), .ZN(n4657) );
  INV_X1 U3105 ( .A(n2392), .ZN(n2393) );
  OR2_X1 U3106 ( .A1(n2366), .A2(n2393), .ZN(n2395) );
  NAND2_X1 U3107 ( .A1(n2395), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  MUX2_X1 U3108 ( .A(n2394), .B(IR_REG_31__SCAN_IN), .S(n2396), .Z(n2398) );
  INV_X1 U3109 ( .A(n2395), .ZN(n2397) );
  NAND2_X1 U3110 ( .A1(n2397), .A2(n2396), .ZN(n2411) );
  NAND2_X1 U3111 ( .A1(n2398), .A2(n2411), .ZN(n2829) );
  MUX2_X1 U3112 ( .A(n4657), .B(n2829), .S(n3419), .Z(n3149) );
  NAND2_X1 U3113 ( .A1(n3137), .A2(n3149), .ZN(n2399) );
  NAND2_X1 U3114 ( .A1(n3049), .A2(n2400), .ZN(n2402) );
  INV_X1 U3115 ( .A(n3137), .ZN(n3858) );
  NAND2_X1 U3116 ( .A1(n3858), .A2(n3084), .ZN(n2401) );
  NOR2_X1 U3117 ( .A1(n2403), .A2(REG3_REG_6__SCAN_IN), .ZN(n2404) );
  NOR2_X1 U3118 ( .A1(n2415), .A2(n2404), .ZN(n3141) );
  NAND2_X1 U3119 ( .A1(n2633), .A2(n3141), .ZN(n2410) );
  NAND2_X1 U3120 ( .A1(n2549), .A2(REG1_REG_6__SCAN_IN), .ZN(n2409) );
  INV_X1 U3121 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2405) );
  OR2_X1 U3122 ( .A1(n2341), .A2(n2405), .ZN(n2408) );
  INV_X1 U3123 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2406) );
  OR2_X1 U3124 ( .A1(n2347), .A2(n2406), .ZN(n2407) );
  NAND4_X1 U3125 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), .ZN(n3857)
         );
  NAND2_X1 U3126 ( .A1(n2411), .A2(IR_REG_31__SCAN_IN), .ZN(n2412) );
  XNOR2_X1 U3127 ( .A(n2412), .B(IR_REG_6__SCAN_IN), .ZN(n4360) );
  MUX2_X1 U3128 ( .A(DATAI_6_), .B(n4360), .S(n3419), .Z(n3110) );
  AND2_X1 U3129 ( .A1(n3857), .A2(n3110), .ZN(n2413) );
  NAND2_X1 U3130 ( .A1(n2353), .A2(REG0_REG_7__SCAN_IN), .ZN(n2420) );
  INV_X1 U3131 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2414) );
  OR2_X1 U3132 ( .A1(n2341), .A2(n2414), .ZN(n2419) );
  OAI21_X1 U3133 ( .B1(n2415), .B2(REG3_REG_7__SCAN_IN), .A(n2440), .ZN(n3193)
         );
  OR2_X1 U3134 ( .A1(n2337), .A2(n3193), .ZN(n2418) );
  INV_X1 U3135 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2416) );
  OR2_X1 U3136 ( .A1(n3418), .A2(n2416), .ZN(n2417) );
  AND2_X1 U3137 ( .A1(n2421), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3138 ( .A1(n2422), .A2(IR_REG_7__SCAN_IN), .ZN(n2425) );
  INV_X1 U3139 ( .A(n2422), .ZN(n2424) );
  NAND2_X1 U3140 ( .A1(n2424), .A2(n2423), .ZN(n2431) );
  MUX2_X1 U3141 ( .A(DATAI_7_), .B(n4359), .S(n3419), .Z(n3074) );
  NAND2_X1 U3142 ( .A1(n3216), .A2(n3074), .ZN(n2650) );
  INV_X1 U3143 ( .A(n3074), .ZN(n3188) );
  NAND2_X1 U3144 ( .A1(n3855), .A2(n3188), .ZN(n3531) );
  NAND2_X1 U3145 ( .A1(n3855), .A2(n3074), .ZN(n2426) );
  NAND2_X1 U3146 ( .A1(n3080), .A2(n2426), .ZN(n3165) );
  NAND2_X1 U3147 ( .A1(n2353), .A2(REG0_REG_8__SCAN_IN), .ZN(n2430) );
  INV_X1 U31480 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3927) );
  OR2_X1 U31490 ( .A1(n3418), .A2(n3927), .ZN(n2429) );
  INV_X1 U3150 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2439) );
  XNOR2_X1 U3151 ( .A(n2440), .B(n2439), .ZN(n4471) );
  OR2_X1 U3152 ( .A1(n2337), .A2(n4471), .ZN(n2428) );
  INV_X1 U3153 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4472) );
  OR2_X1 U3154 ( .A1(n2341), .A2(n4472), .ZN(n2427) );
  INV_X1 U3155 ( .A(DATAI_8_), .ZN(n2434) );
  NAND2_X1 U3156 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  XNOR2_X1 U3157 ( .A(n2433), .B(n2432), .ZN(n4358) );
  MUX2_X1 U3158 ( .A(n2434), .B(n4358), .S(n3419), .Z(n3217) );
  NAND2_X1 U3159 ( .A1(n3231), .A2(n3217), .ZN(n2435) );
  NAND2_X1 U3160 ( .A1(n3165), .A2(n2435), .ZN(n2437) );
  NAND2_X1 U3161 ( .A1(n3854), .A2(n3175), .ZN(n2436) );
  NAND2_X1 U3162 ( .A1(n2437), .A2(n2436), .ZN(n3162) );
  INV_X1 U3163 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2438) );
  OAI21_X1 U3164 ( .B1(n2440), .B2(n2439), .A(n2438), .ZN(n2441) );
  NAND2_X1 U3165 ( .A1(n2441), .A2(n2453), .ZN(n3236) );
  OR2_X1 U3166 ( .A1(n2337), .A2(n3236), .ZN(n2447) );
  INV_X1 U3167 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2442) );
  OR2_X1 U3168 ( .A1(n3418), .A2(n2442), .ZN(n2446) );
  NAND2_X1 U3169 ( .A1(n2353), .A2(REG0_REG_9__SCAN_IN), .ZN(n2445) );
  INV_X1 U3170 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2443) );
  OR2_X1 U3171 ( .A1(n2341), .A2(n2443), .ZN(n2444) );
  NAND4_X1 U3172 ( .A1(n2447), .A2(n2446), .A3(n2445), .A4(n2444), .ZN(n3853)
         );
  NOR2_X1 U3173 ( .A1(n2299), .A2(n2775), .ZN(n2448) );
  MUX2_X1 U3174 ( .A(n2775), .B(n2448), .S(IR_REG_9__SCAN_IN), .Z(n2449) );
  INV_X1 U3175 ( .A(n2449), .ZN(n2450) );
  MUX2_X1 U3176 ( .A(DATAI_9_), .B(n3923), .S(n3419), .Z(n3226) );
  NAND2_X1 U3177 ( .A1(n3259), .A2(n3232), .ZN(n2451) );
  INV_X1 U3178 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3271) );
  OR2_X1 U3179 ( .A1(n3418), .A2(n3271), .ZN(n2458) );
  INV_X1 U3180 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3181 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  NAND2_X1 U3182 ( .A1(n2461), .A2(n2454), .ZN(n3264) );
  OR2_X1 U3183 ( .A1(n2337), .A2(n3264), .ZN(n2457) );
  NAND2_X1 U3184 ( .A1(n2353), .A2(REG0_REG_10__SCAN_IN), .ZN(n2456) );
  INV_X1 U3185 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3240) );
  OR2_X1 U3186 ( .A1(n2341), .A2(n3240), .ZN(n2455) );
  NAND2_X1 U3187 ( .A1(n2467), .A2(IR_REG_31__SCAN_IN), .ZN(n2459) );
  XNOR2_X1 U3188 ( .A(n2459), .B(IR_REG_10__SCAN_IN), .ZN(n3930) );
  MUX2_X1 U3189 ( .A(DATAI_10_), .B(n3930), .S(n3419), .Z(n3252) );
  NAND2_X1 U3190 ( .A1(n2353), .A2(REG0_REG_11__SCAN_IN), .ZN(n2466) );
  INV_X1 U3191 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3306) );
  OR2_X1 U3192 ( .A1(n3418), .A2(n3306), .ZN(n2465) );
  NAND2_X1 U3193 ( .A1(n2461), .A2(n2460), .ZN(n2462) );
  NAND2_X1 U3194 ( .A1(n2475), .A2(n2462), .ZN(n3580) );
  OR2_X1 U3195 ( .A1(n2337), .A2(n3580), .ZN(n2464) );
  INV_X1 U3196 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3581) );
  OR2_X1 U3197 ( .A1(n2341), .A2(n3581), .ZN(n2463) );
  OR2_X1 U3198 ( .A1(n2467), .A2(IR_REG_10__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3199 ( .A1(n2469), .A2(IR_REG_11__SCAN_IN), .ZN(n2472) );
  INV_X1 U3200 ( .A(n2469), .ZN(n2471) );
  INV_X1 U3201 ( .A(IR_REG_11__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3202 ( .A1(n2471), .A2(n2470), .ZN(n2482) );
  MUX2_X1 U3203 ( .A(DATAI_11_), .B(n3922), .S(n3419), .Z(n3297) );
  NAND2_X1 U3204 ( .A1(n3376), .A2(n3297), .ZN(n3284) );
  NAND2_X1 U3205 ( .A1(n3851), .A2(n3317), .ZN(n3286) );
  NAND2_X1 U3206 ( .A1(n3376), .A2(n3317), .ZN(n2473) );
  NAND2_X1 U3207 ( .A1(n3295), .A2(n2473), .ZN(n3277) );
  NAND2_X1 U3208 ( .A1(n2353), .A2(REG0_REG_12__SCAN_IN), .ZN(n2481) );
  INV_X1 U3209 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3279) );
  OR2_X1 U32100 ( .A1(n2341), .A2(n3279), .ZN(n2480) );
  NAND2_X1 U32110 ( .A1(n2475), .A2(n2474), .ZN(n2476) );
  NAND2_X1 U32120 ( .A1(n2477), .A2(n2476), .ZN(n3375) );
  OR2_X1 U32130 ( .A1(n2337), .A2(n3375), .ZN(n2479) );
  INV_X1 U32140 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3361) );
  OR2_X1 U32150 ( .A1(n3418), .A2(n3361), .ZN(n2478) );
  INV_X1 U32160 ( .A(DATAI_12_), .ZN(n2484) );
  NAND2_X1 U32170 ( .A1(n2482), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  XNOR2_X1 U32180 ( .A(n2483), .B(IR_REG_12__SCAN_IN), .ZN(n3934) );
  MUX2_X1 U32190 ( .A(n2484), .B(n4491), .S(n3419), .Z(n3377) );
  NAND2_X1 U32200 ( .A1(n3277), .A2(n2284), .ZN(n2486) );
  INV_X1 U32210 ( .A(n3793), .ZN(n2487) );
  NAND2_X1 U32220 ( .A1(n2353), .A2(REG0_REG_14__SCAN_IN), .ZN(n2495) );
  INV_X1 U32230 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3404) );
  OR2_X1 U32240 ( .A1(n3418), .A2(n3404), .ZN(n2494) );
  INV_X1 U32250 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U32260 ( .A1(n2489), .A2(n4652), .ZN(n2490) );
  NAND2_X1 U32270 ( .A1(n2500), .A2(n2490), .ZN(n3326) );
  OR2_X1 U32280 ( .A1(n2337), .A2(n3326), .ZN(n2493) );
  INV_X1 U32290 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2491) );
  OR2_X1 U32300 ( .A1(n2341), .A2(n2491), .ZN(n2492) );
  OR2_X1 U32310 ( .A1(n2496), .A2(n2775), .ZN(n2497) );
  XNOR2_X1 U32320 ( .A(n2497), .B(IR_REG_14__SCAN_IN), .ZN(n3938) );
  MUX2_X1 U32330 ( .A(DATAI_14_), .B(n3938), .S(n3419), .Z(n3324) );
  NAND2_X1 U32340 ( .A1(n4294), .A2(n3324), .ZN(n3430) );
  NAND2_X1 U32350 ( .A1(n3848), .A2(n3712), .ZN(n3505) );
  NAND2_X1 U32360 ( .A1(n3430), .A2(n3505), .ZN(n3322) );
  NAND2_X1 U32370 ( .A1(n2353), .A2(REG0_REG_15__SCAN_IN), .ZN(n2506) );
  INV_X1 U32380 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2499) );
  OR2_X1 U32390 ( .A1(n2341), .A2(n2499), .ZN(n2505) );
  NAND2_X1 U32400 ( .A1(n2500), .A2(n3834), .ZN(n2501) );
  NAND2_X1 U32410 ( .A1(n2502), .A2(n2501), .ZN(n3842) );
  OR2_X1 U32420 ( .A1(n2337), .A2(n3842), .ZN(n2504) );
  INV_X1 U32430 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4297) );
  OR2_X1 U32440 ( .A1(n3418), .A2(n4297), .ZN(n2503) );
  INV_X1 U32450 ( .A(DATAI_15_), .ZN(n4641) );
  OR2_X1 U32460 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  MUX2_X1 U32470 ( .A(n4641), .B(n4489), .S(n3419), .Z(n3836) );
  NAND2_X1 U32480 ( .A1(n3386), .A2(n2280), .ZN(n2512) );
  NAND2_X1 U32490 ( .A1(n2512), .A2(n2511), .ZN(n4175) );
  NAND2_X1 U32500 ( .A1(n4268), .A2(n4178), .ZN(n3439) );
  NAND2_X1 U32510 ( .A1(n4290), .A2(n4273), .ZN(n3506) );
  NAND2_X1 U32520 ( .A1(n2353), .A2(REG0_REG_17__SCAN_IN), .ZN(n2520) );
  INV_X1 U32530 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4271) );
  OR2_X1 U32540 ( .A1(n3418), .A2(n4271), .ZN(n2519) );
  INV_X1 U32550 ( .A(n2528), .ZN(n2530) );
  NAND2_X1 U32560 ( .A1(n2514), .A2(n2513), .ZN(n2515) );
  NAND2_X1 U32570 ( .A1(n2530), .A2(n2515), .ZN(n4162) );
  OR2_X1 U32580 ( .A1(n2337), .A2(n4162), .ZN(n2518) );
  INV_X1 U32590 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2516) );
  OR2_X1 U32600 ( .A1(n2341), .A2(n2516), .ZN(n2517) );
  INV_X1 U32610 ( .A(DATAI_17_), .ZN(n2523) );
  OR2_X1 U32620 ( .A1(n2521), .A2(n2775), .ZN(n2522) );
  XNOR2_X1 U32630 ( .A(n2522), .B(IR_REG_17__SCAN_IN), .ZN(n3945) );
  MUX2_X1 U32640 ( .A(n2523), .B(n4487), .S(n3419), .Z(n4166) );
  INV_X1 U32650 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3947) );
  OR2_X1 U32660 ( .A1(n3418), .A2(n3947), .ZN(n2527) );
  INV_X1 U32670 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2525) );
  OR2_X1 U32680 ( .A1(n2347), .A2(n2525), .ZN(n2526) );
  AND2_X1 U32690 ( .A1(n2527), .A2(n2526), .ZN(n2534) );
  INV_X1 U32700 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32710 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  NAND2_X1 U32720 ( .A1(n2539), .A2(n2531), .ZN(n4149) );
  OR2_X1 U32730 ( .A1(n4149), .A2(n2337), .ZN(n2533) );
  NAND2_X1 U32740 ( .A1(n3415), .A2(REG2_REG_18__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32750 ( .A1(n2544), .A2(IR_REG_31__SCAN_IN), .ZN(n2536) );
  XNOR2_X1 U32760 ( .A(n2536), .B(IR_REG_18__SCAN_IN), .ZN(n3919) );
  MUX2_X1 U32770 ( .A(DATAI_18_), .B(n3919), .S(n3419), .Z(n4140) );
  NAND2_X1 U32780 ( .A1(n4119), .A2(n4140), .ZN(n4114) );
  NAND2_X1 U32790 ( .A1(n4265), .A2(n4147), .ZN(n4115) );
  NAND2_X1 U32800 ( .A1(n4114), .A2(n4115), .ZN(n4139) );
  NAND2_X1 U32810 ( .A1(n4136), .A2(n4139), .ZN(n4135) );
  NAND2_X1 U32820 ( .A1(n4135), .A2(n2537), .ZN(n4111) );
  INV_X1 U32830 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32840 ( .A1(n2539), .A2(n2538), .ZN(n2540) );
  AND2_X1 U32850 ( .A1(n2547), .A2(n2540), .ZN(n4128) );
  NAND2_X1 U32860 ( .A1(n4128), .A2(n2633), .ZN(n2543) );
  AOI22_X1 U32870 ( .A1(n3415), .A2(REG2_REG_19__SCAN_IN), .B1(n2353), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2542) );
  INV_X1 U32880 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4258) );
  OR2_X1 U32890 ( .A1(n3418), .A2(n4258), .ZN(n2541) );
  INV_X1 U32900 ( .A(n2643), .ZN(n2545) );
  MUX2_X1 U32910 ( .A(DATAI_19_), .B(n4357), .S(n3419), .Z(n2716) );
  NAND2_X1 U32920 ( .A1(n4141), .A2(n2716), .ZN(n2546) );
  AOI21_X1 U32930 ( .B1(n4111), .B2(n2546), .A(n2080), .ZN(n4088) );
  INV_X1 U32940 ( .A(n2553), .ZN(n2554) );
  NAND2_X1 U32950 ( .A1(n2547), .A2(n4520), .ZN(n2548) );
  NAND2_X1 U32960 ( .A1(n2554), .A2(n2548), .ZN(n3781) );
  OR2_X1 U32970 ( .A1(n3781), .A2(n2337), .ZN(n2552) );
  AOI22_X1 U32980 ( .A1(n3415), .A2(REG2_REG_20__SCAN_IN), .B1(n2353), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32990 ( .A1(n2549), .A2(REG1_REG_20__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U33000 ( .A1(n3739), .A2(n4104), .ZN(n3458) );
  INV_X1 U33010 ( .A(n2563), .ZN(n2564) );
  INV_X1 U33020 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3738) );
  NAND2_X1 U33030 ( .A1(n2554), .A2(n3738), .ZN(n2555) );
  NAND2_X1 U33040 ( .A1(n4079), .A2(n2633), .ZN(n2560) );
  INV_X1 U33050 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4250) );
  NAND2_X1 U33060 ( .A1(n2353), .A2(REG0_REG_21__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U33070 ( .A1(n3415), .A2(REG2_REG_21__SCAN_IN), .ZN(n2556) );
  OAI211_X1 U33080 ( .C1(n3418), .C2(n4250), .A(n2557), .B(n2556), .ZN(n2558)
         );
  INV_X1 U33090 ( .A(n2558), .ZN(n2559) );
  INV_X1 U33100 ( .A(n4096), .ZN(n3847) );
  INV_X1 U33110 ( .A(DATAI_21_), .ZN(n2561) );
  NAND2_X1 U33120 ( .A1(n3847), .A2(n4242), .ZN(n2562) );
  INV_X1 U33130 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U33140 ( .A1(n2564), .A2(n3801), .ZN(n2565) );
  NAND2_X1 U33150 ( .A1(n2573), .A2(n2565), .ZN(n3800) );
  OR2_X1 U33160 ( .A1(n3800), .A2(n2337), .ZN(n2570) );
  INV_X1 U33170 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U33180 ( .A1(n2353), .A2(REG0_REG_22__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U33190 ( .A1(n3415), .A2(REG2_REG_22__SCAN_IN), .ZN(n2566) );
  OAI211_X1 U33200 ( .C1(n3418), .C2(n4240), .A(n2567), .B(n2566), .ZN(n2568)
         );
  INV_X1 U33210 ( .A(n2568), .ZN(n2569) );
  INV_X1 U33220 ( .A(DATAI_22_), .ZN(n2571) );
  NOR2_X1 U33230 ( .A1(n3419), .A2(n2571), .ZN(n2572) );
  NAND2_X1 U33240 ( .A1(n4247), .A2(n2572), .ZN(n4042) );
  INV_X1 U33250 ( .A(n4247), .ZN(n4078) );
  NAND2_X1 U33260 ( .A1(n4078), .A2(n4060), .ZN(n2663) );
  NAND2_X1 U33270 ( .A1(n4042), .A2(n2663), .ZN(n4065) );
  INV_X1 U33280 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U33290 ( .A1(n2573), .A2(n3723), .ZN(n2574) );
  AND2_X1 U33300 ( .A1(n2583), .A2(n2574), .ZN(n4051) );
  NAND2_X1 U33310 ( .A1(n4051), .A2(n2633), .ZN(n2579) );
  INV_X1 U33320 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U33330 ( .A1(n3415), .A2(REG2_REG_23__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U33340 ( .A1(n2353), .A2(REG0_REG_23__SCAN_IN), .ZN(n2575) );
  OAI211_X1 U33350 ( .C1(n4234), .C2(n3418), .A(n2576), .B(n2575), .ZN(n2577)
         );
  INV_X1 U33360 ( .A(n2577), .ZN(n2578) );
  INV_X1 U33370 ( .A(DATAI_23_), .ZN(n2580) );
  NAND2_X1 U33380 ( .A1(n4224), .A2(n3647), .ZN(n2581) );
  INV_X1 U33390 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U33400 ( .A1(n2583), .A2(n4654), .ZN(n2584) );
  NAND2_X1 U33410 ( .A1(n4030), .A2(n2633), .ZN(n2589) );
  INV_X1 U33420 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U33430 ( .A1(n3415), .A2(REG2_REG_24__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U33440 ( .A1(n2353), .A2(REG0_REG_24__SCAN_IN), .ZN(n2585) );
  OAI211_X1 U33450 ( .C1(n4230), .C2(n3418), .A(n2586), .B(n2585), .ZN(n2587)
         );
  INV_X1 U33460 ( .A(n2587), .ZN(n2588) );
  NAND2_X1 U33470 ( .A1(n2308), .A2(DATAI_24_), .ZN(n4033) );
  NAND2_X1 U33480 ( .A1(n3747), .A2(n4033), .ZN(n2590) );
  XNOR2_X1 U33490 ( .A(n2599), .B(REG3_REG_25__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U33500 ( .A1(n4013), .A2(n2633), .ZN(n2595) );
  INV_X1 U33510 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4221) );
  NAND2_X1 U33520 ( .A1(n3415), .A2(REG2_REG_25__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U3353 ( .A1(n2353), .A2(REG0_REG_25__SCAN_IN), .ZN(n2591) );
  OAI211_X1 U33540 ( .C1(n4221), .C2(n3418), .A(n2592), .B(n2591), .ZN(n2593)
         );
  INV_X1 U3355 ( .A(n2593), .ZN(n2594) );
  INV_X1 U3356 ( .A(DATAI_25_), .ZN(n4534) );
  NOR2_X1 U3357 ( .A1(n4029), .A2(n4214), .ZN(n2597) );
  NAND2_X1 U3358 ( .A1(n4029), .A2(n4214), .ZN(n2596) );
  NAND2_X1 U3359 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2598) );
  INV_X1 U3360 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4668) );
  INV_X1 U3361 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3821) );
  OAI21_X1 U3362 ( .B1(n2599), .B2(n4668), .A(n3821), .ZN(n2600) );
  NAND2_X1 U3363 ( .A1(n3999), .A2(n2633), .ZN(n2605) );
  INV_X1 U3364 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U3365 ( .A1(n3415), .A2(REG2_REG_26__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3366 ( .A1(n2353), .A2(REG0_REG_26__SCAN_IN), .ZN(n2601) );
  OAI211_X1 U3367 ( .C1(n4212), .C2(n3418), .A(n2602), .B(n2601), .ZN(n2603)
         );
  INV_X1 U3368 ( .A(n2603), .ZN(n2604) );
  NAND2_X1 U3369 ( .A1(n2308), .A2(DATAI_26_), .ZN(n3998) );
  NOR2_X1 U3370 ( .A1(n4218), .A2(n3998), .ZN(n2606) );
  INV_X1 U3371 ( .A(n2608), .ZN(n2607) );
  NAND2_X1 U3372 ( .A1(n2607), .A2(REG3_REG_27__SCAN_IN), .ZN(n2619) );
  INV_X1 U3373 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U3374 ( .A1(n2608), .A2(n4573), .ZN(n2609) );
  NAND2_X1 U3375 ( .A1(n2619), .A2(n2609), .ZN(n3975) );
  INV_X1 U3376 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U3377 ( .A1(n3415), .A2(REG2_REG_27__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U3378 ( .A1(n2353), .A2(REG0_REG_27__SCAN_IN), .ZN(n2610) );
  OAI211_X1 U3379 ( .C1(n2612), .C2(n3418), .A(n2611), .B(n2610), .ZN(n2613)
         );
  INV_X1 U3380 ( .A(n2613), .ZN(n2614) );
  NAND2_X1 U3381 ( .A1(n2308), .A2(DATAI_27_), .ZN(n4204) );
  NAND2_X1 U3382 ( .A1(n3993), .A2(n4204), .ZN(n2616) );
  NAND2_X1 U3383 ( .A1(n3973), .A2(n2616), .ZN(n2618) );
  NAND2_X1 U3384 ( .A1(n3846), .A2(n3974), .ZN(n2617) );
  NAND2_X1 U3385 ( .A1(n2618), .A2(n2617), .ZN(n2729) );
  INV_X1 U3386 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U3387 ( .A1(n2619), .A2(n3690), .ZN(n2620) );
  NAND2_X1 U3388 ( .A1(n3695), .A2(n2633), .ZN(n2626) );
  INV_X1 U3389 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3390 ( .A1(n3415), .A2(REG2_REG_28__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U3391 ( .A1(n2353), .A2(REG0_REG_28__SCAN_IN), .ZN(n2621) );
  OAI211_X1 U3392 ( .C1(n2623), .C2(n3418), .A(n2622), .B(n2621), .ZN(n2624)
         );
  INV_X1 U3393 ( .A(n2624), .ZN(n2625) );
  INV_X1 U3394 ( .A(DATAI_28_), .ZN(n2627) );
  NOR2_X1 U3395 ( .A1(n3419), .A2(n2627), .ZN(n2717) );
  NAND2_X1 U3396 ( .A1(n3684), .A2(n2717), .ZN(n3424) );
  INV_X1 U3397 ( .A(n2717), .ZN(n3691) );
  NAND2_X1 U3398 ( .A1(n4207), .A2(n3691), .ZN(n3421) );
  NAND2_X1 U3399 ( .A1(n3424), .A2(n3421), .ZN(n2731) );
  NOR2_X1 U3400 ( .A1(n3684), .A2(n3691), .ZN(n2628) );
  NAND2_X1 U3401 ( .A1(n2308), .A2(DATAI_29_), .ZN(n3968) );
  INV_X1 U3402 ( .A(n2629), .ZN(n3963) );
  NAND2_X1 U3403 ( .A1(n3415), .A2(REG2_REG_29__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3404 ( .A1(n2353), .A2(REG0_REG_29__SCAN_IN), .ZN(n2630) );
  OAI211_X1 U3405 ( .C1(n2715), .C2(n3418), .A(n2631), .B(n2630), .ZN(n2632)
         );
  AOI21_X1 U3406 ( .B1(n3963), .B2(n2633), .A(n2632), .ZN(n3692) );
  XOR2_X1 U3407 ( .A(n3968), .B(n3692), .Z(n3496) );
  INV_X1 U3408 ( .A(n2642), .ZN(n2635) );
  NAND2_X1 U3409 ( .A1(n2688), .A2(IR_REG_31__SCAN_IN), .ZN(n2636) );
  INV_X1 U3410 ( .A(IR_REG_19__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U3411 ( .A1(n2638), .A2(n2637), .ZN(n2639) );
  NAND2_X1 U3412 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  XNOR2_X1 U3413 ( .A(n4355), .B(n2910), .ZN(n2646) );
  NAND2_X1 U3414 ( .A1(n2646), .A2(n3952), .ZN(n4100) );
  AND2_X1 U3415 ( .A1(n2647), .A2(n4357), .ZN(n2906) );
  NAND2_X1 U3416 ( .A1(n2906), .A2(n2882), .ZN(n4497) );
  NAND2_X1 U3417 ( .A1(n2882), .A2(n3466), .ZN(n2886) );
  NAND2_X1 U3418 ( .A1(n2745), .A2(n3515), .ZN(n2992) );
  NAND2_X1 U3419 ( .A1(n3099), .A2(n2994), .ZN(n3520) );
  NAND2_X1 U3420 ( .A1(n3860), .A2(n3038), .ZN(n3517) );
  AND2_X1 U3421 ( .A1(n3520), .A2(n3517), .ZN(n3483) );
  NAND2_X1 U3422 ( .A1(n2992), .A2(n3483), .ZN(n2991) );
  INV_X1 U3423 ( .A(n3521), .ZN(n2648) );
  AND2_X1 U3424 ( .A1(n3858), .A2(n3149), .ZN(n3045) );
  NAND2_X1 U3425 ( .A1(n3137), .A2(n3084), .ZN(n3499) );
  NAND2_X1 U3426 ( .A1(n3857), .A2(n3138), .ZN(n3523) );
  NAND2_X1 U3427 ( .A1(n3066), .A2(n3523), .ZN(n2649) );
  NAND2_X1 U3428 ( .A1(n3187), .A2(n3110), .ZN(n3527) );
  INV_X1 U3429 ( .A(n2650), .ZN(n2651) );
  NAND2_X1 U3430 ( .A1(n3231), .A2(n3175), .ZN(n3533) );
  NAND2_X1 U3431 ( .A1(n3854), .A2(n3217), .ZN(n3530) );
  AND2_X1 U3432 ( .A1(n3853), .A2(n3232), .ZN(n3155) );
  NAND2_X1 U3433 ( .A1(n3259), .A2(n3226), .ZN(n3534) );
  NAND2_X1 U3434 ( .A1(n3852), .A2(n3265), .ZN(n3498) );
  NAND2_X1 U3435 ( .A1(n3244), .A2(n3498), .ZN(n2652) );
  NAND2_X1 U3436 ( .A1(n3316), .A2(n3252), .ZN(n3503) );
  NAND2_X1 U3437 ( .A1(n3850), .A2(n3377), .ZN(n3335) );
  NAND2_X1 U3438 ( .A1(n3849), .A2(n3793), .ZN(n2653) );
  NAND2_X1 U3439 ( .A1(n3335), .A2(n2653), .ZN(n3538) );
  INV_X1 U3440 ( .A(n3286), .ZN(n3541) );
  NOR2_X1 U3441 ( .A1(n3538), .A2(n3541), .ZN(n2654) );
  NAND2_X1 U3442 ( .A1(n3792), .A2(n3281), .ZN(n3337) );
  NAND2_X1 U3443 ( .A1(n3284), .A2(n3337), .ZN(n2657) );
  INV_X1 U3444 ( .A(n3538), .ZN(n2656) );
  NOR2_X1 U3445 ( .A1(n3849), .A2(n3793), .ZN(n2655) );
  AOI21_X1 U3446 ( .B1(n2657), .B2(n2656), .A(n2655), .ZN(n3542) );
  NAND2_X1 U3447 ( .A1(n2658), .A2(n3430), .ZN(n3383) );
  NAND2_X1 U3448 ( .A1(n4277), .A2(n4288), .ZN(n3437) );
  NAND2_X1 U3449 ( .A1(n4184), .A2(n3836), .ZN(n3504) );
  NAND2_X1 U3450 ( .A1(n3437), .A2(n3504), .ZN(n3485) );
  AND2_X1 U3451 ( .A1(n4182), .A2(n4166), .ZN(n3432) );
  NAND2_X1 U3452 ( .A1(n4141), .A2(n4125), .ZN(n3463) );
  NAND2_X1 U3453 ( .A1(n3463), .A2(n4115), .ZN(n3431) );
  NAND2_X1 U3454 ( .A1(n4244), .A2(n4104), .ZN(n3433) );
  NAND2_X1 U3455 ( .A1(n4091), .A2(n3433), .ZN(n2662) );
  NAND2_X1 U3456 ( .A1(n4276), .A2(n4264), .ZN(n4112) );
  AND2_X1 U3457 ( .A1(n4114), .A2(n4112), .ZN(n2659) );
  OR2_X1 U34580 ( .A1(n4141), .A2(n4125), .ZN(n3464) );
  OAI21_X1 U34590 ( .B1(n3431), .B2(n2659), .A(n3464), .ZN(n4090) );
  NOR2_X1 U3460 ( .A1(n4244), .A2(n4104), .ZN(n2660) );
  OR2_X1 U3461 ( .A1(n4090), .A2(n2660), .ZN(n2661) );
  NAND2_X1 U3462 ( .A1(n2661), .A2(n3433), .ZN(n3549) );
  NAND2_X1 U3463 ( .A1(n4096), .A2(n4242), .ZN(n3456) );
  AND2_X1 U3464 ( .A1(n4042), .A2(n3456), .ZN(n3550) );
  INV_X1 U3465 ( .A(n3550), .ZN(n2665) );
  INV_X1 U3466 ( .A(n3647), .ZN(n4049) );
  NAND2_X1 U34670 ( .A1(n4224), .A2(n4049), .ZN(n3460) );
  NAND2_X1 U3468 ( .A1(n3460), .A2(n2663), .ZN(n3497) );
  NOR2_X1 U34690 ( .A1(n4096), .A2(n4242), .ZN(n4039) );
  AND2_X1 U3470 ( .A1(n4039), .A2(n4042), .ZN(n2664) );
  NOR2_X1 U34710 ( .A1(n3497), .A2(n2664), .ZN(n3441) );
  INV_X1 U3472 ( .A(n3998), .ZN(n2667) );
  NAND2_X1 U34730 ( .A1(n4218), .A2(n2667), .ZN(n2668) );
  INV_X1 U3474 ( .A(n4029), .ZN(n4227) );
  NAND2_X1 U34750 ( .A1(n4227), .A2(n4214), .ZN(n3987) );
  NAND2_X1 U3476 ( .A1(n2668), .A2(n3987), .ZN(n3552) );
  INV_X1 U34770 ( .A(n3552), .ZN(n2669) );
  NAND2_X1 U3478 ( .A1(n4029), .A2(n4016), .ZN(n3454) );
  NAND2_X1 U34790 ( .A1(n4215), .A2(n4033), .ZN(n4004) );
  NAND2_X1 U3480 ( .A1(n3454), .A2(n4004), .ZN(n3988) );
  INV_X1 U34810 ( .A(n4218), .ZN(n4012) );
  AND2_X1 U3482 ( .A1(n4012), .A2(n3998), .ZN(n3422) );
  AOI21_X1 U34830 ( .B1(n2669), .B2(n3988), .A(n3422), .ZN(n3558) );
  XNOR2_X1 U3484 ( .A(n3846), .B(n4204), .ZN(n3980) );
  NAND2_X1 U34850 ( .A1(n3993), .A2(n3974), .ZN(n3423) );
  INV_X1 U3486 ( .A(n3424), .ZN(n2670) );
  XNOR2_X1 U34870 ( .A(n2671), .B(n3496), .ZN(n2682) );
  NAND2_X1 U3488 ( .A1(n4355), .A2(n4357), .ZN(n2672) );
  INV_X1 U34890 ( .A(n2647), .ZN(n2768) );
  NAND2_X1 U3490 ( .A1(n4356), .A2(n2768), .ZN(n3451) );
  NOR2_X1 U34910 ( .A1(n2674), .A2(n2673), .ZN(n2857) );
  NOR2_X1 U3492 ( .A1(n2306), .A2(n2775), .ZN(n2675) );
  MUX2_X1 U34930 ( .A(n2775), .B(n2675), .S(IR_REG_28__SCAN_IN), .Z(n2678) );
  INV_X1 U3494 ( .A(n2676), .ZN(n2677) );
  NAND2_X1 U34950 ( .A1(n4355), .A2(n4356), .ZN(n2887) );
  INV_X1 U3496 ( .A(n2887), .ZN(n2788) );
  NAND2_X1 U34970 ( .A1(n2897), .A2(n2788), .ZN(n4275) );
  AOI21_X1 U3498 ( .B1(B_REG_SCAN_IN), .B2(n2857), .A(n4275), .ZN(n3957) );
  INV_X1 U34990 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3500 ( .A1(n3415), .A2(REG2_REG_30__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U35010 ( .A1(n2353), .A2(REG0_REG_30__SCAN_IN), .ZN(n2679) );
  OAI211_X1 U3502 ( .C1(n3418), .C2(n2681), .A(n2680), .B(n2679), .ZN(n3844)
         );
  NOR2_X2 U35030 ( .A1(n2897), .A2(n2887), .ZN(n4243) );
  NAND2_X1 U3504 ( .A1(n4207), .A2(n4243), .ZN(n2683) );
  NAND2_X1 U35050 ( .A1(n2684), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  MUX2_X1 U35060 ( .A(IR_REG_31__SCAN_IN), .B(n2685), .S(IR_REG_25__SCAN_IN), 
        .Z(n2687) );
  NAND2_X1 U35070 ( .A1(n2687), .A2(n2686), .ZN(n2765) );
  NAND2_X1 U35080 ( .A1(n2765), .A2(B_REG_SCAN_IN), .ZN(n2691) );
  NAND2_X1 U35090 ( .A1(n2697), .A2(n2698), .ZN(n2689) );
  MUX2_X1 U35100 ( .A(n2691), .B(B_REG_SCAN_IN), .S(n2696), .Z(n2694) );
  NAND2_X1 U35110 ( .A1(n2686), .A2(IR_REG_31__SCAN_IN), .ZN(n2692) );
  MUX2_X1 U35120 ( .A(IR_REG_31__SCAN_IN), .B(n2692), .S(IR_REG_26__SCAN_IN), 
        .Z(n2693) );
  NAND2_X1 U35130 ( .A1(n2783), .A2(n2765), .ZN(n2780) );
  NAND2_X1 U35140 ( .A1(n2879), .A2(n2780), .ZN(n2712) );
  XNOR2_X1 U35150 ( .A(n2697), .B(n2698), .ZN(n2787) );
  OR2_X1 U35160 ( .A1(n4497), .A2(n4356), .ZN(n2754) );
  AND2_X1 U35170 ( .A1(n2647), .A2(n3952), .ZN(n2885) );
  OR2_X1 U35180 ( .A1(n2887), .A2(n2885), .ZN(n2890) );
  NAND2_X1 U35190 ( .A1(n2754), .A2(n2890), .ZN(n2699) );
  NOR2_X1 U35200 ( .A1(n2895), .A2(n2699), .ZN(n2711) );
  NOR4_X1 U35210 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2703) );
  NOR4_X1 U35220 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2702) );
  NOR4_X1 U35230 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2701) );
  NOR4_X1 U35240 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2700) );
  NAND4_X1 U35250 ( .A1(n2703), .A2(n2702), .A3(n2701), .A4(n2700), .ZN(n2709)
         );
  NOR2_X1 U35260 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2707) );
  NOR4_X1 U35270 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2706) );
  NOR4_X1 U35280 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2705) );
  NOR4_X1 U35290 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2704) );
  NAND4_X1 U35300 ( .A1(n2707), .A2(n2706), .A3(n2705), .A4(n2704), .ZN(n2708)
         );
  NOR2_X1 U35310 ( .A1(n2709), .A2(n2708), .ZN(n2710) );
  NAND3_X1 U35320 ( .A1(n2712), .A2(n2711), .A3(n2750), .ZN(n2724) );
  NAND2_X1 U35330 ( .A1(n2784), .A2(n2783), .ZN(n2713) );
  MUX2_X1 U35340 ( .A(n2715), .B(n2725), .S(n4518), .Z(n2723) );
  NAND2_X1 U35350 ( .A1(n2915), .A2(n2903), .ZN(n2954) );
  NOR2_X1 U35360 ( .A1(n2954), .A2(n2961), .ZN(n2989) );
  NAND2_X1 U35370 ( .A1(n2989), .A2(n3038), .ZN(n3027) );
  NOR2_X2 U35380 ( .A1(n3051), .A2(n3084), .ZN(n3060) );
  NAND2_X1 U35390 ( .A1(n3060), .A2(n3138), .ZN(n3075) );
  OR2_X2 U35400 ( .A1(n4145), .A2(n2716), .ZN(n4124) );
  NOR2_X4 U35410 ( .A1(n4124), .A2(n4094), .ZN(n4102) );
  INV_X1 U35420 ( .A(n4033), .ZN(n4223) );
  INV_X1 U35430 ( .A(n2718), .ZN(n2736) );
  INV_X1 U35440 ( .A(n3968), .ZN(n3426) );
  NAND2_X1 U35450 ( .A1(n2736), .A2(n3426), .ZN(n2719) );
  NAND2_X1 U35460 ( .A1(n4199), .A2(n2719), .ZN(n3966) );
  INV_X1 U35470 ( .A(n2886), .ZN(n2904) );
  NAND2_X1 U35480 ( .A1(n2723), .A2(n2722), .ZN(U3547) );
  INV_X1 U35490 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2726) );
  XNOR2_X1 U35500 ( .A(n2729), .B(n2731), .ZN(n3597) );
  INV_X1 U35510 ( .A(n4506), .ZN(n4262) );
  INV_X1 U35520 ( .A(n3692), .ZN(n3845) );
  OAI22_X1 U35530 ( .A1(n3993), .A2(n4293), .B1(n4274), .B2(n3691), .ZN(n2730)
         );
  AOI21_X1 U35540 ( .B1(n4289), .B2(n3845), .A(n2730), .ZN(n2734) );
  INV_X1 U35550 ( .A(n2731), .ZN(n3453) );
  XNOR2_X1 U35560 ( .A(n2732), .B(n3453), .ZN(n2733) );
  NAND2_X1 U35570 ( .A1(n2733), .A2(n4171), .ZN(n3592) );
  OAI211_X1 U35580 ( .C1(n3597), .C2(n4262), .A(n2734), .B(n3592), .ZN(n2738)
         );
  MUX2_X1 U35590 ( .A(REG1_REG_28__SCAN_IN), .B(n2738), .S(n4518), .Z(n2735)
         );
  INV_X1 U35600 ( .A(n2735), .ZN(n2737) );
  OAI21_X1 U35610 ( .B1(n2050), .B2(n3691), .A(n2736), .ZN(n3589) );
  NAND2_X1 U35620 ( .A1(n2737), .A2(n2283), .ZN(U3546) );
  MUX2_X1 U35630 ( .A(REG0_REG_28__SCAN_IN), .B(n2738), .S(n4513), .Z(n2739)
         );
  INV_X1 U35640 ( .A(n2739), .ZN(n2740) );
  NAND2_X1 U35650 ( .A1(n2740), .A2(n2285), .ZN(U3514) );
  INV_X1 U35660 ( .A(n4484), .ZN(n2741) );
  INV_X2 U35670 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U35680 ( .A1(n2742), .A2(n3476), .ZN(n2743) );
  NAND2_X1 U35690 ( .A1(n2744), .A2(n2743), .ZN(n2965) );
  INV_X1 U35700 ( .A(n4100), .ZN(n3171) );
  NAND2_X1 U35710 ( .A1(n2965), .A2(n3171), .ZN(n2749) );
  OAI21_X1 U35720 ( .B1(n3476), .B2(n2746), .A(n2745), .ZN(n2747) );
  NAND2_X1 U35730 ( .A1(n2747), .A2(n4171), .ZN(n2748) );
  NAND2_X1 U35740 ( .A1(n2749), .A2(n2748), .ZN(n2963) );
  INV_X1 U35750 ( .A(n2890), .ZN(n2751) );
  NOR2_X1 U35760 ( .A1(n2895), .A2(n2751), .ZN(n2753) );
  NAND4_X1 U35770 ( .A1(n2880), .A2(n2753), .A3(n2752), .A4(n2879), .ZN(n2755)
         );
  MUX2_X1 U35780 ( .A(n2963), .B(REG2_REG_2__SCAN_IN), .S(n4482), .Z(n2763) );
  INV_X1 U35790 ( .A(n2910), .ZN(n2849) );
  NAND2_X1 U35800 ( .A1(n2849), .A2(n4357), .ZN(n3033) );
  INV_X1 U35810 ( .A(n3033), .ZN(n2756) );
  AND2_X1 U3582 ( .A1(n4473), .A2(n2756), .ZN(n4477) );
  NOR2_X1 U3583 ( .A1(n4470), .A2(n3874), .ZN(n2757) );
  AOI21_X1 U3584 ( .B1(n2965), .B2(n4477), .A(n2757), .ZN(n2761) );
  NAND2_X1 U3585 ( .A1(n4473), .A2(n4287), .ZN(n4190) );
  INV_X1 U3586 ( .A(n4190), .ZN(n3325) );
  AOI22_X1 U3587 ( .A1(n3325), .A2(n2961), .B1(n4183), .B2(n3860), .ZN(n2760)
         );
  NAND2_X1 U3588 ( .A1(n4473), .A2(n3952), .ZN(n4148) );
  INV_X1 U3589 ( .A(n4146), .ZN(n4283) );
  XNOR2_X1 U3590 ( .A(n2954), .B(n2931), .ZN(n2967) );
  NAND2_X1 U3591 ( .A1(n4476), .A2(n2967), .ZN(n2759) );
  NAND2_X1 U3592 ( .A1(n4185), .A2(n3862), .ZN(n2758) );
  NAND4_X1 U3593 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n2762)
         );
  OR2_X1 U3594 ( .A1(n2763), .A2(n2762), .ZN(U3288) );
  NAND2_X1 U3595 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2764) );
  OAI21_X1 U3596 ( .B1(n2765), .B2(U3149), .A(n2764), .ZN(U3327) );
  INV_X1 U3597 ( .A(DATAI_26_), .ZN(n4610) );
  NAND2_X1 U3598 ( .A1(n2766), .A2(STATE_REG_SCAN_IN), .ZN(n2767) );
  OAI21_X1 U3599 ( .B1(STATE_REG_SCAN_IN), .B2(n4610), .A(n2767), .ZN(U3326)
         );
  INV_X1 U3600 ( .A(DATAI_20_), .ZN(n4680) );
  NAND2_X1 U3601 ( .A1(n2768), .A2(STATE_REG_SCAN_IN), .ZN(n2769) );
  OAI21_X1 U3602 ( .B1(STATE_REG_SCAN_IN), .B2(n4680), .A(n2769), .ZN(U3332)
         );
  INV_X1 U3603 ( .A(DATAI_24_), .ZN(n4542) );
  NAND2_X1 U3604 ( .A1(n2696), .A2(STATE_REG_SCAN_IN), .ZN(n2770) );
  OAI21_X1 U3605 ( .B1(STATE_REG_SCAN_IN), .B2(n4542), .A(n2770), .ZN(U3328)
         );
  INV_X1 U3606 ( .A(DATAI_27_), .ZN(n4681) );
  NAND2_X1 U3607 ( .A1(n2857), .A2(STATE_REG_SCAN_IN), .ZN(n2771) );
  OAI21_X1 U3608 ( .B1(STATE_REG_SCAN_IN), .B2(n4681), .A(n2771), .ZN(U3325)
         );
  INV_X1 U3609 ( .A(DATAI_29_), .ZN(n4643) );
  NAND2_X1 U3610 ( .A1(n2772), .A2(STATE_REG_SCAN_IN), .ZN(n2773) );
  OAI21_X1 U3611 ( .B1(STATE_REG_SCAN_IN), .B2(n4643), .A(n2773), .ZN(U3323)
         );
  INV_X1 U3612 ( .A(n2897), .ZN(n2920) );
  NAND2_X1 U3613 ( .A1(n2920), .A2(STATE_REG_SCAN_IN), .ZN(n2774) );
  OAI21_X1 U3614 ( .B1(STATE_REG_SCAN_IN), .B2(n2627), .A(n2774), .ZN(U3324)
         );
  INV_X1 U3615 ( .A(DATAI_31_), .ZN(n4530) );
  OR4_X1 U3616 ( .A1(n2776), .A2(IR_REG_30__SCAN_IN), .A3(n2775), .A4(U3149), 
        .ZN(n2777) );
  OAI21_X1 U3617 ( .B1(STATE_REG_SCAN_IN), .B2(n4530), .A(n2777), .ZN(U3321)
         );
  INV_X1 U3618 ( .A(n2895), .ZN(n2778) );
  INV_X1 U3619 ( .A(D_REG_1__SCAN_IN), .ZN(n2782) );
  INV_X1 U3620 ( .A(n2780), .ZN(n2781) );
  AOI22_X1 U3621 ( .A1(n4483), .A2(n2782), .B1(n2781), .B2(n4484), .ZN(U3459)
         );
  INV_X1 U3622 ( .A(D_REG_0__SCAN_IN), .ZN(n2786) );
  AND2_X1 U3623 ( .A1(n4484), .A2(n2783), .ZN(n2785) );
  AOI22_X1 U3624 ( .A1(n4483), .A2(n2786), .B1(n2785), .B2(n2784), .ZN(U3458)
         );
  OR2_X1 U3625 ( .A1(n2787), .A2(U3149), .ZN(n3577) );
  NAND2_X1 U3626 ( .A1(n2895), .A2(n3577), .ZN(n2791) );
  AOI21_X1 U3627 ( .B1(n2788), .B2(n2787), .A(n3419), .ZN(n2790) );
  INV_X1 U3628 ( .A(n2790), .ZN(n2789) );
  AND2_X1 U3629 ( .A1(n2791), .A2(n2790), .ZN(n2809) );
  INV_X1 U3630 ( .A(n2809), .ZN(n2795) );
  INV_X1 U3631 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2792) );
  AOI21_X1 U3632 ( .B1(n2857), .B2(n2792), .A(n2897), .ZN(n2859) );
  OAI21_X1 U3633 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2857), .A(n2859), .ZN(n2793)
         );
  MUX2_X1 U3634 ( .A(n2793), .B(n2859), .S(IR_REG_0__SCAN_IN), .Z(n2794) );
  OAI22_X1 U3635 ( .A1(n2795), .A2(n2794), .B1(STATE_REG_SCAN_IN), .B2(n2902), 
        .ZN(n2796) );
  AOI21_X1 U3636 ( .B1(n4463), .B2(ADDR_REG_0__SCAN_IN), .A(n2796), .ZN(n2798)
         );
  INV_X1 U3637 ( .A(n2857), .ZN(n2806) );
  NAND3_X1 U3638 ( .A1(n4465), .A2(IR_REG_0__SCAN_IN), .A3(n2346), .ZN(n2797)
         );
  NAND2_X1 U3639 ( .A1(n2798), .A2(n2797), .ZN(U3240) );
  INV_X1 U3640 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3879) );
  INV_X1 U3641 ( .A(n4364), .ZN(n3877) );
  MUX2_X1 U3642 ( .A(REG2_REG_2__SCAN_IN), .B(n3879), .S(n4364), .Z(n2802) );
  INV_X1 U3643 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2799) );
  AND2_X1 U3644 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2800)
         );
  NAND2_X1 U3645 ( .A1(n4365), .A2(REG2_REG_1__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U3646 ( .A1(n3881), .A2(n3880), .ZN(n2801) );
  INV_X1 U3647 ( .A(n4363), .ZN(n2816) );
  XNOR2_X1 U3648 ( .A(n2803), .B(n2865), .ZN(n2860) );
  INV_X1 U3649 ( .A(n2860), .ZN(n2805) );
  INV_X1 U3650 ( .A(n2803), .ZN(n2804) );
  MUX2_X1 U3651 ( .A(REG2_REG_5__SCAN_IN), .B(n2387), .S(n2829), .Z(n2807) );
  NOR2_X1 U3652 ( .A1(n2897), .A2(n2806), .ZN(n3573) );
  AOI211_X1 U3653 ( .C1(n2808), .C2(n2807), .A(n2825), .B(n4459), .ZN(n2812)
         );
  NOR2_X1 U3654 ( .A1(STATE_REG_SCAN_IN), .A2(n2383), .ZN(n3151) );
  AOI21_X1 U3655 ( .B1(n4463), .B2(ADDR_REG_5__SCAN_IN), .A(n3151), .ZN(n2810)
         );
  OAI21_X1 U3656 ( .B1(n4469), .B2(n2829), .A(n2810), .ZN(n2811) );
  NOR2_X1 U3657 ( .A1(n2812), .A2(n2811), .ZN(n2824) );
  XNOR2_X1 U3658 ( .A(n2829), .B(REG1_REG_5__SCAN_IN), .ZN(n2822) );
  XNOR2_X1 U3659 ( .A(n4364), .B(n2813), .ZN(n3887) );
  XNOR2_X1 U3660 ( .A(n4365), .B(n2338), .ZN(n3867) );
  AND2_X1 U3661 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U3662 ( .A1(n3867), .A2(n3866), .ZN(n3865) );
  NAND2_X1 U3663 ( .A1(n4365), .A2(REG1_REG_1__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U3664 ( .A1(n3865), .A2(n2814), .ZN(n3886) );
  NAND2_X1 U3665 ( .A1(n3887), .A2(n3886), .ZN(n3885) );
  NAND2_X1 U3666 ( .A1(n4364), .A2(REG1_REG_2__SCAN_IN), .ZN(n2815) );
  NAND2_X1 U3667 ( .A1(n3885), .A2(n2815), .ZN(n2817) );
  XNOR2_X1 U3668 ( .A(n2817), .B(n2816), .ZN(n3894) );
  NAND2_X1 U3669 ( .A1(n3894), .A2(REG1_REG_3__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U3670 ( .A1(n2817), .A2(n4363), .ZN(n2818) );
  NAND2_X1 U3671 ( .A1(n3893), .A2(n2818), .ZN(n2819) );
  INV_X1 U3672 ( .A(n2819), .ZN(n2820) );
  XNOR2_X1 U3673 ( .A(n2819), .B(n2865), .ZN(n2862) );
  NAND2_X1 U3674 ( .A1(n2862), .A2(REG1_REG_4__SCAN_IN), .ZN(n2861) );
  OAI21_X1 U3675 ( .B1(n2820), .B2(n2865), .A(n2861), .ZN(n2821) );
  NAND2_X1 U3676 ( .A1(n2821), .A2(n2822), .ZN(n2827) );
  OAI211_X1 U3677 ( .C1(n2822), .C2(n2821), .A(n4465), .B(n2827), .ZN(n2823)
         );
  NAND2_X1 U3678 ( .A1(n2824), .A2(n2823), .ZN(U3245) );
  INV_X1 U3679 ( .A(n2829), .ZN(n4361) );
  XNOR2_X1 U3680 ( .A(n2840), .B(REG2_REG_6__SCAN_IN), .ZN(n2835) );
  INV_X1 U3681 ( .A(n4469), .ZN(n3892) );
  NAND2_X1 U3682 ( .A1(n4463), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U3683 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3684 ( .A1(n2826), .A2(n3136), .ZN(n2833) );
  OAI21_X1 U3685 ( .B1(n2829), .B2(n2828), .A(n2827), .ZN(n2837) );
  XNOR2_X1 U3686 ( .A(n2837), .B(n4360), .ZN(n2831) );
  INV_X1 U3687 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3118) );
  NOR2_X1 U3688 ( .A1(n2831), .A2(n3118), .ZN(n2836) );
  INV_X1 U3689 ( .A(n4465), .ZN(n2830) );
  AOI211_X1 U3690 ( .C1(n2831), .C2(n3118), .A(n2836), .B(n2830), .ZN(n2832)
         );
  AOI211_X1 U3691 ( .C1(n3892), .C2(n4360), .A(n2833), .B(n2832), .ZN(n2834)
         );
  OAI21_X1 U3692 ( .B1(n2835), .B2(n4459), .A(n2834), .ZN(U3246) );
  NOR2_X1 U3693 ( .A1(n4463), .A2(n3856), .ZN(U3148) );
  MUX2_X1 U3694 ( .A(REG1_REG_7__SCAN_IN), .B(n2416), .S(n4359), .Z(n2838) );
  XNOR2_X1 U3695 ( .A(n2871), .B(n2838), .ZN(n2845) );
  INV_X1 U3696 ( .A(n4359), .ZN(n2869) );
  INV_X1 U3697 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4660) );
  NOR2_X1 U3698 ( .A1(STATE_REG_SCAN_IN), .A2(n4660), .ZN(n3190) );
  AOI21_X1 U3699 ( .B1(n4463), .B2(ADDR_REG_7__SCAN_IN), .A(n3190), .ZN(n2839)
         );
  OAI21_X1 U3700 ( .B1(n4469), .B2(n2869), .A(n2839), .ZN(n2844) );
  MUX2_X1 U3701 ( .A(n2414), .B(REG2_REG_7__SCAN_IN), .S(n4359), .Z(n2841) );
  NOR2_X1 U3702 ( .A1(n2842), .A2(n2841), .ZN(n2873) );
  AOI211_X1 U3703 ( .C1(n2842), .C2(n2841), .A(n4459), .B(n2873), .ZN(n2843)
         );
  AOI211_X1 U3704 ( .C1(n4465), .C2(n2845), .A(n2844), .B(n2843), .ZN(n2846)
         );
  INV_X1 U3705 ( .A(n2846), .ZN(U3247) );
  OR2_X4 U3706 ( .A1(n3681), .A2(n4146), .ZN(n3683) );
  INV_X1 U3707 ( .A(n3683), .ZN(n2848) );
  NAND2_X1 U3708 ( .A1(n2851), .A2(n2850), .ZN(n2855) );
  NAND2_X1 U3709 ( .A1(n2979), .A2(REG1_REG_0__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U3710 ( .A1(n2912), .A2(n2852), .ZN(n2854) );
  INV_X1 U3711 ( .A(n2913), .ZN(n2853) );
  OAI21_X1 U3712 ( .B1(n2855), .B2(n2854), .A(n2853), .ZN(n2899) );
  NAND2_X1 U3713 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3868) );
  AOI21_X1 U3714 ( .B1(n2857), .B2(n3868), .A(n2897), .ZN(n2856) );
  OAI21_X1 U3715 ( .B1(n2899), .B2(n2857), .A(n2856), .ZN(n2858) );
  OAI211_X1 U3716 ( .C1(IR_REG_0__SCAN_IN), .C2(n2859), .A(n2858), .B(U4043), 
        .ZN(n3891) );
  XNOR2_X1 U3717 ( .A(n2860), .B(REG2_REG_4__SCAN_IN), .ZN(n2867) );
  OAI211_X1 U3718 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2862), .A(n4465), .B(n2861), 
        .ZN(n2864) );
  AND2_X1 U3719 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3102) );
  AOI21_X1 U3720 ( .B1(n4463), .B2(ADDR_REG_4__SCAN_IN), .A(n3102), .ZN(n2863)
         );
  OAI211_X1 U3721 ( .C1(n4469), .C2(n2865), .A(n2864), .B(n2863), .ZN(n2866)
         );
  AOI21_X1 U3722 ( .B1(n4411), .B2(n2867), .A(n2866), .ZN(n2868) );
  NAND2_X1 U3723 ( .A1(n3891), .A2(n2868), .ZN(U3244) );
  NOR2_X1 U3724 ( .A1(n4359), .A2(REG1_REG_7__SCAN_IN), .ZN(n2870) );
  XOR2_X1 U3725 ( .A(REG1_REG_8__SCAN_IN), .B(n3924), .Z(n2872) );
  NAND2_X1 U3726 ( .A1(n2872), .A2(n4465), .ZN(n2878) );
  AOI21_X1 U3727 ( .B1(n4359), .B2(REG2_REG_7__SCAN_IN), .A(n2873), .ZN(n3904)
         );
  XNOR2_X1 U3728 ( .A(REG2_REG_8__SCAN_IN), .B(n3905), .ZN(n2874) );
  NAND2_X1 U3729 ( .A1(n4411), .A2(n2874), .ZN(n2875) );
  NAND2_X1 U3730 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3215) );
  NAND2_X1 U3731 ( .A1(n2875), .A2(n3215), .ZN(n2876) );
  AOI21_X1 U3732 ( .B1(n4463), .B2(ADDR_REG_8__SCAN_IN), .A(n2876), .ZN(n2877)
         );
  OAI211_X1 U3733 ( .C1(n4469), .C2(n4358), .A(n2878), .B(n2877), .ZN(U3248)
         );
  NAND3_X1 U3734 ( .A1(n2881), .A2(n2880), .A3(n2879), .ZN(n2922) );
  INV_X1 U3735 ( .A(n2911), .ZN(n2883) );
  NAND2_X1 U3736 ( .A1(n4484), .A2(n2883), .ZN(n2884) );
  NAND2_X1 U3737 ( .A1(n2922), .A2(n3574), .ZN(n2981) );
  INV_X1 U3738 ( .A(n2981), .ZN(n2892) );
  OR2_X1 U3739 ( .A1(n2886), .A2(n2885), .ZN(n2888) );
  NAND2_X1 U3740 ( .A1(n2888), .A2(n2887), .ZN(n2894) );
  NAND2_X1 U3741 ( .A1(n2894), .A2(n4274), .ZN(n2889) );
  NAND2_X1 U3742 ( .A1(n2922), .A2(n2889), .ZN(n2891) );
  NAND2_X1 U3743 ( .A1(n2891), .A2(n2890), .ZN(n2980) );
  NOR3_X1 U3744 ( .A1(n2892), .A2(n2980), .A3(n2895), .ZN(n2941) );
  NOR3_X1 U3745 ( .A1(n2922), .A2(n2895), .A3(n4274), .ZN(n2893) );
  OR2_X1 U3746 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  NAND2_X1 U3747 ( .A1(n3574), .A2(n2897), .ZN(n2898) );
  OAI22_X1 U3748 ( .A1(n2899), .A2(n3827), .B1(n2916), .B2(n3822), .ZN(n2900)
         );
  AOI21_X1 U3749 ( .B1(n3098), .B2(n2952), .A(n2900), .ZN(n2901) );
  OAI21_X1 U3750 ( .B1(n2941), .B2(n2902), .A(n2901), .ZN(U3229) );
  NAND2_X1 U3751 ( .A1(n3864), .A2(n2903), .ZN(n3512) );
  AND2_X1 U3752 ( .A1(n3510), .A2(n3512), .ZN(n4498) );
  INV_X1 U3753 ( .A(n4477), .ZN(n3587) );
  NAND2_X1 U3754 ( .A1(n2952), .A2(n2904), .ZN(n4495) );
  AOI21_X1 U3755 ( .B1(n4122), .B2(n4100), .A(n4498), .ZN(n2905) );
  AOI21_X1 U3756 ( .B1(n4289), .B2(n3862), .A(n2905), .ZN(n4496) );
  OAI21_X1 U3757 ( .B1(n2906), .B2(n4495), .A(n4496), .ZN(n2907) );
  AOI22_X1 U3758 ( .A1(n2907), .A2(n4473), .B1(REG3_REG_0__SCAN_IN), .B2(n4186), .ZN(n2909) );
  NAND2_X1 U3759 ( .A1(n4087), .A2(REG2_REG_0__SCAN_IN), .ZN(n2908) );
  OAI211_X1 U3760 ( .C1(n4498), .C2(n3587), .A(n2909), .B(n2908), .ZN(U3290)
         );
  INV_X2 U3761 ( .A(n3666), .ZN(n2972) );
  OAI22_X1 U3762 ( .A1(n2916), .A2(n3683), .B1(n3656), .B2(n2915), .ZN(n2927)
         );
  AOI211_X1 U3763 ( .C1(n2918), .C2(n2917), .A(n3827), .B(n2929), .ZN(n2919)
         );
  INV_X1 U3764 ( .A(n2919), .ZN(n2925) );
  NAND2_X1 U3765 ( .A1(n3574), .A2(n2920), .ZN(n2921) );
  NOR2_X1 U3766 ( .A1(n2922), .A2(n2921), .ZN(n3700) );
  INV_X2 U3767 ( .A(n3700), .ZN(n3835) );
  OAI22_X1 U3768 ( .A1(n2946), .A2(n3835), .B1(n3822), .B2(n2932), .ZN(n2923)
         );
  AOI21_X1 U3769 ( .B1(n3098), .B2(n3008), .A(n2923), .ZN(n2924) );
  OAI211_X1 U3770 ( .C1(n2941), .C2(n3004), .A(n2925), .B(n2924), .ZN(U3219)
         );
  AND2_X1 U3771 ( .A1(n2927), .A2(n2926), .ZN(n2928) );
  OAI22_X1 U3772 ( .A1(n2932), .A2(n3683), .B1(n3645), .B2(n2931), .ZN(n2975)
         );
  XNOR2_X1 U3773 ( .A(n2974), .B(n2933), .ZN(n2934) );
  NOR2_X1 U3774 ( .A1(n2935), .A2(n2934), .ZN(n2937) );
  OAI21_X1 U3775 ( .B1(n2937), .B2(n2936), .A(n3832), .ZN(n2940) );
  OAI22_X1 U3776 ( .A1(n3099), .A2(n3822), .B1(n3835), .B2(n2916), .ZN(n2938)
         );
  AOI21_X1 U3777 ( .B1(n3098), .B2(n2961), .A(n2938), .ZN(n2939) );
  OAI211_X1 U3778 ( .C1(n2941), .C2(n3874), .A(n2940), .B(n2939), .ZN(U3234)
         );
  INV_X1 U3779 ( .A(n4497), .ZN(n4504) );
  OR2_X1 U3780 ( .A1(n2942), .A2(n3475), .ZN(n2943) );
  NAND2_X1 U3781 ( .A1(n2944), .A2(n2943), .ZN(n2949) );
  INV_X1 U3782 ( .A(n2949), .ZN(n3002) );
  AOI22_X1 U3783 ( .A1(n3861), .A2(n4289), .B1(n4287), .B2(n3008), .ZN(n2945)
         );
  OAI21_X1 U3784 ( .B1(n2946), .B2(n4293), .A(n2945), .ZN(n2951) );
  INV_X1 U3785 ( .A(n2947), .ZN(n2948) );
  AOI21_X1 U3786 ( .B1(n3475), .B2(n3510), .A(n2948), .ZN(n2950) );
  OAI22_X1 U3787 ( .A1(n2950), .A2(n4122), .B1(n4100), .B2(n2949), .ZN(n3005)
         );
  AOI211_X1 U3788 ( .C1(n4504), .C2(n3002), .A(n2951), .B(n3005), .ZN(n2960)
         );
  NAND2_X1 U3789 ( .A1(n3008), .A2(n2952), .ZN(n2953) );
  NAND2_X1 U3790 ( .A1(n2954), .A2(n2953), .ZN(n3011) );
  INV_X1 U3791 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2955) );
  OAI22_X1 U3792 ( .A1(n4347), .A2(n3011), .B1(n4513), .B2(n2955), .ZN(n2956)
         );
  INV_X1 U3793 ( .A(n2956), .ZN(n2957) );
  OAI21_X1 U3794 ( .B1(n2960), .B2(n4511), .A(n2957), .ZN(U3469) );
  OAI22_X1 U3795 ( .A1(n4299), .A2(n3011), .B1(n4518), .B2(n2338), .ZN(n2958)
         );
  INV_X1 U3796 ( .A(n2958), .ZN(n2959) );
  OAI21_X1 U3797 ( .B1(n2960), .B2(n4516), .A(n2959), .ZN(U3519) );
  AOI22_X1 U3798 ( .A1(n3860), .A2(n4289), .B1(n2961), .B2(n4287), .ZN(n2962)
         );
  OAI21_X1 U3799 ( .B1(n2916), .B2(n4293), .A(n2962), .ZN(n2964) );
  AOI211_X1 U3800 ( .C1(n4504), .C2(n2965), .A(n2964), .B(n2963), .ZN(n2969)
         );
  AOI22_X1 U3801 ( .A1(n2727), .A2(n2967), .B1(REG0_REG_2__SCAN_IN), .B2(n4511), .ZN(n2966) );
  OAI21_X1 U3802 ( .B1(n2969), .B2(n4511), .A(n2966), .ZN(U3471) );
  AOI22_X1 U3803 ( .A1(n2720), .A2(n2967), .B1(REG1_REG_2__SCAN_IN), .B2(n4516), .ZN(n2968) );
  OAI21_X1 U3804 ( .B1(n2969), .B2(n4516), .A(n2968), .ZN(U3520) );
  NAND2_X1 U3805 ( .A1(n3860), .A2(n3662), .ZN(n2971) );
  NAND2_X1 U3806 ( .A1(n3663), .A2(n2994), .ZN(n2970) );
  NAND2_X1 U3807 ( .A1(n2971), .A2(n2970), .ZN(n2973) );
  XNOR2_X1 U3808 ( .A(n2973), .B(n2972), .ZN(n3092) );
  OAI22_X1 U3809 ( .A1(n3099), .A2(n3683), .B1(n3656), .B2(n3038), .ZN(n3091)
         );
  XNOR2_X1 U3810 ( .A(n3092), .B(n3091), .ZN(n3093) );
  INV_X1 U3811 ( .A(n2974), .ZN(n2976) );
  XOR2_X1 U3812 ( .A(n3093), .B(n3094), .Z(n2988) );
  OAI22_X1 U3813 ( .A1(n2932), .A2(n3835), .B1(n3822), .B2(n3148), .ZN(n2986)
         );
  OAI21_X1 U3814 ( .B1(n2980), .B2(n2979), .A(STATE_REG_SCAN_IN), .ZN(n2983)
         );
  MUX2_X1 U3815 ( .A(U3149), .B(n3825), .S(n2984), .Z(n2985) );
  AOI211_X1 U3816 ( .C1(n2994), .C2(n3098), .A(n2986), .B(n2985), .ZN(n2987)
         );
  OAI21_X1 U3817 ( .B1(n2988), .B2(n3827), .A(n2987), .ZN(U3215) );
  OR2_X1 U3818 ( .A1(n2989), .A2(n3038), .ZN(n2990) );
  NAND2_X1 U3819 ( .A1(n2990), .A2(n3027), .ZN(n3035) );
  XNOR2_X1 U3820 ( .A(n3013), .B(n3483), .ZN(n3044) );
  OAI21_X1 U3821 ( .B1(n3483), .B2(n2992), .A(n2991), .ZN(n2993) );
  AOI22_X1 U3822 ( .A1(n2993), .A2(n4171), .B1(n4243), .B2(n3861), .ZN(n3039)
         );
  AOI22_X1 U3823 ( .A1(n3859), .A2(n4289), .B1(n4287), .B2(n2994), .ZN(n2995)
         );
  OAI211_X1 U3824 ( .C1(n4262), .C2(n3044), .A(n3039), .B(n2995), .ZN(n3000)
         );
  NAND2_X1 U3825 ( .A1(n3000), .A2(n4518), .ZN(n2997) );
  NAND2_X1 U3826 ( .A1(n4516), .A2(REG1_REG_3__SCAN_IN), .ZN(n2996) );
  OAI211_X1 U3827 ( .C1(n4299), .C2(n3035), .A(n2997), .B(n2996), .ZN(U3521)
         );
  OAI22_X1 U3828 ( .A1(n4347), .A2(n3035), .B1(n4513), .B2(n2998), .ZN(n2999)
         );
  AOI21_X1 U3829 ( .B1(n3000), .B2(n4513), .A(n2999), .ZN(n3001) );
  INV_X1 U3830 ( .A(n3001), .ZN(U3473) );
  NAND2_X1 U3831 ( .A1(n4477), .A2(n3002), .ZN(n3003) );
  OAI21_X1 U3832 ( .B1(n4470), .B2(n3004), .A(n3003), .ZN(n3007) );
  MUX2_X1 U3833 ( .A(REG2_REG_1__SCAN_IN), .B(n3005), .S(n4473), .Z(n3006) );
  AOI211_X1 U3834 ( .C1(n4185), .C2(n3864), .A(n3007), .B(n3006), .ZN(n3010)
         );
  AOI22_X1 U3835 ( .A1(n3325), .A2(n3008), .B1(n4183), .B2(n3861), .ZN(n3009)
         );
  OAI211_X1 U3836 ( .C1(n4127), .C2(n3011), .A(n3010), .B(n3009), .ZN(U3289)
         );
  NAND2_X1 U3837 ( .A1(n3013), .A2(n3012), .ZN(n3016) );
  NAND2_X1 U3838 ( .A1(n3016), .A2(n3014), .ZN(n3020) );
  NAND2_X1 U3839 ( .A1(n3016), .A2(n3015), .ZN(n3018) );
  INV_X1 U3840 ( .A(n3017), .ZN(n3477) );
  NAND2_X1 U3841 ( .A1(n3018), .A2(n3477), .ZN(n3019) );
  INV_X1 U3842 ( .A(n4505), .ZN(n3032) );
  XOR2_X1 U3843 ( .A(n3477), .B(n3021), .Z(n3026) );
  AOI22_X1 U3844 ( .A1(n3860), .A2(n4243), .B1(n3022), .B2(n4287), .ZN(n3023)
         );
  OAI21_X1 U3845 ( .B1(n3137), .B2(n4275), .A(n3023), .ZN(n3024) );
  AOI21_X1 U3846 ( .B1(n4505), .B2(n3171), .A(n3024), .ZN(n3025) );
  OAI21_X1 U3847 ( .B1(n3026), .B2(n4122), .A(n3025), .ZN(n4502) );
  INV_X1 U3848 ( .A(n3027), .ZN(n3028) );
  OAI211_X1 U3849 ( .C1(n3028), .C2(n3100), .A(n4146), .B(n3051), .ZN(n4501)
         );
  OAI22_X1 U3850 ( .A1(n4501), .A2(n4357), .B1(n4470), .B2(n3105), .ZN(n3029)
         );
  OAI21_X1 U3851 ( .B1(n4502), .B2(n3029), .A(n4473), .ZN(n3031) );
  NAND2_X1 U3852 ( .A1(n4087), .A2(REG2_REG_4__SCAN_IN), .ZN(n3030) );
  OAI211_X1 U3853 ( .C1(n3032), .C2(n3587), .A(n3031), .B(n3030), .ZN(U3286)
         );
  NAND2_X1 U3854 ( .A1(n4100), .A2(n3033), .ZN(n3034) );
  INV_X1 U3855 ( .A(n3035), .ZN(n3042) );
  OAI22_X1 U3856 ( .A1(n4473), .A2(n3895), .B1(REG3_REG_3__SCAN_IN), .B2(n4470), .ZN(n3036) );
  AOI21_X1 U3857 ( .B1(n4183), .B2(n3859), .A(n3036), .ZN(n3037) );
  OAI21_X1 U3858 ( .B1(n3038), .B2(n4190), .A(n3037), .ZN(n3041) );
  NOR2_X1 U3859 ( .A1(n3039), .A2(n4482), .ZN(n3040) );
  AOI211_X1 U3860 ( .C1(n3042), .C2(n4476), .A(n3041), .B(n3040), .ZN(n3043)
         );
  OAI21_X1 U3861 ( .B1(n4154), .B2(n3044), .A(n3043), .ZN(U3287) );
  INV_X1 U3862 ( .A(n3045), .ZN(n3524) );
  AND2_X1 U3863 ( .A1(n3524), .A2(n3499), .ZN(n3471) );
  XOR2_X1 U3864 ( .A(n3471), .B(n3046), .Z(n3047) );
  NAND2_X1 U3865 ( .A1(n3047), .A2(n4171), .ZN(n3086) );
  AND2_X1 U3866 ( .A1(n3049), .A2(n3048), .ZN(n3050) );
  XNOR2_X1 U3867 ( .A(n3050), .B(n3471), .ZN(n3088) );
  AND2_X1 U3868 ( .A1(n3051), .A2(n3084), .ZN(n3052) );
  NOR2_X1 U3869 ( .A1(n3060), .A2(n3052), .ZN(n3106) );
  INV_X1 U3870 ( .A(n3106), .ZN(n3056) );
  AOI22_X1 U3871 ( .A1(n4185), .A2(n3859), .B1(n4183), .B2(n3857), .ZN(n3055)
         );
  OAI22_X1 U3872 ( .A1(n4473), .A2(n2387), .B1(n3154), .B2(n4470), .ZN(n3053)
         );
  AOI21_X1 U3873 ( .B1(n3084), .B2(n3325), .A(n3053), .ZN(n3054) );
  OAI211_X1 U3874 ( .C1(n4127), .C2(n3056), .A(n3055), .B(n3054), .ZN(n3057)
         );
  AOI21_X1 U3875 ( .B1(n3088), .B2(n4177), .A(n3057), .ZN(n3058) );
  OAI21_X1 U3876 ( .B1(n3086), .B2(n4482), .A(n3058), .ZN(U3285) );
  AND2_X1 U3877 ( .A1(n3527), .A2(n3523), .ZN(n3481) );
  XOR2_X1 U3878 ( .A(n3481), .B(n3059), .Z(n3115) );
  OR2_X1 U3879 ( .A1(n3060), .A2(n3138), .ZN(n3061) );
  NAND2_X1 U3880 ( .A1(n3075), .A2(n3061), .ZN(n3119) );
  INV_X1 U3881 ( .A(n3119), .ZN(n3065) );
  INV_X1 U3882 ( .A(n4185), .ZN(n3329) );
  AOI22_X1 U3883 ( .A1(n3325), .A2(n3110), .B1(n4183), .B2(n3855), .ZN(n3063)
         );
  AOI22_X1 U3884 ( .A1(n4087), .A2(REG2_REG_6__SCAN_IN), .B1(n3141), .B2(n4186), .ZN(n3062) );
  OAI211_X1 U3885 ( .C1(n3137), .C2(n3329), .A(n3063), .B(n3062), .ZN(n3064)
         );
  AOI21_X1 U3886 ( .B1(n4476), .B2(n3065), .A(n3064), .ZN(n3069) );
  XNOR2_X1 U3887 ( .A(n3066), .B(n3481), .ZN(n3113) );
  NAND2_X1 U3888 ( .A1(n4473), .A2(n4171), .ZN(n3334) );
  INV_X1 U3889 ( .A(n3334), .ZN(n3067) );
  NAND2_X1 U3890 ( .A1(n3113), .A2(n3067), .ZN(n3068) );
  OAI211_X1 U3891 ( .C1(n3115), .C2(n4154), .A(n3069), .B(n3068), .ZN(U3284)
         );
  XNOR2_X1 U3892 ( .A(n3070), .B(n3528), .ZN(n3073) );
  AOI22_X1 U3893 ( .A1(n3854), .A2(n4289), .B1(n4287), .B2(n3074), .ZN(n3071)
         );
  OAI21_X1 U3894 ( .B1(n3187), .B2(n4293), .A(n3071), .ZN(n3072) );
  AOI21_X1 U3895 ( .B1(n3073), .B2(n4171), .A(n3072), .ZN(n4510) );
  AOI21_X1 U3896 ( .B1(n3075), .B2(n3074), .A(n4283), .ZN(n3076) );
  NAND2_X1 U3897 ( .A1(n3076), .A2(n3174), .ZN(n4509) );
  INV_X1 U3898 ( .A(n4509), .ZN(n3079) );
  INV_X1 U3899 ( .A(n4148), .ZN(n3078) );
  OAI22_X1 U3900 ( .A1(n4473), .A2(n2414), .B1(n3193), .B2(n4470), .ZN(n3077)
         );
  AOI21_X1 U3901 ( .B1(n3079), .B2(n3078), .A(n3077), .ZN(n3083) );
  NAND2_X1 U3902 ( .A1(n3081), .A2(n3528), .ZN(n4507) );
  NAND3_X1 U3903 ( .A1(n3080), .A2(n4507), .A3(n4177), .ZN(n3082) );
  OAI211_X1 U3904 ( .C1(n4510), .C2(n4087), .A(n3083), .B(n3082), .ZN(U3283)
         );
  AOI22_X1 U3905 ( .A1(n3857), .A2(n4289), .B1(n4287), .B2(n3084), .ZN(n3085)
         );
  OAI211_X1 U3906 ( .C1(n3148), .C2(n4293), .A(n3086), .B(n3085), .ZN(n3087)
         );
  AOI21_X1 U3907 ( .B1(n3088), .B2(n4506), .A(n3087), .ZN(n3109) );
  AOI22_X1 U3908 ( .A1(n2727), .A2(n3106), .B1(REG0_REG_5__SCAN_IN), .B2(n4511), .ZN(n3089) );
  OAI21_X1 U3909 ( .B1(n3109), .B2(n4511), .A(n3089), .ZN(U3477) );
  OAI22_X1 U3910 ( .A1(n3148), .A2(n3682), .B1(n3681), .B2(n3100), .ZN(n3090)
         );
  XNOR2_X1 U3911 ( .A(n3090), .B(n2972), .ZN(n3124) );
  OAI22_X1 U3912 ( .A1(n3148), .A2(n3683), .B1(n3645), .B2(n3100), .ZN(n3123)
         );
  XNOR2_X1 U3913 ( .A(n3124), .B(n3123), .ZN(n3096) );
  AOI211_X1 U3914 ( .C1(n3096), .C2(n3095), .A(n3827), .B(n3125), .ZN(n3097)
         );
  INV_X1 U3915 ( .A(n3097), .ZN(n3104) );
  INV_X1 U3916 ( .A(n3822), .ZN(n3839) );
  OAI22_X1 U3917 ( .A1(n3837), .A2(n3100), .B1(n3099), .B2(n3835), .ZN(n3101)
         );
  AOI211_X1 U3918 ( .C1(n3839), .C2(n3858), .A(n3102), .B(n3101), .ZN(n3103)
         );
  OAI211_X1 U3919 ( .C1(n3843), .C2(n3105), .A(n3104), .B(n3103), .ZN(U3227)
         );
  NAND2_X1 U3920 ( .A1(n4516), .A2(REG1_REG_5__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U3921 ( .A1(n2720), .A2(n3106), .ZN(n3107) );
  OAI211_X1 U3922 ( .C1(n3109), .C2(n4516), .A(n3108), .B(n3107), .ZN(U3523)
         );
  AOI22_X1 U3923 ( .A1(n3855), .A2(n4289), .B1(n3110), .B2(n4287), .ZN(n3111)
         );
  OAI21_X1 U3924 ( .B1(n3137), .B2(n4293), .A(n3111), .ZN(n3112) );
  AOI21_X1 U3925 ( .B1(n3113), .B2(n4171), .A(n3112), .ZN(n3114) );
  OAI21_X1 U3926 ( .B1(n3115), .B2(n4262), .A(n3114), .ZN(n3121) );
  OAI22_X1 U3927 ( .A1(n4347), .A2(n3119), .B1(n4513), .B2(n2406), .ZN(n3116)
         );
  AOI21_X1 U3928 ( .B1(n3121), .B2(n4513), .A(n3116), .ZN(n3117) );
  INV_X1 U3929 ( .A(n3117), .ZN(U3479) );
  OAI22_X1 U3930 ( .A1(n4299), .A2(n3119), .B1(n4518), .B2(n3118), .ZN(n3120)
         );
  AOI21_X1 U3931 ( .B1(n3121), .B2(n4518), .A(n3120), .ZN(n3122) );
  INV_X1 U3932 ( .A(n3122), .ZN(U3524) );
  OAI22_X1 U3933 ( .A1(n3137), .A2(n3645), .B1(n3681), .B2(n3149), .ZN(n3126)
         );
  XNOR2_X1 U3934 ( .A(n3126), .B(n2972), .ZN(n3127) );
  OAI22_X1 U3935 ( .A1(n3137), .A2(n3683), .B1(n3656), .B2(n3149), .ZN(n3128)
         );
  XNOR2_X1 U3936 ( .A(n3127), .B(n3128), .ZN(n3146) );
  INV_X1 U3937 ( .A(n3127), .ZN(n3130) );
  INV_X1 U3938 ( .A(n3128), .ZN(n3129) );
  NOR2_X1 U3939 ( .A1(n3130), .A2(n3129), .ZN(n3131) );
  INV_X1 U3940 ( .A(n3131), .ZN(n3132) );
  OAI22_X1 U3941 ( .A1(n3187), .A2(n3682), .B1(n3681), .B2(n3138), .ZN(n3134)
         );
  XNOR2_X1 U3942 ( .A(n3134), .B(n2972), .ZN(n3182) );
  OAI22_X1 U3943 ( .A1(n3187), .A2(n3683), .B1(n3656), .B2(n3138), .ZN(n3183)
         );
  XNOR2_X1 U3944 ( .A(n3182), .B(n3183), .ZN(n3135) );
  XNOR2_X1 U3945 ( .A(n3184), .B(n3135), .ZN(n3143) );
  OAI21_X1 U3946 ( .B1(n3822), .B2(n3216), .A(n3136), .ZN(n3140) );
  OAI22_X1 U3947 ( .A1(n3837), .A2(n3138), .B1(n3137), .B2(n3835), .ZN(n3139)
         );
  AOI211_X1 U3948 ( .C1(n3141), .C2(n3825), .A(n3140), .B(n3139), .ZN(n3142)
         );
  OAI21_X1 U3949 ( .B1(n3143), .B2(n3827), .A(n3142), .ZN(U3236) );
  AOI211_X1 U3950 ( .C1(n3144), .C2(n3146), .A(n3827), .B(n3145), .ZN(n3147)
         );
  INV_X1 U3951 ( .A(n3147), .ZN(n3153) );
  OAI22_X1 U3952 ( .A1(n3837), .A2(n3149), .B1(n3148), .B2(n3835), .ZN(n3150)
         );
  AOI211_X1 U3953 ( .C1(n3839), .C2(n3857), .A(n3151), .B(n3150), .ZN(n3152)
         );
  OAI211_X1 U3954 ( .C1(n3843), .C2(n3154), .A(n3153), .B(n3152), .ZN(U3224)
         );
  INV_X1 U3955 ( .A(n3155), .ZN(n3507) );
  AND2_X1 U3956 ( .A1(n3507), .A2(n3534), .ZN(n3484) );
  XOR2_X1 U3957 ( .A(n3484), .B(n3156), .Z(n3157) );
  NAND2_X1 U3958 ( .A1(n3157), .A2(n4171), .ZN(n3195) );
  INV_X1 U3959 ( .A(n3173), .ZN(n3158) );
  AOI21_X1 U3960 ( .B1(n3226), .B2(n3158), .A(n3238), .ZN(n3199) );
  AOI22_X1 U3961 ( .A1(n3325), .A2(n3226), .B1(n4183), .B2(n3852), .ZN(n3159)
         );
  OAI21_X1 U3962 ( .B1(n3231), .B2(n3329), .A(n3159), .ZN(n3161) );
  OAI22_X1 U3963 ( .A1(n3236), .A2(n4470), .B1(n2443), .B2(n4473), .ZN(n3160)
         );
  AOI211_X1 U3964 ( .C1(n3199), .C2(n4476), .A(n3161), .B(n3160), .ZN(n3164)
         );
  XNOR2_X1 U3965 ( .A(n3162), .B(n3484), .ZN(n3197) );
  NAND2_X1 U3966 ( .A1(n3197), .A2(n4177), .ZN(n3163) );
  OAI211_X1 U3967 ( .C1(n3195), .C2(n4482), .A(n3164), .B(n3163), .ZN(U3281)
         );
  AND2_X1 U3968 ( .A1(n3533), .A2(n3530), .ZN(n3482) );
  XNOR2_X1 U3969 ( .A(n3165), .B(n3482), .ZN(n4478) );
  INV_X1 U3970 ( .A(n4478), .ZN(n3172) );
  XNOR2_X1 U3971 ( .A(n3166), .B(n3482), .ZN(n3169) );
  OAI22_X1 U3972 ( .A1(n3216), .A2(n4293), .B1(n3217), .B2(n4274), .ZN(n3167)
         );
  AOI21_X1 U3973 ( .B1(n4289), .B2(n3853), .A(n3167), .ZN(n3168) );
  OAI21_X1 U3974 ( .B1(n3169), .B2(n4122), .A(n3168), .ZN(n3170) );
  AOI21_X1 U3975 ( .B1(n3171), .B2(n4478), .A(n3170), .ZN(n4481) );
  OAI21_X1 U3976 ( .B1(n4497), .B2(n3172), .A(n4481), .ZN(n3178) );
  NAND2_X1 U3977 ( .A1(n3178), .A2(n4518), .ZN(n3177) );
  AOI21_X1 U3978 ( .B1(n3175), .B2(n3174), .A(n3173), .ZN(n4475) );
  NAND2_X1 U3979 ( .A1(n4475), .A2(n2720), .ZN(n3176) );
  OAI211_X1 U3980 ( .C1(n4518), .C2(n3927), .A(n3177), .B(n3176), .ZN(U3526)
         );
  INV_X1 U3981 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U3982 ( .A1(n3178), .A2(n4513), .ZN(n3180) );
  NAND2_X1 U3983 ( .A1(n4475), .A2(n2727), .ZN(n3179) );
  OAI211_X1 U3984 ( .C1(n4513), .C2(n3181), .A(n3180), .B(n3179), .ZN(U3483)
         );
  OAI22_X1 U3985 ( .A1(n3216), .A2(n3682), .B1(n3681), .B2(n3188), .ZN(n3185)
         );
  XNOR2_X1 U3986 ( .A(n3185), .B(n3666), .ZN(n3205) );
  OAI22_X1 U3987 ( .A1(n3216), .A2(n3683), .B1(n3645), .B2(n3188), .ZN(n3204)
         );
  XNOR2_X1 U3988 ( .A(n3205), .B(n3204), .ZN(n3202) );
  XOR2_X1 U3989 ( .A(n3203), .B(n3202), .Z(n3186) );
  NAND2_X1 U3990 ( .A1(n3186), .A2(n3832), .ZN(n3192) );
  OAI22_X1 U3991 ( .A1(n3837), .A2(n3188), .B1(n3187), .B2(n3835), .ZN(n3189)
         );
  AOI211_X1 U3992 ( .C1(n3839), .C2(n3854), .A(n3190), .B(n3189), .ZN(n3191)
         );
  OAI211_X1 U3993 ( .C1(n3843), .C2(n3193), .A(n3192), .B(n3191), .ZN(U3210)
         );
  AOI22_X1 U3994 ( .A1(n3852), .A2(n4289), .B1(n4287), .B2(n3226), .ZN(n3194)
         );
  OAI211_X1 U3995 ( .C1(n3231), .C2(n4293), .A(n3195), .B(n3194), .ZN(n3196)
         );
  AOI21_X1 U3996 ( .B1(n3197), .B2(n4506), .A(n3196), .ZN(n3201) );
  AOI22_X1 U3997 ( .A1(n3199), .A2(n2727), .B1(REG0_REG_9__SCAN_IN), .B2(n4511), .ZN(n3198) );
  OAI21_X1 U3998 ( .B1(n3201), .B2(n4511), .A(n3198), .ZN(U3485) );
  AOI22_X1 U3999 ( .A1(n3199), .A2(n2720), .B1(REG1_REG_9__SCAN_IN), .B2(n4516), .ZN(n3200) );
  OAI21_X1 U4000 ( .B1(n3201), .B2(n4516), .A(n3200), .ZN(U3527) );
  INV_X1 U4001 ( .A(n3204), .ZN(n3206) );
  OAI22_X1 U4002 ( .A1(n3231), .A2(n3645), .B1(n3681), .B2(n3217), .ZN(n3208)
         );
  XNOR2_X1 U4003 ( .A(n3208), .B(n2972), .ZN(n3212) );
  INV_X1 U4004 ( .A(n3212), .ZN(n3210) );
  OAI22_X1 U4005 ( .A1(n3231), .A2(n3683), .B1(n3645), .B2(n3217), .ZN(n3211)
         );
  INV_X1 U4006 ( .A(n3211), .ZN(n3209) );
  NAND2_X1 U4007 ( .A1(n3210), .A2(n3209), .ZN(n3223) );
  INV_X1 U4008 ( .A(n3223), .ZN(n3213) );
  AND2_X1 U4009 ( .A1(n3212), .A2(n3211), .ZN(n3224) );
  NOR2_X1 U4010 ( .A1(n3213), .A2(n3224), .ZN(n3214) );
  XNOR2_X1 U4011 ( .A(n3225), .B(n3214), .ZN(n3222) );
  INV_X1 U4012 ( .A(n4471), .ZN(n3220) );
  OAI21_X1 U4013 ( .B1(n3822), .B2(n3259), .A(n3215), .ZN(n3219) );
  OAI22_X1 U4014 ( .A1(n3837), .A2(n3217), .B1(n3216), .B2(n3835), .ZN(n3218)
         );
  AOI211_X1 U4015 ( .C1(n3220), .C2(n3825), .A(n3219), .B(n3218), .ZN(n3221)
         );
  OAI21_X1 U4016 ( .B1(n3222), .B2(n3827), .A(n3221), .ZN(U3218) );
  OAI22_X1 U4017 ( .A1(n3259), .A2(n3683), .B1(n3645), .B2(n3232), .ZN(n3248)
         );
  NAND2_X1 U4018 ( .A1(n3853), .A2(n3662), .ZN(n3228) );
  NAND2_X1 U4019 ( .A1(n3663), .A2(n3226), .ZN(n3227) );
  NAND2_X1 U4020 ( .A1(n3228), .A2(n3227), .ZN(n3229) );
  XNOR2_X1 U4021 ( .A(n3229), .B(n2972), .ZN(n3249) );
  XOR2_X1 U4022 ( .A(n3248), .B(n3249), .Z(n3250) );
  XNOR2_X1 U4023 ( .A(n3251), .B(n3250), .ZN(n3230) );
  NAND2_X1 U4024 ( .A1(n3230), .A2(n3832), .ZN(n3235) );
  AND2_X1 U4025 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4378) );
  OAI22_X1 U4026 ( .A1(n3837), .A2(n3232), .B1(n3231), .B2(n3835), .ZN(n3233)
         );
  AOI211_X1 U4027 ( .C1(n3839), .C2(n3852), .A(n4378), .B(n3233), .ZN(n3234)
         );
  OAI211_X1 U4028 ( .C1(n3843), .C2(n3236), .A(n3235), .B(n3234), .ZN(U3228)
         );
  AND2_X1 U4029 ( .A1(n3503), .A2(n3498), .ZN(n3472) );
  XOR2_X1 U4030 ( .A(n3472), .B(n3237), .Z(n3270) );
  OR2_X1 U4031 ( .A1(n3238), .A2(n3265), .ZN(n3239) );
  NAND2_X1 U4032 ( .A1(n3292), .A2(n3239), .ZN(n3276) );
  OAI22_X1 U4033 ( .A1(n4473), .A2(n3240), .B1(n3264), .B2(n4470), .ZN(n3241)
         );
  AOI21_X1 U4034 ( .B1(n4185), .B2(n3853), .A(n3241), .ZN(n3243) );
  AOI22_X1 U4035 ( .A1(n3325), .A2(n3252), .B1(n4183), .B2(n3851), .ZN(n3242)
         );
  OAI211_X1 U4036 ( .C1(n3276), .C2(n4127), .A(n3243), .B(n3242), .ZN(n3246)
         );
  XOR2_X1 U4037 ( .A(n3472), .B(n3244), .Z(n3268) );
  NOR2_X1 U4038 ( .A1(n3268), .A2(n3334), .ZN(n3245) );
  AOI211_X1 U4039 ( .C1(n4177), .C2(n3270), .A(n3246), .B(n3245), .ZN(n3247)
         );
  INV_X1 U4040 ( .A(n3247), .ZN(U3280) );
  NAND2_X1 U4041 ( .A1(n3852), .A2(n3662), .ZN(n3254) );
  NAND2_X1 U4042 ( .A1(n3663), .A2(n3252), .ZN(n3253) );
  NAND2_X1 U40430 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  XNOR2_X1 U4044 ( .A(n3255), .B(n2972), .ZN(n3310) );
  NOR2_X1 U4045 ( .A1(n3645), .A2(n3265), .ZN(n3256) );
  AOI21_X1 U4046 ( .B1(n2848), .B2(n3852), .A(n3256), .ZN(n3308) );
  XNOR2_X1 U4047 ( .A(n3310), .B(n3308), .ZN(n3257) );
  NAND2_X1 U4048 ( .A1(n3258), .A2(n3257), .ZN(n3312) );
  OAI211_X1 U4049 ( .C1(n3258), .C2(n3257), .A(n3312), .B(n3832), .ZN(n3263)
         );
  NAND2_X1 U4050 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4382) );
  INV_X1 U4051 ( .A(n4382), .ZN(n3261) );
  OAI22_X1 U4052 ( .A1(n3837), .A2(n3265), .B1(n3259), .B2(n3835), .ZN(n3260)
         );
  AOI211_X1 U4053 ( .C1(n3839), .C2(n3851), .A(n3261), .B(n3260), .ZN(n3262)
         );
  OAI211_X1 U4054 ( .C1(n3843), .C2(n3264), .A(n3263), .B(n3262), .ZN(U3214)
         );
  OAI22_X1 U4055 ( .A1(n3376), .A2(n4275), .B1(n4274), .B2(n3265), .ZN(n3266)
         );
  AOI21_X1 U4056 ( .B1(n4243), .B2(n3853), .A(n3266), .ZN(n3267) );
  OAI21_X1 U4057 ( .B1(n3268), .B2(n4122), .A(n3267), .ZN(n3269) );
  AOI21_X1 U4058 ( .B1(n4506), .B2(n3270), .A(n3269), .ZN(n3273) );
  MUX2_X1 U4059 ( .A(n3271), .B(n3273), .S(n4518), .Z(n3272) );
  OAI21_X1 U4060 ( .B1(n4299), .B2(n3276), .A(n3272), .ZN(U3528) );
  INV_X1 U4061 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3274) );
  MUX2_X1 U4062 ( .A(n3274), .B(n3273), .S(n4513), .Z(n3275) );
  OAI21_X1 U4063 ( .B1(n3276), .B2(n4347), .A(n3275), .ZN(U3487) );
  AND2_X1 U4064 ( .A1(n3337), .A2(n3335), .ZN(n3473) );
  INV_X1 U4065 ( .A(n3473), .ZN(n3287) );
  XNOR2_X1 U4066 ( .A(n3277), .B(n3287), .ZN(n3352) );
  AND2_X1 U4067 ( .A1(n3293), .A2(n3281), .ZN(n3278) );
  OR2_X1 U4068 ( .A1(n3278), .A2(n3344), .ZN(n3363) );
  OAI22_X1 U4069 ( .A1(n4473), .A2(n3279), .B1(n3375), .B2(n4470), .ZN(n3280)
         );
  AOI21_X1 U4070 ( .B1(n3281), .B2(n3325), .A(n3280), .ZN(n3283) );
  AOI22_X1 U4071 ( .A1(n4185), .A2(n3851), .B1(n4183), .B2(n3849), .ZN(n3282)
         );
  OAI211_X1 U4072 ( .C1(n3363), .C2(n4127), .A(n3283), .B(n3282), .ZN(n3290)
         );
  INV_X1 U4073 ( .A(n3284), .ZN(n3285) );
  AOI21_X1 U4074 ( .B1(n3298), .B2(n3286), .A(n3285), .ZN(n3338) );
  XNOR2_X1 U4075 ( .A(n3338), .B(n3287), .ZN(n3288) );
  NAND2_X1 U4076 ( .A1(n3288), .A2(n4171), .ZN(n3355) );
  NOR2_X1 U4077 ( .A1(n3355), .A2(n4482), .ZN(n3289) );
  AOI211_X1 U4078 ( .C1(n4177), .C2(n3352), .A(n3290), .B(n3289), .ZN(n3291)
         );
  INV_X1 U4079 ( .A(n3291), .ZN(U3278) );
  OAI21_X1 U4080 ( .B1(n2109), .B2(n3317), .A(n3293), .ZN(n3582) );
  INV_X1 U4081 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3303) );
  INV_X1 U4082 ( .A(n3295), .ZN(n3296) );
  AOI21_X1 U4083 ( .B1(n3486), .B2(n3294), .A(n3296), .ZN(n3588) );
  AOI22_X1 U4084 ( .A1(n3850), .A2(n4289), .B1(n4287), .B2(n3297), .ZN(n3301)
         );
  XNOR2_X1 U4085 ( .A(n3298), .B(n3486), .ZN(n3299) );
  NAND2_X1 U4086 ( .A1(n3299), .A2(n4171), .ZN(n3300) );
  OAI211_X1 U4087 ( .C1(n3588), .C2(n4100), .A(n3301), .B(n3300), .ZN(n3579)
         );
  OAI22_X1 U4088 ( .A1(n3588), .A2(n4497), .B1(n3316), .B2(n4293), .ZN(n3302)
         );
  NOR2_X1 U4089 ( .A1(n3579), .A2(n3302), .ZN(n3305) );
  MUX2_X1 U4090 ( .A(n3303), .B(n3305), .S(n4513), .Z(n3304) );
  OAI21_X1 U4091 ( .B1(n3582), .B2(n4347), .A(n3304), .ZN(U3489) );
  MUX2_X1 U4092 ( .A(n3306), .B(n3305), .S(n4518), .Z(n3307) );
  OAI21_X1 U4093 ( .B1(n4299), .B2(n3582), .A(n3307), .ZN(U3529) );
  INV_X1 U4094 ( .A(n3308), .ZN(n3309) );
  NAND2_X1 U4095 ( .A1(n3310), .A2(n3309), .ZN(n3311) );
  NAND2_X1 U4096 ( .A1(n3312), .A2(n3311), .ZN(n3366) );
  OAI22_X1 U4097 ( .A1(n3376), .A2(n3645), .B1(n3681), .B2(n3317), .ZN(n3313)
         );
  XNOR2_X1 U4098 ( .A(n3313), .B(n2972), .ZN(n3364) );
  OAI22_X1 U4099 ( .A1(n3376), .A2(n3683), .B1(n3645), .B2(n3317), .ZN(n3365)
         );
  XNOR2_X1 U4100 ( .A(n3364), .B(n3365), .ZN(n3314) );
  XNOR2_X1 U4101 ( .A(n3366), .B(n3314), .ZN(n3315) );
  NAND2_X1 U4102 ( .A1(n3315), .A2(n3832), .ZN(n3320) );
  AND2_X1 U4103 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4398) );
  OAI22_X1 U4104 ( .A1(n3837), .A2(n3317), .B1(n3316), .B2(n3835), .ZN(n3318)
         );
  AOI211_X1 U4105 ( .C1(n3839), .C2(n3850), .A(n4398), .B(n3318), .ZN(n3319)
         );
  OAI211_X1 U4106 ( .C1(n3843), .C2(n3580), .A(n3320), .B(n3319), .ZN(U3233)
         );
  XNOR2_X1 U4107 ( .A(n3438), .B(n3322), .ZN(n3398) );
  OAI21_X1 U4108 ( .B1(n3323), .B2(n3322), .A(n3321), .ZN(n3400) );
  NAND2_X1 U4109 ( .A1(n3400), .A2(n4177), .ZN(n3333) );
  OAI21_X1 U4110 ( .B1(n3346), .B2(n3712), .A(n3387), .ZN(n3406) );
  INV_X1 U4111 ( .A(n3406), .ZN(n3331) );
  AOI22_X1 U4112 ( .A1(n3325), .A2(n3324), .B1(n4183), .B2(n4184), .ZN(n3328)
         );
  INV_X1 U4113 ( .A(n3326), .ZN(n3715) );
  AOI22_X1 U4114 ( .A1(n4087), .A2(REG2_REG_14__SCAN_IN), .B1(n3715), .B2(
        n4186), .ZN(n3327) );
  OAI211_X1 U4115 ( .C1(n3711), .C2(n3329), .A(n3328), .B(n3327), .ZN(n3330)
         );
  AOI21_X1 U4116 ( .B1(n3331), .B2(n4476), .A(n3330), .ZN(n3332) );
  OAI211_X1 U4117 ( .C1(n3398), .C2(n3334), .A(n3333), .B(n3332), .ZN(U3276)
         );
  XNOR2_X1 U4118 ( .A(n3711), .B(n3793), .ZN(n3469) );
  INV_X1 U4119 ( .A(n3335), .ZN(n3336) );
  AOI21_X1 U4120 ( .B1(n3338), .B2(n3337), .A(n3336), .ZN(n3339) );
  XOR2_X1 U4121 ( .A(n3469), .B(n3339), .Z(n3342) );
  OAI22_X1 U4122 ( .A1(n4294), .A2(n4275), .B1(n4274), .B2(n3793), .ZN(n3340)
         );
  AOI21_X1 U4123 ( .B1(n4243), .B2(n3850), .A(n3340), .ZN(n3341) );
  OAI21_X1 U4124 ( .B1(n3342), .B2(n4122), .A(n3341), .ZN(n3407) );
  INV_X1 U4125 ( .A(n3407), .ZN(n3351) );
  XOR2_X1 U4126 ( .A(n3469), .B(n3343), .Z(n3408) );
  NOR2_X1 U4127 ( .A1(n3344), .A2(n3793), .ZN(n3345) );
  OR2_X1 U4128 ( .A1(n3346), .A2(n3345), .ZN(n3414) );
  INV_X1 U4129 ( .A(n3797), .ZN(n3347) );
  AOI22_X1 U4130 ( .A1(n4482), .A2(REG2_REG_13__SCAN_IN), .B1(n3347), .B2(
        n4186), .ZN(n3348) );
  OAI21_X1 U4131 ( .B1(n3414), .B2(n4127), .A(n3348), .ZN(n3349) );
  AOI21_X1 U4132 ( .B1(n3408), .B2(n4177), .A(n3349), .ZN(n3350) );
  OAI21_X1 U4133 ( .B1(n4087), .B2(n3351), .A(n3350), .ZN(U3277) );
  INV_X1 U4134 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4135 ( .A1(n3352), .A2(n4506), .ZN(n3357) );
  OAI22_X1 U4136 ( .A1(n3711), .A2(n4275), .B1(n4274), .B2(n3377), .ZN(n3354)
         );
  NOR2_X1 U4137 ( .A1(n3376), .A2(n4293), .ZN(n3353) );
  NOR2_X1 U4138 ( .A1(n3354), .A2(n3353), .ZN(n3356) );
  MUX2_X1 U4139 ( .A(n3358), .B(n3360), .S(n4513), .Z(n3359) );
  OAI21_X1 U4140 ( .B1(n3363), .B2(n4347), .A(n3359), .ZN(U3491) );
  MUX2_X1 U4141 ( .A(n3361), .B(n3360), .S(n4518), .Z(n3362) );
  OAI21_X1 U4142 ( .B1(n4299), .B2(n3363), .A(n3362), .ZN(U3530) );
  OAI21_X1 U4143 ( .B1(n3366), .B2(n3365), .A(n3364), .ZN(n3368) );
  NAND2_X1 U4144 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  AND2_X1 U4145 ( .A1(n3368), .A2(n3367), .ZN(n3600) );
  OAI22_X1 U4146 ( .A1(n3792), .A2(n3645), .B1(n3681), .B2(n3377), .ZN(n3369)
         );
  XNOR2_X1 U4147 ( .A(n3369), .B(n2972), .ZN(n3370) );
  OAI22_X1 U4148 ( .A1(n3792), .A2(n3683), .B1(n3645), .B2(n3377), .ZN(n3371)
         );
  NAND2_X1 U4149 ( .A1(n3370), .A2(n3371), .ZN(n3599) );
  INV_X1 U4150 ( .A(n3370), .ZN(n3373) );
  INV_X1 U4151 ( .A(n3371), .ZN(n3372) );
  NAND2_X1 U4152 ( .A1(n3373), .A2(n3372), .ZN(n3601) );
  NAND2_X1 U4153 ( .A1(n3599), .A2(n3601), .ZN(n3374) );
  XNOR2_X1 U4154 ( .A(n3600), .B(n3374), .ZN(n3382) );
  INV_X1 U4155 ( .A(n3375), .ZN(n3380) );
  NAND2_X1 U4156 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4402) );
  OAI21_X1 U4157 ( .B1(n3822), .B2(n3711), .A(n4402), .ZN(n3379) );
  OAI22_X1 U4158 ( .A1(n3837), .A2(n3377), .B1(n3376), .B2(n3835), .ZN(n3378)
         );
  AOI211_X1 U4159 ( .C1(n3380), .C2(n3825), .A(n3379), .B(n3378), .ZN(n3381)
         );
  OAI21_X1 U4160 ( .B1(n3382), .B2(n3827), .A(n3381), .ZN(U3221) );
  AOI21_X1 U4161 ( .B1(n3383), .B2(n3485), .A(n4122), .ZN(n3385) );
  NAND2_X1 U4162 ( .A1(n3385), .A2(n3384), .ZN(n4292) );
  XNOR2_X1 U4163 ( .A(n3386), .B(n3485), .ZN(n4296) );
  NAND2_X1 U4164 ( .A1(n4296), .A2(n4177), .ZN(n3395) );
  INV_X1 U4165 ( .A(n3387), .ZN(n3388) );
  OAI21_X1 U4166 ( .B1(n3388), .B2(n3836), .A(n4179), .ZN(n4353) );
  INV_X1 U4167 ( .A(n4353), .ZN(n3393) );
  AOI22_X1 U4168 ( .A1(n4183), .A2(n4290), .B1(n4185), .B2(n3848), .ZN(n3391)
         );
  INV_X1 U4169 ( .A(n3842), .ZN(n3389) );
  AOI22_X1 U4170 ( .A1(n4087), .A2(REG2_REG_15__SCAN_IN), .B1(n3389), .B2(
        n4186), .ZN(n3390) );
  OAI211_X1 U4171 ( .C1(n3836), .C2(n4190), .A(n3391), .B(n3390), .ZN(n3392)
         );
  AOI21_X1 U4172 ( .B1(n3393), .B2(n4476), .A(n3392), .ZN(n3394) );
  OAI211_X1 U4173 ( .C1(n4482), .C2(n4292), .A(n3395), .B(n3394), .ZN(U3275)
         );
  INV_X1 U4174 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3401) );
  OAI22_X1 U4175 ( .A1(n4277), .A2(n4275), .B1(n4274), .B2(n3712), .ZN(n3396)
         );
  AOI21_X1 U4176 ( .B1(n4243), .B2(n3849), .A(n3396), .ZN(n3397) );
  OAI21_X1 U4177 ( .B1(n3398), .B2(n4122), .A(n3397), .ZN(n3399) );
  AOI21_X1 U4178 ( .B1(n3400), .B2(n4506), .A(n3399), .ZN(n3403) );
  MUX2_X1 U4179 ( .A(n3401), .B(n3403), .S(n4513), .Z(n3402) );
  OAI21_X1 U4180 ( .B1(n3406), .B2(n4347), .A(n3402), .ZN(U3495) );
  MUX2_X1 U4181 ( .A(n3404), .B(n3403), .S(n4518), .Z(n3405) );
  OAI21_X1 U4182 ( .B1(n4299), .B2(n3406), .A(n3405), .ZN(U3532) );
  AOI21_X1 U4183 ( .B1(n4506), .B2(n3408), .A(n3407), .ZN(n3411) );
  MUX2_X1 U4184 ( .A(n3409), .B(n3411), .S(n4518), .Z(n3410) );
  OAI21_X1 U4185 ( .B1(n4299), .B2(n3414), .A(n3410), .ZN(U3531) );
  INV_X1 U4186 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3412) );
  MUX2_X1 U4187 ( .A(n3412), .B(n3411), .S(n4513), .Z(n3413) );
  OAI21_X1 U4188 ( .B1(n3414), .B2(n4347), .A(n3413), .ZN(U3493) );
  INV_X1 U4189 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U4190 ( .A1(n3415), .A2(REG2_REG_31__SCAN_IN), .ZN(n3417) );
  NAND2_X1 U4191 ( .A1(n2353), .A2(REG0_REG_31__SCAN_IN), .ZN(n3416) );
  OAI211_X1 U4192 ( .C1(n3418), .C2(n4195), .A(n3417), .B(n3416), .ZN(n3958)
         );
  INV_X1 U4193 ( .A(DATAI_30_), .ZN(n4642) );
  NOR2_X1 U4194 ( .A1(n3419), .A2(n4642), .ZN(n4202) );
  INV_X1 U4195 ( .A(n4202), .ZN(n3450) );
  OR2_X1 U4196 ( .A1(n3692), .A2(n3426), .ZN(n3420) );
  AND2_X1 U4197 ( .A1(n3421), .A2(n3420), .ZN(n3425) );
  INV_X1 U4198 ( .A(n3425), .ZN(n3557) );
  NOR3_X1 U4199 ( .A1(n3557), .A2(n3980), .A3(n3422), .ZN(n3448) );
  NAND2_X1 U4200 ( .A1(n3424), .A2(n3423), .ZN(n3444) );
  NAND2_X1 U4201 ( .A1(n3425), .A2(n3444), .ZN(n3429) );
  NAND2_X1 U4202 ( .A1(n3692), .A2(n3426), .ZN(n3427) );
  NAND2_X1 U4203 ( .A1(n2308), .A2(DATAI_31_), .ZN(n3959) );
  NAND2_X1 U4204 ( .A1(n3958), .A2(n3959), .ZN(n3564) );
  OAI211_X1 U4205 ( .C1(n3450), .C2(n3844), .A(n3427), .B(n3564), .ZN(n3443)
         );
  INV_X1 U4206 ( .A(n3443), .ZN(n3428) );
  NAND2_X1 U4207 ( .A1(n3429), .A2(n3428), .ZN(n3560) );
  NAND2_X1 U4208 ( .A1(n3430), .A2(n3437), .ZN(n3544) );
  NAND2_X1 U4209 ( .A1(n3504), .A2(n3505), .ZN(n3436) );
  INV_X1 U4210 ( .A(n3506), .ZN(n3435) );
  INV_X1 U4211 ( .A(n3431), .ZN(n3434) );
  INV_X1 U4212 ( .A(n3432), .ZN(n3465) );
  NAND3_X1 U4213 ( .A1(n3434), .A2(n3433), .A3(n3465), .ZN(n3509) );
  AOI211_X1 U4214 ( .C1(n3437), .C2(n3436), .A(n3435), .B(n3509), .ZN(n3543)
         );
  OAI21_X1 U4215 ( .B1(n3438), .B2(n3544), .A(n3543), .ZN(n3440) );
  OR2_X1 U4216 ( .A1(n3509), .A2(n3439), .ZN(n3548) );
  NAND4_X1 U4217 ( .A1(n3440), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3442)
         );
  NAND2_X1 U4218 ( .A1(n3455), .A2(n3461), .ZN(n3553) );
  AOI21_X1 U4219 ( .B1(n3442), .B2(n3441), .A(n3553), .ZN(n3446) );
  NOR3_X1 U4220 ( .A1(n3444), .A2(n3443), .A3(n3552), .ZN(n3445) );
  OAI21_X1 U4221 ( .B1(n3446), .B2(n3988), .A(n3445), .ZN(n3447) );
  OAI21_X1 U4222 ( .B1(n3448), .B2(n3560), .A(n3447), .ZN(n3449) );
  OAI21_X1 U4223 ( .B1(n3958), .B2(n3450), .A(n3449), .ZN(n3571) );
  NAND2_X1 U4224 ( .A1(n3844), .A2(n3450), .ZN(n3561) );
  AOI21_X1 U4225 ( .B1(n3561), .B2(n3958), .A(n3959), .ZN(n3452) );
  NOR2_X1 U4226 ( .A1(n3452), .A2(n3451), .ZN(n3570) );
  XNOR2_X1 U4227 ( .A(n4218), .B(n3998), .ZN(n3990) );
  NAND3_X1 U4228 ( .A1(n3453), .A2(n2174), .A3(n3990), .ZN(n3495) );
  NAND2_X1 U4229 ( .A1(n3987), .A2(n3454), .ZN(n4009) );
  NAND2_X1 U4230 ( .A1(n3455), .A2(n4004), .ZN(n4025) );
  INV_X1 U4231 ( .A(n3456), .ZN(n4040) );
  OR2_X1 U4232 ( .A1(n4039), .A2(n4040), .ZN(n4074) );
  INV_X1 U4233 ( .A(n4074), .ZN(n4071) );
  INV_X1 U4234 ( .A(n3457), .ZN(n3459) );
  NAND2_X1 U4235 ( .A1(n3459), .A2(n3458), .ZN(n4093) );
  NAND3_X1 U4236 ( .A1(n4071), .A2(n4498), .A3(n4093), .ZN(n3462) );
  NAND2_X1 U4237 ( .A1(n3461), .A2(n3460), .ZN(n4043) );
  NOR4_X1 U4238 ( .A1(n4025), .A2(n3462), .A3(n4065), .A4(n4043), .ZN(n3493)
         );
  NAND2_X1 U4239 ( .A1(n3464), .A2(n3463), .ZN(n4118) );
  NAND2_X1 U4240 ( .A1(n3465), .A2(n4112), .ZN(n4157) );
  NOR2_X1 U4241 ( .A1(n4118), .A2(n4157), .ZN(n3470) );
  XNOR2_X1 U4242 ( .A(n3844), .B(n4202), .ZN(n3468) );
  OR2_X1 U4243 ( .A1(n3958), .A2(n3959), .ZN(n3562) );
  AND3_X1 U4244 ( .A1(n3562), .A2(n3564), .A3(n3466), .ZN(n3467) );
  AND4_X1 U4245 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3492)
         );
  INV_X1 U4246 ( .A(n4139), .ZN(n3474) );
  NAND4_X1 U4247 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3480)
         );
  INV_X1 U4248 ( .A(n3475), .ZN(n3478) );
  NAND4_X1 U4249 ( .A1(n2211), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3479)
         );
  NOR2_X1 U4250 ( .A1(n3480), .A2(n3479), .ZN(n3491) );
  NAND4_X1 U4251 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3489)
         );
  INV_X1 U4252 ( .A(n3485), .ZN(n3487) );
  NAND4_X1 U4253 ( .A1(n3487), .A2(n4176), .A3(n3486), .A4(n3528), .ZN(n3488)
         );
  NOR2_X1 U4254 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  NAND4_X1 U4255 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3494)
         );
  NOR4_X1 U4256 ( .A1(n3496), .A2(n3495), .A3(n4009), .A4(n3494), .ZN(n3568)
         );
  INV_X1 U4257 ( .A(n3497), .ZN(n3555) );
  INV_X1 U4258 ( .A(n3498), .ZN(n3540) );
  INV_X1 U4259 ( .A(n3531), .ZN(n3500) );
  NOR2_X1 U4260 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  NAND4_X1 U4261 ( .A1(n3501), .A2(n3507), .A3(n3530), .A4(n3523), .ZN(n3502)
         );
  NAND2_X1 U4262 ( .A1(n3503), .A2(n3502), .ZN(n3537) );
  NAND4_X1 U4263 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(n3508)
         );
  NOR2_X1 U4264 ( .A1(n3509), .A2(n3508), .ZN(n3536) );
  OAI211_X1 U4265 ( .C1(n4356), .C2(n2096), .A(n3512), .B(n3511), .ZN(n3513)
         );
  NAND3_X1 U4266 ( .A1(n3515), .A2(n3514), .A3(n3513), .ZN(n3516) );
  NAND3_X1 U4267 ( .A1(n3518), .A2(n3517), .A3(n3516), .ZN(n3519) );
  NAND3_X1 U4268 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3522) );
  NAND4_X1 U4269 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3526)
         );
  NAND3_X1 U4270 ( .A1(n3528), .A2(n3527), .A3(n3526), .ZN(n3529) );
  NAND3_X1 U4271 ( .A1(n3531), .A2(n3530), .A3(n3529), .ZN(n3532) );
  NAND3_X1 U4272 ( .A1(n3534), .A2(n3533), .A3(n3532), .ZN(n3535) );
  AOI22_X1 U4273 ( .A1(n3543), .A2(n3537), .B1(n3536), .B2(n3535), .ZN(n3539)
         );
  OR4_X1 U4274 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3547) );
  INV_X1 U4275 ( .A(n3542), .ZN(n3545) );
  OAI21_X1 U4276 ( .B1(n3545), .B2(n3544), .A(n3543), .ZN(n3546) );
  AND4_X1 U4277 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3551)
         );
  OAI21_X1 U4278 ( .B1(n4039), .B2(n3551), .A(n3550), .ZN(n3554) );
  AOI211_X1 U4279 ( .C1(n3555), .C2(n3554), .A(n3553), .B(n3552), .ZN(n3556)
         );
  AOI211_X1 U4280 ( .C1(n3846), .C2(n4204), .A(n3557), .B(n3556), .ZN(n3559)
         );
  NAND2_X1 U4281 ( .A1(n3559), .A2(n3558), .ZN(n3566) );
  INV_X1 U4282 ( .A(n3560), .ZN(n3565) );
  NAND2_X1 U4283 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  AOI22_X1 U4284 ( .A1(n3566), .A2(n3565), .B1(n3564), .B2(n3563), .ZN(n3567)
         );
  MUX2_X1 U4285 ( .A(n3568), .B(n3567), .S(n2647), .Z(n3569) );
  AOI21_X1 U4286 ( .B1(n3571), .B2(n3570), .A(n3569), .ZN(n3572) );
  XNOR2_X1 U4287 ( .A(n3572), .B(n3952), .ZN(n3578) );
  NAND2_X1 U4288 ( .A1(n3574), .A2(n3573), .ZN(n3575) );
  OAI211_X1 U4289 ( .C1(n4355), .C2(n3577), .A(n3575), .B(B_REG_SCAN_IN), .ZN(
        n3576) );
  OAI21_X1 U4290 ( .B1(n3578), .B2(n3577), .A(n3576), .ZN(U3239) );
  NAND2_X1 U4291 ( .A1(n3579), .A2(n4473), .ZN(n3586) );
  OAI22_X1 U4292 ( .A1(n4473), .A2(n3581), .B1(n3580), .B2(n4470), .ZN(n3584)
         );
  NOR2_X1 U4293 ( .A1(n3582), .A2(n4127), .ZN(n3583) );
  AOI211_X1 U4294 ( .C1(n4185), .C2(n3852), .A(n3584), .B(n3583), .ZN(n3585)
         );
  OAI211_X1 U4295 ( .C1(n3588), .C2(n3587), .A(n3586), .B(n3585), .ZN(U3279)
         );
  INV_X1 U4296 ( .A(n3589), .ZN(n3595) );
  AOI22_X1 U4297 ( .A1(n3845), .A2(n4183), .B1(n3846), .B2(n4185), .ZN(n3591)
         );
  AOI22_X1 U4298 ( .A1(n3695), .A2(n4186), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4087), .ZN(n3590) );
  OAI211_X1 U4299 ( .C1(n3691), .C2(n4190), .A(n3591), .B(n3590), .ZN(n3594)
         );
  NOR2_X1 U4300 ( .A1(n3592), .A2(n4087), .ZN(n3593) );
  AOI211_X1 U4301 ( .C1(n4476), .C2(n3595), .A(n3594), .B(n3593), .ZN(n3596)
         );
  OAI21_X1 U4302 ( .B1(n3597), .B2(n4154), .A(n3596), .ZN(U3262) );
  OAI22_X1 U4303 ( .A1(n4218), .A2(n3682), .B1(n3681), .B2(n3998), .ZN(n3598)
         );
  XNOR2_X1 U4304 ( .A(n3598), .B(n2972), .ZN(n3671) );
  OAI22_X1 U4305 ( .A1(n4218), .A2(n3683), .B1(n3656), .B2(n3998), .ZN(n3672)
         );
  NAND2_X1 U4306 ( .A1(n3671), .A2(n3672), .ZN(n3817) );
  NAND2_X1 U4307 ( .A1(n3600), .A2(n3599), .ZN(n3602) );
  NAND2_X1 U4308 ( .A1(n3602), .A2(n3601), .ZN(n3787) );
  OAI22_X1 U4309 ( .A1(n3711), .A2(n3645), .B1(n3681), .B2(n3793), .ZN(n3603)
         );
  XOR2_X1 U4310 ( .A(n2972), .B(n3603), .Z(n3789) );
  NAND2_X1 U4311 ( .A1(n3787), .A2(n3789), .ZN(n3606) );
  OAI22_X1 U4312 ( .A1(n3711), .A2(n3683), .B1(n3645), .B2(n3793), .ZN(n3788)
         );
  INV_X1 U4313 ( .A(n3787), .ZN(n3605) );
  INV_X1 U4314 ( .A(n3789), .ZN(n3604) );
  OAI22_X1 U4315 ( .A1(n4294), .A2(n3645), .B1(n3681), .B2(n3712), .ZN(n3607)
         );
  XNOR2_X1 U4316 ( .A(n3607), .B(n2972), .ZN(n3609) );
  OAI22_X1 U4317 ( .A1(n4294), .A2(n3683), .B1(n3645), .B2(n3712), .ZN(n3608)
         );
  NAND2_X1 U4318 ( .A1(n3609), .A2(n3608), .ZN(n3707) );
  NAND2_X1 U4319 ( .A1(n3706), .A2(n3707), .ZN(n3610) );
  OR2_X1 U4320 ( .A1(n3609), .A2(n3608), .ZN(n3708) );
  NAND2_X1 U4321 ( .A1(n3610), .A2(n3708), .ZN(n3612) );
  OAI22_X1 U4322 ( .A1(n4277), .A2(n3645), .B1(n3681), .B2(n3836), .ZN(n3611)
         );
  XOR2_X1 U4323 ( .A(n2972), .B(n3611), .Z(n3613) );
  NAND2_X1 U4324 ( .A1(n3612), .A2(n3613), .ZN(n3752) );
  OAI22_X1 U4325 ( .A1(n4277), .A2(n3683), .B1(n3682), .B2(n3836), .ZN(n3830)
         );
  INV_X1 U4326 ( .A(n3612), .ZN(n3615) );
  OAI22_X1 U4327 ( .A1(n4268), .A2(n3683), .B1(n3645), .B2(n4273), .ZN(n3619)
         );
  OAI22_X1 U4328 ( .A1(n4268), .A2(n3645), .B1(n3681), .B2(n4273), .ZN(n3616)
         );
  XNOR2_X1 U4329 ( .A(n3616), .B(n2972), .ZN(n3618) );
  XOR2_X1 U4330 ( .A(n3619), .B(n3618), .Z(n3755) );
  INV_X1 U4331 ( .A(n3618), .ZN(n3621) );
  INV_X1 U4332 ( .A(n3619), .ZN(n3620) );
  NAND2_X1 U4333 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  OAI22_X1 U4334 ( .A1(n4276), .A2(n3645), .B1(n3681), .B2(n4166), .ZN(n3623)
         );
  XNOR2_X1 U4335 ( .A(n3623), .B(n2972), .ZN(n3762) );
  OAI22_X1 U4336 ( .A1(n4276), .A2(n3683), .B1(n3645), .B2(n4166), .ZN(n3763)
         );
  NAND2_X1 U4337 ( .A1(n3762), .A2(n3763), .ZN(n3624) );
  OAI22_X1 U4338 ( .A1(n4119), .A2(n3645), .B1(n3681), .B2(n4147), .ZN(n3625)
         );
  XNOR2_X1 U4339 ( .A(n3625), .B(n2972), .ZN(n3626) );
  OAI22_X1 U4340 ( .A1(n4119), .A2(n3683), .B1(n3656), .B2(n4147), .ZN(n3627)
         );
  AND2_X1 U4341 ( .A1(n3626), .A2(n3627), .ZN(n3807) );
  INV_X1 U4342 ( .A(n3626), .ZN(n3629) );
  INV_X1 U4343 ( .A(n3627), .ZN(n3628) );
  NAND2_X1 U4344 ( .A1(n3629), .A2(n3628), .ZN(n3808) );
  OAI22_X1 U4345 ( .A1(n3782), .A2(n3683), .B1(n3656), .B2(n4125), .ZN(n3632)
         );
  OAI22_X1 U4346 ( .A1(n3782), .A2(n3645), .B1(n3681), .B2(n4125), .ZN(n3630)
         );
  XNOR2_X1 U4347 ( .A(n3630), .B(n2972), .ZN(n3631) );
  XOR2_X1 U4348 ( .A(n3632), .B(n3631), .Z(n3729) );
  OAI22_X1 U4349 ( .A1(n3739), .A2(n3645), .B1(n3681), .B2(n4104), .ZN(n3636)
         );
  XNOR2_X1 U4350 ( .A(n3636), .B(n2972), .ZN(n3637) );
  OAI22_X1 U4351 ( .A1(n3739), .A2(n3683), .B1(n3656), .B2(n4104), .ZN(n3638)
         );
  NAND2_X1 U4352 ( .A1(n3637), .A2(n3638), .ZN(n3778) );
  INV_X1 U4353 ( .A(n3637), .ZN(n3640) );
  INV_X1 U4354 ( .A(n3638), .ZN(n3639) );
  NAND2_X1 U4355 ( .A1(n3640), .A2(n3639), .ZN(n3780) );
  OAI22_X1 U4356 ( .A1(n4096), .A2(n3645), .B1(n3681), .B2(n4082), .ZN(n3641)
         );
  XNOR2_X1 U4357 ( .A(n3641), .B(n2972), .ZN(n3735) );
  OAI22_X1 U4358 ( .A1(n4096), .A2(n3683), .B1(n3656), .B2(n4082), .ZN(n3734)
         );
  NOR2_X1 U4359 ( .A1(n3735), .A2(n3734), .ZN(n3644) );
  INV_X1 U4360 ( .A(n3735), .ZN(n3643) );
  INV_X1 U4361 ( .A(n3734), .ZN(n3642) );
  OAI22_X1 U4362 ( .A1(n4247), .A2(n3645), .B1(n3681), .B2(n4060), .ZN(n3646)
         );
  XNOR2_X1 U4363 ( .A(n3646), .B(n2972), .ZN(n3653) );
  OAI22_X1 U4364 ( .A1(n4247), .A2(n3683), .B1(n3656), .B2(n4060), .ZN(n3652)
         );
  XNOR2_X1 U4365 ( .A(n3653), .B(n3652), .ZN(n3799) );
  NAND2_X1 U4366 ( .A1(n4224), .A2(n3662), .ZN(n3649) );
  NAND2_X1 U4367 ( .A1(n3663), .A2(n3647), .ZN(n3648) );
  NAND2_X1 U4368 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  XNOR2_X1 U4369 ( .A(n3650), .B(n3666), .ZN(n3655) );
  NOR2_X1 U4370 ( .A1(n3645), .A2(n4049), .ZN(n3651) );
  AOI21_X1 U4371 ( .B1(n4224), .B2(n2848), .A(n3651), .ZN(n3654) );
  XNOR2_X1 U4372 ( .A(n3655), .B(n3654), .ZN(n3720) );
  NOR2_X1 U4373 ( .A1(n3653), .A2(n3652), .ZN(n3721) );
  NOR2_X1 U4374 ( .A1(n3655), .A2(n3654), .ZN(n3657) );
  OAI22_X1 U4375 ( .A1(n3747), .A2(n3683), .B1(n3656), .B2(n4033), .ZN(n3658)
         );
  INV_X1 U4376 ( .A(n3657), .ZN(n3659) );
  NAND2_X1 U4377 ( .A1(n3659), .A2(n2278), .ZN(n3660) );
  OAI22_X1 U4378 ( .A1(n3747), .A2(n3682), .B1(n3681), .B2(n4033), .ZN(n3661)
         );
  XNOR2_X1 U4379 ( .A(n3661), .B(n2972), .ZN(n3772) );
  NAND2_X1 U4380 ( .A1(n4029), .A2(n3662), .ZN(n3665) );
  NAND2_X1 U4381 ( .A1(n3663), .A2(n4214), .ZN(n3664) );
  NAND2_X1 U4382 ( .A1(n3665), .A2(n3664), .ZN(n3667) );
  XNOR2_X1 U4383 ( .A(n3667), .B(n3666), .ZN(n3670) );
  NOR2_X1 U4384 ( .A1(n3656), .A2(n4016), .ZN(n3668) );
  AOI21_X1 U4385 ( .B1(n4029), .B2(n2848), .A(n3668), .ZN(n3669) );
  NOR2_X1 U4386 ( .A1(n3670), .A2(n3669), .ZN(n3744) );
  NAND2_X1 U4387 ( .A1(n3817), .A2(n3816), .ZN(n3675) );
  INV_X1 U4388 ( .A(n3671), .ZN(n3674) );
  INV_X1 U4389 ( .A(n3672), .ZN(n3673) );
  NAND2_X1 U4390 ( .A1(n3674), .A2(n3673), .ZN(n3818) );
  NAND2_X1 U4391 ( .A1(n3675), .A2(n3818), .ZN(n3698) );
  OAI22_X1 U4392 ( .A1(n3993), .A2(n3682), .B1(n4204), .B2(n3681), .ZN(n3676)
         );
  XNOR2_X1 U4393 ( .A(n3676), .B(n2972), .ZN(n3678) );
  OAI22_X1 U4394 ( .A1(n3993), .A2(n3683), .B1(n4204), .B2(n3656), .ZN(n3677)
         );
  XNOR2_X1 U4395 ( .A(n3678), .B(n3677), .ZN(n3699) );
  INV_X1 U4396 ( .A(n3677), .ZN(n3680) );
  INV_X1 U4397 ( .A(n3678), .ZN(n3679) );
  OAI22_X1 U4398 ( .A1(n3698), .A2(n3699), .B1(n3680), .B2(n3679), .ZN(n3689)
         );
  OAI22_X1 U4399 ( .A1(n3684), .A2(n3682), .B1(n3681), .B2(n3691), .ZN(n3687)
         );
  OAI22_X1 U4400 ( .A1(n3684), .A2(n3683), .B1(n3645), .B2(n3691), .ZN(n3685)
         );
  XNOR2_X1 U4401 ( .A(n3685), .B(n2972), .ZN(n3686) );
  XOR2_X1 U4402 ( .A(n3687), .B(n3686), .Z(n3688) );
  XNOR2_X1 U4403 ( .A(n3689), .B(n3688), .ZN(n3697) );
  OAI22_X1 U4404 ( .A1(n3993), .A2(n3835), .B1(STATE_REG_SCAN_IN), .B2(n3690), 
        .ZN(n3694) );
  OAI22_X1 U4405 ( .A1(n3692), .A2(n3822), .B1(n3820), .B2(n3691), .ZN(n3693)
         );
  AOI211_X1 U4406 ( .C1(n3695), .C2(n3825), .A(n3694), .B(n3693), .ZN(n3696)
         );
  OAI21_X1 U4407 ( .B1(n3697), .B2(n3827), .A(n3696), .ZN(U3217) );
  XNOR2_X1 U4408 ( .A(n3698), .B(n3699), .ZN(n3705) );
  NOR2_X1 U4409 ( .A1(n3843), .A2(n3975), .ZN(n3703) );
  AOI22_X1 U4410 ( .A1(n4012), .A2(n3700), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3701) );
  OAI21_X1 U4411 ( .B1(n3837), .B2(n4204), .A(n3701), .ZN(n3702) );
  AOI211_X1 U4412 ( .C1(n3839), .C2(n4207), .A(n3703), .B(n3702), .ZN(n3704)
         );
  OAI21_X1 U4413 ( .B1(n3705), .B2(n3827), .A(n3704), .ZN(U3211) );
  NAND2_X1 U4414 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  XNOR2_X1 U4415 ( .A(n3706), .B(n3709), .ZN(n3717) );
  NOR2_X1 U4416 ( .A1(n4652), .A2(STATE_REG_SCAN_IN), .ZN(n4425) );
  INV_X1 U4417 ( .A(n4425), .ZN(n3710) );
  OAI21_X1 U4418 ( .B1(n3822), .B2(n4277), .A(n3710), .ZN(n3714) );
  OAI22_X1 U4419 ( .A1(n3820), .A2(n3712), .B1(n3711), .B2(n3835), .ZN(n3713)
         );
  AOI211_X1 U4420 ( .C1(n3715), .C2(n3825), .A(n3714), .B(n3713), .ZN(n3716)
         );
  OAI21_X1 U4421 ( .B1(n3717), .B2(n3827), .A(n3716), .ZN(U3212) );
  OAI21_X1 U4422 ( .B1(n3719), .B2(n3721), .A(n3720), .ZN(n3722) );
  NAND3_X1 U4423 ( .A1(n2274), .A2(n3722), .A3(n3832), .ZN(n3727) );
  OAI22_X1 U4424 ( .A1(n4247), .A2(n3835), .B1(STATE_REG_SCAN_IN), .B2(n3723), 
        .ZN(n3725) );
  OAI22_X1 U4425 ( .A1(n3747), .A2(n3822), .B1(n3837), .B2(n4049), .ZN(n3724)
         );
  AOI211_X1 U4426 ( .C1(n4051), .C2(n3825), .A(n3725), .B(n3724), .ZN(n3726)
         );
  NAND2_X1 U4427 ( .A1(n3727), .A2(n3726), .ZN(U3213) );
  XOR2_X1 U4428 ( .A(n3729), .B(n3728), .Z(n3733) );
  NAND2_X1 U4429 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3951) );
  OAI21_X1 U4430 ( .B1(n3822), .B2(n3739), .A(n3951), .ZN(n3731) );
  OAI22_X1 U4431 ( .A1(n3820), .A2(n4125), .B1(n4119), .B2(n3835), .ZN(n3730)
         );
  AOI211_X1 U4432 ( .C1(n4128), .C2(n3825), .A(n3731), .B(n3730), .ZN(n3732)
         );
  OAI21_X1 U4433 ( .B1(n3733), .B2(n3827), .A(n3732), .ZN(U3216) );
  XNOR2_X1 U4434 ( .A(n3735), .B(n3734), .ZN(n3736) );
  XNOR2_X1 U4435 ( .A(n3737), .B(n3736), .ZN(n3743) );
  OAI22_X1 U4436 ( .A1(n4247), .A2(n3822), .B1(STATE_REG_SCAN_IN), .B2(n3738), 
        .ZN(n3741) );
  OAI22_X1 U4437 ( .A1(n3820), .A2(n4082), .B1(n3739), .B2(n3835), .ZN(n3740)
         );
  AOI211_X1 U4438 ( .C1(n4079), .C2(n3825), .A(n3741), .B(n3740), .ZN(n3742)
         );
  OAI21_X1 U4439 ( .B1(n3743), .B2(n3827), .A(n3742), .ZN(U3220) );
  NOR2_X1 U4440 ( .A1(n3744), .A2(n2069), .ZN(n3745) );
  XNOR2_X1 U4441 ( .A(n3746), .B(n3745), .ZN(n3751) );
  OAI22_X1 U4442 ( .A1(n3747), .A2(n3835), .B1(n3820), .B2(n4016), .ZN(n3749)
         );
  OAI22_X1 U4443 ( .A1(n4218), .A2(n3822), .B1(STATE_REG_SCAN_IN), .B2(n4668), 
        .ZN(n3748) );
  AOI211_X1 U4444 ( .C1(n4013), .C2(n3825), .A(n3749), .B(n3748), .ZN(n3750)
         );
  OAI21_X1 U4445 ( .B1(n3751), .B2(n3827), .A(n3750), .ZN(U3222) );
  INV_X1 U4446 ( .A(n3829), .ZN(n3753) );
  OAI21_X1 U4447 ( .B1(n3753), .B2(n3830), .A(n3752), .ZN(n3754) );
  XOR2_X1 U4448 ( .A(n3755), .B(n3754), .Z(n3760) );
  INV_X1 U4449 ( .A(n3756), .ZN(n4187) );
  NAND2_X1 U4450 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4440) );
  OAI21_X1 U4451 ( .B1(n3822), .B2(n4276), .A(n4440), .ZN(n3758) );
  OAI22_X1 U4452 ( .A1(n3820), .A2(n4273), .B1(n4277), .B2(n3835), .ZN(n3757)
         );
  AOI211_X1 U4453 ( .C1(n4187), .C2(n3825), .A(n3758), .B(n3757), .ZN(n3759)
         );
  OAI21_X1 U4454 ( .B1(n3760), .B2(n3827), .A(n3759), .ZN(U3223) );
  XOR2_X1 U4455 ( .A(n3763), .B(n3762), .Z(n3764) );
  XNOR2_X1 U4456 ( .A(n3761), .B(n3764), .ZN(n3765) );
  NAND2_X1 U4457 ( .A1(n3765), .A2(n3832), .ZN(n3768) );
  NOR2_X1 U4458 ( .A1(STATE_REG_SCAN_IN), .A2(n2513), .ZN(n4453) );
  OAI22_X1 U4459 ( .A1(n3837), .A2(n4166), .B1(n4268), .B2(n3835), .ZN(n3766)
         );
  AOI211_X1 U4460 ( .C1(n3839), .C2(n4265), .A(n4453), .B(n3766), .ZN(n3767)
         );
  OAI211_X1 U4461 ( .C1(n3843), .C2(n4162), .A(n3768), .B(n3767), .ZN(U3225)
         );
  NAND2_X1 U4462 ( .A1(n3770), .A2(n3769), .ZN(n3771) );
  XOR2_X1 U4463 ( .A(n3772), .B(n3771), .Z(n3776) );
  INV_X1 U4464 ( .A(n4224), .ZN(n3802) );
  OAI22_X1 U4465 ( .A1(n3802), .A2(n3835), .B1(STATE_REG_SCAN_IN), .B2(n4654), 
        .ZN(n3774) );
  OAI22_X1 U4466 ( .A1(n4227), .A2(n3822), .B1(n3820), .B2(n4033), .ZN(n3773)
         );
  AOI211_X1 U4467 ( .C1(n4030), .C2(n3825), .A(n3774), .B(n3773), .ZN(n3775)
         );
  OAI21_X1 U4468 ( .B1(n3776), .B2(n3827), .A(n3775), .ZN(U3226) );
  AOI21_X1 U4469 ( .B1(n3780), .B2(n3778), .A(n3777), .ZN(n3779) );
  AOI21_X1 U4470 ( .B1(n2055), .B2(n3780), .A(n3779), .ZN(n3786) );
  INV_X1 U4471 ( .A(n3781), .ZN(n4106) );
  OAI22_X1 U4472 ( .A1(n3822), .A2(n4096), .B1(STATE_REG_SCAN_IN), .B2(n4520), 
        .ZN(n3784) );
  OAI22_X1 U4473 ( .A1(n3837), .A2(n4104), .B1(n3782), .B2(n3835), .ZN(n3783)
         );
  AOI211_X1 U4474 ( .C1(n4106), .C2(n3825), .A(n3784), .B(n3783), .ZN(n3785)
         );
  OAI21_X1 U4475 ( .B1(n3786), .B2(n3827), .A(n3785), .ZN(U3230) );
  XNOR2_X1 U4476 ( .A(n3789), .B(n3788), .ZN(n3790) );
  XNOR2_X1 U4477 ( .A(n3787), .B(n3790), .ZN(n3791) );
  NAND2_X1 U4478 ( .A1(n3791), .A2(n3832), .ZN(n3796) );
  AND2_X1 U4479 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4415) );
  OAI22_X1 U4480 ( .A1(n3837), .A2(n3793), .B1(n3792), .B2(n3835), .ZN(n3794)
         );
  AOI211_X1 U4481 ( .C1(n3839), .C2(n3848), .A(n4415), .B(n3794), .ZN(n3795)
         );
  OAI211_X1 U4482 ( .C1(n3843), .C2(n3797), .A(n3796), .B(n3795), .ZN(U3231)
         );
  AOI21_X1 U4483 ( .B1(n3799), .B2(n3798), .A(n3719), .ZN(n3806) );
  INV_X1 U4484 ( .A(n3800), .ZN(n4063) );
  OAI22_X1 U4485 ( .A1(n3835), .A2(n4096), .B1(STATE_REG_SCAN_IN), .B2(n3801), 
        .ZN(n3804) );
  OAI22_X1 U4486 ( .A1(n3837), .A2(n4060), .B1(n3802), .B2(n3822), .ZN(n3803)
         );
  AOI211_X1 U4487 ( .C1(n4063), .C2(n3825), .A(n3804), .B(n3803), .ZN(n3805)
         );
  OAI21_X1 U4488 ( .B1(n3806), .B2(n3827), .A(n3805), .ZN(U3232) );
  INV_X1 U4489 ( .A(n3807), .ZN(n3809) );
  NAND2_X1 U4490 ( .A1(n3809), .A2(n3808), .ZN(n3810) );
  XNOR2_X1 U4491 ( .A(n3811), .B(n3810), .ZN(n3812) );
  NAND2_X1 U4492 ( .A1(n3812), .A2(n3832), .ZN(n3815) );
  AND2_X1 U4493 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4462) );
  OAI22_X1 U4494 ( .A1(n3837), .A2(n4147), .B1(n4276), .B2(n3835), .ZN(n3813)
         );
  AOI211_X1 U4495 ( .C1(n3839), .C2(n4141), .A(n4462), .B(n3813), .ZN(n3814)
         );
  OAI211_X1 U4496 ( .C1(n3843), .C2(n4149), .A(n3815), .B(n3814), .ZN(U3235)
         );
  NAND2_X1 U4497 ( .A1(n3818), .A2(n3817), .ZN(n3819) );
  XNOR2_X1 U4498 ( .A(n3816), .B(n3819), .ZN(n3828) );
  OAI22_X1 U4499 ( .A1(n4227), .A2(n3835), .B1(n3820), .B2(n3998), .ZN(n3824)
         );
  OAI22_X1 U4500 ( .A1(n3993), .A2(n3822), .B1(STATE_REG_SCAN_IN), .B2(n3821), 
        .ZN(n3823) );
  AOI211_X1 U4501 ( .C1(n3999), .C2(n3825), .A(n3824), .B(n3823), .ZN(n3826)
         );
  OAI21_X1 U4502 ( .B1(n3828), .B2(n3827), .A(n3826), .ZN(U3237) );
  NAND2_X1 U4503 ( .A1(n3829), .A2(n3752), .ZN(n3831) );
  XNOR2_X1 U4504 ( .A(n3831), .B(n3830), .ZN(n3833) );
  NAND2_X1 U4505 ( .A1(n3833), .A2(n3832), .ZN(n3841) );
  NOR2_X1 U4506 ( .A1(n3834), .A2(STATE_REG_SCAN_IN), .ZN(n4434) );
  OAI22_X1 U4507 ( .A1(n3837), .A2(n3836), .B1(n4294), .B2(n3835), .ZN(n3838)
         );
  AOI211_X1 U4508 ( .C1(n3839), .C2(n4290), .A(n4434), .B(n3838), .ZN(n3840)
         );
  OAI211_X1 U4509 ( .C1(n3843), .C2(n3842), .A(n3841), .B(n3840), .ZN(U3238)
         );
  MUX2_X1 U4510 ( .A(DATAO_REG_31__SCAN_IN), .B(n3958), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4511 ( .A(DATAO_REG_30__SCAN_IN), .B(n3844), .S(n3856), .Z(U3580)
         );
  MUX2_X1 U4512 ( .A(DATAO_REG_29__SCAN_IN), .B(n3845), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4513 ( .A(DATAO_REG_28__SCAN_IN), .B(n4207), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4514 ( .A(DATAO_REG_27__SCAN_IN), .B(n3846), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4515 ( .A(DATAO_REG_26__SCAN_IN), .B(n4012), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4516 ( .A(DATAO_REG_25__SCAN_IN), .B(n4029), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4517 ( .A(DATAO_REG_24__SCAN_IN), .B(n4215), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4518 ( .A(DATAO_REG_23__SCAN_IN), .B(n4224), .S(n3856), .Z(U3573)
         );
  MUX2_X1 U4519 ( .A(DATAO_REG_22__SCAN_IN), .B(n4078), .S(n3856), .Z(U3572)
         );
  MUX2_X1 U4520 ( .A(DATAO_REG_21__SCAN_IN), .B(n3847), .S(n3856), .Z(U3571)
         );
  MUX2_X1 U4521 ( .A(DATAO_REG_20__SCAN_IN), .B(n4244), .S(n3856), .Z(U3570)
         );
  MUX2_X1 U4522 ( .A(DATAO_REG_19__SCAN_IN), .B(n4141), .S(n3856), .Z(U3569)
         );
  MUX2_X1 U4523 ( .A(DATAO_REG_18__SCAN_IN), .B(n4265), .S(n3856), .Z(U3568)
         );
  MUX2_X1 U4524 ( .A(DATAO_REG_17__SCAN_IN), .B(n4182), .S(n3856), .Z(U3567)
         );
  MUX2_X1 U4525 ( .A(DATAO_REG_16__SCAN_IN), .B(n4290), .S(n3856), .Z(U3566)
         );
  MUX2_X1 U4526 ( .A(DATAO_REG_15__SCAN_IN), .B(n4184), .S(n3856), .Z(U3565)
         );
  MUX2_X1 U4527 ( .A(DATAO_REG_14__SCAN_IN), .B(n3848), .S(n3856), .Z(U3564)
         );
  MUX2_X1 U4528 ( .A(DATAO_REG_13__SCAN_IN), .B(n3849), .S(n3856), .Z(U3563)
         );
  MUX2_X1 U4529 ( .A(DATAO_REG_12__SCAN_IN), .B(n3850), .S(n3856), .Z(U3562)
         );
  MUX2_X1 U4530 ( .A(DATAO_REG_11__SCAN_IN), .B(n3851), .S(n3856), .Z(U3561)
         );
  MUX2_X1 U4531 ( .A(DATAO_REG_10__SCAN_IN), .B(n3852), .S(n3856), .Z(U3560)
         );
  MUX2_X1 U4532 ( .A(DATAO_REG_9__SCAN_IN), .B(n3853), .S(U4043), .Z(U3559) );
  MUX2_X1 U4533 ( .A(DATAO_REG_8__SCAN_IN), .B(n3854), .S(n3856), .Z(U3558) );
  MUX2_X1 U4534 ( .A(DATAO_REG_7__SCAN_IN), .B(n3855), .S(n3856), .Z(U3557) );
  MUX2_X1 U4535 ( .A(DATAO_REG_6__SCAN_IN), .B(n3857), .S(n3856), .Z(U3556) );
  MUX2_X1 U4536 ( .A(DATAO_REG_5__SCAN_IN), .B(n3858), .S(U4043), .Z(U3555) );
  MUX2_X1 U4537 ( .A(DATAO_REG_4__SCAN_IN), .B(n3859), .S(U4043), .Z(U3554) );
  MUX2_X1 U4538 ( .A(DATAO_REG_3__SCAN_IN), .B(n3860), .S(U4043), .Z(U3553) );
  MUX2_X1 U4539 ( .A(DATAO_REG_2__SCAN_IN), .B(n3861), .S(U4043), .Z(U3552) );
  MUX2_X1 U4540 ( .A(DATAO_REG_1__SCAN_IN), .B(n3862), .S(U4043), .Z(U3551) );
  MUX2_X1 U4541 ( .A(DATAO_REG_0__SCAN_IN), .B(n3864), .S(U4043), .Z(U3550) );
  NAND2_X1 U4542 ( .A1(n3892), .A2(n4365), .ZN(n3873) );
  OAI211_X1 U4543 ( .C1(n3867), .C2(n3866), .A(n4465), .B(n3865), .ZN(n3872)
         );
  OAI211_X1 U4544 ( .C1(n2800), .C2(n3869), .A(n4411), .B(n3881), .ZN(n3871)
         );
  AOI22_X1 U4545 ( .A1(n4463), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3870) );
  NAND4_X1 U4546 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(U3241)
         );
  NOR2_X1 U4547 ( .A1(n3874), .A2(STATE_REG_SCAN_IN), .ZN(n3875) );
  AOI21_X1 U4548 ( .B1(n4463), .B2(ADDR_REG_2__SCAN_IN), .A(n3875), .ZN(n3876)
         );
  OAI21_X1 U4549 ( .B1(n4469), .B2(n3877), .A(n3876), .ZN(n3878) );
  INV_X1 U4550 ( .A(n3878), .ZN(n3890) );
  MUX2_X1 U4551 ( .A(n3879), .B(REG2_REG_2__SCAN_IN), .S(n4364), .Z(n3882) );
  NAND3_X1 U4552 ( .A1(n3882), .A2(n3881), .A3(n3880), .ZN(n3883) );
  NAND3_X1 U4553 ( .A1(n4411), .A2(n3884), .A3(n3883), .ZN(n3889) );
  OAI211_X1 U4554 ( .C1(n3887), .C2(n3886), .A(n4465), .B(n3885), .ZN(n3888)
         );
  NAND4_X1 U4555 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(U3242)
         );
  NAND2_X1 U4556 ( .A1(n3892), .A2(n4363), .ZN(n3901) );
  OAI211_X1 U4557 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3894), .A(n4465), .B(n3893), 
        .ZN(n3900) );
  AOI22_X1 U4558 ( .A1(n4463), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3899) );
  XNOR2_X1 U4559 ( .A(n3896), .B(n3895), .ZN(n3897) );
  NAND2_X1 U4560 ( .A1(n4411), .A2(n3897), .ZN(n3898) );
  NAND4_X1 U4561 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(U3243)
         );
  MUX2_X1 U4562 ( .A(REG2_REG_19__SCAN_IN), .B(n4130), .S(n4357), .Z(n3918) );
  INV_X1 U4563 ( .A(n3919), .ZN(n4486) );
  INV_X1 U4564 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4565 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4486), .B1(n3919), .B2(
        n3902), .ZN(n4461) );
  NOR2_X1 U4566 ( .A1(n3945), .A2(REG2_REG_17__SCAN_IN), .ZN(n3903) );
  AOI21_X1 U4567 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3945), .A(n3903), .ZN(n4451) );
  NOR2_X1 U4568 ( .A1(n4410), .A2(n4490), .ZN(n4409) );
  NAND2_X1 U4569 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3922), .ZN(n3909) );
  INV_X1 U4570 ( .A(n3922), .ZN(n4492) );
  AOI22_X1 U4571 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3922), .B1(n4492), .B2(
        n3581), .ZN(n4394) );
  NAND2_X1 U4572 ( .A1(n3923), .A2(REG2_REG_9__SCAN_IN), .ZN(n3906) );
  INV_X1 U4573 ( .A(n3923), .ZN(n4494) );
  AOI22_X1 U4574 ( .A1(n3923), .A2(REG2_REG_9__SCAN_IN), .B1(n2443), .B2(n4494), .ZN(n4374) );
  NAND2_X1 U4575 ( .A1(n3930), .A2(n3907), .ZN(n3908) );
  INV_X1 U4576 ( .A(n3930), .ZN(n4493) );
  XNOR2_X1 U4577 ( .A(n3907), .B(n4493), .ZN(n4381) );
  NAND2_X1 U4578 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4381), .ZN(n4380) );
  NAND2_X1 U4579 ( .A1(n3934), .A2(n3910), .ZN(n3911) );
  NOR2_X1 U4580 ( .A1(n2179), .A2(n3912), .ZN(n3913) );
  NOR2_X1 U4581 ( .A1(n2491), .A2(n4423), .ZN(n4422) );
  NOR2_X1 U4582 ( .A1(n3913), .A2(n4422), .ZN(n4432) );
  NAND2_X1 U4583 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3920), .ZN(n3914) );
  OAI21_X1 U4584 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3920), .A(n3914), .ZN(n4431) );
  NOR2_X1 U4585 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  INV_X1 U4586 ( .A(n3942), .ZN(n4488) );
  NAND2_X1 U4587 ( .A1(n3915), .A2(n4488), .ZN(n3916) );
  AOI21_X1 U4588 ( .B1(n3919), .B2(REG2_REG_18__SCAN_IN), .A(n4460), .ZN(n3917) );
  XOR2_X1 U4589 ( .A(n3918), .B(n3917), .Z(n3956) );
  AOI22_X1 U4590 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3919), .B1(n4486), .B2(
        n3947), .ZN(n4466) );
  NOR2_X1 U4591 ( .A1(n3945), .A2(REG1_REG_17__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4592 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3920), .ZN(n3941) );
  AOI22_X1 U4593 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3920), .B1(n4489), .B2(
        n4297), .ZN(n4437) );
  NAND2_X1 U4594 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3921), .ZN(n3937) );
  AOI22_X1 U4595 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3921), .B1(n4490), .B2(
        n3409), .ZN(n4419) );
  NAND2_X1 U4596 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3922), .ZN(n3933) );
  AOI22_X1 U4597 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3922), .B1(n4492), .B2(
        n3306), .ZN(n4391) );
  NAND2_X1 U4598 ( .A1(n3923), .A2(REG1_REG_9__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4599 ( .A1(n3923), .A2(REG1_REG_9__SCAN_IN), .B1(n2442), .B2(n4494), .ZN(n4371) );
  INV_X1 U4600 ( .A(n3925), .ZN(n3926) );
  OAI22_X1 U4601 ( .A1(n3928), .A2(n3927), .B1(n3926), .B2(n4358), .ZN(n4370)
         );
  NAND2_X1 U4602 ( .A1(n4371), .A2(n4370), .ZN(n4369) );
  NAND2_X1 U4603 ( .A1(n3929), .A2(n4369), .ZN(n3931) );
  NAND2_X1 U4604 ( .A1(n3930), .A2(n3931), .ZN(n3932) );
  XNOR2_X1 U4605 ( .A(n3931), .B(n4493), .ZN(n4386) );
  NAND2_X1 U4606 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4386), .ZN(n4385) );
  NAND2_X1 U4607 ( .A1(n3934), .A2(n3935), .ZN(n3936) );
  NAND2_X1 U4608 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4406), .ZN(n4405) );
  NAND2_X1 U4609 ( .A1(n3936), .A2(n4405), .ZN(n4418) );
  NAND2_X1 U4610 ( .A1(n4419), .A2(n4418), .ZN(n4417) );
  NAND2_X1 U4611 ( .A1(n3937), .A2(n4417), .ZN(n3939) );
  NAND2_X1 U4612 ( .A1(n3938), .A2(n3939), .ZN(n3940) );
  XNOR2_X1 U4613 ( .A(n3939), .B(n2179), .ZN(n4427) );
  NAND2_X1 U4614 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4427), .ZN(n4426) );
  NOR2_X1 U4615 ( .A1(n3942), .A2(n3943), .ZN(n3944) );
  AOI22_X1 U4616 ( .A1(n3945), .A2(n4271), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4487), .ZN(n4454) );
  OAI21_X1 U4617 ( .B1(n3947), .B2(n4486), .A(n4464), .ZN(n3949) );
  MUX2_X1 U4618 ( .A(n4258), .B(REG1_REG_19__SCAN_IN), .S(n4357), .Z(n3948) );
  XNOR2_X1 U4619 ( .A(n3949), .B(n3948), .ZN(n3954) );
  NAND2_X1 U4620 ( .A1(n4463), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3950) );
  OAI211_X1 U4621 ( .C1(n4469), .C2(n3952), .A(n3951), .B(n3950), .ZN(n3953)
         );
  AOI21_X1 U4622 ( .B1(n3954), .B2(n4465), .A(n3953), .ZN(n3955) );
  OAI21_X1 U4623 ( .B1(n3956), .B2(n4459), .A(n3955), .ZN(U3259) );
  NOR2_X2 U4624 ( .A1(n4199), .A2(n4202), .ZN(n4198) );
  XNOR2_X1 U4625 ( .A(n4198), .B(n3959), .ZN(n4303) );
  NAND2_X1 U4626 ( .A1(n3958), .A2(n3957), .ZN(n4200) );
  OAI21_X1 U4627 ( .B1(n3959), .B2(n4274), .A(n4200), .ZN(n4300) );
  NAND2_X1 U4628 ( .A1(n4473), .A2(n4300), .ZN(n3961) );
  NAND2_X1 U4629 ( .A1(n4087), .A2(REG2_REG_31__SCAN_IN), .ZN(n3960) );
  OAI211_X1 U4630 ( .C1(n4303), .C2(n4127), .A(n3961), .B(n3960), .ZN(U3260)
         );
  INV_X1 U4631 ( .A(n3962), .ZN(n3972) );
  NAND2_X1 U4632 ( .A1(n3963), .A2(n4186), .ZN(n3964) );
  OAI211_X1 U4633 ( .C1(n3966), .C2(n4127), .A(n3965), .B(n3964), .ZN(n3970)
         );
  AOI22_X1 U4634 ( .A1(n4207), .A2(n4185), .B1(n4087), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n3967) );
  OAI21_X1 U4635 ( .B1(n3968), .B2(n4190), .A(n3967), .ZN(n3969) );
  AOI21_X1 U4636 ( .B1(n3970), .B2(n4473), .A(n3969), .ZN(n3971) );
  OAI21_X1 U4637 ( .B1(n3972), .B2(n4154), .A(n3971), .ZN(U3354) );
  XNOR2_X1 U4638 ( .A(n3973), .B(n3980), .ZN(n4208) );
  AOI21_X1 U4639 ( .B1(n3974), .B2(n3997), .A(n2050), .ZN(n4309) );
  AOI22_X1 U4640 ( .A1(n4207), .A2(n4183), .B1(n4185), .B2(n4012), .ZN(n3978)
         );
  INV_X1 U4641 ( .A(n3975), .ZN(n3976) );
  AOI22_X1 U4642 ( .A1(n3976), .A2(n4186), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4482), .ZN(n3977) );
  OAI211_X1 U4643 ( .C1(n4204), .C2(n4190), .A(n3978), .B(n3977), .ZN(n3979)
         );
  AOI21_X1 U4644 ( .B1(n4309), .B2(n4476), .A(n3979), .ZN(n3985) );
  NAND2_X1 U4645 ( .A1(n3981), .A2(n3980), .ZN(n3982) );
  AOI21_X1 U4646 ( .B1(n3983), .B2(n3982), .A(n4122), .ZN(n4205) );
  NAND2_X1 U4647 ( .A1(n4205), .A2(n4473), .ZN(n3984) );
  OAI211_X1 U4648 ( .C1(n4208), .C2(n4154), .A(n3985), .B(n3984), .ZN(U3263)
         );
  XNOR2_X1 U4649 ( .A(n3986), .B(n3990), .ZN(n4211) );
  INV_X1 U4650 ( .A(n4211), .ZN(n4003) );
  INV_X1 U4651 ( .A(n4005), .ZN(n3989) );
  OAI21_X1 U4652 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n3992) );
  INV_X1 U4653 ( .A(n3990), .ZN(n3991) );
  XNOR2_X1 U4654 ( .A(n3992), .B(n3991), .ZN(n3996) );
  OAI22_X1 U4655 ( .A1(n3993), .A2(n4275), .B1(n4274), .B2(n3998), .ZN(n3994)
         );
  AOI21_X1 U4656 ( .B1(n4243), .B2(n4029), .A(n3994), .ZN(n3995) );
  OAI21_X1 U4657 ( .B1(n3996), .B2(n4122), .A(n3995), .ZN(n4210) );
  OAI21_X1 U4658 ( .B1(n4011), .B2(n3998), .A(n3997), .ZN(n4314) );
  AOI22_X1 U4659 ( .A1(n3999), .A2(n4186), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4482), .ZN(n4000) );
  OAI21_X1 U4660 ( .B1(n4314), .B2(n4127), .A(n4000), .ZN(n4001) );
  AOI21_X1 U4661 ( .B1(n4210), .B2(n4473), .A(n4001), .ZN(n4002) );
  OAI21_X1 U4662 ( .B1(n4003), .B2(n4154), .A(n4002), .ZN(U3264) );
  NAND2_X1 U4663 ( .A1(n4005), .A2(n4004), .ZN(n4006) );
  XNOR2_X1 U4664 ( .A(n4006), .B(n4009), .ZN(n4007) );
  NAND2_X1 U4665 ( .A1(n4007), .A2(n4171), .ZN(n4217) );
  XNOR2_X1 U4666 ( .A(n4008), .B(n4009), .ZN(n4220) );
  NAND2_X1 U4667 ( .A1(n4220), .A2(n4177), .ZN(n4020) );
  NOR2_X1 U4668 ( .A1(n4026), .A2(n4016), .ZN(n4010) );
  OR2_X1 U4669 ( .A1(n4011), .A2(n4010), .ZN(n4318) );
  INV_X1 U4670 ( .A(n4318), .ZN(n4018) );
  AOI22_X1 U4671 ( .A1(n4012), .A2(n4183), .B1(n4185), .B2(n4215), .ZN(n4015)
         );
  AOI22_X1 U4672 ( .A1(n4013), .A2(n4186), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4482), .ZN(n4014) );
  OAI211_X1 U4673 ( .C1(n4016), .C2(n4190), .A(n4015), .B(n4014), .ZN(n4017)
         );
  AOI21_X1 U4674 ( .B1(n4018), .B2(n4476), .A(n4017), .ZN(n4019) );
  OAI211_X1 U4675 ( .C1(n4482), .C2(n4217), .A(n4020), .B(n4019), .ZN(U3265)
         );
  INV_X1 U4676 ( .A(n4025), .ZN(n4021) );
  XNOR2_X1 U4677 ( .A(n4022), .B(n4021), .ZN(n4023) );
  NAND2_X1 U4678 ( .A1(n4023), .A2(n4171), .ZN(n4226) );
  XOR2_X1 U4679 ( .A(n4025), .B(n4024), .Z(n4229) );
  NAND2_X1 U4680 ( .A1(n4229), .A2(n4177), .ZN(n4037) );
  INV_X1 U4681 ( .A(n4048), .ZN(n4028) );
  INV_X1 U4682 ( .A(n4026), .ZN(n4027) );
  OAI21_X1 U4683 ( .B1(n4028), .B2(n4033), .A(n4027), .ZN(n4322) );
  INV_X1 U4684 ( .A(n4322), .ZN(n4035) );
  AOI22_X1 U4685 ( .A1(n4029), .A2(n4183), .B1(n4185), .B2(n4224), .ZN(n4032)
         );
  AOI22_X1 U4686 ( .A1(n4030), .A2(n4186), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4482), .ZN(n4031) );
  OAI211_X1 U4687 ( .C1(n4033), .C2(n4190), .A(n4032), .B(n4031), .ZN(n4034)
         );
  AOI21_X1 U4688 ( .B1(n4035), .B2(n4476), .A(n4034), .ZN(n4036) );
  OAI211_X1 U4689 ( .C1(n4482), .C2(n4226), .A(n4037), .B(n4036), .ZN(U3266)
         );
  XOR2_X1 U4690 ( .A(n4043), .B(n4038), .Z(n4233) );
  INV_X1 U4691 ( .A(n4233), .ZN(n4055) );
  INV_X1 U4692 ( .A(n4039), .ZN(n4041) );
  AOI21_X1 U4693 ( .B1(n4072), .B2(n4041), .A(n4040), .ZN(n4056) );
  OAI21_X1 U4694 ( .B1(n4056), .B2(n4065), .A(n4042), .ZN(n4044) );
  XNOR2_X1 U4695 ( .A(n4044), .B(n4043), .ZN(n4047) );
  OAI22_X1 U4696 ( .A1(n4247), .A2(n4293), .B1(n4274), .B2(n4049), .ZN(n4045)
         );
  AOI21_X1 U4697 ( .B1(n4215), .B2(n4289), .A(n4045), .ZN(n4046) );
  OAI21_X1 U4698 ( .B1(n4047), .B2(n4122), .A(n4046), .ZN(n4232) );
  INV_X1 U4699 ( .A(n4062), .ZN(n4050) );
  OAI21_X1 U4700 ( .B1(n4050), .B2(n4049), .A(n4048), .ZN(n4326) );
  AOI22_X1 U4701 ( .A1(REG2_REG_23__SCAN_IN), .A2(n4482), .B1(n4051), .B2(
        n4186), .ZN(n4052) );
  OAI21_X1 U4702 ( .B1(n4326), .B2(n4127), .A(n4052), .ZN(n4053) );
  AOI21_X1 U4703 ( .B1(n4232), .B2(n4473), .A(n4053), .ZN(n4054) );
  OAI21_X1 U4704 ( .B1(n4055), .B2(n4154), .A(n4054), .ZN(U3267) );
  XOR2_X1 U4705 ( .A(n4065), .B(n4056), .Z(n4059) );
  OAI22_X1 U4706 ( .A1(n4096), .A2(n4293), .B1(n4060), .B2(n4274), .ZN(n4057)
         );
  AOI21_X1 U4707 ( .B1(n4224), .B2(n4289), .A(n4057), .ZN(n4058) );
  OAI21_X1 U4708 ( .B1(n4059), .B2(n4122), .A(n4058), .ZN(n4237) );
  OR2_X1 U4709 ( .A1(n4076), .A2(n4060), .ZN(n4061) );
  NAND2_X1 U4710 ( .A1(n4062), .A2(n4061), .ZN(n4330) );
  AOI22_X1 U4711 ( .A1(n4087), .A2(REG2_REG_22__SCAN_IN), .B1(n4063), .B2(
        n4186), .ZN(n4064) );
  OAI21_X1 U4712 ( .B1(n4330), .B2(n4127), .A(n4064), .ZN(n4069) );
  NOR2_X1 U4713 ( .A1(n4066), .A2(n4065), .ZN(n4236) );
  INV_X1 U4714 ( .A(n4238), .ZN(n4067) );
  NOR3_X1 U4715 ( .A1(n4236), .A2(n4067), .A3(n4154), .ZN(n4068) );
  AOI211_X1 U4716 ( .C1(n4473), .C2(n4237), .A(n4069), .B(n4068), .ZN(n4070)
         );
  INV_X1 U4717 ( .A(n4070), .ZN(U3268) );
  XNOR2_X1 U4718 ( .A(n4072), .B(n4071), .ZN(n4073) );
  NAND2_X1 U4719 ( .A1(n4073), .A2(n4171), .ZN(n4246) );
  XNOR2_X1 U4720 ( .A(n4075), .B(n4074), .ZN(n4249) );
  NAND2_X1 U4721 ( .A1(n4249), .A2(n4177), .ZN(n4086) );
  INV_X1 U4722 ( .A(n4076), .ZN(n4077) );
  OAI21_X1 U4723 ( .B1(n4102), .B2(n4082), .A(n4077), .ZN(n4334) );
  INV_X1 U4724 ( .A(n4334), .ZN(n4084) );
  AOI22_X1 U4725 ( .A1(n4078), .A2(n4183), .B1(n4185), .B2(n4244), .ZN(n4081)
         );
  AOI22_X1 U4726 ( .A1(n4482), .A2(REG2_REG_21__SCAN_IN), .B1(n4079), .B2(
        n4186), .ZN(n4080) );
  OAI211_X1 U4727 ( .C1(n4082), .C2(n4190), .A(n4081), .B(n4080), .ZN(n4083)
         );
  AOI21_X1 U4728 ( .B1(n4084), .B2(n4476), .A(n4083), .ZN(n4085) );
  OAI211_X1 U4729 ( .C1(n4087), .C2(n4246), .A(n4086), .B(n4085), .ZN(U3269)
         );
  XOR2_X1 U4730 ( .A(n4093), .B(n4089), .Z(n4101) );
  NOR2_X1 U4731 ( .A1(n4091), .A2(n4090), .ZN(n4092) );
  XOR2_X1 U4732 ( .A(n4093), .B(n4092), .Z(n4098) );
  AOI22_X1 U4733 ( .A1(n4141), .A2(n4243), .B1(n4094), .B2(n4287), .ZN(n4095)
         );
  OAI21_X1 U4734 ( .B1(n4096), .B2(n4275), .A(n4095), .ZN(n4097) );
  AOI21_X1 U4735 ( .B1(n4098), .B2(n4171), .A(n4097), .ZN(n4099) );
  OAI21_X1 U4736 ( .B1(n4101), .B2(n4100), .A(n4099), .ZN(n4252) );
  INV_X1 U4737 ( .A(n4252), .ZN(n4110) );
  INV_X1 U4738 ( .A(n4101), .ZN(n4253) );
  INV_X1 U4739 ( .A(n4124), .ZN(n4105) );
  INV_X1 U4740 ( .A(n4102), .ZN(n4103) );
  OAI21_X1 U4741 ( .B1(n4105), .B2(n4104), .A(n4103), .ZN(n4338) );
  AOI22_X1 U4742 ( .A1(n4482), .A2(REG2_REG_20__SCAN_IN), .B1(n4106), .B2(
        n4186), .ZN(n4107) );
  OAI21_X1 U4743 ( .B1(n4338), .B2(n4127), .A(n4107), .ZN(n4108) );
  AOI21_X1 U4744 ( .B1(n4253), .B2(n4477), .A(n4108), .ZN(n4109) );
  OAI21_X1 U4745 ( .B1(n4110), .B2(n4482), .A(n4109), .ZN(U3270) );
  XNOR2_X1 U4746 ( .A(n4111), .B(n4118), .ZN(n4257) );
  INV_X1 U4747 ( .A(n4257), .ZN(n4134) );
  NAND2_X1 U4748 ( .A1(n4113), .A2(n4112), .ZN(n4138) );
  INV_X1 U4749 ( .A(n4114), .ZN(n4116) );
  OAI21_X1 U4750 ( .B1(n4138), .B2(n4116), .A(n4115), .ZN(n4117) );
  XOR2_X1 U4751 ( .A(n4118), .B(n4117), .Z(n4123) );
  OAI22_X1 U4752 ( .A1(n4119), .A2(n4293), .B1(n4274), .B2(n4125), .ZN(n4120)
         );
  AOI21_X1 U4753 ( .B1(n4244), .B2(n4289), .A(n4120), .ZN(n4121) );
  OAI21_X1 U4754 ( .B1(n4123), .B2(n4122), .A(n4121), .ZN(n4256) );
  INV_X1 U4755 ( .A(n4145), .ZN(n4126) );
  OAI21_X1 U4756 ( .B1(n4126), .B2(n4125), .A(n4124), .ZN(n4342) );
  NOR2_X1 U4757 ( .A1(n4342), .A2(n4127), .ZN(n4132) );
  INV_X1 U4758 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4130) );
  INV_X1 U4759 ( .A(n4128), .ZN(n4129) );
  OAI22_X1 U4760 ( .A1(n4473), .A2(n4130), .B1(n4129), .B2(n4470), .ZN(n4131)
         );
  AOI211_X1 U4761 ( .C1(n4256), .C2(n4473), .A(n4132), .B(n4131), .ZN(n4133)
         );
  OAI21_X1 U4762 ( .B1(n4134), .B2(n4154), .A(n4133), .ZN(U3271) );
  OAI21_X1 U4763 ( .B1(n4136), .B2(n4139), .A(n4135), .ZN(n4137) );
  INV_X1 U4764 ( .A(n4137), .ZN(n4263) );
  XOR2_X1 U4765 ( .A(n4139), .B(n4138), .Z(n4144) );
  AOI22_X1 U4766 ( .A1(n4141), .A2(n4289), .B1(n4140), .B2(n4287), .ZN(n4142)
         );
  OAI21_X1 U4767 ( .B1(n4276), .B2(n4293), .A(n4142), .ZN(n4143) );
  AOI21_X1 U4768 ( .B1(n4144), .B2(n4171), .A(n4143), .ZN(n4261) );
  INV_X1 U4769 ( .A(n4261), .ZN(n4152) );
  OAI211_X1 U4770 ( .C1(n4159), .C2(n4147), .A(n4146), .B(n4145), .ZN(n4260)
         );
  NOR2_X1 U4771 ( .A1(n4260), .A2(n4148), .ZN(n4151) );
  OAI22_X1 U4772 ( .A1(n4473), .A2(n3902), .B1(n4149), .B2(n4470), .ZN(n4150)
         );
  AOI211_X1 U4773 ( .C1(n4152), .C2(n4473), .A(n4151), .B(n4150), .ZN(n4153)
         );
  OAI21_X1 U4774 ( .B1(n4263), .B2(n4154), .A(n4153), .ZN(U3272) );
  XNOR2_X1 U4775 ( .A(n4155), .B(n4157), .ZN(n4156) );
  NAND2_X1 U4776 ( .A1(n4156), .A2(n4171), .ZN(n4267) );
  XNOR2_X1 U4777 ( .A(n4158), .B(n4157), .ZN(n4270) );
  NAND2_X1 U4778 ( .A1(n4270), .A2(n4177), .ZN(n4170) );
  INV_X1 U4779 ( .A(n4181), .ZN(n4161) );
  INV_X1 U4780 ( .A(n4159), .ZN(n4160) );
  OAI21_X1 U4781 ( .B1(n4161), .B2(n4166), .A(n4160), .ZN(n4348) );
  INV_X1 U4782 ( .A(n4348), .ZN(n4168) );
  AOI22_X1 U4783 ( .A1(n4185), .A2(n4290), .B1(n4183), .B2(n4265), .ZN(n4165)
         );
  INV_X1 U4784 ( .A(n4162), .ZN(n4163) );
  AOI22_X1 U4785 ( .A1(n4482), .A2(REG2_REG_17__SCAN_IN), .B1(n4163), .B2(
        n4186), .ZN(n4164) );
  OAI211_X1 U4786 ( .C1(n4166), .C2(n4190), .A(n4165), .B(n4164), .ZN(n4167)
         );
  AOI21_X1 U4787 ( .B1(n4168), .B2(n4476), .A(n4167), .ZN(n4169) );
  OAI211_X1 U4788 ( .C1(n4482), .C2(n4267), .A(n4170), .B(n4169), .ZN(U3273)
         );
  OAI211_X1 U4789 ( .C1(n4173), .C2(n4176), .A(n4172), .B(n4171), .ZN(n4281)
         );
  AOI21_X1 U4790 ( .B1(n4176), .B2(n4175), .A(n4174), .ZN(n4285) );
  NAND2_X1 U4791 ( .A1(n4285), .A2(n4177), .ZN(n4194) );
  NAND2_X1 U4792 ( .A1(n4179), .A2(n4178), .ZN(n4180) );
  NAND2_X1 U4793 ( .A1(n4181), .A2(n4180), .ZN(n4282) );
  INV_X1 U4794 ( .A(n4282), .ZN(n4192) );
  AOI22_X1 U4795 ( .A1(n4185), .A2(n4184), .B1(n4183), .B2(n4182), .ZN(n4189)
         );
  AOI22_X1 U4796 ( .A1(n4482), .A2(REG2_REG_16__SCAN_IN), .B1(n4187), .B2(
        n4186), .ZN(n4188) );
  OAI211_X1 U4797 ( .C1(n4273), .C2(n4190), .A(n4189), .B(n4188), .ZN(n4191)
         );
  AOI21_X1 U4798 ( .B1(n4192), .B2(n4476), .A(n4191), .ZN(n4193) );
  OAI211_X1 U4799 ( .C1(n4482), .C2(n4281), .A(n4194), .B(n4193), .ZN(U3274)
         );
  NOR2_X1 U4800 ( .A1(n4518), .A2(n4195), .ZN(n4196) );
  AOI21_X1 U4801 ( .B1(n4518), .B2(n4300), .A(n4196), .ZN(n4197) );
  OAI21_X1 U4802 ( .B1(n4303), .B2(n4299), .A(n4197), .ZN(U3549) );
  AOI21_X1 U4803 ( .B1(n4202), .B2(n4199), .A(n4198), .ZN(n4366) );
  INV_X1 U4804 ( .A(n4366), .ZN(n4306) );
  INV_X1 U4805 ( .A(n4200), .ZN(n4201) );
  AOI21_X1 U4806 ( .B1(n4202), .B2(n4287), .A(n4201), .ZN(n4368) );
  MUX2_X1 U4807 ( .A(n4368), .B(n2681), .S(n4516), .Z(n4203) );
  OAI21_X1 U4808 ( .B1(n4306), .B2(n4299), .A(n4203), .ZN(U3548) );
  OAI22_X1 U4809 ( .A1(n4218), .A2(n4293), .B1(n4204), .B2(n4274), .ZN(n4206)
         );
  INV_X1 U4810 ( .A(n4209), .ZN(U3545) );
  AOI21_X1 U4811 ( .B1(n4211), .B2(n4506), .A(n4210), .ZN(n4311) );
  MUX2_X1 U4812 ( .A(n4212), .B(n4311), .S(n4518), .Z(n4213) );
  OAI21_X1 U4813 ( .B1(n4299), .B2(n4314), .A(n4213), .ZN(U3544) );
  AOI22_X1 U4814 ( .A1(n4215), .A2(n4243), .B1(n4214), .B2(n4287), .ZN(n4216)
         );
  OAI211_X1 U4815 ( .C1(n4218), .C2(n4275), .A(n4217), .B(n4216), .ZN(n4219)
         );
  AOI21_X1 U4816 ( .B1(n4220), .B2(n4506), .A(n4219), .ZN(n4315) );
  MUX2_X1 U4817 ( .A(n4221), .B(n4315), .S(n4518), .Z(n4222) );
  OAI21_X1 U4818 ( .B1(n4299), .B2(n4318), .A(n4222), .ZN(U3543) );
  AOI22_X1 U4819 ( .A1(n4224), .A2(n4243), .B1(n4287), .B2(n4223), .ZN(n4225)
         );
  OAI211_X1 U4820 ( .C1(n4227), .C2(n4275), .A(n4226), .B(n4225), .ZN(n4228)
         );
  AOI21_X1 U4821 ( .B1(n4229), .B2(n4506), .A(n4228), .ZN(n4319) );
  MUX2_X1 U4822 ( .A(n4230), .B(n4319), .S(n4518), .Z(n4231) );
  OAI21_X1 U4823 ( .B1(n4299), .B2(n4322), .A(n4231), .ZN(U3542) );
  AOI21_X1 U4824 ( .B1(n4233), .B2(n4506), .A(n4232), .ZN(n4323) );
  MUX2_X1 U4825 ( .A(n4234), .B(n4323), .S(n4518), .Z(n4235) );
  OAI21_X1 U4826 ( .B1(n4299), .B2(n4326), .A(n4235), .ZN(U3541) );
  NOR2_X1 U4827 ( .A1(n4236), .A2(n4262), .ZN(n4239) );
  AOI21_X1 U4828 ( .B1(n4239), .B2(n4238), .A(n4237), .ZN(n4327) );
  MUX2_X1 U4829 ( .A(n4240), .B(n4327), .S(n4518), .Z(n4241) );
  OAI21_X1 U4830 ( .B1(n4299), .B2(n4330), .A(n4241), .ZN(U3540) );
  AOI22_X1 U4831 ( .A1(n4244), .A2(n4243), .B1(n4242), .B2(n4287), .ZN(n4245)
         );
  OAI211_X1 U4832 ( .C1(n4247), .C2(n4275), .A(n4246), .B(n4245), .ZN(n4248)
         );
  AOI21_X1 U4833 ( .B1(n4249), .B2(n4506), .A(n4248), .ZN(n4331) );
  MUX2_X1 U4834 ( .A(n4250), .B(n4331), .S(n4518), .Z(n4251) );
  OAI21_X1 U4835 ( .B1(n4299), .B2(n4334), .A(n4251), .ZN(U3539) );
  INV_X1 U4836 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4254) );
  AOI21_X1 U4837 ( .B1(n4504), .B2(n4253), .A(n4252), .ZN(n4335) );
  MUX2_X1 U4838 ( .A(n4254), .B(n4335), .S(n4518), .Z(n4255) );
  OAI21_X1 U4839 ( .B1(n4299), .B2(n4338), .A(n4255), .ZN(U3538) );
  AOI21_X1 U4840 ( .B1(n4257), .B2(n4506), .A(n4256), .ZN(n4339) );
  MUX2_X1 U4841 ( .A(n4258), .B(n4339), .S(n4518), .Z(n4259) );
  OAI21_X1 U4842 ( .B1(n4299), .B2(n4342), .A(n4259), .ZN(U3537) );
  OAI211_X1 U4843 ( .C1(n4263), .C2(n4262), .A(n4261), .B(n4260), .ZN(n4343)
         );
  MUX2_X1 U4844 ( .A(REG1_REG_18__SCAN_IN), .B(n4343), .S(n4518), .Z(U3536) );
  AOI22_X1 U4845 ( .A1(n4265), .A2(n4289), .B1(n4287), .B2(n4264), .ZN(n4266)
         );
  OAI211_X1 U4846 ( .C1(n4268), .C2(n4293), .A(n4267), .B(n4266), .ZN(n4269)
         );
  AOI21_X1 U4847 ( .B1(n4270), .B2(n4506), .A(n4269), .ZN(n4344) );
  MUX2_X1 U4848 ( .A(n4271), .B(n4344), .S(n4518), .Z(n4272) );
  OAI21_X1 U4849 ( .B1(n4299), .B2(n4348), .A(n4272), .ZN(U3535) );
  OAI22_X1 U4850 ( .A1(n4276), .A2(n4275), .B1(n4274), .B2(n4273), .ZN(n4279)
         );
  NOR2_X1 U4851 ( .A1(n4277), .A2(n4293), .ZN(n4278) );
  NOR2_X1 U4852 ( .A1(n4279), .A2(n4278), .ZN(n4280) );
  OAI211_X1 U4853 ( .C1(n4283), .C2(n4282), .A(n4281), .B(n4280), .ZN(n4284)
         );
  AOI21_X1 U4854 ( .B1(n4285), .B2(n4506), .A(n4284), .ZN(n4286) );
  INV_X1 U4855 ( .A(n4286), .ZN(n4349) );
  MUX2_X1 U4856 ( .A(REG1_REG_16__SCAN_IN), .B(n4349), .S(n4518), .Z(U3534) );
  AOI22_X1 U4857 ( .A1(n4290), .A2(n4289), .B1(n4288), .B2(n4287), .ZN(n4291)
         );
  OAI211_X1 U4858 ( .C1(n4294), .C2(n4293), .A(n4292), .B(n4291), .ZN(n4295)
         );
  AOI21_X1 U4859 ( .B1(n4296), .B2(n4506), .A(n4295), .ZN(n4350) );
  MUX2_X1 U4860 ( .A(n4297), .B(n4350), .S(n4518), .Z(n4298) );
  OAI21_X1 U4861 ( .B1(n4299), .B2(n4353), .A(n4298), .ZN(U3533) );
  NAND2_X1 U4862 ( .A1(n4513), .A2(n4300), .ZN(n4302) );
  NAND2_X1 U4863 ( .A1(n4511), .A2(REG0_REG_31__SCAN_IN), .ZN(n4301) );
  OAI211_X1 U4864 ( .C1(n4303), .C2(n4347), .A(n4302), .B(n4301), .ZN(U3517)
         );
  INV_X1 U4865 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4304) );
  MUX2_X1 U4866 ( .A(n4368), .B(n4304), .S(n4511), .Z(n4305) );
  OAI21_X1 U4867 ( .B1(n4306), .B2(n4347), .A(n4305), .ZN(U3516) );
  MUX2_X1 U4868 ( .A(REG0_REG_27__SCAN_IN), .B(n4307), .S(n4513), .Z(n4308) );
  AOI21_X1 U4869 ( .B1(n4309), .B2(n2727), .A(n4308), .ZN(n4310) );
  INV_X1 U4870 ( .A(n4310), .ZN(U3513) );
  INV_X1 U4871 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4312) );
  MUX2_X1 U4872 ( .A(n4312), .B(n4311), .S(n4513), .Z(n4313) );
  OAI21_X1 U4873 ( .B1(n4314), .B2(n4347), .A(n4313), .ZN(U3512) );
  INV_X1 U4874 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4316) );
  MUX2_X1 U4875 ( .A(n4316), .B(n4315), .S(n4513), .Z(n4317) );
  OAI21_X1 U4876 ( .B1(n4318), .B2(n4347), .A(n4317), .ZN(U3511) );
  INV_X1 U4877 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4320) );
  MUX2_X1 U4878 ( .A(n4320), .B(n4319), .S(n4513), .Z(n4321) );
  OAI21_X1 U4879 ( .B1(n4322), .B2(n4347), .A(n4321), .ZN(U3510) );
  INV_X1 U4880 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4324) );
  MUX2_X1 U4881 ( .A(n4324), .B(n4323), .S(n4513), .Z(n4325) );
  OAI21_X1 U4882 ( .B1(n4326), .B2(n4347), .A(n4325), .ZN(U3509) );
  INV_X1 U4883 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4328) );
  MUX2_X1 U4884 ( .A(n4328), .B(n4327), .S(n4513), .Z(n4329) );
  OAI21_X1 U4885 ( .B1(n4330), .B2(n4347), .A(n4329), .ZN(U3508) );
  INV_X1 U4886 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4332) );
  MUX2_X1 U4887 ( .A(n4332), .B(n4331), .S(n4513), .Z(n4333) );
  OAI21_X1 U4888 ( .B1(n4334), .B2(n4347), .A(n4333), .ZN(U3507) );
  INV_X1 U4889 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4336) );
  MUX2_X1 U4890 ( .A(n4336), .B(n4335), .S(n4513), .Z(n4337) );
  OAI21_X1 U4891 ( .B1(n4338), .B2(n4347), .A(n4337), .ZN(U3506) );
  INV_X1 U4892 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4340) );
  MUX2_X1 U4893 ( .A(n4340), .B(n4339), .S(n4513), .Z(n4341) );
  OAI21_X1 U4894 ( .B1(n4342), .B2(n4347), .A(n4341), .ZN(U3505) );
  MUX2_X1 U4895 ( .A(REG0_REG_18__SCAN_IN), .B(n4343), .S(n4513), .Z(U3503) );
  INV_X1 U4896 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4345) );
  MUX2_X1 U4897 ( .A(n4345), .B(n4344), .S(n4513), .Z(n4346) );
  OAI21_X1 U4898 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(U3501) );
  MUX2_X1 U4899 ( .A(REG0_REG_16__SCAN_IN), .B(n4349), .S(n4513), .Z(U3499) );
  INV_X1 U4900 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4351) );
  MUX2_X1 U4901 ( .A(n4351), .B(n4350), .S(n4513), .Z(n4352) );
  OAI21_X1 U4902 ( .B1(n4353), .B2(n4347), .A(n4352), .ZN(U3497) );
  MUX2_X1 U4903 ( .A(DATAI_30_), .B(n4354), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4904 ( .A(DATAI_22_), .B(n4355), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4905 ( .A(n4356), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4906 ( .A(n4357), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4907 ( .A(DATAI_8_), .B(n2147), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4908 ( .A(n4359), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4909 ( .A(DATAI_6_), .B(n4360), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U4910 ( .A(n4361), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4911 ( .A(DATAI_4_), .B(n4362), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4912 ( .A(n4363), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4913 ( .A(n4364), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4914 ( .A(n4365), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4915 ( .A1(n4366), .A2(n4476), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4482), .ZN(n4367) );
  OAI21_X1 U4916 ( .B1(n4482), .B2(n4368), .A(n4367), .ZN(U3261) );
  OAI211_X1 U4917 ( .C1(n4371), .C2(n4370), .A(n4465), .B(n4369), .ZN(n4376)
         );
  OAI211_X1 U4918 ( .C1(n4374), .C2(n4373), .A(n4411), .B(n4372), .ZN(n4375)
         );
  OAI211_X1 U4919 ( .C1(n4469), .C2(n4494), .A(n4376), .B(n4375), .ZN(n4377)
         );
  AOI211_X1 U4920 ( .C1(n4463), .C2(ADDR_REG_9__SCAN_IN), .A(n4378), .B(n4377), 
        .ZN(n4379) );
  INV_X1 U4921 ( .A(n4379), .ZN(U3249) );
  OAI211_X1 U4922 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4381), .A(n4411), .B(n4380), .ZN(n4383) );
  NAND2_X1 U4923 ( .A1(n4383), .A2(n4382), .ZN(n4384) );
  AOI21_X1 U4924 ( .B1(n4463), .B2(ADDR_REG_10__SCAN_IN), .A(n4384), .ZN(n4388) );
  OAI211_X1 U4925 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4386), .A(n4465), .B(n4385), .ZN(n4387) );
  OAI211_X1 U4926 ( .C1(n4469), .C2(n4493), .A(n4388), .B(n4387), .ZN(U3250)
         );
  OAI211_X1 U4927 ( .C1(n4391), .C2(n4390), .A(n4465), .B(n4389), .ZN(n4396)
         );
  OAI211_X1 U4928 ( .C1(n4394), .C2(n4393), .A(n4411), .B(n4392), .ZN(n4395)
         );
  OAI211_X1 U4929 ( .C1(n4469), .C2(n4492), .A(n4396), .B(n4395), .ZN(n4397)
         );
  AOI211_X1 U4930 ( .C1(n4463), .C2(ADDR_REG_11__SCAN_IN), .A(n4398), .B(n4397), .ZN(n4399) );
  INV_X1 U4931 ( .A(n4399), .ZN(U3251) );
  OAI211_X1 U4932 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4401), .A(n4411), .B(n4400), .ZN(n4403) );
  NAND2_X1 U4933 ( .A1(n4403), .A2(n4402), .ZN(n4404) );
  AOI21_X1 U4934 ( .B1(n4463), .B2(ADDR_REG_12__SCAN_IN), .A(n4404), .ZN(n4408) );
  OAI211_X1 U4935 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4406), .A(n4465), .B(n4405), .ZN(n4407) );
  OAI211_X1 U4936 ( .C1(n4469), .C2(n4491), .A(n4408), .B(n4407), .ZN(U3252)
         );
  AOI21_X1 U4937 ( .B1(n4410), .B2(n4490), .A(n4409), .ZN(n4414) );
  OAI21_X1 U4938 ( .B1(n4414), .B2(n4413), .A(n4411), .ZN(n4412) );
  AOI21_X1 U4939 ( .B1(n4414), .B2(n4413), .A(n4412), .ZN(n4416) );
  AOI211_X1 U4940 ( .C1(n4463), .C2(ADDR_REG_13__SCAN_IN), .A(n4416), .B(n4415), .ZN(n4421) );
  OAI211_X1 U4941 ( .C1(n4419), .C2(n4418), .A(n4465), .B(n4417), .ZN(n4420)
         );
  OAI211_X1 U4942 ( .C1(n4469), .C2(n4490), .A(n4421), .B(n4420), .ZN(U3253)
         );
  AOI211_X1 U4943 ( .C1(n2491), .C2(n4423), .A(n4422), .B(n4459), .ZN(n4424)
         );
  AOI211_X1 U4944 ( .C1(n4463), .C2(ADDR_REG_14__SCAN_IN), .A(n4425), .B(n4424), .ZN(n4429) );
  OAI211_X1 U4945 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4427), .A(n4465), .B(n4426), .ZN(n4428) );
  OAI211_X1 U4946 ( .C1(n4469), .C2(n2179), .A(n4429), .B(n4428), .ZN(U3254)
         );
  AOI211_X1 U4947 ( .C1(n4432), .C2(n4431), .A(n4430), .B(n4459), .ZN(n4433)
         );
  AOI211_X1 U4948 ( .C1(n4463), .C2(ADDR_REG_15__SCAN_IN), .A(n4434), .B(n4433), .ZN(n4439) );
  OAI211_X1 U4949 ( .C1(n4437), .C2(n4436), .A(n4465), .B(n4435), .ZN(n4438)
         );
  OAI211_X1 U4950 ( .C1(n4469), .C2(n4489), .A(n4439), .B(n4438), .ZN(U3255)
         );
  INV_X1 U4951 ( .A(n4440), .ZN(n4444) );
  AOI221_X1 U4952 ( .B1(n4442), .B2(n4441), .C1(n2313), .C2(n4441), .A(n4459), 
        .ZN(n4443) );
  AOI211_X1 U4953 ( .C1(n4463), .C2(ADDR_REG_16__SCAN_IN), .A(n4444), .B(n4443), .ZN(n4448) );
  OAI221_X1 U4954 ( .B1(n4446), .B2(REG1_REG_16__SCAN_IN), .C1(n4446), .C2(
        n4445), .A(n4465), .ZN(n4447) );
  OAI211_X1 U4955 ( .C1(n4469), .C2(n4488), .A(n4448), .B(n4447), .ZN(U3256)
         );
  AOI221_X1 U4956 ( .B1(n4451), .B2(n4450), .C1(n4449), .C2(n4450), .A(n4459), 
        .ZN(n4452) );
  AOI211_X1 U4957 ( .C1(n4463), .C2(ADDR_REG_17__SCAN_IN), .A(n4453), .B(n4452), .ZN(n4458) );
  OAI221_X1 U4958 ( .B1(n4456), .B2(n4455), .C1(n4456), .C2(n4454), .A(n4465), 
        .ZN(n4457) );
  OAI211_X1 U4959 ( .C1(n4469), .C2(n4487), .A(n4458), .B(n4457), .ZN(U3257)
         );
  OAI211_X1 U4960 ( .C1(n4466), .C2(n2066), .A(n4465), .B(n4464), .ZN(n4467)
         );
  OAI211_X1 U4961 ( .C1(n4469), .C2(n4486), .A(n4468), .B(n4467), .ZN(U3258)
         );
  OAI22_X1 U4962 ( .A1(n4473), .A2(n4472), .B1(n4471), .B2(n4470), .ZN(n4474)
         );
  INV_X1 U4963 ( .A(n4474), .ZN(n4480) );
  AOI22_X1 U4964 ( .A1(n4478), .A2(n4477), .B1(n4476), .B2(n4475), .ZN(n4479)
         );
  OAI211_X1 U4965 ( .C1(n4482), .C2(n4481), .A(n4480), .B(n4479), .ZN(U3282)
         );
  AND2_X1 U4966 ( .A1(D_REG_31__SCAN_IN), .A2(n4483), .ZN(U3291) );
  AND2_X1 U4967 ( .A1(D_REG_30__SCAN_IN), .A2(n4483), .ZN(U3292) );
  AND2_X1 U4968 ( .A1(D_REG_29__SCAN_IN), .A2(n4483), .ZN(U3293) );
  AND2_X1 U4969 ( .A1(D_REG_28__SCAN_IN), .A2(n4483), .ZN(U3294) );
  AND2_X1 U4970 ( .A1(D_REG_27__SCAN_IN), .A2(n4483), .ZN(U3295) );
  AND2_X1 U4971 ( .A1(D_REG_26__SCAN_IN), .A2(n4483), .ZN(U3296) );
  AND2_X1 U4972 ( .A1(D_REG_25__SCAN_IN), .A2(n4483), .ZN(U3297) );
  AND2_X1 U4973 ( .A1(D_REG_24__SCAN_IN), .A2(n4483), .ZN(U3298) );
  AND2_X1 U4974 ( .A1(D_REG_23__SCAN_IN), .A2(n4483), .ZN(U3299) );
  AND2_X1 U4975 ( .A1(D_REG_22__SCAN_IN), .A2(n4483), .ZN(U3300) );
  AND2_X1 U4976 ( .A1(D_REG_21__SCAN_IN), .A2(n4483), .ZN(U3301) );
  AND2_X1 U4977 ( .A1(D_REG_20__SCAN_IN), .A2(n4483), .ZN(U3302) );
  AND2_X1 U4978 ( .A1(D_REG_19__SCAN_IN), .A2(n4483), .ZN(U3303) );
  AND2_X1 U4979 ( .A1(D_REG_18__SCAN_IN), .A2(n4483), .ZN(U3304) );
  AND2_X1 U4980 ( .A1(D_REG_17__SCAN_IN), .A2(n4483), .ZN(U3305) );
  AND2_X1 U4981 ( .A1(D_REG_16__SCAN_IN), .A2(n4483), .ZN(U3306) );
  AND2_X1 U4982 ( .A1(D_REG_15__SCAN_IN), .A2(n4483), .ZN(U3307) );
  AND2_X1 U4983 ( .A1(D_REG_14__SCAN_IN), .A2(n4483), .ZN(U3308) );
  AND2_X1 U4984 ( .A1(D_REG_13__SCAN_IN), .A2(n4483), .ZN(U3309) );
  AND2_X1 U4985 ( .A1(D_REG_12__SCAN_IN), .A2(n4483), .ZN(U3310) );
  AND2_X1 U4986 ( .A1(D_REG_11__SCAN_IN), .A2(n4483), .ZN(U3311) );
  AND2_X1 U4987 ( .A1(D_REG_10__SCAN_IN), .A2(n4483), .ZN(U3312) );
  AND2_X1 U4988 ( .A1(D_REG_9__SCAN_IN), .A2(n4483), .ZN(U3313) );
  AND2_X1 U4989 ( .A1(D_REG_8__SCAN_IN), .A2(n4483), .ZN(U3314) );
  AND2_X1 U4990 ( .A1(D_REG_7__SCAN_IN), .A2(n4483), .ZN(U3315) );
  AND2_X1 U4991 ( .A1(D_REG_6__SCAN_IN), .A2(n4483), .ZN(U3316) );
  AND2_X1 U4992 ( .A1(D_REG_5__SCAN_IN), .A2(n4483), .ZN(U3317) );
  AND2_X1 U4993 ( .A1(D_REG_4__SCAN_IN), .A2(n4483), .ZN(U3318) );
  AND2_X1 U4994 ( .A1(D_REG_3__SCAN_IN), .A2(n4483), .ZN(U3319) );
  AND2_X1 U4995 ( .A1(D_REG_2__SCAN_IN), .A2(n4483), .ZN(U3320) );
  AOI21_X1 U4996 ( .B1(U3149), .B2(n2580), .A(n4484), .ZN(U3329) );
  INV_X1 U4997 ( .A(DATAI_18_), .ZN(n4485) );
  AOI22_X1 U4998 ( .A1(STATE_REG_SCAN_IN), .A2(n4486), .B1(n4485), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n4487), .B1(n2523), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5000 ( .A(DATAI_16_), .ZN(n4656) );
  AOI22_X1 U5001 ( .A1(STATE_REG_SCAN_IN), .A2(n4488), .B1(n4656), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5002 ( .A1(STATE_REG_SCAN_IN), .A2(n4489), .B1(n4641), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5003 ( .A(DATAI_14_), .ZN(n4666) );
  AOI22_X1 U5004 ( .A1(STATE_REG_SCAN_IN), .A2(n2179), .B1(n4666), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5005 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .B1(n2336), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5006 ( .A1(STATE_REG_SCAN_IN), .A2(n4491), .B1(n2484), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5007 ( .A(DATAI_11_), .ZN(n4639) );
  AOI22_X1 U5008 ( .A1(STATE_REG_SCAN_IN), .A2(n4492), .B1(n4639), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5009 ( .A(DATAI_10_), .ZN(n4551) );
  AOI22_X1 U5010 ( .A1(STATE_REG_SCAN_IN), .A2(n4493), .B1(n4551), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5011 ( .A(DATAI_9_), .ZN(n4659) );
  AOI22_X1 U5012 ( .A1(STATE_REG_SCAN_IN), .A2(n4494), .B1(n4659), .B2(U3149), 
        .ZN(U3343) );
  OAI211_X1 U5013 ( .C1(n4498), .C2(n4497), .A(n4496), .B(n4495), .ZN(n4499)
         );
  INV_X1 U5014 ( .A(n4499), .ZN(n4514) );
  INV_X1 U5015 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5016 ( .A1(n4513), .A2(n4514), .B1(n4500), .B2(n4511), .ZN(U3467)
         );
  INV_X1 U5017 ( .A(n4501), .ZN(n4503) );
  AOI211_X1 U5018 ( .C1(n4505), .C2(n4504), .A(n4503), .B(n4502), .ZN(n4515)
         );
  AOI22_X1 U5019 ( .A1(n4513), .A2(n4515), .B1(n2369), .B2(n4511), .ZN(U3475)
         );
  NAND3_X1 U5020 ( .A1(n3080), .A2(n4507), .A3(n4506), .ZN(n4508) );
  INV_X1 U5021 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5022 ( .A1(n4513), .A2(n4517), .B1(n4512), .B2(n4511), .ZN(U3481)
         );
  AOI22_X1 U5023 ( .A1(n4518), .A2(n4514), .B1(n2346), .B2(n4516), .ZN(U3518)
         );
  AOI22_X1 U5024 ( .A1(n4518), .A2(n4515), .B1(n2373), .B2(n4516), .ZN(U3522)
         );
  AOI22_X1 U5025 ( .A1(n4518), .A2(n4517), .B1(n2416), .B2(n4516), .ZN(U3525)
         );
  AOI22_X1 U5026 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4702) );
  AOI22_X1 U5027 ( .A1(n4520), .A2(keyinput_g53), .B1(keyinput_g20), .B2(n4639), .ZN(n4519) );
  OAI221_X1 U5028 ( .B1(n4520), .B2(keyinput_g53), .C1(n4639), .C2(
        keyinput_g20), .A(n4519), .ZN(n4528) );
  XNOR2_X1 U5029 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4524) );
  XNOR2_X1 U5030 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4523) );
  XNOR2_X1 U5031 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_g42), .ZN(n4522) );
  XNOR2_X1 U5032 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4521) );
  NAND4_X1 U5033 ( .A1(n4524), .A2(n4523), .A3(n4522), .A4(n4521), .ZN(n4527)
         );
  XNOR2_X1 U5034 ( .A(keyinput_g2), .B(n4643), .ZN(n4526) );
  XNOR2_X1 U5035 ( .A(keyinput_g3), .B(n2627), .ZN(n4525) );
  NOR4_X1 U5036 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(n4563)
         );
  AOI22_X1 U5037 ( .A1(n4530), .A2(keyinput_g0), .B1(n4652), .B2(keyinput_g35), 
        .ZN(n4529) );
  OAI221_X1 U5038 ( .B1(n4530), .B2(keyinput_g0), .C1(n4652), .C2(keyinput_g35), .A(n4529), .ZN(n4538) );
  AOI22_X1 U5039 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(REG3_REG_10__SCAN_IN), 
        .B2(keyinput_g37), .ZN(n4531) );
  OAI221_X1 U5040 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(REG3_REG_10__SCAN_IN), .C2(keyinput_g37), .A(n4531), .ZN(n4537) );
  AOI22_X1 U5041 ( .A1(n4657), .A2(keyinput_g26), .B1(n4656), .B2(keyinput_g15), .ZN(n4532) );
  OAI221_X1 U5042 ( .B1(n4657), .B2(keyinput_g26), .C1(n4656), .C2(
        keyinput_g15), .A(n4532), .ZN(n4536) );
  AOI22_X1 U5043 ( .A1(n4534), .A2(keyinput_g6), .B1(n4660), .B2(keyinput_g33), 
        .ZN(n4533) );
  OAI221_X1 U5044 ( .B1(n4534), .B2(keyinput_g6), .C1(n4660), .C2(keyinput_g33), .A(n4533), .ZN(n4535) );
  NOR4_X1 U5045 ( .A1(n4538), .A2(n4537), .A3(n4536), .A4(n4535), .ZN(n4562)
         );
  AOI22_X1 U5046 ( .A1(n2580), .A2(keyinput_g8), .B1(n2513), .B2(keyinput_g48), 
        .ZN(n4539) );
  OAI221_X1 U5047 ( .B1(n2580), .B2(keyinput_g8), .C1(n2513), .C2(keyinput_g48), .A(n4539), .ZN(n4549) );
  INV_X1 U5048 ( .A(DATAI_19_), .ZN(n4541) );
  AOI22_X1 U5049 ( .A1(n4668), .A2(keyinput_g45), .B1(keyinput_g12), .B2(n4541), .ZN(n4540) );
  OAI221_X1 U5050 ( .B1(n4668), .B2(keyinput_g45), .C1(n4541), .C2(
        keyinput_g12), .A(n4540), .ZN(n4548) );
  XOR2_X1 U5051 ( .A(n3690), .B(keyinput_g40), .Z(n4546) );
  XOR2_X1 U5052 ( .A(n4542), .B(keyinput_g7), .Z(n4545) );
  XNOR2_X1 U5053 ( .A(DATAI_3_), .B(keyinput_g28), .ZN(n4544) );
  XNOR2_X1 U5054 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_g62), .ZN(n4543) );
  NAND4_X1 U5055 ( .A1(n4546), .A2(n4545), .A3(n4544), .A4(n4543), .ZN(n4547)
         );
  NOR3_X1 U5056 ( .A1(n4549), .A2(n4548), .A3(n4547), .ZN(n4561) );
  AOI22_X1 U5057 ( .A1(n4551), .A2(keyinput_g21), .B1(n3738), .B2(keyinput_g43), .ZN(n4550) );
  OAI221_X1 U5058 ( .B1(n4551), .B2(keyinput_g21), .C1(n3738), .C2(
        keyinput_g43), .A(n4550), .ZN(n4559) );
  XNOR2_X1 U5059 ( .A(n4618), .B(keyinput_g58), .ZN(n4558) );
  XNOR2_X1 U5060 ( .A(keyinput_g18), .B(n2336), .ZN(n4557) );
  XNOR2_X1 U5061 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_g36), .ZN(n4555) );
  XNOR2_X1 U5062 ( .A(DATAI_1_), .B(keyinput_g30), .ZN(n4554) );
  XNOR2_X1 U5063 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_g49), .ZN(n4553) );
  XNOR2_X1 U5064 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4552) );
  NAND4_X1 U5065 ( .A1(n4555), .A2(n4554), .A3(n4553), .A4(n4552), .ZN(n4556)
         );
  NOR4_X1 U5066 ( .A1(n4559), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4560)
         );
  NAND4_X1 U5067 ( .A1(n4563), .A2(n4562), .A3(n4561), .A4(n4560), .ZN(n4700)
         );
  AOI22_X1 U5068 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_26_), .B2(
        keyinput_g5), .ZN(n4564) );
  OAI221_X1 U5069 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_26_), .C2(
        keyinput_g5), .A(n4564), .ZN(n4571) );
  AOI22_X1 U5070 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(DATAI_27_), .B2(
        keyinput_g4), .ZN(n4565) );
  OAI221_X1 U5071 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(DATAI_27_), .C2(
        keyinput_g4), .A(n4565), .ZN(n4570) );
  AOI22_X1 U5072 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_g51), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_g55), .ZN(n4566) );
  OAI221_X1 U5073 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_g55), .A(n4566), .ZN(n4569) );
  AOI22_X1 U5074 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .ZN(n4567) );
  OAI221_X1 U5075 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_g44), .A(n4567), .ZN(n4568) );
  NOR4_X1 U5076 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4599)
         );
  XNOR2_X1 U5077 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_g41), .ZN(n4579) );
  AOI22_X1 U5078 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(n4573), 
        .B2(keyinput_g34), .ZN(n4572) );
  OAI221_X1 U5079 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(n4573), 
        .C2(keyinput_g34), .A(n4572), .ZN(n4578) );
  AOI22_X1 U5080 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(DATAI_21_), .B2(
        keyinput_g10), .ZN(n4574) );
  OAI221_X1 U5081 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(DATAI_21_), .C2(
        keyinput_g10), .A(n4574), .ZN(n4577) );
  AOI22_X1 U5082 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput_g32), .ZN(n4575) );
  OAI221_X1 U5083 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_g32), .A(n4575), .ZN(n4576) );
  NOR4_X1 U5084 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4598)
         );
  AOI22_X1 U5085 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(REG3_REG_5__SCAN_IN), 
        .B2(keyinput_g47), .ZN(n4580) );
  OAI221_X1 U5086 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(REG3_REG_5__SCAN_IN), 
        .C2(keyinput_g47), .A(n4580), .ZN(n4587) );
  AOI22_X1 U5087 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_g59), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_g60), .ZN(n4581) );
  OAI221_X1 U5088 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_g59), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_g60), .A(n4581), .ZN(n4586) );
  AOI22_X1 U5089 ( .A1(DATAI_30_), .A2(keyinput_g1), .B1(DATAI_20_), .B2(
        keyinput_g11), .ZN(n4582) );
  OAI221_X1 U5090 ( .B1(DATAI_30_), .B2(keyinput_g1), .C1(DATAI_20_), .C2(
        keyinput_g11), .A(n4582), .ZN(n4585) );
  AOI22_X1 U5091 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_g46), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_g63), .ZN(n4583) );
  OAI221_X1 U5092 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_g63), .A(n4583), .ZN(n4584) );
  NOR4_X1 U5093 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4597)
         );
  AOI22_X1 U5094 ( .A1(DATAI_12_), .A2(keyinput_g19), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n4588) );
  OAI221_X1 U5095 ( .B1(DATAI_12_), .B2(keyinput_g19), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n4588), .ZN(n4595) );
  AOI22_X1 U5096 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .ZN(n4589) );
  OAI221_X1 U5097 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_g54), .A(n4589), .ZN(n4594) );
  AOI22_X1 U5098 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput_g56), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_g57), .ZN(n4590) );
  OAI221_X1 U5099 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_g56), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_g57), .A(n4590), .ZN(n4593) );
  AOI22_X1 U5100 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(IR_REG_6__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n4591) );
  OAI221_X1 U5101 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(IR_REG_6__SCAN_IN), 
        .C2(keyinput_g61), .A(n4591), .ZN(n4592) );
  NOR4_X1 U5102 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NAND4_X1 U5103 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4699)
         );
  AOI22_X1 U5104 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n4600) );
  OAI221_X1 U5105 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_25_), .C2(
        keyinput_f6), .A(n4600), .ZN(n4607) );
  AOI22_X1 U5106 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n4601) );
  OAI221_X1 U5107 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4601), .ZN(n4606) );
  AOI22_X1 U5108 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n4602) );
  OAI221_X1 U5109 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(REG3_REG_3__SCAN_IN), .C2(keyinput_f38), .A(n4602), .ZN(n4605) );
  AOI22_X1 U5110 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(DATAI_23_), .B2(
        keyinput_f8), .ZN(n4603) );
  OAI221_X1 U5111 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_23_), .C2(
        keyinput_f8), .A(n4603), .ZN(n4604) );
  NOR4_X1 U5112 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4637)
         );
  INV_X1 U5113 ( .A(DATAI_2_), .ZN(n4608) );
  XOR2_X1 U5114 ( .A(n4608), .B(keyinput_f29), .Z(n4616) );
  AOI22_X1 U5115 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(n4610), .B2(
        keyinput_f5), .ZN(n4609) );
  OAI221_X1 U5116 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(n4610), .C2(
        keyinput_f5), .A(n4609), .ZN(n4615) );
  AOI22_X1 U5117 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .ZN(n4611) );
  OAI221_X1 U5118 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4611), .ZN(n4614) );
  AOI22_X1 U5119 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n4612) );
  OAI221_X1 U5120 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n4612), .ZN(n4613) );
  NOR4_X1 U5121 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), .ZN(n4636)
         );
  AOI22_X1 U5122 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_f50), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_f60), .ZN(n4617) );
  OAI221_X1 U5123 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_f50), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_f60), .A(n4617), .ZN(n4625) );
  AOI22_X1 U5124 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_f57), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_f58), .ZN(n4619) );
  OAI221_X1 U5125 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_f57), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_f58), .A(n4619), .ZN(n4624) );
  AOI22_X1 U5126 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_f41), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4620) );
  OAI221_X1 U5127 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_f41), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4620), .ZN(n4623) );
  AOI22_X1 U5128 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .ZN(n4621) );
  OAI221_X1 U5129 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4621), .ZN(n4622) );
  NOR4_X1 U5130 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(n4635)
         );
  AOI22_X1 U5131 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .ZN(n4626) );
  OAI221_X1 U5132 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_f54), .A(n4626), .ZN(n4633) );
  AOI22_X1 U5133 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4627) );
  OAI221_X1 U5134 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4627), .ZN(n4632) );
  AOI22_X1 U5135 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(IR_REG_6__SCAN_IN), 
        .B2(keyinput_f61), .ZN(n4628) );
  OAI221_X1 U5136 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(IR_REG_6__SCAN_IN), 
        .C2(keyinput_f61), .A(n4628), .ZN(n4631) );
  AOI22_X1 U5137 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n4629) );
  OAI221_X1 U5138 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_f62), .A(n4629), .ZN(n4630) );
  NOR4_X1 U5139 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4634)
         );
  NAND4_X1 U5140 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4693)
         );
  AOI22_X1 U5141 ( .A1(n2627), .A2(keyinput_f3), .B1(keyinput_f20), .B2(n4639), 
        .ZN(n4638) );
  OAI221_X1 U5142 ( .B1(n2627), .B2(keyinput_f3), .C1(n4639), .C2(keyinput_f20), .A(n4638), .ZN(n4650) );
  AOI22_X1 U5143 ( .A1(n4642), .A2(keyinput_f1), .B1(n4641), .B2(keyinput_f16), 
        .ZN(n4640) );
  OAI221_X1 U5144 ( .B1(n4642), .B2(keyinput_f1), .C1(n4641), .C2(keyinput_f16), .A(n4640), .ZN(n4649) );
  XOR2_X1 U5145 ( .A(n4643), .B(keyinput_f2), .Z(n4647) );
  XNOR2_X1 U5146 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n4646) );
  XNOR2_X1 U5147 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_f37), .ZN(n4645) );
  XNOR2_X1 U5148 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4644) );
  NAND4_X1 U5149 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4648)
         );
  NOR3_X1 U5150 ( .A1(n4650), .A2(n4649), .A3(n4648), .ZN(n4691) );
  AOI22_X1 U5151 ( .A1(n2523), .A2(keyinput_f14), .B1(n4652), .B2(keyinput_f35), .ZN(n4651) );
  OAI221_X1 U5152 ( .B1(n2523), .B2(keyinput_f14), .C1(n4652), .C2(
        keyinput_f35), .A(n4651), .ZN(n4664) );
  AOI22_X1 U5153 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(n4654), .B2(
        keyinput_f49), .ZN(n4653) );
  OAI221_X1 U5154 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(n4654), .C2(
        keyinput_f49), .A(n4653), .ZN(n4663) );
  AOI22_X1 U5155 ( .A1(n4657), .A2(keyinput_f26), .B1(n4656), .B2(keyinput_f15), .ZN(n4655) );
  OAI221_X1 U5156 ( .B1(n4657), .B2(keyinput_f26), .C1(n4656), .C2(
        keyinput_f15), .A(n4655), .ZN(n4662) );
  AOI22_X1 U5157 ( .A1(n4660), .A2(keyinput_f33), .B1(keyinput_f22), .B2(n4659), .ZN(n4658) );
  OAI221_X1 U5158 ( .B1(n4660), .B2(keyinput_f33), .C1(n4659), .C2(
        keyinput_f22), .A(n4658), .ZN(n4661) );
  NOR4_X1 U5159 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), .ZN(n4690)
         );
  AOI22_X1 U5160 ( .A1(n4666), .A2(keyinput_f17), .B1(keyinput_f18), .B2(n2336), .ZN(n4665) );
  OAI221_X1 U5161 ( .B1(n4666), .B2(keyinput_f17), .C1(n2336), .C2(
        keyinput_f18), .A(n4665), .ZN(n4675) );
  AOI22_X1 U5162 ( .A1(n2513), .A2(keyinput_f48), .B1(n4668), .B2(keyinput_f45), .ZN(n4667) );
  OAI221_X1 U5163 ( .B1(n2513), .B2(keyinput_f48), .C1(n4668), .C2(
        keyinput_f45), .A(n4667), .ZN(n4674) );
  XOR2_X1 U5164 ( .A(n2484), .B(keyinput_f19), .Z(n4672) );
  XNOR2_X1 U5165 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4671) );
  XNOR2_X1 U5166 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_f39), .ZN(n4670) );
  XNOR2_X1 U5167 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n4669) );
  NAND4_X1 U5168 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4673)
         );
  NOR3_X1 U5169 ( .A1(n4675), .A2(n4674), .A3(n4673), .ZN(n4689) );
  AOI22_X1 U5170 ( .A1(n2434), .A2(keyinput_f23), .B1(n2383), .B2(keyinput_f47), .ZN(n4676) );
  OAI221_X1 U5171 ( .B1(n2434), .B2(keyinput_f23), .C1(n2383), .C2(
        keyinput_f47), .A(n4676), .ZN(n4687) );
  INV_X1 U5172 ( .A(DATAI_6_), .ZN(n4678) );
  AOI22_X1 U5173 ( .A1(n3738), .A2(keyinput_f43), .B1(keyinput_f25), .B2(n4678), .ZN(n4677) );
  OAI221_X1 U5174 ( .B1(n3738), .B2(keyinput_f43), .C1(n4678), .C2(
        keyinput_f25), .A(n4677), .ZN(n4686) );
  AOI22_X1 U5175 ( .A1(n4680), .A2(keyinput_f11), .B1(U3149), .B2(keyinput_f32), .ZN(n4679) );
  OAI221_X1 U5176 ( .B1(n4680), .B2(keyinput_f11), .C1(U3149), .C2(
        keyinput_f32), .A(n4679), .ZN(n4685) );
  XOR2_X1 U5177 ( .A(n4681), .B(keyinput_f4), .Z(n4683) );
  XNOR2_X1 U5178 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_f63), .ZN(n4682) );
  NAND2_X1 U5179 ( .A1(n4683), .A2(n4682), .ZN(n4684) );
  NOR4_X1 U5180 ( .A1(n4687), .A2(n4686), .A3(n4685), .A4(n4684), .ZN(n4688)
         );
  NAND4_X1 U5181 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4692)
         );
  OAI22_X1 U5182 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(n4693), .B2(n4692), 
        .ZN(n4695) );
  INV_X1 U5183 ( .A(keyinput_g24), .ZN(n4694) );
  NAND2_X1 U5184 ( .A1(n4695), .A2(n4694), .ZN(n4697) );
  OAI211_X1 U5185 ( .C1(n4695), .C2(keyinput_f24), .A(DATAI_7_), .B(
        keyinput_g24), .ZN(n4696) );
  OAI21_X1 U5186 ( .B1(DATAI_7_), .B2(n4697), .A(n4696), .ZN(n4698) );
  OAI21_X1 U5187 ( .B1(n4700), .B2(n4699), .A(n4698), .ZN(n4701) );
  XOR2_X1 U5188 ( .A(n4702), .B(n4701), .Z(U3352) );
endmodule

