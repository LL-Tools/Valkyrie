

module b20_C_AntiSAT_k_128_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157;

  INV_X1 U4852 ( .A(n6248), .ZN(n5707) );
  CLKBUF_X3 U4853 ( .A(n6308), .Z(n8261) );
  INV_X1 U4854 ( .A(n8056), .ZN(n8052) );
  AND2_X1 U4855 ( .A1(n6188), .A2(n8254), .ZN(n8246) );
  INV_X2 U4856 ( .A(n7975), .ZN(n8973) );
  INV_X1 U4858 ( .A(n6091), .ZN(n7059) );
  AND2_X1 U4859 ( .A1(n5078), .A2(n8270), .ZN(n5428) );
  NOR2_X1 U4860 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5193) );
  NAND2_X1 U4861 ( .A1(n9318), .A2(n4800), .ZN(n9304) );
  INV_X1 U4862 ( .A(n8977), .ZN(n7977) );
  NAND2_X1 U4863 ( .A1(n9333), .A2(n4802), .ZN(n9318) );
  INV_X1 U4864 ( .A(n8798), .ZN(n8604) );
  AND2_X1 U4865 ( .A1(n5634), .A2(n6258), .ZN(n9268) );
  NAND2_X1 U4866 ( .A1(n5438), .A2(n6373), .ZN(n5442) );
  INV_X1 U4867 ( .A(n5442), .ZN(n5457) );
  INV_X1 U4868 ( .A(n6934), .ZN(n9693) );
  BUF_X1 U4869 ( .A(n5438), .Z(n6397) );
  NAND2_X1 U4870 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U4871 ( .A1(n4889), .A2(n4890), .ZN(n4891) );
  NAND2_X2 U4872 ( .A1(n6133), .A2(n6134), .ZN(n5768) );
  INV_X1 U4873 ( .A(n8549), .ZN(n8478) );
  NOR2_X1 U4874 ( .A1(n9236), .A2(n9418), .ZN(n9457) );
  AOI21_X2 U4875 ( .B1(n5050), .B2(P1_IR_REG_29__SCAN_IN), .A(n5049), .ZN(
        n5078) );
  AND2_X1 U4876 ( .A1(n5738), .A2(n5739), .ZN(n4346) );
  AND4_X1 U4877 ( .A1(n5193), .A2(n5031), .A3(n5030), .A4(n5029), .ZN(n4347)
         );
  NAND2_X2 U4878 ( .A1(n5696), .A2(n5695), .ZN(n5438) );
  OAI21_X2 U4879 ( .B1(n8358), .B2(n4659), .A(n4658), .ZN(n4666) );
  NOR2_X2 U4880 ( .A1(n7507), .A2(n5864), .ZN(n7578) );
  NAND2_X2 U4881 ( .A1(n7637), .A2(n6225), .ZN(n6227) );
  OAI21_X2 U4882 ( .B1(n8947), .B2(n8950), .A(n8948), .ZN(n9036) );
  NOR2_X2 U4883 ( .A1(n9054), .A2(n7960), .ZN(n8947) );
  XNOR2_X1 U4884 ( .A(n5756), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9760) );
  NOR2_X2 U4885 ( .A1(n6850), .A2(n6940), .ZN(n6839) );
  OAI21_X2 U4886 ( .B1(n6380), .B2(n5442), .A(n4539), .ZN(n6940) );
  AND2_X1 U4887 ( .A1(n8791), .A2(n4416), .ZN(n4815) );
  XNOR2_X1 U4888 ( .A(n6244), .B(n6260), .ZN(n8289) );
  NOR3_X1 U4889 ( .A1(n8232), .A2(n8230), .A3(n8231), .ZN(n8238) );
  AND2_X1 U4890 ( .A1(n8298), .A2(n8350), .ZN(n8033) );
  OR4_X2 U4891 ( .A1(n8092), .A2(n8582), .A3(n8594), .A4(n8091), .ZN(n8094) );
  NOR2_X1 U4892 ( .A1(n4559), .A2(n8214), .ZN(n4555) );
  INV_X1 U4893 ( .A(n4558), .ZN(n4557) );
  INV_X1 U4894 ( .A(n8182), .ZN(n8643) );
  NAND2_X1 U4895 ( .A1(n7840), .A2(n4393), .ZN(n7839) );
  AOI21_X1 U4896 ( .B1(n7553), .B2(n6337), .A(n6336), .ZN(n7750) );
  OAI21_X1 U4897 ( .B1(n6993), .B2(n4740), .A(n4738), .ZN(n7204) );
  AND4_X2 U4898 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n8592)
         );
  AND4_X1 U4899 ( .A1(n7063), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n8581)
         );
  OR2_X1 U4900 ( .A1(n7453), .A2(n7235), .ZN(n7659) );
  NAND2_X1 U4901 ( .A1(n6076), .A2(n6075), .ZN(n8798) );
  CLKBUF_X2 U4902 ( .A(n8571), .Z(n4348) );
  NAND2_X1 U4903 ( .A1(n5263), .A2(n5262), .ZN(n7729) );
  XNOR2_X1 U4904 ( .A(n7021), .B(n8973), .ZN(n7247) );
  AND3_X1 U4905 ( .A1(n4498), .A2(P2_REG2_REG_7__SCAN_IN), .A3(n7272), .ZN(
        n7273) );
  NAND2_X1 U4906 ( .A1(n5326), .A2(n5325), .ZN(n9445) );
  AND2_X1 U4907 ( .A1(n4461), .A2(n4460), .ZN(n4934) );
  INV_X1 U4908 ( .A(n8429), .ZN(n7146) );
  NAND2_X2 U4909 ( .A1(n8104), .A2(n8099), .ZN(n8105) );
  NAND2_X1 U4910 ( .A1(n4680), .A2(n4487), .ZN(n8444) );
  INV_X1 U4911 ( .A(n8246), .ZN(n8227) );
  OR2_X1 U4912 ( .A1(n8431), .A2(n6979), .ZN(n8104) );
  INV_X1 U4913 ( .A(n6304), .ZN(n6984) );
  NAND4_X1 U4914 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n9130)
         );
  AND4_X1 U4915 ( .A1(n5765), .A2(n5764), .A3(n5762), .A4(n5763), .ZN(n7159)
         );
  INV_X2 U4916 ( .A(n4346), .ZN(n6090) );
  NAND2_X1 U4917 ( .A1(n5760), .A2(n5759), .ZN(n9812) );
  CLKBUF_X1 U4918 ( .A(n4346), .Z(n6070) );
  INV_X8 U4919 ( .A(n7984), .ZN(n8975) );
  INV_X4 U4921 ( .A(n7965), .ZN(n7984) );
  NAND2_X1 U4922 ( .A1(n4478), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6682) );
  MUX2_X1 U4923 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6104), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6105) );
  NAND2_X1 U4924 ( .A1(n5195), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U4925 ( .A1(n4370), .A2(n6680), .ZN(n6649) );
  OR2_X1 U4926 ( .A1(n7890), .A2(n4505), .ZN(n5733) );
  AND2_X1 U4927 ( .A1(n6100), .A2(n6107), .ZN(n6102) );
  NAND2_X1 U4928 ( .A1(n5734), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5748) );
  XNOR2_X1 U4929 ( .A(n4792), .B(n5037), .ZN(n5696) );
  NAND2_X1 U4930 ( .A1(n4353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U4931 ( .B1(n6373), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n4892), .ZN(
        n5439) );
  OR2_X1 U4932 ( .A1(n5701), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5699) );
  NAND4_X1 U4933 ( .A1(n4692), .A2(n4694), .A3(n4882), .A4(n4347), .ZN(n5701)
         );
  INV_X4 U4934 ( .A(n4891), .ZN(n6373) );
  AND2_X1 U4936 ( .A1(n5033), .A2(n5187), .ZN(n4692) );
  NOR2_X1 U4937 ( .A1(n4798), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4694) );
  AND2_X1 U4938 ( .A1(n4824), .A2(n4820), .ZN(n4819) );
  AND3_X1 U4939 ( .A1(n5032), .A2(n5188), .A3(n5189), .ZN(n5033) );
  AND2_X2 U4940 ( .A1(n5380), .A2(n5381), .ZN(n5187) );
  AND2_X1 U4941 ( .A1(n4507), .A2(n5718), .ZN(n4667) );
  AND2_X1 U4942 ( .A1(n5814), .A2(n5800), .ZN(n4824) );
  AND2_X1 U4943 ( .A1(n5721), .A2(n4677), .ZN(n4676) );
  INV_X1 U4944 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5946) );
  NOR2_X1 U4945 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5030) );
  INV_X1 U4946 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5718) );
  INV_X1 U4947 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5194) );
  NOR2_X1 U4948 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4542) );
  INV_X1 U4949 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5381) );
  INV_X4 U4950 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U4951 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  OAI21_X2 U4952 ( .B1(n7856), .B2(n5519), .A(n5595), .ZN(n9414) );
  NAND2_X2 U4953 ( .A1(n6480), .A2(n7435), .ZN(n6479) );
  XNOR2_X2 U4954 ( .A(n6587), .B(n6585), .ZN(n6614) );
  NOR2_X2 U4955 ( .A1(n9419), .A2(n9420), .ZN(n9417) );
  NOR2_X2 U4956 ( .A1(n4368), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5954) );
  OR2_X2 U4957 ( .A1(n5926), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4368) );
  NOR2_X2 U4958 ( .A1(n8958), .A2(n8962), .ZN(n9048) );
  NOR2_X2 U4959 ( .A1(n8959), .A2(n8960), .ZN(n8958) );
  OR2_X2 U4960 ( .A1(n6068), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n4369) );
  OR2_X2 U4961 ( .A1(n6090), .A2(n8578), .ZN(n6083) );
  NOR4_X2 U4962 ( .A1(n8233), .A2(n8247), .A3(n8094), .A4(n8093), .ZN(n8096)
         );
  NOR2_X1 U4963 ( .A1(n4755), .A2(n6237), .ZN(n4754) );
  INV_X1 U4964 ( .A(n4758), .ZN(n4755) );
  AND2_X1 U4965 ( .A1(n4627), .A2(n4460), .ZN(n4459) );
  OR2_X1 U4966 ( .A1(n9486), .A2(n7966), .ZN(n6254) );
  NAND2_X1 U4967 ( .A1(n7931), .A2(n7930), .ZN(n4727) );
  NAND2_X1 U4968 ( .A1(n8939), .A2(n5738), .ZN(n5779) );
  NAND2_X1 U4969 ( .A1(n4512), .A2(n4511), .ZN(n7762) );
  INV_X1 U4970 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5971) );
  AND2_X1 U4972 ( .A1(n5859), .A2(n5858), .ZN(n6332) );
  NOR2_X1 U4973 ( .A1(n9546), .A2(n9238), .ZN(n5706) );
  NAND2_X1 U4974 ( .A1(n5486), .A2(n5485), .ZN(n5688) );
  INV_X1 U4975 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5485) );
  AND2_X1 U4976 ( .A1(n5152), .A2(n5151), .ZN(n9058) );
  INV_X1 U4977 ( .A(n5430), .ZN(n5373) );
  XNOR2_X1 U4978 ( .A(n5359), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U4979 ( .A(n8517), .B(n8524), .ZN(n8500) );
  AND2_X1 U4980 ( .A1(n8732), .A2(n8166), .ZN(n4441) );
  AND2_X1 U4981 ( .A1(n4676), .A2(n5907), .ZN(n4675) );
  INV_X1 U4982 ( .A(n5217), .ZN(n4959) );
  INV_X1 U4983 ( .A(n4954), .ZN(n4457) );
  OR2_X1 U4984 ( .A1(n6701), .A2(n6745), .ZN(n4680) );
  OR2_X1 U4985 ( .A1(n6126), .A2(n8811), .ZN(n8207) );
  NOR2_X1 U4986 ( .A1(n8743), .A2(n4831), .ZN(n4830) );
  INV_X1 U4987 ( .A(n5920), .ZN(n4831) );
  AND2_X1 U4988 ( .A1(n5720), .A2(n4574), .ZN(n4573) );
  INV_X1 U4989 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5720) );
  AND2_X1 U4990 ( .A1(n9022), .A2(n9117), .ZN(n6228) );
  XNOR2_X1 U4991 ( .A(n5017), .B(n5016), .ZN(n5063) );
  OAI21_X1 U4992 ( .B1(n5163), .B2(n4849), .A(n4846), .ZN(n4992) );
  INV_X1 U4993 ( .A(n4850), .ZN(n4849) );
  AOI21_X1 U4994 ( .B1(n4850), .B2(n4848), .A(n4847), .ZN(n4846) );
  AOI21_X1 U4995 ( .B1(n4863), .B2(n4862), .A(n5258), .ZN(n4861) );
  OAI21_X1 U4996 ( .B1(n6373), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n4440), .ZN(
        n4918) );
  NAND2_X1 U4997 ( .A1(n6373), .A2(n6382), .ZN(n4440) );
  INV_X1 U4998 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U4999 ( .A1(n6701), .A2(n6745), .ZN(n8442) );
  NAND2_X1 U5000 ( .A1(n7506), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U5001 ( .A1(n4496), .A2(n7816), .ZN(n4492) );
  NOR2_X1 U5002 ( .A1(n8552), .A2(n8530), .ZN(n8533) );
  AND2_X1 U5003 ( .A1(n6079), .A2(n6078), .ZN(n8236) );
  AOI21_X1 U5004 ( .B1(n8599), .B2(n6065), .A(n4449), .ZN(n8587) );
  AND2_X1 U5005 ( .A1(n8799), .A2(n8588), .ZN(n4449) );
  AOI21_X1 U5006 ( .B1(n4557), .B2(n4555), .A(n8213), .ZN(n4554) );
  AOI22_X1 U5007 ( .A1(n8611), .A2(n8616), .B1(n8889), .B2(n8623), .ZN(n8599)
         );
  AOI21_X1 U5008 ( .B1(n4811), .B2(n4810), .A(n4809), .ZN(n8621) );
  NAND2_X1 U5009 ( .A1(n8897), .A2(n8818), .ZN(n4810) );
  AND2_X1 U5010 ( .A1(n8639), .A2(n8417), .ZN(n4809) );
  INV_X1 U5011 ( .A(n8633), .ZN(n4811) );
  OR2_X1 U5012 ( .A1(n8690), .A2(n6120), .ZN(n6123) );
  AND4_X1 U5013 ( .A1(n5942), .A2(n5941), .A3(n5940), .A4(n5939), .ZN(n8745)
         );
  AND4_X1 U5014 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n8746)
         );
  INV_X1 U5015 ( .A(n8055), .ZN(n5996) );
  NOR2_X1 U5016 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  NAND2_X1 U5017 ( .A1(n5788), .A2(n6982), .ZN(n4806) );
  NAND2_X1 U5018 ( .A1(n5768), .A2(n6376), .ZN(n8056) );
  NAND2_X1 U5019 ( .A1(n5748), .A2(n5735), .ZN(n5737) );
  INV_X1 U5020 ( .A(n6134), .ZN(n8549) );
  INV_X1 U5021 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4656) );
  AOI21_X1 U5022 ( .B1(n5984), .B2(n5973), .A(n4505), .ZN(n4657) );
  AND3_X1 U5023 ( .A1(n4823), .A2(n4819), .A3(n4574), .ZN(n5856) );
  NAND2_X1 U5024 ( .A1(n5073), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5167) );
  INV_X1 U5025 ( .A(n5178), .ZN(n5073) );
  NOR2_X1 U5026 ( .A1(n9026), .A2(n4737), .ZN(n4736) );
  NOR2_X1 U5027 ( .A1(n9016), .A2(n4350), .ZN(n4737) );
  AND4_X1 U5028 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n8965)
         );
  NOR2_X1 U5030 ( .A1(n9301), .A2(n4801), .ZN(n4800) );
  INV_X1 U5031 ( .A(n6254), .ZN(n4801) );
  AOI21_X1 U5032 ( .B1(n4754), .B2(n4760), .A(n4395), .ZN(n4752) );
  NAND2_X1 U5033 ( .A1(n4723), .A2(n4727), .ZN(n4719) );
  NAND2_X1 U5034 ( .A1(n4718), .A2(n4727), .ZN(n4717) );
  INV_X1 U5035 ( .A(n4721), .ZN(n4718) );
  AOI21_X1 U5036 ( .B1(n4723), .B2(n4722), .A(n4391), .ZN(n4721) );
  OR2_X1 U5037 ( .A1(n9532), .A2(n9118), .ZN(n6225) );
  NAND2_X1 U5038 ( .A1(n7039), .A2(n7206), .ZN(n4740) );
  NAND2_X1 U5039 ( .A1(n4739), .A2(n7206), .ZN(n4738) );
  INV_X1 U5040 ( .A(n4741), .ZN(n4739) );
  INV_X1 U5041 ( .A(n9344), .ZN(n9491) );
  INV_X1 U5042 ( .A(n6397), .ZN(n5459) );
  NAND2_X1 U5043 ( .A1(n4513), .A2(n4367), .ZN(n4512) );
  NAND2_X1 U5044 ( .A1(n8521), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U5045 ( .A1(n8519), .A2(n8521), .ZN(n4685) );
  NOR2_X1 U5046 ( .A1(n4470), .A2(n9797), .ZN(n4468) );
  NOR2_X1 U5047 ( .A1(n4471), .A2(n4474), .ZN(n4470) );
  NOR2_X1 U5048 ( .A1(n6099), .A2(n4366), .ZN(n4474) );
  OR2_X1 U5049 ( .A1(n6087), .A2(n4469), .ZN(n4467) );
  NAND2_X1 U5050 ( .A1(n4472), .A2(n8726), .ZN(n4469) );
  NAND2_X1 U5051 ( .A1(n4473), .A2(n8092), .ZN(n4472) );
  AOI21_X1 U5052 ( .B1(n5649), .B2(n6262), .A(n4356), .ZN(n4536) );
  NOR2_X1 U5053 ( .A1(n5553), .A2(n5707), .ZN(n4519) );
  NAND2_X1 U5054 ( .A1(n7037), .A2(n5707), .ZN(n4521) );
  NAND2_X1 U5055 ( .A1(n5553), .A2(n6248), .ZN(n4522) );
  NAND2_X1 U5056 ( .A1(n6998), .A2(n4517), .ZN(n4516) );
  NOR2_X1 U5057 ( .A1(n7037), .A2(n6248), .ZN(n4517) );
  NAND2_X1 U5058 ( .A1(n5599), .A2(n5676), .ZN(n4530) );
  AOI21_X1 U5059 ( .B1(n5599), .B2(n5598), .A(n5678), .ZN(n4532) );
  MUX2_X1 U5060 ( .A(n8203), .B(n8202), .S(n8227), .Z(n8209) );
  OAI22_X1 U5061 ( .A1(n5615), .A2(n9357), .B1(n5614), .B2(n6248), .ZN(n4534)
         );
  NAND2_X1 U5062 ( .A1(n8523), .A2(n4595), .ZN(n8529) );
  NAND2_X1 U5063 ( .A1(n8525), .A2(n8524), .ZN(n4595) );
  AND3_X1 U5064 ( .A1(n5907), .A2(n5946), .A3(n5973), .ZN(n5726) );
  INV_X1 U5065 ( .A(n5633), .ZN(n4527) );
  NAND2_X1 U5066 ( .A1(n4528), .A2(n5637), .ZN(n4524) );
  NAND2_X1 U5067 ( .A1(n6258), .A2(n6259), .ZN(n5635) );
  INV_X1 U5068 ( .A(n6258), .ZN(n4785) );
  NOR2_X1 U5069 ( .A1(n5455), .A2(n4422), .ZN(n4857) );
  INV_X1 U5070 ( .A(n5230), .ZN(n4956) );
  INV_X1 U5071 ( .A(SI_15_), .ZN(n4955) );
  NAND2_X1 U5072 ( .A1(n5283), .A2(n4944), .ZN(n4865) );
  NAND2_X1 U5073 ( .A1(n4614), .A2(n4392), .ZN(n4461) );
  NAND2_X1 U5074 ( .A1(n4647), .A2(n8588), .ZN(n4645) );
  AOI21_X1 U5075 ( .B1(n4660), .B2(n4665), .A(n4408), .ZN(n4658) );
  INV_X1 U5076 ( .A(n4660), .ZN(n4659) );
  NAND2_X1 U5077 ( .A1(n4633), .A2(n4632), .ZN(n9769) );
  INV_X1 U5078 ( .A(n9771), .ZN(n4633) );
  INV_X1 U5079 ( .A(n9772), .ZN(n4632) );
  NOR2_X1 U5080 ( .A1(n6699), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U5081 ( .A1(n8436), .A2(n4418), .ZN(n7287) );
  NAND2_X1 U5082 ( .A1(n7765), .A2(n7766), .ZN(n7817) );
  INV_X1 U5083 ( .A(n4414), .ZN(n4583) );
  XNOR2_X1 U5084 ( .A(n8817), .B(n8418), .ZN(n8182) );
  OR2_X1 U5085 ( .A1(n8908), .A2(n8656), .ZN(n8196) );
  OR2_X1 U5086 ( .A1(n8385), .A2(n8706), .ZN(n8189) );
  OR2_X1 U5087 ( .A1(n8708), .A2(n8716), .ZN(n8188) );
  INV_X1 U5088 ( .A(n6111), .ZN(n4545) );
  OR2_X1 U5089 ( .A1(n6549), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U5090 ( .A1(n6162), .A2(n6550), .ZN(n6195) );
  OR2_X1 U5091 ( .A1(n6549), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U5092 ( .A1(n6188), .A2(n8095), .ZN(n6300) );
  AND2_X1 U5093 ( .A1(n8165), .A2(n8164), .ZN(n8743) );
  OR2_X1 U5094 ( .A1(n6195), .A2(n6194), .ZN(n6975) );
  OR3_X1 U5095 ( .A1(n7864), .A2(n7872), .A3(n7810), .ZN(n6346) );
  INV_X1 U5096 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10039) );
  INV_X1 U5097 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U5098 ( .A1(n5722), .A2(n4827), .ZN(n6158) );
  NOR3_X1 U5099 ( .A1(n5727), .A2(n4351), .A3(P2_IR_REG_10__SCAN_IN), .ZN(
        n4827) );
  AND2_X1 U5100 ( .A1(n4675), .A2(n5948), .ZN(n4674) );
  INV_X2 U5101 ( .A(n5877), .ZN(n5722) );
  INV_X1 U5102 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4822) );
  OR2_X1 U5103 ( .A1(n7247), .A2(n4446), .ZN(n7181) );
  NAND2_X1 U5104 ( .A1(n4630), .A2(n7216), .ZN(n7219) );
  NAND2_X1 U5105 ( .A1(n7463), .A2(n8975), .ZN(n4630) );
  AOI21_X1 U5106 ( .B1(n4783), .B2(n4785), .A(n4782), .ZN(n4781) );
  INV_X1 U5107 ( .A(n6259), .ZN(n4782) );
  OR2_X1 U5108 ( .A1(n9258), .A2(n8978), .ZN(n5633) );
  OR2_X1 U5109 ( .A1(n9491), .A2(n9058), .ZN(n5618) );
  INV_X1 U5110 ( .A(n4789), .ZN(n4788) );
  NOR2_X1 U5111 ( .A1(n9400), .A2(n4790), .ZN(n4789) );
  INV_X1 U5112 ( .A(n5600), .ZN(n4790) );
  OR2_X1 U5113 ( .A1(n5241), .A2(n5224), .ZN(n5466) );
  AND2_X1 U5114 ( .A1(n6222), .A2(n4767), .ZN(n4766) );
  NAND2_X1 U5115 ( .A1(n4768), .A2(n4770), .ZN(n4767) );
  INV_X1 U5116 ( .A(n4771), .ZN(n4768) );
  OR2_X1 U5117 ( .A1(n7729), .A2(n7545), .ZN(n5666) );
  NAND2_X1 U5118 ( .A1(n5662), .A2(n7200), .ZN(n4797) );
  INV_X1 U5119 ( .A(n9432), .ZN(n4699) );
  CLKBUF_X1 U5120 ( .A(n6205), .Z(n7101) );
  INV_X1 U5121 ( .A(n9581), .ZN(n9420) );
  OR2_X1 U5122 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  OR2_X1 U5123 ( .A1(n5442), .A2(n6392), .ZN(n5443) );
  NOR2_X1 U5124 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5192) );
  NOR2_X1 U5125 ( .A1(n4948), .A2(n4867), .ZN(n4866) );
  INV_X1 U5126 ( .A(n4944), .ZN(n4867) );
  OAI21_X1 U5127 ( .B1(P1_RD_REG_SCAN_IN), .B2(P1_ADDR_REG_19__SCAN_IN), .A(
        n4886), .ZN(n4890) );
  INV_X1 U5128 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U5129 ( .A1(n4647), .A2(n8588), .ZN(n4646) );
  INV_X1 U5130 ( .A(n4645), .ZN(n4644) );
  INV_X1 U5131 ( .A(n4652), .ZN(n4651) );
  OAI21_X1 U5132 ( .B1(n4655), .B2(n4653), .A(n8388), .ZN(n4652) );
  NAND2_X1 U5133 ( .A1(n4642), .A2(n4644), .ZN(n4639) );
  AND2_X1 U5134 ( .A1(n8042), .A2(n4643), .ZN(n4642) );
  NAND2_X1 U5135 ( .A1(n4646), .A2(n4645), .ZN(n4643) );
  AND2_X1 U5136 ( .A1(n4364), .A2(n8012), .ZN(n4655) );
  NAND2_X1 U5137 ( .A1(n4364), .A2(n4415), .ZN(n4654) );
  OAI21_X1 U5138 ( .B1(n8333), .B2(n4653), .A(n4651), .ZN(n8386) );
  INV_X1 U5139 ( .A(n8428), .ZN(n7242) );
  NAND2_X1 U5140 ( .A1(n8245), .A2(n8780), .ZN(n4579) );
  NAND2_X1 U5141 ( .A1(n8248), .A2(n8249), .ZN(n4439) );
  NOR2_X1 U5142 ( .A1(n8247), .A2(n8095), .ZN(n4438) );
  NAND2_X1 U5143 ( .A1(n9774), .A2(n9775), .ZN(n9773) );
  NAND2_X1 U5144 ( .A1(n6682), .A2(n6680), .ZN(n6678) );
  XNOR2_X1 U5145 ( .A(n7287), .B(n4499), .ZN(n6760) );
  NAND2_X1 U5146 ( .A1(n6760), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7289) );
  NOR2_X1 U5147 ( .A1(n7279), .A2(n7280), .ZN(n7281) );
  OR2_X1 U5148 ( .A1(n7281), .A2(n7282), .ZN(n4592) );
  NAND2_X1 U5149 ( .A1(n7508), .A2(n4419), .ZN(n7583) );
  AND2_X1 U5150 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  NAND2_X1 U5151 ( .A1(n7734), .A2(n7678), .ZN(n7680) );
  NAND2_X1 U5152 ( .A1(n7680), .A2(n7679), .ZN(n7765) );
  XNOR2_X1 U5153 ( .A(n7817), .B(n7812), .ZN(n7767) );
  NAND2_X1 U5154 ( .A1(n4683), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5155 ( .A1(n4586), .A2(n4589), .ZN(n4585) );
  INV_X1 U5156 ( .A(n4587), .ZN(n4586) );
  AOI21_X1 U5157 ( .B1(n7772), .B2(n7773), .A(n4588), .ZN(n4587) );
  INV_X1 U5158 ( .A(n7829), .ZN(n4588) );
  OR2_X1 U5159 ( .A1(n4511), .A2(n4510), .ZN(n4509) );
  NAND2_X1 U5160 ( .A1(n4513), .A2(n4382), .ZN(n4508) );
  NOR2_X1 U5161 ( .A1(n8452), .A2(n4495), .ZN(n8469) );
  NOR2_X1 U5162 ( .A1(n7824), .A2(n7823), .ZN(n4495) );
  NAND2_X1 U5163 ( .A1(n8503), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8539) );
  INV_X1 U5164 ( .A(n8598), .ZN(n8605) );
  INV_X1 U5165 ( .A(n8632), .ZN(n4552) );
  AND2_X1 U5166 ( .A1(n8066), .A2(n8217), .ZN(n8598) );
  NAND2_X1 U5167 ( .A1(n4808), .A2(n6046), .ZN(n8611) );
  NAND2_X1 U5168 ( .A1(n8893), .A2(n8811), .ZN(n6046) );
  NAND2_X1 U5169 ( .A1(n8621), .A2(n4868), .ZN(n4808) );
  INV_X1 U5170 ( .A(n8208), .ZN(n4559) );
  OAI21_X1 U5171 ( .B1(n8208), .B2(n8204), .A(n8207), .ZN(n4558) );
  AND2_X1 U5172 ( .A1(n8207), .A2(n8205), .ZN(n8629) );
  OAI21_X1 U5173 ( .B1(n8642), .B2(n8643), .A(n8185), .ZN(n8632) );
  OAI22_X1 U5174 ( .A1(n8644), .A2(n8182), .B1(n8418), .B2(n8817), .ZN(n8633)
         );
  AOI21_X1 U5175 ( .B1(n6123), .B2(n4567), .A(n4566), .ZN(n8642) );
  OAI21_X1 U5176 ( .B1(n4568), .B2(n4569), .A(n8179), .ZN(n4566) );
  NOR2_X1 U5177 ( .A1(n4568), .A2(n4572), .ZN(n4567) );
  INV_X1 U5178 ( .A(n8200), .ZN(n4568) );
  AOI21_X1 U5179 ( .B1(n8655), .B2(n8654), .A(n6030), .ZN(n8644) );
  NOR2_X1 U5180 ( .A1(n8662), .A2(n6029), .ZN(n6030) );
  AND2_X1 U5181 ( .A1(n8196), .A2(n8195), .ZN(n4569) );
  NAND2_X1 U5182 ( .A1(n6123), .A2(n4571), .ZN(n4570) );
  BUF_X1 U5183 ( .A(n5804), .Z(n7058) );
  AND2_X1 U5184 ( .A1(n8195), .A2(n8192), .ZN(n8668) );
  INV_X1 U5185 ( .A(n8674), .ZN(n8706) );
  INV_X1 U5186 ( .A(n4564), .ZN(n4563) );
  OAI21_X1 U5187 ( .B1(n8168), .B2(n8190), .A(n8175), .ZN(n4564) );
  NAND2_X1 U5188 ( .A1(n5919), .A2(n5918), .ZN(n8762) );
  AND4_X1 U5189 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n8767)
         );
  OR2_X1 U5190 ( .A1(n9793), .A2(n9795), .ZN(n9791) );
  AND2_X1 U5191 ( .A1(n8112), .A2(n8118), .ZN(n8109) );
  AND2_X1 U5192 ( .A1(n6360), .A2(n8246), .ZN(n8728) );
  AND2_X1 U5193 ( .A1(n8117), .A2(n8111), .ZN(n6908) );
  NAND2_X1 U5194 ( .A1(n5770), .A2(n5769), .ZN(n6982) );
  INV_X1 U5195 ( .A(n8728), .ZN(n9794) );
  NAND2_X1 U5196 ( .A1(n6981), .A2(n6970), .ZN(n6969) );
  NAND2_X1 U5197 ( .A1(n7159), .A2(n8872), .ZN(n8070) );
  INV_X1 U5198 ( .A(n5779), .ZN(n5804) );
  OR2_X1 U5199 ( .A1(n6549), .A2(n6173), .ZN(n6973) );
  NAND2_X1 U5200 ( .A1(n5975), .A2(n5974), .ZN(n5983) );
  INV_X1 U5201 ( .A(n9813), .ZN(n9842) );
  NOR2_X1 U5202 ( .A1(n6191), .A2(n6180), .ZN(n6358) );
  NOR2_X1 U5203 ( .A1(n6975), .A2(n6180), .ZN(n6353) );
  AND2_X1 U5204 ( .A1(n6346), .A2(n6554), .ZN(n6974) );
  NAND2_X1 U5205 ( .A1(n4667), .A2(n4542), .ZN(n5799) );
  INV_X1 U5206 ( .A(n4596), .ZN(n4445) );
  INV_X1 U5207 ( .A(n6486), .ZN(n6570) );
  NAND2_X1 U5208 ( .A1(n5068), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U5209 ( .A1(n7050), .A2(n8970), .ZN(n4762) );
  AOI21_X1 U5210 ( .B1(n4736), .B2(n4350), .A(n4396), .ZN(n4735) );
  INV_X1 U5211 ( .A(n5464), .ZN(n5149) );
  AND2_X1 U5212 ( .A1(n5113), .A2(n5112), .ZN(n9294) );
  NAND2_X1 U5213 ( .A1(n4751), .A2(n4750), .ZN(n9300) );
  AOI21_X1 U5214 ( .B1(n4406), .B2(n4752), .A(n4359), .ZN(n4750) );
  AND2_X1 U5215 ( .A1(n9319), .A2(n6253), .ZN(n4802) );
  INV_X1 U5216 ( .A(n4754), .ZN(n4753) );
  AND2_X1 U5217 ( .A1(n6254), .A2(n5620), .ZN(n9319) );
  AOI21_X1 U5218 ( .B1(n4759), .B2(n6236), .A(n4403), .ZN(n4758) );
  NAND2_X1 U5219 ( .A1(n5520), .A2(n4789), .ZN(n9397) );
  NAND2_X1 U5220 ( .A1(n9414), .A2(n9413), .ZN(n5520) );
  OR2_X1 U5221 ( .A1(n9420), .A2(n8965), .ZN(n5600) );
  AOI21_X1 U5222 ( .B1(n4713), .B2(n4387), .A(n4714), .ZN(n9396) );
  AND2_X1 U5223 ( .A1(n5600), .A2(n5597), .ZN(n9413) );
  NAND2_X1 U5224 ( .A1(n7839), .A2(n5671), .ZN(n7856) );
  INV_X1 U5225 ( .A(n5519), .ZN(n7855) );
  NOR2_X1 U5226 ( .A1(n6228), .A2(n4726), .ZN(n4725) );
  INV_X1 U5227 ( .A(n4871), .ZN(n4726) );
  INV_X1 U5228 ( .A(n6228), .ZN(n4724) );
  NAND2_X1 U5229 ( .A1(n4772), .A2(n6219), .ZN(n4771) );
  NAND2_X1 U5230 ( .A1(n7463), .A2(n9122), .ZN(n4770) );
  AND2_X1 U5231 ( .A1(n7652), .A2(n5568), .ZN(n7495) );
  NAND2_X1 U5232 ( .A1(n5514), .A2(n4796), .ZN(n7455) );
  INV_X1 U5233 ( .A(n4797), .ZN(n4796) );
  AOI21_X1 U5234 ( .B1(n7039), .B2(n4742), .A(n4397), .ZN(n4741) );
  INV_X1 U5235 ( .A(n6215), .ZN(n4742) );
  NAND2_X1 U5236 ( .A1(n6209), .A2(n6964), .ZN(n6210) );
  NAND2_X1 U5237 ( .A1(n6875), .A2(n6208), .ZN(n4712) );
  NAND2_X1 U5238 ( .A1(n6582), .A2(n6207), .ZN(n6208) );
  XNOR2_X1 U5239 ( .A(n9131), .B(n6582), .ZN(n6881) );
  AND2_X1 U5240 ( .A1(n9720), .A2(n7435), .ZN(n9242) );
  NAND2_X1 U5241 ( .A1(n6600), .A2(n6599), .ZN(n9441) );
  NAND2_X1 U5242 ( .A1(n5239), .A2(n5238), .ZN(n9532) );
  INV_X1 U5243 ( .A(n5446), .ZN(n5460) );
  AND2_X1 U5244 ( .A1(n6248), .A2(n7435), .ZN(n9726) );
  OR2_X1 U5245 ( .A1(n6956), .A2(n6288), .ZN(n6293) );
  INV_X1 U5246 ( .A(n9391), .ZN(n9715) );
  AND2_X1 U5247 ( .A1(n6605), .A2(n6297), .ZN(n6600) );
  NAND2_X1 U5248 ( .A1(n6274), .A2(n6273), .ZN(n6591) );
  OAI21_X1 U5249 ( .B1(n5063), .B2(n5019), .A(n5018), .ZN(n5057) );
  OR2_X1 U5250 ( .A1(n5017), .A2(n5016), .ZN(n5018) );
  NAND2_X1 U5251 ( .A1(n5051), .A2(n5048), .ZN(n5049) );
  AND2_X1 U5252 ( .A1(n5044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U5253 ( .A1(n5047), .A2(n7886), .ZN(n5048) );
  OAI21_X1 U5254 ( .B1(n5004), .B2(n4837), .A(n4832), .ZN(n5085) );
  AND2_X1 U5255 ( .A1(n4833), .A2(n4835), .ZN(n4832) );
  NAND2_X1 U5256 ( .A1(n4434), .A2(n5098), .ZN(n4835) );
  NAND2_X1 U5257 ( .A1(n4836), .A2(n4834), .ZN(n4833) );
  AND2_X1 U5258 ( .A1(n5096), .A2(n5008), .ZN(n5107) );
  NOR2_X1 U5259 ( .A1(n5153), .A2(n4853), .ZN(n4852) );
  INV_X1 U5260 ( .A(n4980), .ZN(n4853) );
  AOI21_X1 U5261 ( .B1(n4852), .B2(n4981), .A(n4851), .ZN(n4850) );
  INV_X1 U5262 ( .A(n4986), .ZN(n4851) );
  NAND2_X1 U5263 ( .A1(n4978), .A2(n4977), .ZN(n5163) );
  OAI21_X1 U5264 ( .B1(n5171), .B2(n5172), .A(n4976), .ZN(n4978) );
  XNOR2_X1 U5265 ( .A(n5690), .B(n5689), .ZN(n6395) );
  INV_X1 U5266 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5689) );
  XNOR2_X1 U5267 ( .A(n5154), .B(n5153), .ZN(n7572) );
  OAI21_X1 U5268 ( .B1(n5163), .B2(n4981), .A(n4980), .ZN(n5154) );
  XNOR2_X1 U5269 ( .A(n5171), .B(n5174), .ZN(n7364) );
  AOI21_X1 U5270 ( .B1(n4453), .B2(n4454), .A(n4422), .ZN(n4452) );
  NAND2_X1 U5271 ( .A1(n5285), .A2(n4944), .ZN(n5271) );
  OAI21_X1 U5272 ( .B1(n4463), .B2(n4462), .A(n4928), .ZN(n5317) );
  NAND2_X1 U5273 ( .A1(n4616), .A2(n4376), .ZN(n4462) );
  INV_X1 U5274 ( .A(n4614), .ZN(n4463) );
  NOR2_X1 U5275 ( .A1(n4841), .A2(n4844), .ZN(n4447) );
  INV_X1 U5276 ( .A(n5370), .ZN(n4841) );
  AOI21_X1 U5277 ( .B1(n5413), .B2(n4843), .A(n4405), .ZN(n4842) );
  INV_X1 U5278 ( .A(n4917), .ZN(n4843) );
  XNOR2_X1 U5279 ( .A(n4915), .B(SI_5_), .ZN(n5370) );
  NAND2_X1 U5280 ( .A1(n4914), .A2(n4913), .ZN(n5371) );
  INV_X1 U5281 ( .A(n5768), .ZN(n6371) );
  NAND2_X1 U5282 ( .A1(n4669), .A2(n4668), .ZN(n8290) );
  OR2_X1 U5283 ( .A1(n4670), .A2(n8368), .ZN(n4668) );
  AOI21_X1 U5284 ( .B1(n4672), .B2(n4671), .A(n4433), .ZN(n4670) );
  OR2_X1 U5285 ( .A1(n8010), .A2(n8745), .ZN(n4874) );
  AND4_X1 U5286 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n8689)
         );
  INV_X1 U5287 ( .A(n10138), .ZN(n8400) );
  INV_X1 U5288 ( .A(n8818), .ZN(n8417) );
  INV_X1 U5289 ( .A(n7611), .ZN(n10122) );
  OR2_X1 U5290 ( .A1(n6090), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5782) );
  XNOR2_X1 U5291 ( .A(n6633), .B(n4590), .ZN(n9761) );
  NOR2_X1 U5292 ( .A1(n6702), .A2(n4436), .ZN(n6704) );
  NAND2_X1 U5293 ( .A1(n4482), .A2(n4479), .ZN(n7507) );
  NOR2_X1 U5294 ( .A1(n4481), .A2(n4690), .ZN(n4480) );
  OR2_X1 U5295 ( .A1(n7582), .A2(n7581), .ZN(n7669) );
  XNOR2_X1 U5296 ( .A(n7670), .B(n7742), .ZN(n7733) );
  OR2_X1 U5297 ( .A1(n7762), .A2(n7812), .ZN(n4682) );
  NAND2_X1 U5298 ( .A1(n7762), .A2(n4431), .ZN(n4681) );
  NOR2_X1 U5299 ( .A1(n8500), .A2(n8710), .ZN(n8518) );
  OAI21_X1 U5300 ( .B1(n8533), .B2(n4365), .A(n4594), .ZN(n4593) );
  AOI21_X1 U5301 ( .B1(n8555), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8536), .ZN(
        n4594) );
  INV_X1 U5302 ( .A(n9779), .ZN(n8542) );
  OR2_X1 U5303 ( .A1(n8567), .A2(n9778), .ZN(n4635) );
  AOI21_X1 U5304 ( .B1(n8566), .B2(n9788), .A(n8565), .ZN(n4634) );
  INV_X1 U5305 ( .A(n8236), .ZN(n8787) );
  AND2_X1 U5306 ( .A1(n6355), .A2(n6974), .ZN(n9804) );
  INV_X1 U5307 ( .A(n6354), .ZN(n6355) );
  INV_X1 U5308 ( .A(n8721), .ZN(n9802) );
  XNOR2_X1 U5309 ( .A(n8582), .B(n8577), .ZN(n4818) );
  AOI21_X1 U5310 ( .B1(n4815), .B2(n9797), .A(n9894), .ZN(n4813) );
  NOR2_X1 U5311 ( .A1(n4373), .A2(n6143), .ZN(n4465) );
  AND2_X1 U5312 ( .A1(n5751), .A2(n5750), .ZN(n8897) );
  OR2_X1 U5313 ( .A1(n9878), .A2(n9865), .ZN(n8935) );
  NOR2_X1 U5314 ( .A1(n4609), .A2(n7996), .ZN(n4608) );
  INV_X1 U5315 ( .A(n7983), .ZN(n4609) );
  NAND2_X1 U5316 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  INV_X1 U5317 ( .A(n7997), .ZN(n4606) );
  INV_X1 U5318 ( .A(n7996), .ZN(n4607) );
  NAND2_X1 U5319 ( .A1(n9278), .A2(n9088), .ZN(n4610) );
  NAND2_X1 U5320 ( .A1(n4613), .A2(n7917), .ZN(n4612) );
  INV_X1 U5321 ( .A(n9386), .ZN(n9505) );
  INV_X1 U5322 ( .A(n5709), .ZN(n5714) );
  NAND2_X1 U5323 ( .A1(n4839), .A2(n6597), .ZN(n4535) );
  NAND2_X1 U5324 ( .A1(n5650), .A2(n9699), .ZN(n4839) );
  AND2_X1 U5325 ( .A1(n5487), .A2(n5688), .ZN(n6478) );
  AND3_X1 U5326 ( .A1(n5170), .A2(n5169), .A3(n5168), .ZN(n9057) );
  INV_X1 U5327 ( .A(n7947), .ZN(n9113) );
  AND2_X1 U5328 ( .A1(n5143), .A2(n5142), .ZN(n9344) );
  NOR2_X1 U5329 ( .A1(n6293), .A2(n6953), .ZN(n9509) );
  OR2_X1 U5330 ( .A1(n5043), .A2(n5459), .ZN(n9546) );
  AND3_X1 U5331 ( .A1(n5349), .A2(n5348), .A3(n5347), .ZN(n7096) );
  NAND2_X1 U5332 ( .A1(n9738), .A2(n9722), .ZN(n9586) );
  OR2_X1 U5333 ( .A1(n6395), .A2(P1_U3086), .ZN(n7621) );
  CLKBUF_X1 U5334 ( .A(n6480), .Z(n9699) );
  AND2_X1 U5335 ( .A1(n4518), .A2(n4516), .ZN(n4515) );
  NAND2_X1 U5336 ( .A1(n4520), .A2(n4519), .ZN(n4518) );
  MUX2_X1 U5337 ( .A(n8131), .B(n8130), .S(n8227), .Z(n8140) );
  OAI21_X1 U5338 ( .B1(n8174), .B2(n8173), .A(n8172), .ZN(n8191) );
  NAND2_X1 U5339 ( .A1(n4531), .A2(n4529), .ZN(n5613) );
  OAI21_X1 U5340 ( .B1(n4532), .B2(n5602), .A(n5707), .ZN(n4531) );
  AOI21_X1 U5341 ( .B1(n4530), .B2(n4386), .A(n4354), .ZN(n4529) );
  OAI21_X1 U5342 ( .B1(n4533), .B2(n5619), .A(n5621), .ZN(n5631) );
  AOI21_X1 U5343 ( .B1(n4534), .B2(n5618), .A(n5617), .ZN(n4533) );
  NOR2_X1 U5344 ( .A1(n4380), .A2(n4352), .ZN(n4525) );
  NAND2_X1 U5345 ( .A1(n8088), .A2(n4476), .ZN(n6012) );
  INV_X1 U5346 ( .A(n7899), .ZN(n4476) );
  INV_X1 U5347 ( .A(n4852), .ZN(n4848) );
  INV_X1 U5348 ( .A(n5140), .ZN(n4847) );
  INV_X1 U5349 ( .A(SI_17_), .ZN(n4960) );
  INV_X1 U5350 ( .A(n4866), .ZN(n4862) );
  NAND2_X1 U5351 ( .A1(n4879), .A2(n4464), .ZN(n4460) );
  INV_X1 U5352 ( .A(n4928), .ZN(n4464) );
  INV_X1 U5353 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4887) );
  INV_X1 U5354 ( .A(n7828), .ZN(n4589) );
  INV_X1 U5355 ( .A(n7673), .ZN(n4511) );
  INV_X1 U5356 ( .A(n7761), .ZN(n4510) );
  NAND2_X1 U5357 ( .A1(n8455), .A2(n8456), .ZN(n8488) );
  INV_X1 U5358 ( .A(n8529), .ZN(n8526) );
  OR2_X1 U5359 ( .A1(n6098), .A2(n8581), .ZN(n8241) );
  AND2_X1 U5360 ( .A1(n8048), .A2(n8798), .ZN(n8222) );
  AND2_X1 U5361 ( .A1(n6012), .A2(n8717), .ZN(n6011) );
  NAND2_X1 U5362 ( .A1(n8667), .A2(n8672), .ZN(n4477) );
  NOR2_X1 U5363 ( .A1(n8190), .A2(n4562), .ZN(n4561) );
  INV_X1 U5364 ( .A(n8169), .ZN(n4562) );
  NAND2_X1 U5365 ( .A1(n5793), .A2(n4412), .ZN(n4803) );
  NAND2_X1 U5366 ( .A1(n6304), .A2(n9812), .ZN(n8071) );
  OR2_X1 U5367 ( .A1(n7563), .A2(n7562), .ZN(n7566) );
  INV_X1 U5368 ( .A(n6973), .ZN(n6180) );
  NAND2_X1 U5369 ( .A1(n6158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U5370 ( .A1(n6145), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6175) );
  INV_X1 U5371 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6174) );
  INV_X1 U5372 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5947) );
  AND2_X1 U5373 ( .A1(n5722), .A2(n4675), .ZN(n5949) );
  INV_X1 U5374 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4677) );
  NOR2_X1 U5375 ( .A1(n4736), .A2(n7939), .ZN(n4732) );
  NOR2_X1 U5376 ( .A1(n7938), .A2(n7937), .ZN(n4731) );
  INV_X1 U5377 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5310) );
  OR2_X1 U5378 ( .A1(n8997), .A2(n4621), .ZN(n4620) );
  INV_X1 U5379 ( .A(n4877), .ZN(n4621) );
  NAND2_X1 U5380 ( .A1(n5637), .A2(n4527), .ZN(n4526) );
  INV_X1 U5381 ( .A(n5635), .ZN(n5624) );
  NOR2_X1 U5382 ( .A1(n9505), .A2(n9512), .ZN(n4705) );
  INV_X1 U5383 ( .A(n6229), .ZN(n4715) );
  INV_X1 U5384 ( .A(n4719), .ZN(n4716) );
  INV_X1 U5385 ( .A(n4725), .ZN(n4722) );
  INV_X1 U5386 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U5387 ( .A1(n4711), .A2(n9106), .ZN(n4710) );
  NOR2_X1 U5388 ( .A1(n9538), .A2(n7729), .ZN(n4711) );
  OR2_X1 U5389 ( .A1(n5329), .A2(n5310), .ZN(n5312) );
  NOR2_X1 U5390 ( .A1(n9445), .A2(n9679), .ZN(n4700) );
  NOR2_X1 U5391 ( .A1(n7112), .A2(n7050), .ZN(n6860) );
  NAND2_X1 U5392 ( .A1(n9291), .A2(n9558), .ZN(n9275) );
  AND2_X1 U5393 ( .A1(n9308), .A2(n9562), .ZN(n9291) );
  AND2_X1 U5394 ( .A1(n9329), .A2(n9339), .ZN(n9323) );
  AND2_X1 U5395 ( .A1(n9344), .A2(n9348), .ZN(n9339) );
  NOR2_X1 U5396 ( .A1(n7659), .A2(n7729), .ZN(n7713) );
  NAND2_X1 U5397 ( .A1(n5015), .A2(n5014), .ZN(n5017) );
  INV_X1 U5398 ( .A(n5003), .ZN(n4834) );
  NAND2_X1 U5399 ( .A1(n5034), .A2(n4799), .ZN(n4798) );
  INV_X1 U5400 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4799) );
  AND2_X1 U5401 ( .A1(n5003), .A2(n5002), .ZN(n5120) );
  AND2_X1 U5402 ( .A1(n4997), .A2(n4996), .ZN(n5129) );
  INV_X1 U5403 ( .A(SI_20_), .ZN(n5172) );
  INV_X1 U5404 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U5405 ( .A1(n4859), .A2(n4967), .ZN(n5186) );
  NAND2_X1 U5406 ( .A1(n4854), .A2(n4417), .ZN(n4859) );
  AOI21_X1 U5407 ( .B1(n4858), .B2(n4857), .A(n4856), .ZN(n4855) );
  INV_X1 U5408 ( .A(n4964), .ZN(n4856) );
  AOI21_X1 U5409 ( .B1(n5246), .B2(n4456), .A(n4424), .ZN(n4454) );
  NOR2_X1 U5410 ( .A1(n4456), .A2(n4858), .ZN(n4453) );
  INV_X1 U5411 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4958) );
  NOR2_X1 U5412 ( .A1(n4939), .A2(n4628), .ZN(n4627) );
  INV_X1 U5413 ( .A(n4933), .ZN(n4628) );
  NAND2_X1 U5414 ( .A1(n4626), .A2(n4625), .ZN(n5285) );
  NOR2_X1 U5415 ( .A1(n5283), .A2(n4624), .ZN(n4625) );
  NOR2_X2 U5416 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5380) );
  OAI21_X1 U5417 ( .B1(n6376), .B2(n4538), .A(n4537), .ZN(n4904) );
  NAND2_X1 U5418 ( .A1(n4891), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4537) );
  OR2_X1 U5419 ( .A1(n4891), .A2(n4894), .ZN(n4895) );
  XNOR2_X1 U5420 ( .A(n8261), .B(n7170), .ZN(n6318) );
  NOR2_X1 U5421 ( .A1(n5988), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5976) );
  NOR2_X1 U5422 ( .A1(n8004), .A2(n8423), .ZN(n4672) );
  NAND2_X1 U5423 ( .A1(n8004), .A2(n8423), .ZN(n4671) );
  NOR2_X1 U5424 ( .A1(n8377), .A2(n4661), .ZN(n4660) );
  INV_X1 U5425 ( .A(n4662), .ZN(n4661) );
  NAND2_X1 U5426 ( .A1(n8023), .A2(n8314), .ZN(n4662) );
  NAND2_X1 U5427 ( .A1(n8358), .A2(n4664), .ZN(n4663) );
  XNOR2_X1 U5428 ( .A(n6308), .B(n9812), .ZN(n6305) );
  OR2_X1 U5429 ( .A1(n6000), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5988) );
  OR2_X1 U5430 ( .A1(n6057), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6068) );
  AND2_X1 U5431 ( .A1(n6361), .A2(n6360), .ZN(n8409) );
  NAND2_X1 U5432 ( .A1(n6156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U5433 ( .A1(n4500), .A2(n4503), .ZN(n9775) );
  NAND2_X1 U5434 ( .A1(n6658), .A2(n6642), .ZN(n4500) );
  NAND2_X1 U5435 ( .A1(n9769), .A2(n4390), .ZN(n6672) );
  NAND2_X1 U5436 ( .A1(n4680), .A2(n8442), .ZN(n4679) );
  OAI21_X1 U5437 ( .B1(n6700), .B2(n4486), .A(n4484), .ZN(n4488) );
  NOR2_X1 U5438 ( .A1(n4485), .A2(n6703), .ZN(n4484) );
  NAND2_X1 U5439 ( .A1(n7289), .A2(n7290), .ZN(n7293) );
  NAND2_X1 U5440 ( .A1(n7514), .A2(n7515), .ZN(n7596) );
  NAND2_X1 U5441 ( .A1(n4592), .A2(n4591), .ZN(n7514) );
  INV_X1 U5442 ( .A(n7513), .ZN(n4591) );
  NAND2_X1 U5443 ( .A1(n7584), .A2(n7585), .ZN(n7587) );
  OAI21_X1 U5444 ( .B1(n7774), .B2(n7773), .A(n7772), .ZN(n7830) );
  NAND2_X1 U5445 ( .A1(n7819), .A2(n7820), .ZN(n7822) );
  NAND2_X1 U5446 ( .A1(n7822), .A2(n7821), .ZN(n8455) );
  INV_X1 U5447 ( .A(n4582), .ZN(n4581) );
  AOI21_X1 U5448 ( .B1(n4362), .B2(n4583), .A(n8459), .ZN(n4582) );
  NAND2_X1 U5449 ( .A1(n7774), .A2(n4414), .ZN(n4584) );
  XNOR2_X1 U5450 ( .A(n8488), .B(n8477), .ZN(n8457) );
  NAND2_X1 U5451 ( .A1(n8492), .A2(n8493), .ZN(n8501) );
  NAND2_X1 U5452 ( .A1(n8507), .A2(n8508), .ZN(n8523) );
  AOI21_X1 U5453 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8499), .A(n8498), .ZN(
        n8517) );
  XNOR2_X1 U5454 ( .A(n8537), .B(n8524), .ZN(n8503) );
  NAND2_X1 U5455 ( .A1(n8501), .A2(n4631), .ZN(n8537) );
  NAND2_X1 U5456 ( .A1(n8499), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4631) );
  INV_X1 U5457 ( .A(n4473), .ZN(n4471) );
  NAND2_X1 U5458 ( .A1(n6099), .A2(n4366), .ZN(n4473) );
  NAND2_X1 U5459 ( .A1(n4548), .A2(n4549), .ZN(n8593) );
  AOI21_X1 U5460 ( .B1(n4349), .B2(n4556), .A(n8218), .ZN(n4549) );
  OR2_X1 U5461 ( .A1(n8222), .A2(n8223), .ZN(n8594) );
  OR2_X1 U5462 ( .A1(n8184), .A2(n8626), .ZN(n8634) );
  NAND2_X1 U5463 ( .A1(n4477), .A2(n6014), .ZN(n7899) );
  INV_X1 U5464 ( .A(n4477), .ZN(n8669) );
  NAND2_X1 U5465 ( .A1(n8692), .A2(n8188), .ZN(n8707) );
  INV_X1 U5466 ( .A(n8163), .ZN(n8732) );
  AND2_X1 U5467 ( .A1(n8160), .A2(n8159), .ZN(n8772) );
  OR2_X1 U5468 ( .A1(n5888), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U5469 ( .A1(n5898), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U5470 ( .A1(n9791), .A2(n4575), .ZN(n6113) );
  AND2_X1 U5471 ( .A1(n4880), .A2(n8134), .ZN(n4575) );
  OR2_X1 U5472 ( .A1(n5871), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5888) );
  AOI21_X1 U5473 ( .B1(n7562), .B2(n5855), .A(n4400), .ZN(n4826) );
  NAND2_X1 U5474 ( .A1(n7566), .A2(n5855), .ZN(n9796) );
  AND2_X1 U5475 ( .A1(n5844), .A2(n7276), .ZN(n5862) );
  NOR2_X1 U5476 ( .A1(n5833), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5844) );
  AND4_X1 U5477 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n10130)
         );
  OR2_X1 U5478 ( .A1(n5820), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5833) );
  AOI21_X1 U5479 ( .B1(n4545), .B2(n8119), .A(n4544), .ZN(n4543) );
  INV_X1 U5480 ( .A(n8122), .ZN(n4544) );
  NAND2_X1 U5481 ( .A1(n4804), .A2(n4805), .ZN(n7346) );
  AND2_X1 U5482 ( .A1(n4803), .A2(n4381), .ZN(n4804) );
  NOR2_X1 U5483 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5807) );
  INV_X1 U5484 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5806) );
  OR2_X1 U5485 ( .A1(n6090), .A2(n6949), .ZN(n5795) );
  OAI21_X1 U5486 ( .B1(n7157), .B2(n8070), .A(n8068), .ZN(n6970) );
  NAND2_X1 U5487 ( .A1(n8071), .A2(n8068), .ZN(n7157) );
  NAND2_X1 U5488 ( .A1(n6977), .A2(n6976), .ZN(n7139) );
  AND4_X1 U5489 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n6976)
         );
  AOI21_X1 U5490 ( .B1(n8587), .B2(n6077), .A(n4448), .ZN(n8576) );
  NOR2_X1 U5491 ( .A1(n8794), .A2(n8798), .ZN(n4448) );
  OR2_X1 U5492 ( .A1(n9859), .A2(n6188), .ZN(n6354) );
  NAND2_X1 U5493 ( .A1(n5986), .A2(n5985), .ZN(n8385) );
  NAND2_X1 U5494 ( .A1(n8762), .A2(n5920), .ZN(n8744) );
  OR2_X1 U5495 ( .A1(n6989), .A2(n8254), .ZN(n9859) );
  NAND2_X1 U5496 ( .A1(n6141), .A2(n8246), .ZN(n9813) );
  AND2_X1 U5497 ( .A1(n9859), .A2(n7615), .ZN(n9872) );
  NAND2_X1 U5498 ( .A1(n6160), .A2(n6161), .ZN(n6549) );
  NOR3_X1 U5499 ( .A1(n5727), .A2(n4351), .A3(n4829), .ZN(n4828) );
  NAND2_X1 U5500 ( .A1(n5721), .A2(n10039), .ZN(n4829) );
  INV_X1 U5501 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5736) );
  INV_X1 U5502 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5747) );
  INV_X1 U5503 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U5504 ( .A1(n6146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U5505 ( .A1(n6175), .A2(n6174), .ZN(n6146) );
  INV_X1 U5506 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U5507 ( .A1(n6148), .A2(n6153), .ZN(n6150) );
  NAND2_X1 U5508 ( .A1(n6102), .A2(n6101), .ZN(n6156) );
  INV_X1 U5509 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6101) );
  INV_X1 U5510 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6107) );
  AND2_X1 U5511 ( .A1(n4822), .A2(n5719), .ZN(n4820) );
  AND2_X1 U5512 ( .A1(n4824), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U5513 ( .A1(n4505), .A2(n4507), .ZN(n4504) );
  OR2_X1 U5514 ( .A1(n4541), .A2(n4506), .ZN(n4501) );
  NAND2_X1 U5515 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4506) );
  NAND2_X1 U5516 ( .A1(n7544), .A2(n7542), .ZN(n7539) );
  OAI21_X1 U5517 ( .B1(n9015), .B2(n4733), .A(n4730), .ZN(n8959) );
  NAND2_X1 U5518 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  AOI21_X1 U5519 ( .B1(n4732), .B2(n4735), .A(n4731), .ZN(n4730) );
  INV_X1 U5520 ( .A(n7939), .ZN(n4734) );
  INV_X1 U5521 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5327) );
  OR2_X1 U5522 ( .A1(n5336), .A2(n5327), .ZN(n5329) );
  AND2_X1 U5523 ( .A1(n4746), .A2(n7185), .ZN(n4745) );
  INV_X1 U5524 ( .A(n7224), .ZN(n4746) );
  NAND2_X1 U5525 ( .A1(n7019), .A2(n4375), .ZN(n4747) );
  NAND2_X1 U5526 ( .A1(n6570), .A2(n6487), .ZN(n6492) );
  INV_X1 U5527 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U5528 ( .A1(n5069), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5278) );
  INV_X1 U5529 ( .A(n5293), .ZN(n5069) );
  INV_X1 U5530 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7393) );
  INV_X1 U5531 ( .A(n7219), .ZN(n7308) );
  OR2_X1 U5532 ( .A1(n5305), .A2(n7314), .ZN(n5293) );
  INV_X1 U5533 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7314) );
  OAI21_X1 U5534 ( .B1(n7971), .B2(n9724), .A(n6573), .ZN(n6574) );
  NAND2_X1 U5535 ( .A1(n9035), .A2(n7970), .ZN(n9005) );
  NAND2_X1 U5536 ( .A1(n5070), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5241) );
  INV_X1 U5537 ( .A(n5685), .ZN(n5711) );
  NOR4_X1 U5538 ( .A1(n5483), .A2(n5523), .A3(n5685), .A4(n5482), .ZN(n5648)
         );
  AND2_X1 U5539 ( .A1(n9546), .A2(n9238), .ZN(n5685) );
  NOR2_X1 U5540 ( .A1(n5184), .A2(n5183), .ZN(n7947) );
  AND4_X1 U5541 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n7545)
         );
  AND4_X1 U5542 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n9123)
         );
  AND4_X1 U5543 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n7192)
         );
  AND4_X1 U5544 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n6830)
         );
  AND2_X1 U5545 ( .A1(n6260), .A2(n4783), .ZN(n4777) );
  OAI21_X1 U5546 ( .B1(n6260), .B2(n4358), .A(n4779), .ZN(n4778) );
  NAND2_X1 U5547 ( .A1(n6260), .A2(n4781), .ZN(n4779) );
  NAND2_X1 U5548 ( .A1(n6261), .A2(n4781), .ZN(n4780) );
  AND2_X1 U5549 ( .A1(n5628), .A2(n6256), .ZN(n9286) );
  AND2_X1 U5550 ( .A1(n5124), .A2(n5123), .ZN(n9311) );
  NAND2_X1 U5551 ( .A1(n9318), .A2(n6254), .ZN(n9302) );
  NAND2_X1 U5552 ( .A1(n5074), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5158) );
  OR2_X1 U5553 ( .A1(n5158), .A2(n8953), .ZN(n5145) );
  AND2_X1 U5554 ( .A1(n6249), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U5555 ( .A1(n4788), .A2(n5677), .ZN(n4787) );
  AND2_X1 U5556 ( .A1(n9417), .A2(n4702), .ZN(n9348) );
  NOR2_X1 U5557 ( .A1(n4704), .A2(n9349), .ZN(n4702) );
  NAND2_X1 U5558 ( .A1(n9397), .A2(n5677), .ZN(n9389) );
  NAND2_X1 U5559 ( .A1(n9417), .A2(n9409), .ZN(n9403) );
  NAND2_X1 U5560 ( .A1(n9417), .A2(n4705), .ZN(n9381) );
  NAND2_X1 U5561 ( .A1(n5071), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5468) );
  INV_X1 U5562 ( .A(n5466), .ZN(n5071) );
  NOR2_X1 U5563 ( .A1(n7659), .A2(n4709), .ZN(n7714) );
  INV_X1 U5564 ( .A(n4711), .ZN(n4709) );
  OR2_X1 U5565 ( .A1(n5278), .A2(n7393), .ZN(n5265) );
  OR2_X1 U5566 ( .A1(n5265), .A2(n5251), .ZN(n5253) );
  AOI21_X1 U5567 ( .B1(n4766), .B2(n4769), .A(n4394), .ZN(n4764) );
  INV_X1 U5568 ( .A(n4770), .ZN(n4769) );
  INV_X1 U5569 ( .A(n5557), .ZN(n4795) );
  AND2_X1 U5570 ( .A1(n7083), .A2(n4696), .ZN(n7452) );
  NOR2_X1 U5571 ( .A1(n7264), .A2(n4698), .ZN(n4696) );
  NAND2_X1 U5572 ( .A1(n7083), .A2(n4700), .ZN(n7032) );
  OR2_X1 U5573 ( .A1(n5404), .A2(n6813), .ZN(n5336) );
  NAND2_X1 U5574 ( .A1(n7083), .A2(n7096), .ZN(n7084) );
  OR2_X1 U5575 ( .A1(n6861), .A2(n6937), .ZN(n6850) );
  NAND2_X1 U5576 ( .A1(n9724), .A2(n6206), .ZN(n4775) );
  NAND2_X1 U5577 ( .A1(n5504), .A2(n5503), .ZN(n6883) );
  NAND2_X1 U5578 ( .A1(n9724), .A2(n7113), .ZN(n7112) );
  CLKBUF_X1 U5579 ( .A(n7101), .Z(n7109) );
  INV_X1 U5580 ( .A(n9080), .ZN(n9069) );
  NAND2_X1 U5581 ( .A1(n5059), .A2(n5058), .ZN(n5642) );
  NAND2_X1 U5582 ( .A1(n5065), .A2(n5064), .ZN(n6291) );
  NAND2_X1 U5583 ( .A1(n5131), .A2(n5130), .ZN(n9486) );
  AND2_X1 U5584 ( .A1(n7574), .A2(n7490), .ZN(n9720) );
  NOR2_X1 U5585 ( .A1(n9446), .A2(n9726), .ZN(n9716) );
  XNOR2_X1 U5586 ( .A(n5057), .B(n5056), .ZN(n8269) );
  XNOR2_X1 U5587 ( .A(n5700), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U5588 ( .A1(n5699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5700) );
  XNOR2_X1 U5589 ( .A(n5702), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6271) );
  XNOR2_X1 U5590 ( .A(n5186), .B(n5185), .ZN(n7154) );
  NAND2_X1 U5591 ( .A1(n4444), .A2(n4377), .ZN(n5220) );
  INV_X1 U5592 ( .A(n5322), .ZN(n4444) );
  NAND2_X1 U5593 ( .A1(n4458), .A2(n4954), .ZN(n5232) );
  NAND2_X1 U5594 ( .A1(n5247), .A2(n4952), .ZN(n4458) );
  NAND2_X1 U5595 ( .A1(n4860), .A2(n4863), .ZN(n5259) );
  NAND2_X1 U5596 ( .A1(n5285), .A2(n4629), .ZN(n6411) );
  OAI21_X1 U5597 ( .B1(n4934), .B2(n4624), .A(n4622), .ZN(n4629) );
  INV_X1 U5598 ( .A(n4623), .ZN(n4622) );
  OAI21_X1 U5599 ( .B1(n4627), .B2(n4624), .A(n5283), .ZN(n4623) );
  NAND2_X1 U5600 ( .A1(n4615), .A2(n5371), .ZN(n4614) );
  AND2_X1 U5601 ( .A1(n4447), .A2(n5341), .ZN(n4615) );
  INV_X1 U5602 ( .A(n4617), .ZN(n4616) );
  OAI21_X1 U5603 ( .B1(n4842), .B2(n4618), .A(n4922), .ZN(n4617) );
  XNOR2_X1 U5604 ( .A(n4907), .B(SI_3_), .ZN(n5378) );
  INV_X1 U5605 ( .A(n4640), .ZN(n8043) );
  INV_X1 U5606 ( .A(n4646), .ZN(n4641) );
  OAI21_X1 U5607 ( .B1(n8396), .B2(n4644), .A(n4642), .ZN(n8260) );
  NAND2_X1 U5608 ( .A1(n6313), .A2(n6312), .ZN(n6821) );
  AOI21_X1 U5609 ( .B1(n4651), .B2(n4653), .A(n4425), .ZN(n4649) );
  AOI21_X1 U5610 ( .B1(n8396), .B2(n4642), .A(n4638), .ZN(n4637) );
  NAND2_X1 U5611 ( .A1(n4639), .A2(n8259), .ZN(n4638) );
  AND4_X1 U5612 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n7611)
         );
  AND4_X1 U5613 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(n7564)
         );
  XNOR2_X1 U5614 ( .A(n6305), .B(n6304), .ZN(n6895) );
  NAND2_X1 U5615 ( .A1(n4346), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U5616 ( .A1(n8333), .A2(n8012), .ZN(n8342) );
  NAND2_X1 U5617 ( .A1(n4450), .A2(n5997), .ZN(n8708) );
  NAND2_X1 U5618 ( .A1(n6871), .A2(n8052), .ZN(n4450) );
  OAI21_X1 U5619 ( .B1(n8005), .B2(n4672), .A(n4671), .ZN(n8370) );
  NAND2_X1 U5620 ( .A1(n4663), .A2(n4662), .ZN(n8378) );
  INV_X1 U5621 ( .A(n8425), .ZN(n10129) );
  AND4_X1 U5622 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n8716)
         );
  NAND2_X1 U5623 ( .A1(n4650), .A2(n4654), .ZN(n8387) );
  NAND2_X1 U5624 ( .A1(n8333), .A2(n4655), .ZN(n4650) );
  AND2_X1 U5625 ( .A1(n6056), .A2(n6055), .ZN(n8404) );
  INV_X1 U5626 ( .A(n10134), .ZN(n8403) );
  AOI21_X1 U5627 ( .B1(n8615), .B2(n6070), .A(n6054), .ZN(n8623) );
  AND2_X1 U5628 ( .A1(n6352), .A2(n6351), .ZN(n10138) );
  AOI21_X1 U5629 ( .B1(n8290), .B2(n8291), .A(n4873), .ZN(n8407) );
  INV_X1 U5630 ( .A(n8383), .ZN(n10126) );
  OAI21_X1 U5631 ( .B1(n8063), .B2(n4578), .A(n4374), .ZN(n4577) );
  NAND2_X1 U5632 ( .A1(n4439), .A2(n4438), .ZN(n8250) );
  NAND2_X1 U5633 ( .A1(n4579), .A2(n6188), .ZN(n4578) );
  XNOR2_X1 U5634 ( .A(n6144), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8254) );
  OR2_X1 U5635 ( .A1(n6631), .A2(P2_U3151), .ZN(n8532) );
  OAI22_X1 U5636 ( .A1(n6634), .A2(n9760), .B1(n9762), .B2(n9761), .ZN(n9785)
         );
  INV_X1 U5637 ( .A(n4592), .ZN(n7512) );
  XNOR2_X1 U5638 ( .A(n7583), .B(n7577), .ZN(n7510) );
  NAND2_X1 U5639 ( .A1(n7510), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7584) );
  NOR2_X1 U5640 ( .A1(n7578), .A2(n7579), .ZN(n7582) );
  OR2_X1 U5641 ( .A1(n7761), .A2(n7812), .ZN(n4683) );
  NAND2_X1 U5642 ( .A1(n4427), .A2(n4682), .ZN(n4684) );
  INV_X1 U5643 ( .A(n4496), .ZN(n4491) );
  INV_X1 U5644 ( .A(n7814), .ZN(n4493) );
  NAND2_X1 U5645 ( .A1(n4490), .A2(n4489), .ZN(n8452) );
  NAND2_X1 U5646 ( .A1(n7814), .A2(n4494), .ZN(n4489) );
  NAND2_X1 U5647 ( .A1(n4407), .A2(n4682), .ZN(n4490) );
  INV_X1 U5648 ( .A(n9788), .ZN(n8534) );
  XNOR2_X1 U5649 ( .A(n8469), .B(n8477), .ZN(n8453) );
  NOR2_X1 U5650 ( .A1(n8453), .A2(n8735), .ZN(n8470) );
  OAI21_X1 U5651 ( .B1(n8453), .B2(n4688), .A(n4687), .ZN(n8498) );
  NAND2_X1 U5652 ( .A1(n4689), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U5653 ( .A1(n8471), .A2(n4689), .ZN(n4687) );
  INV_X1 U5654 ( .A(n8473), .ZN(n4689) );
  NAND2_X1 U5655 ( .A1(n4550), .A2(n4554), .ZN(n8606) );
  NAND2_X1 U5656 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  INV_X1 U5657 ( .A(n8404), .ZN(n8799) );
  NAND2_X1 U5658 ( .A1(n6048), .A2(n6047), .ZN(n8614) );
  NAND2_X1 U5659 ( .A1(n4553), .A2(n4557), .ZN(n8617) );
  NAND2_X1 U5660 ( .A1(n8632), .A2(n4559), .ZN(n4553) );
  NOR2_X1 U5661 ( .A1(n8632), .A2(n8184), .ZN(n8627) );
  AOI21_X1 U5662 ( .B1(n8625), .B2(n6070), .A(n6045), .ZN(n8811) );
  INV_X1 U5663 ( .A(n8897), .ZN(n8639) );
  AND2_X1 U5664 ( .A1(n5746), .A2(n5745), .ZN(n8818) );
  NAND2_X1 U5665 ( .A1(n6032), .A2(n6031), .ZN(n8817) );
  NAND2_X1 U5666 ( .A1(n7572), .A2(n8052), .ZN(n6032) );
  NAND2_X1 U5667 ( .A1(n4570), .A2(n4569), .ZN(n8652) );
  NAND2_X1 U5668 ( .A1(n6022), .A2(n6021), .ZN(n8662) );
  AND2_X1 U5669 ( .A1(n4570), .A2(n8195), .ZN(n7906) );
  AND2_X1 U5670 ( .A1(n6123), .A2(n6122), .ZN(n8665) );
  NAND2_X1 U5671 ( .A1(n4565), .A2(n8168), .ZN(n8718) );
  NAND2_X1 U5672 ( .A1(n9791), .A2(n8134), .ZN(n7609) );
  INV_X1 U5673 ( .A(n6332), .ZN(n10135) );
  INV_X1 U5674 ( .A(n7557), .ZN(n9851) );
  INV_X1 U5675 ( .A(n10130), .ZN(n10120) );
  NAND2_X1 U5676 ( .A1(n4547), .A2(n6111), .ZN(n7342) );
  NAND2_X1 U5677 ( .A1(n6110), .A2(n6913), .ZN(n4547) );
  INV_X1 U5678 ( .A(n5793), .ZN(n4807) );
  INV_X2 U5679 ( .A(n9807), .ZN(n9808) );
  NAND2_X1 U5680 ( .A1(n6299), .A2(n7365), .ZN(n6989) );
  INV_X1 U5681 ( .A(n8614), .ZN(n8889) );
  AND2_X1 U5682 ( .A1(n6039), .A2(n6038), .ZN(n8893) );
  NAND2_X1 U5683 ( .A1(n5962), .A2(n5961), .ZN(n8908) );
  INV_X1 U5684 ( .A(n5983), .ZN(n8914) );
  INV_X1 U5685 ( .A(n8385), .ZN(n8918) );
  INV_X2 U5686 ( .A(n9878), .ZN(n9880) );
  NAND2_X1 U5687 ( .A1(n6974), .A2(n6549), .ZN(n6561) );
  INV_X1 U5688 ( .A(n6161), .ZN(n7872) );
  XNOR2_X1 U5689 ( .A(n6147), .B(n6152), .ZN(n7864) );
  NAND2_X1 U5690 ( .A1(n6150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U5691 ( .A1(n6150), .A2(n6149), .ZN(n7810) );
  OR2_X1 U5692 ( .A1(n6148), .A2(n6153), .ZN(n6149) );
  INV_X1 U5693 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9963) );
  INV_X1 U5694 ( .A(n8254), .ZN(n7573) );
  INV_X1 U5695 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7492) );
  INV_X1 U5696 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7155) );
  INV_X1 U5697 ( .A(n6299), .ZN(n8558) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6924) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6872) );
  INV_X1 U5700 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6714) );
  INV_X1 U5701 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6414) );
  INV_X1 U5702 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6410) );
  INV_X1 U5703 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6406) );
  INV_X1 U5704 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6379) );
  NOR2_X1 U5705 ( .A1(n5799), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5813) );
  INV_X1 U5706 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6390) );
  AND2_X1 U5707 ( .A1(n6395), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6297) );
  INV_X1 U5708 ( .A(n7957), .ZN(n7959) );
  AND2_X1 U5709 ( .A1(n7990), .A2(n7989), .ZN(n8991) );
  NAND2_X1 U5710 ( .A1(n5087), .A2(n5086), .ZN(n9258) );
  NOR2_X1 U5711 ( .A1(n9046), .A2(n4877), .ZN(n8998) );
  NAND2_X1 U5712 ( .A1(n4744), .A2(n7223), .ZN(n7386) );
  NAND2_X1 U5713 ( .A1(n4747), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U5714 ( .A1(n5275), .A2(n5274), .ZN(n7235) );
  NAND2_X1 U5715 ( .A1(n5223), .A2(n5222), .ZN(n9022) );
  AOI21_X1 U5716 ( .B1(n9015), .B2(n9016), .A(n4350), .ZN(n9025) );
  NAND2_X1 U5717 ( .A1(n5462), .A2(n5461), .ZN(n9521) );
  NOR2_X1 U5718 ( .A1(n9048), .A2(n9047), .ZN(n9046) );
  XNOR2_X1 U5719 ( .A(n7957), .B(n4728), .ZN(n9056) );
  INV_X1 U5720 ( .A(n7958), .ZN(n4728) );
  NAND2_X1 U5721 ( .A1(n9015), .A2(n4736), .ZN(n4729) );
  NAND2_X1 U5722 ( .A1(n5110), .A2(n5109), .ZN(n9293) );
  INV_X1 U5723 ( .A(n9059), .ZN(n9098) );
  INV_X1 U5724 ( .A(n9061), .ZN(n9101) );
  NAND2_X1 U5725 ( .A1(n5118), .A2(n5117), .ZN(n9109) );
  NAND4_X1 U5726 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n9129)
         );
  NAND4_X1 U5727 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5417), .ZN(n9131)
         );
  INV_X2 U5728 ( .A(P1_U3973), .ZN(n9132) );
  INV_X1 U5729 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U5730 ( .A1(n9255), .A2(n9254), .ZN(n9464) );
  AND2_X1 U5731 ( .A1(n9333), .A2(n6253), .ZN(n9320) );
  NAND2_X1 U5732 ( .A1(n4749), .A2(n4752), .ZN(n9317) );
  OR2_X1 U5733 ( .A1(n9363), .A2(n4753), .ZN(n4749) );
  NAND2_X1 U5734 ( .A1(n4756), .A2(n4758), .ZN(n9332) );
  NAND2_X1 U5735 ( .A1(n9363), .A2(n4759), .ZN(n4756) );
  NAND2_X1 U5736 ( .A1(n4757), .A2(n6235), .ZN(n9347) );
  OR2_X1 U5737 ( .A1(n9363), .A2(n6236), .ZN(n4757) );
  AND2_X1 U5738 ( .A1(n5176), .A2(n5175), .ZN(n9386) );
  NAND2_X1 U5739 ( .A1(n5520), .A2(n5600), .ZN(n9399) );
  OAI21_X1 U5740 ( .B1(n6227), .B2(n4719), .A(n4717), .ZN(n9412) );
  NAND2_X1 U5741 ( .A1(n4720), .A2(n4723), .ZN(n7851) );
  NAND2_X1 U5742 ( .A1(n6227), .A2(n4725), .ZN(n4720) );
  NAND2_X1 U5743 ( .A1(n6227), .A2(n4871), .ZN(n7838) );
  INV_X1 U5744 ( .A(n9532), .ZN(n9106) );
  INV_X1 U5745 ( .A(n7235), .ZN(n6221) );
  NAND2_X1 U5746 ( .A1(n4765), .A2(n4770), .ZN(n7493) );
  NAND2_X1 U5747 ( .A1(n6218), .A2(n4771), .ZN(n4765) );
  NAND2_X1 U5748 ( .A1(n7455), .A2(n5516), .ZN(n7459) );
  NAND2_X1 U5749 ( .A1(n7031), .A2(n7039), .ZN(n7030) );
  NAND2_X1 U5750 ( .A1(n6993), .A2(n6215), .ZN(n7031) );
  INV_X1 U5751 ( .A(n9247), .ZN(n9450) );
  INV_X1 U5752 ( .A(n9724), .ZN(n7117) );
  OR2_X1 U5753 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  INV_X1 U5754 ( .A(n4540), .ZN(n4539) );
  OAI21_X1 U5755 ( .B1(n6397), .B2(n6445), .A(n5372), .ZN(n4540) );
  INV_X1 U5756 ( .A(n9530), .ZN(n7728) );
  INV_X1 U5758 ( .A(n5642), .ZN(n9550) );
  INV_X1 U5759 ( .A(n9293), .ZN(n9562) );
  AND2_X1 U5760 ( .A1(n5122), .A2(n5121), .ZN(n9566) );
  AND2_X1 U5761 ( .A1(n5212), .A2(n5211), .ZN(n9581) );
  NAND2_X1 U5762 ( .A1(n5320), .A2(n5319), .ZN(n9432) );
  INV_X2 U5763 ( .A(n7727), .ZN(n9738) );
  OAI21_X1 U5764 ( .B1(n5057), .B2(n5056), .A(n5024), .ZN(n5027) );
  INV_X1 U5765 ( .A(n5078), .ZN(n7883) );
  XNOR2_X1 U5766 ( .A(n5085), .B(n5084), .ZN(n8942) );
  INV_X1 U5767 ( .A(n5042), .ZN(n4791) );
  XNOR2_X1 U5768 ( .A(n5101), .B(n5100), .ZN(n8049) );
  NAND2_X1 U5769 ( .A1(n5108), .A2(n5107), .ZN(n5097) );
  OAI21_X1 U5770 ( .B1(n5701), .B2(n5036), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4792) );
  INV_X1 U5771 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5035) );
  INV_X1 U5772 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5697) );
  OAI21_X2 U5773 ( .B1(n5699), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5698) );
  INV_X1 U5774 ( .A(n6270), .ZN(n7867) );
  INV_X1 U5775 ( .A(n6271), .ZN(n7807) );
  NAND2_X1 U5776 ( .A1(n4845), .A2(n4850), .ZN(n5141) );
  INV_X1 U5777 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7576) );
  INV_X1 U5778 ( .A(n6478), .ZN(n7574) );
  INV_X1 U5779 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7489) );
  INV_X1 U5780 ( .A(n6262), .ZN(n7490) );
  NAND2_X1 U5781 ( .A1(n4347), .A2(n4882), .ZN(n4695) );
  INV_X1 U5782 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8276) );
  INV_X1 U5783 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6874) );
  INV_X1 U5784 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U5785 ( .A1(n4619), .A2(n4842), .ZN(n5342) );
  NAND2_X1 U5786 ( .A1(n5371), .A2(n4447), .ZN(n4619) );
  NAND2_X1 U5787 ( .A1(n4840), .A2(n4917), .ZN(n5414) );
  INV_X1 U5788 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6381) );
  XNOR2_X1 U5789 ( .A(n5371), .B(n5370), .ZN(n6380) );
  INV_X1 U5790 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6375) );
  CLKBUF_X1 U5791 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9596) );
  INV_X1 U5792 ( .A(n4513), .ZN(n7732) );
  INV_X1 U5793 ( .A(n4512), .ZN(n7674) );
  AOI21_X1 U5794 ( .B1(n8535), .B2(n8541), .A(n4593), .ZN(n8545) );
  OAI21_X1 U5795 ( .B1(n4636), .B2(n9779), .A(n4399), .ZN(P2_U3201) );
  XNOR2_X1 U5796 ( .A(n8564), .B(n8563), .ZN(n4636) );
  AND3_X1 U5797 ( .A1(n4467), .A2(n4466), .A3(n4475), .ZN(n7876) );
  AND2_X1 U5798 ( .A1(n4816), .A2(n4416), .ZN(n8792) );
  NOR2_X1 U5799 ( .A1(n6199), .A2(n6201), .ZN(n6202) );
  NAND2_X1 U5800 ( .A1(n9894), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4817) );
  OAI21_X1 U5801 ( .B1(n4818), .B2(n4814), .A(n4813), .ZN(n4812) );
  INV_X1 U5802 ( .A(n4815), .ZN(n4814) );
  OAI21_X1 U5803 ( .B1(n6198), .B2(n8935), .A(n6184), .ZN(n6185) );
  NAND2_X1 U5804 ( .A1(n4816), .A2(n4815), .ZN(n8883) );
  AOI21_X1 U5805 ( .B1(n9077), .B2(n4603), .A(n4426), .ZN(n4602) );
  OAI21_X1 U5806 ( .B1(n4536), .B2(n4535), .A(n5694), .ZN(n4838) );
  NAND2_X1 U5807 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  INV_X1 U5808 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9234) );
  MUX2_X1 U5809 ( .A(n9458), .B(n9543), .S(n9509), .Z(n9459) );
  MUX2_X1 U5810 ( .A(n9544), .B(n9543), .S(n9738), .Z(n9545) );
  AND2_X1 U5811 ( .A1(n5639), .A2(n5638), .ZN(n6260) );
  AND2_X1 U5812 ( .A1(n4554), .A2(n8066), .ZN(n4349) );
  AND2_X1 U5813 ( .A1(n7926), .A2(n7925), .ZN(n4350) );
  NAND4_X1 U5814 ( .A1(n5730), .A2(n5729), .A3(n5728), .A4(n6154), .ZN(n4351)
         );
  NAND2_X1 U5815 ( .A1(n5291), .A2(n5290), .ZN(n7463) );
  AND3_X1 U5816 ( .A1(n5634), .A2(n9267), .A3(n6248), .ZN(n4352) );
  OR2_X1 U5817 ( .A1(n5358), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4353) );
  AND2_X1 U5818 ( .A1(n5605), .A2(n6248), .ZN(n4354) );
  OR2_X1 U5819 ( .A1(n8428), .A2(n9830), .ZN(n4355) );
  INV_X1 U5820 ( .A(n9130), .ZN(n6209) );
  OR2_X1 U5821 ( .A1(n5648), .A2(n9699), .ZN(n4356) );
  AND2_X1 U5822 ( .A1(n5677), .A2(n6248), .ZN(n4357) );
  AND2_X1 U5823 ( .A1(n4781), .A2(n4784), .ZN(n4358) );
  INV_X1 U5824 ( .A(n4760), .ZN(n4759) );
  NAND2_X1 U5825 ( .A1(n4379), .A2(n6235), .ZN(n4760) );
  INV_X1 U5826 ( .A(n4665), .ZN(n4664) );
  INV_X1 U5827 ( .A(n4556), .ZN(n4551) );
  NAND2_X1 U5828 ( .A1(n4557), .A2(n6127), .ZN(n4556) );
  INV_X1 U5829 ( .A(n9349), .ZN(n9571) );
  NAND2_X1 U5830 ( .A1(n5156), .A2(n5155), .ZN(n9349) );
  AND2_X1 U5831 ( .A1(n9486), .A2(n9110), .ZN(n4359) );
  OAI21_X1 U5832 ( .B1(n4717), .B2(n4715), .A(n4423), .ZN(n4714) );
  OR2_X1 U5833 ( .A1(n9047), .A2(n8997), .ZN(n4360) );
  NAND2_X1 U5834 ( .A1(n5165), .A2(n5164), .ZN(n9372) );
  INV_X1 U5835 ( .A(n9372), .ZN(n9575) );
  AND2_X1 U5836 ( .A1(n4504), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4361) );
  AND2_X1 U5837 ( .A1(n4585), .A2(n8458), .ZN(n4362) );
  OR2_X1 U5838 ( .A1(n4959), .A2(SI_16_), .ZN(n4363) );
  NAND2_X1 U5839 ( .A1(n8013), .A2(n8420), .ZN(n4364) );
  INV_X1 U5840 ( .A(n8794), .ZN(n8048) );
  NAND2_X1 U5841 ( .A1(n6067), .A2(n6066), .ZN(n8794) );
  INV_X1 U5842 ( .A(n9278), .ZN(n9558) );
  NAND2_X1 U5843 ( .A1(n5103), .A2(n5102), .ZN(n9278) );
  INV_X1 U5844 ( .A(n7577), .ZN(n4690) );
  OAI21_X1 U5845 ( .B1(n5923), .B2(n5946), .A(n5933), .ZN(n8454) );
  OR2_X1 U5846 ( .A1(n8534), .A2(n8541), .ZN(n4365) );
  INV_X1 U5847 ( .A(n8502), .ZN(n8499) );
  INV_X1 U5848 ( .A(n6745), .ZN(n4486) );
  AND2_X1 U5850 ( .A1(n8787), .A2(n8793), .ZN(n4366) );
  OR2_X1 U5851 ( .A1(n7742), .A2(n7670), .ZN(n4367) );
  INV_X1 U5852 ( .A(n5799), .ZN(n4823) );
  AND2_X1 U5853 ( .A1(n9229), .A2(n7574), .ZN(n6248) );
  NAND4_X1 U5854 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n6204)
         );
  OR2_X1 U5855 ( .A1(n6647), .A2(n6673), .ZN(n4370) );
  NAND4_X1 U5856 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n8429)
         );
  OR2_X1 U5857 ( .A1(n7273), .A2(n7274), .ZN(n4371) );
  OR2_X1 U5858 ( .A1(n9486), .A2(n9110), .ZN(n4372) );
  NOR2_X1 U5859 ( .A1(n7878), .A2(n9859), .ZN(n4373) );
  NOR2_X1 U5860 ( .A1(n8096), .A2(n7365), .ZN(n4374) );
  NOR2_X1 U5861 ( .A1(n7186), .A2(n4748), .ZN(n4375) );
  NAND2_X1 U5862 ( .A1(n5033), .A2(n5187), .ZN(n5233) );
  AND2_X1 U5863 ( .A1(n4928), .A2(n4927), .ZN(n4376) );
  INV_X1 U5864 ( .A(n6582), .ZN(n7050) );
  AND3_X1 U5865 ( .A1(n5427), .A2(n5426), .A3(n5425), .ZN(n6582) );
  XNOR2_X1 U5866 ( .A(n5027), .B(n5026), .ZN(n7885) );
  AND4_X1 U5867 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n4377)
         );
  AND2_X1 U5868 ( .A1(n7996), .A2(n7997), .ZN(n4378) );
  OR2_X1 U5869 ( .A1(n9349), .A2(n9112), .ZN(n4379) );
  AND2_X1 U5870 ( .A1(n5635), .A2(n6248), .ZN(n4380) );
  NOR2_X1 U5871 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5189) );
  OR2_X1 U5872 ( .A1(n5983), .A2(n8689), .ZN(n8195) );
  AND3_X1 U5873 ( .A1(n5400), .A2(n5399), .A3(n5398), .ZN(n7320) );
  INV_X1 U5874 ( .A(n4938), .ZN(n4624) );
  AND3_X1 U5875 ( .A1(n5386), .A2(n5385), .A3(n5384), .ZN(n6964) );
  NAND2_X1 U5876 ( .A1(n7146), .A2(n9825), .ZN(n4381) );
  NAND2_X1 U5877 ( .A1(n4824), .A2(n4823), .ZN(n5826) );
  NAND2_X1 U5878 ( .A1(n5201), .A2(n5200), .ZN(n9512) );
  AND2_X1 U5879 ( .A1(n4367), .A2(n7761), .ZN(n4382) );
  NOR2_X1 U5880 ( .A1(n8470), .A2(n8471), .ZN(n4383) );
  NOR2_X1 U5881 ( .A1(n8518), .A2(n8519), .ZN(n4384) );
  NAND2_X1 U5882 ( .A1(n4823), .A2(n4821), .ZN(n4385) );
  AND4_X1 U5883 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n7041)
         );
  AND2_X1 U5884 ( .A1(n4357), .A2(n5597), .ZN(n4386) );
  AND2_X1 U5885 ( .A1(n4716), .A2(n6229), .ZN(n4387) );
  INV_X1 U5886 ( .A(n9538), .ZN(n7719) );
  NAND2_X1 U5887 ( .A1(n5250), .A2(n5249), .ZN(n9538) );
  INV_X1 U5888 ( .A(n7039), .ZN(n4743) );
  INV_X1 U5889 ( .A(n4784), .ZN(n4783) );
  OAI21_X1 U5890 ( .B1(n9268), .B2(n4785), .A(n9251), .ZN(n4784) );
  AND2_X1 U5891 ( .A1(n4376), .A2(n4879), .ZN(n4388) );
  AND2_X1 U5892 ( .A1(n4663), .A2(n4660), .ZN(n4389) );
  OR2_X1 U5893 ( .A1(n9784), .A2(n9883), .ZN(n4390) );
  AND2_X1 U5894 ( .A1(n8799), .A2(n8613), .ZN(n8219) );
  INV_X1 U5895 ( .A(n6795), .ZN(n9127) );
  AND4_X1 U5896 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n6795)
         );
  AND2_X1 U5897 ( .A1(n9521), .A2(n9116), .ZN(n4391) );
  AND2_X1 U5898 ( .A1(n4616), .A2(n4388), .ZN(n4392) );
  INV_X1 U5899 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7886) );
  AND2_X1 U5900 ( .A1(n5590), .A2(n5671), .ZN(n4393) );
  NOR2_X1 U5901 ( .A1(n6221), .A2(n6220), .ZN(n4394) );
  AND2_X1 U5902 ( .A1(n9344), .A2(n9058), .ZN(n4395) );
  INV_X1 U5903 ( .A(n4704), .ZN(n4703) );
  NAND2_X1 U5904 ( .A1(n4705), .A2(n9575), .ZN(n4704) );
  AND2_X1 U5905 ( .A1(n8897), .A2(n8417), .ZN(n8184) );
  INV_X1 U5906 ( .A(n4666), .ZN(n8030) );
  NOR2_X1 U5907 ( .A1(n7933), .A2(n7932), .ZN(n4396) );
  NOR2_X1 U5908 ( .A1(n9432), .A2(n9124), .ZN(n4397) );
  OR2_X2 U5909 ( .A1(n5040), .A2(n4798), .ZN(n4398) );
  AND2_X1 U5910 ( .A1(n4635), .A2(n4634), .ZN(n4399) );
  AND2_X1 U5911 ( .A1(n6332), .A2(n7611), .ZN(n4400) );
  OR2_X1 U5912 ( .A1(n4695), .A2(n5233), .ZN(n4401) );
  INV_X1 U5913 ( .A(n4572), .ZN(n4571) );
  NAND2_X1 U5914 ( .A1(n6122), .A2(n8668), .ZN(n4572) );
  INV_X1 U5915 ( .A(n4698), .ZN(n4697) );
  NAND2_X1 U5916 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  INV_X1 U5917 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5651) );
  OR2_X1 U5918 ( .A1(n8662), .A2(n8833), .ZN(n8179) );
  AND2_X1 U5919 ( .A1(n4620), .A2(n7955), .ZN(n4402) );
  NOR2_X1 U5920 ( .A1(n9571), .A2(n7956), .ZN(n4403) );
  AND2_X1 U5921 ( .A1(n5041), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4404) );
  INV_X1 U5922 ( .A(n7463), .ZN(n4772) );
  AND2_X1 U5923 ( .A1(n4919), .A2(SI_6_), .ZN(n4405) );
  AND2_X1 U5924 ( .A1(n4753), .A2(n4372), .ZN(n4406) );
  AND2_X1 U5925 ( .A1(n4681), .A2(n4492), .ZN(n4407) );
  AND2_X1 U5926 ( .A1(n7004), .A2(n5350), .ZN(n5554) );
  INV_X1 U5927 ( .A(n5554), .ZN(n4520) );
  AND2_X1 U5928 ( .A1(n8026), .A2(n8824), .ZN(n4408) );
  NAND2_X1 U5929 ( .A1(n9258), .A2(n8978), .ZN(n6259) );
  NAND2_X1 U5930 ( .A1(n4393), .A2(n4724), .ZN(n4723) );
  INV_X1 U5931 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4507) );
  INV_X1 U5932 ( .A(n7180), .ZN(n4446) );
  AND2_X1 U5933 ( .A1(n4752), .A2(n4372), .ZN(n4409) );
  AND3_X1 U5934 ( .A1(n5625), .A2(n5637), .A3(n4525), .ZN(n4410) );
  INV_X1 U5935 ( .A(n5341), .ZN(n4618) );
  OR2_X1 U5936 ( .A1(n8799), .A2(n8613), .ZN(n8217) );
  AND2_X1 U5937 ( .A1(n7505), .A2(n4691), .ZN(n4411) );
  NAND2_X1 U5938 ( .A1(n8429), .A2(n7170), .ZN(n4412) );
  OAI21_X1 U5939 ( .B1(n9048), .B2(n4360), .A(n4402), .ZN(n7957) );
  INV_X1 U5940 ( .A(n4864), .ZN(n4863) );
  OAI21_X1 U5941 ( .B1(n4948), .B2(n4865), .A(n4947), .ZN(n4864) );
  NOR2_X1 U5942 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5188) );
  INV_X1 U5943 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5907) );
  INV_X1 U5944 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5041) );
  XNOR2_X1 U5945 ( .A(n4657), .B(n4656), .ZN(n6299) );
  NOR2_X1 U5946 ( .A1(n5862), .A2(n5845), .ZN(n4413) );
  NAND2_X1 U5947 ( .A1(n4747), .A2(n7185), .ZN(n7225) );
  AND2_X1 U5948 ( .A1(n4589), .A2(n7772), .ZN(n4414) );
  INV_X1 U5949 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U5950 ( .A1(n4729), .A2(n4735), .ZN(n9065) );
  NAND2_X1 U5951 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5984) );
  INV_X1 U5952 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4574) );
  AND2_X1 U5953 ( .A1(n8340), .A2(n8716), .ZN(n4415) );
  NOR2_X1 U5954 ( .A1(n5970), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U5955 ( .A1(n8798), .A2(n8728), .ZN(n4416) );
  NAND3_X1 U5956 ( .A1(n4823), .A2(n4819), .A3(n4573), .ZN(n5877) );
  NAND2_X1 U5957 ( .A1(n7539), .A2(n7540), .ZN(n7918) );
  INV_X1 U5958 ( .A(n7918), .ZN(n4613) );
  NOR3_X1 U5959 ( .A1(n7659), .A2(n9022), .A3(n4710), .ZN(n4707) );
  AND2_X1 U5960 ( .A1(n6064), .A2(n6063), .ZN(n8613) );
  NAND2_X1 U5961 ( .A1(n4823), .A2(n4819), .ZN(n5851) );
  AND2_X1 U5962 ( .A1(n4855), .A2(n5208), .ZN(n4417) );
  INV_X1 U5963 ( .A(n8656), .ZN(n8675) );
  AND3_X1 U5964 ( .A1(n5969), .A2(n5968), .A3(n5967), .ZN(n8656) );
  NAND2_X1 U5965 ( .A1(n9417), .A2(n4703), .ZN(n4706) );
  INV_X1 U5966 ( .A(n4456), .ZN(n4455) );
  NOR2_X1 U5967 ( .A1(n4957), .A2(n4457), .ZN(n4456) );
  NAND2_X1 U5968 ( .A1(n5722), .A2(n4676), .ZN(n4678) );
  OR2_X1 U5969 ( .A1(n8440), .A2(n6759), .ZN(n4418) );
  OR2_X1 U5970 ( .A1(n7509), .A2(n7291), .ZN(n4419) );
  AND2_X1 U5971 ( .A1(n4584), .A2(n4585), .ZN(n4420) );
  AND2_X1 U5972 ( .A1(n4584), .A2(n4362), .ZN(n4421) );
  AND2_X1 U5973 ( .A1(n4959), .A2(SI_16_), .ZN(n4422) );
  OR2_X1 U5974 ( .A1(n9581), .A2(n8965), .ZN(n4423) );
  INV_X1 U5975 ( .A(n4363), .ZN(n4858) );
  AND2_X1 U5976 ( .A1(n4956), .A2(n4955), .ZN(n4424) );
  NAND2_X1 U5977 ( .A1(n8308), .A2(n8306), .ZN(n4425) );
  INV_X1 U5978 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5979 ( .A1(n8003), .A2(n4610), .ZN(n4426) );
  AND2_X1 U5980 ( .A1(n4681), .A2(n4491), .ZN(n4427) );
  OR2_X1 U5981 ( .A1(n9554), .A2(n9586), .ZN(n4428) );
  AND2_X1 U5982 ( .A1(n4454), .A2(n4363), .ZN(n4429) );
  INV_X1 U5983 ( .A(n8368), .ZN(n4673) );
  OR2_X1 U5984 ( .A1(n7733), .A2(n7683), .ZN(n4513) );
  AND2_X1 U5985 ( .A1(n4493), .A2(n4684), .ZN(n4430) );
  AND2_X1 U5986 ( .A1(n7761), .A2(n7812), .ZN(n4431) );
  AND2_X1 U5987 ( .A1(n4807), .A2(n4806), .ZN(n4432) );
  OAI21_X1 U5988 ( .B1(n6993), .B2(n4743), .A(n4741), .ZN(n7203) );
  AND2_X1 U5989 ( .A1(n8006), .A2(n8746), .ZN(n4433) );
  INV_X1 U5990 ( .A(n7816), .ZN(n4494) );
  NAND2_X1 U5991 ( .A1(n7083), .A2(n4697), .ZN(n4701) );
  INV_X1 U5992 ( .A(n4708), .ZN(n7845) );
  NOR2_X1 U5993 ( .A1(n7659), .A2(n4710), .ZN(n4708) );
  INV_X1 U5994 ( .A(n4837), .ZN(n4836) );
  NAND2_X1 U5995 ( .A1(n5098), .A2(n5107), .ZN(n4837) );
  NAND2_X1 U5996 ( .A1(n5096), .A2(n5099), .ZN(n4434) );
  AND2_X1 U5997 ( .A1(n5662), .A2(n5514), .ZN(n4435) );
  XNOR2_X1 U5998 ( .A(n5748), .B(n5747), .ZN(n6133) );
  AND2_X2 U5999 ( .A1(n6196), .A2(n6971), .ZN(n9897) );
  NAND2_X1 U6000 ( .A1(n6109), .A2(n6300), .ZN(n8726) );
  INV_X1 U6001 ( .A(n8726), .ZN(n9797) );
  INV_X1 U6002 ( .A(n9699), .ZN(n9229) );
  AND2_X1 U6003 ( .A1(n4679), .A2(n6703), .ZN(n4436) );
  XNOR2_X1 U6004 ( .A(n5652), .B(n5651), .ZN(n7435) );
  XNOR2_X1 U6005 ( .A(n6108), .B(n6107), .ZN(n7365) );
  NAND2_X1 U6006 ( .A1(n6105), .A2(n6156), .ZN(n8069) );
  INV_X1 U6007 ( .A(n8069), .ZN(n6188) );
  INV_X1 U6008 ( .A(n9760), .ZN(n4590) );
  NAND2_X1 U6009 ( .A1(n6766), .A2(n7288), .ZN(n7272) );
  INV_X1 U6010 ( .A(n7288), .ZN(n4499) );
  NOR2_X2 U6011 ( .A1(n4348), .A2(n6081), .ZN(n8578) );
  NAND2_X1 U6012 ( .A1(n5998), .A2(n8343), .ZN(n6000) );
  NAND2_X1 U6013 ( .A1(n6024), .A2(n6023), .ZN(n6033) );
  NAND2_X1 U6014 ( .A1(n4437), .A2(n4898), .ZN(n4901) );
  INV_X1 U6015 ( .A(n5441), .ZN(n4437) );
  NAND2_X1 U6016 ( .A1(n4897), .A2(SI_0_), .ZN(n5441) );
  NAND2_X1 U6017 ( .A1(n9553), .A2(n4428), .ZN(P1_U3518) );
  NAND2_X1 U6018 ( .A1(n9354), .A2(n6252), .ZN(n9335) );
  NAND2_X1 U6019 ( .A1(n7640), .A2(n5518), .ZN(n7643) );
  NAND2_X1 U6020 ( .A1(n9287), .A2(n9286), .ZN(n9269) );
  OAI21_X1 U6021 ( .B1(n5520), .B2(n5601), .A(n4786), .ZN(n6251) );
  OAI21_X1 U6022 ( .B1(n5514), .B2(n4794), .A(n4793), .ZN(n7494) );
  INV_X1 U6023 ( .A(n5413), .ZN(n4844) );
  AOI211_X1 U6024 ( .C1(n8216), .C2(n8610), .A(n8215), .B(n8605), .ZN(n8221)
         );
  NOR2_X1 U6025 ( .A1(n8225), .A2(n8224), .ZN(n8232) );
  MUX2_X1 U6026 ( .A(n8108), .B(n8107), .S(n8227), .Z(n8110) );
  NAND2_X1 U6027 ( .A1(n4442), .A2(n4441), .ZN(n8167) );
  NAND3_X1 U6028 ( .A1(n8162), .A2(n8161), .A3(n8743), .ZN(n4442) );
  NOR3_X1 U6029 ( .A1(n8133), .A2(n8140), .A3(n8132), .ZN(n8145) );
  AOI211_X1 U6030 ( .C1(n8200), .C2(n8199), .A(n8198), .B(n8643), .ZN(n8201)
         );
  NAND2_X1 U6031 ( .A1(n4577), .A2(n8250), .ZN(n4576) );
  XNOR2_X1 U6032 ( .A(n4576), .B(n8558), .ZN(n8257) );
  NAND2_X1 U6033 ( .A1(n4443), .A2(n6580), .ZN(n6615) );
  NAND2_X1 U6034 ( .A1(n6624), .A2(n6625), .ZN(n4443) );
  NAND2_X2 U6035 ( .A1(n6810), .A2(n6811), .ZN(n7019) );
  OAI21_X2 U6036 ( .B1(n5220), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5458) );
  OR2_X2 U6037 ( .A1(n6479), .A2(n6478), .ZN(n6481) );
  AOI21_X2 U6038 ( .B1(n4599), .B2(n7531), .A(n4445), .ZN(n7538) );
  NAND2_X1 U6039 ( .A1(n6853), .A2(n5655), .ZN(n5550) );
  NAND2_X1 U6040 ( .A1(n6829), .A2(n5535), .ZN(n6997) );
  AOI211_X2 U6041 ( .C1(n9466), .C2(n9735), .A(n9465), .B(n9464), .ZN(n9551)
         );
  NAND2_X1 U6042 ( .A1(n9266), .A2(n6258), .ZN(n9252) );
  NAND2_X2 U6043 ( .A1(n9005), .A2(n9006), .ZN(n9004) );
  OR2_X2 U6044 ( .A1(n6480), .A2(n6483), .ZN(n7049) );
  NOR2_X2 U6045 ( .A1(n9056), .A2(n9055), .ZN(n9054) );
  NOR2_X1 U6046 ( .A1(n4745), .A2(n4598), .ZN(n4597) );
  INV_X2 U6047 ( .A(n7971), .ZN(n8970) );
  NAND2_X1 U6048 ( .A1(n5247), .A2(n4429), .ZN(n4451) );
  OAI21_X1 U6049 ( .B1(n5247), .B2(n4455), .A(n4454), .ZN(n5219) );
  NAND2_X1 U6050 ( .A1(n4451), .A2(n4452), .ZN(n5456) );
  NAND2_X1 U6051 ( .A1(n4461), .A2(n4459), .ZN(n4626) );
  NAND2_X1 U6052 ( .A1(n4614), .A2(n4616), .ZN(n5321) );
  INV_X1 U6053 ( .A(n6143), .ZN(n4475) );
  NAND3_X1 U6054 ( .A1(n4467), .A2(n4466), .A3(n4465), .ZN(n6197) );
  NAND2_X1 U6055 ( .A1(n6087), .A2(n4468), .ZN(n4466) );
  MUX2_X1 U6056 ( .A(n6379), .B(n6381), .S(n6373), .Z(n4915) );
  INV_X1 U6057 ( .A(n6649), .ZN(n4478) );
  NAND2_X1 U6058 ( .A1(n6647), .A2(n6673), .ZN(n6680) );
  AOI21_X1 U6059 ( .B1(n7505), .B2(n4691), .A(n7577), .ZN(n4483) );
  NAND2_X1 U6060 ( .A1(n7505), .A2(n4480), .ZN(n4479) );
  INV_X1 U6061 ( .A(n4691), .ZN(n4481) );
  INV_X1 U6062 ( .A(n4483), .ZN(n4482) );
  NAND2_X1 U6063 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U6064 ( .A1(n8444), .A2(n8442), .ZN(n6763) );
  INV_X1 U6065 ( .A(n4488), .ZN(n4487) );
  NAND2_X1 U6066 ( .A1(n4497), .A2(n4499), .ZN(n4498) );
  INV_X1 U6067 ( .A(n6766), .ZN(n4497) );
  NAND2_X1 U6068 ( .A1(n7272), .A2(n4498), .ZN(n6767) );
  NAND3_X2 U6069 ( .A1(n4501), .A2(n4502), .A3(n4504), .ZN(n6658) );
  NAND3_X1 U6070 ( .A1(n4501), .A2(n4502), .A3(n4361), .ZN(n4503) );
  NAND2_X1 U6071 ( .A1(n4541), .A2(n4507), .ZN(n4502) );
  NAND2_X1 U6072 ( .A1(n4508), .A2(n4509), .ZN(n7811) );
  NAND2_X1 U6073 ( .A1(n4514), .A2(n4515), .ZN(n5565) );
  NAND4_X1 U6074 ( .A1(n5551), .A2(n5552), .A3(n4522), .A4(n4521), .ZN(n4514)
         );
  OAI21_X1 U6075 ( .B1(n5565), .B2(n5564), .A(n5563), .ZN(n5566) );
  INV_X1 U6076 ( .A(n5632), .ZN(n4528) );
  NAND2_X1 U6077 ( .A1(n5626), .A2(n4410), .ZN(n4523) );
  NAND4_X1 U6078 ( .A1(n4524), .A2(n4523), .A3(n4526), .A4(n6260), .ZN(n5641)
         );
  CLKBUF_X1 U6079 ( .A(n4542), .Z(n4541) );
  NAND2_X1 U6080 ( .A1(n4541), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6645) );
  OAI22_X1 U6081 ( .A1(n6657), .A2(n9760), .B1(n4541), .B2(n6656), .ZN(n9755)
         );
  AND2_X1 U6082 ( .A1(n4541), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U6083 ( .A1(n6984), .A2(n5761), .ZN(n8068) );
  NAND2_X1 U6084 ( .A1(n4546), .A2(n4543), .ZN(n7361) );
  NAND3_X1 U6085 ( .A1(n6110), .A2(n8119), .A3(n6913), .ZN(n4546) );
  NAND2_X1 U6086 ( .A1(n4349), .A2(n8632), .ZN(n4548) );
  NAND2_X1 U6087 ( .A1(n8733), .A2(n8169), .ZN(n4565) );
  NAND2_X1 U6088 ( .A1(n4560), .A2(n4563), .ZN(n8690) );
  NAND2_X1 U6089 ( .A1(n8733), .A2(n4561), .ZN(n4560) );
  INV_X1 U6090 ( .A(n7774), .ZN(n4580) );
  AOI21_X1 U6091 ( .B1(n4580), .B2(n4362), .A(n4581), .ZN(n8475) );
  MUX2_X1 U6092 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n8549), .Z(n6633) );
  OR2_X1 U6093 ( .A1(n4599), .A2(n4597), .ZN(n7532) );
  AOI21_X1 U6094 ( .B1(n4597), .B2(n7531), .A(n4884), .ZN(n4596) );
  INV_X1 U6095 ( .A(n7223), .ZN(n4598) );
  NAND2_X1 U6096 ( .A1(n7385), .A2(n4600), .ZN(n4599) );
  NAND3_X1 U6097 ( .A1(n7019), .A2(n7223), .A3(n4375), .ZN(n4600) );
  NAND2_X1 U6098 ( .A1(n4601), .A2(n4605), .ZN(n4611) );
  NAND2_X1 U6099 ( .A1(n9004), .A2(n4608), .ZN(n4601) );
  AND2_X2 U6100 ( .A1(n9077), .A2(n4378), .ZN(n8984) );
  NAND2_X1 U6101 ( .A1(n4604), .A2(n4602), .ZN(P1_U3214) );
  AND2_X1 U6102 ( .A1(n4378), .A2(n9095), .ZN(n4603) );
  NAND2_X1 U6103 ( .A1(n4611), .A2(n9095), .ZN(n4604) );
  NAND2_X2 U6104 ( .A1(n9004), .A2(n7983), .ZN(n9077) );
  NAND2_X2 U6105 ( .A1(n9093), .A2(n4612), .ZN(n9015) );
  NAND2_X2 U6106 ( .A1(n9092), .A2(n9094), .ZN(n9093) );
  XNOR2_X2 U6107 ( .A(n7918), .B(n7917), .ZN(n9092) );
  NAND2_X1 U6108 ( .A1(n4626), .A2(n4938), .ZN(n5284) );
  NAND2_X1 U6109 ( .A1(n4934), .A2(n4933), .ZN(n5299) );
  MUX2_X1 U6110 ( .A(n9883), .B(P2_REG1_REG_2__SCAN_IN), .S(n6658), .Z(n9771)
         );
  AOI21_X1 U6111 ( .B1(n8396), .B2(n4641), .A(n4644), .ZN(n4640) );
  INV_X1 U6112 ( .A(n4637), .ZN(n8263) );
  INV_X1 U6113 ( .A(n8394), .ZN(n4647) );
  NAND2_X1 U6114 ( .A1(n8333), .A2(n4651), .ZN(n4648) );
  NAND2_X1 U6115 ( .A1(n4648), .A2(n4649), .ZN(n8307) );
  AOI21_X1 U6116 ( .B1(n8358), .B2(n8315), .A(n8314), .ZN(n8317) );
  OR2_X1 U6117 ( .A1(n8024), .A2(n8019), .ZN(n4665) );
  NAND3_X1 U6118 ( .A1(n8005), .A2(n4673), .A3(n4671), .ZN(n4669) );
  NAND2_X1 U6119 ( .A1(n5722), .A2(n4674), .ZN(n5970) );
  NAND2_X1 U6120 ( .A1(n5722), .A2(n5721), .ZN(n5884) );
  INV_X1 U6121 ( .A(n4678), .ZN(n5908) );
  NAND2_X1 U6122 ( .A1(n8040), .A2(n8039), .ZN(n8396) );
  NOR2_X1 U6123 ( .A1(n5884), .A2(n5727), .ZN(n6100) );
  NAND3_X1 U6124 ( .A1(n4682), .A2(n4683), .A3(n4681), .ZN(n7763) );
  INV_X1 U6125 ( .A(n4684), .ZN(n7813) );
  OAI21_X1 U6126 ( .B1(n8500), .B2(n4686), .A(n4685), .ZN(n8547) );
  AND2_X1 U6127 ( .A1(n5187), .A2(n5651), .ZN(n4693) );
  NAND4_X1 U6128 ( .A1(n4693), .A2(n4882), .A3(n4347), .A4(n5033), .ZN(n5358)
         );
  INV_X1 U6129 ( .A(n4701), .ZN(n7207) );
  INV_X1 U6130 ( .A(n4706), .ZN(n9371) );
  NOR2_X2 U6131 ( .A1(n9256), .A2(n6291), .ZN(n9243) );
  OR2_X2 U6132 ( .A1(n9275), .A2(n9258), .ZN(n9256) );
  INV_X1 U6133 ( .A(n4707), .ZN(n7853) );
  AND2_X2 U6134 ( .A1(n5448), .A2(n5447), .ZN(n9724) );
  AND2_X1 U6135 ( .A1(n5443), .A2(n5444), .ZN(n5448) );
  OAI21_X1 U6136 ( .B1(n6864), .B2(n4712), .A(n6859), .ZN(n6966) );
  NAND2_X1 U6137 ( .A1(n4712), .A2(n6864), .ZN(n6859) );
  INV_X1 U6138 ( .A(n6227), .ZN(n4713) );
  NAND2_X1 U6139 ( .A1(n7019), .A2(n7018), .ZN(n7187) );
  INV_X1 U6140 ( .A(n7018), .ZN(n4748) );
  NAND2_X1 U6141 ( .A1(n9363), .A2(n4409), .ZN(n4751) );
  XNOR2_X2 U6142 ( .A(n4761), .B(n8973), .ZN(n6587) );
  NAND2_X1 U6143 ( .A1(n6581), .A2(n4762), .ZN(n4761) );
  AND2_X4 U6144 ( .A1(n8977), .A2(n7975), .ZN(n7971) );
  NAND2_X1 U6145 ( .A1(n4763), .A2(n4764), .ZN(n7651) );
  NAND2_X1 U6146 ( .A1(n6218), .A2(n4766), .ZN(n4763) );
  INV_X1 U6147 ( .A(n6218), .ZN(n7451) );
  AOI21_X2 U6148 ( .B1(n6809), .B2(n6808), .A(n6807), .ZN(n6810) );
  NAND2_X2 U6149 ( .A1(n6781), .A2(n6780), .ZN(n6809) );
  OR2_X2 U6150 ( .A1(n6738), .A2(n6737), .ZN(n6781) );
  AND2_X2 U6151 ( .A1(n6731), .A2(n6730), .ZN(n6738) );
  OAI211_X1 U6152 ( .C1(n5448), .C2(n5502), .A(n4774), .B(n4773), .ZN(n6205)
         );
  NAND3_X1 U6153 ( .A1(n5447), .A2(n5448), .A3(n5502), .ZN(n4773) );
  OR2_X1 U6154 ( .A1(n5447), .A2(n5502), .ZN(n4774) );
  NAND2_X1 U6155 ( .A1(n7101), .A2(n7108), .ZN(n7107) );
  NAND2_X1 U6156 ( .A1(n7107), .A2(n4775), .ZN(n6876) );
  NAND2_X1 U6157 ( .A1(n6257), .A2(n4777), .ZN(n4776) );
  OAI211_X1 U6158 ( .C1(n6257), .C2(n4780), .A(n4778), .B(n4776), .ZN(n6265)
         );
  NAND2_X1 U6159 ( .A1(n6257), .A2(n9268), .ZN(n9266) );
  OAI21_X2 U6160 ( .B1(n4791), .B2(n4404), .A(n5044), .ZN(n5695) );
  AOI21_X1 U6161 ( .B1(n5516), .B2(n4797), .A(n4795), .ZN(n4793) );
  INV_X1 U6162 ( .A(n5516), .ZN(n4794) );
  NOR2_X2 U6163 ( .A1(n5358), .A2(n4398), .ZN(n5046) );
  OAI21_X2 U6164 ( .B1(n6841), .B2(n5508), .A(n5657), .ZN(n6829) );
  NAND2_X1 U6165 ( .A1(n5550), .A2(n5534), .ZN(n6841) );
  NAND4_X1 U6166 ( .A1(n4803), .A2(n4355), .A3(n4805), .A4(n4381), .ZN(n5819)
         );
  NAND3_X1 U6167 ( .A1(n6982), .A2(n5788), .A3(n4412), .ZN(n4805) );
  NAND2_X1 U6168 ( .A1(n4812), .A2(n4817), .ZN(P2_U3487) );
  NAND2_X1 U6169 ( .A1(n4818), .A2(n8726), .ZN(n4816) );
  NAND2_X1 U6170 ( .A1(n4825), .A2(n4826), .ZN(n5870) );
  NAND2_X1 U6171 ( .A1(n7563), .A2(n5855), .ZN(n4825) );
  NAND2_X1 U6172 ( .A1(n5722), .A2(n4828), .ZN(n5734) );
  NAND2_X1 U6173 ( .A1(n8762), .A2(n4830), .ZN(n8748) );
  NAND2_X1 U6174 ( .A1(n5004), .A2(n5003), .ZN(n5108) );
  NAND3_X1 U6175 ( .A1(n4838), .A2(n5715), .A3(n5716), .ZN(P1_U3242) );
  NAND2_X1 U6176 ( .A1(n5371), .A2(n5370), .ZN(n4840) );
  NAND2_X1 U6177 ( .A1(n5163), .A2(n4852), .ZN(n4845) );
  NAND2_X1 U6178 ( .A1(n5219), .A2(n4857), .ZN(n4854) );
  NAND2_X1 U6179 ( .A1(n4854), .A2(n4855), .ZN(n5209) );
  NAND2_X1 U6180 ( .A1(n5284), .A2(n4866), .ZN(n4860) );
  OAI21_X1 U6181 ( .B1(n5284), .B2(n4864), .A(n4861), .ZN(n4951) );
  OR2_X1 U6182 ( .A1(n5785), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6183 ( .A1(n6197), .A2(n9880), .ZN(n6187) );
  AND2_X1 U6184 ( .A1(n7729), .A2(n9120), .ZN(n6223) );
  NAND2_X1 U6185 ( .A1(n7494), .A2(n7495), .ZN(n7653) );
  INV_X1 U6186 ( .A(n6091), .ZN(n5778) );
  NOR3_X1 U6187 ( .A1(n8221), .A2(n8220), .A3(n8594), .ZN(n8225) );
  OAI21_X1 U6188 ( .B1(n9285), .B2(n6241), .A(n4875), .ZN(n9265) );
  NAND2_X1 U6189 ( .A1(n5501), .A2(n7100), .ZN(n7103) );
  NAND2_X1 U6190 ( .A1(n4992), .A2(n4991), .ZN(n5128) );
  OR3_X1 U6191 ( .A1(n5635), .A2(n9267), .A3(n6248), .ZN(n5625) );
  NAND2_X2 U6192 ( .A1(n7653), .A2(n5517), .ZN(n7708) );
  OAI21_X1 U6193 ( .B1(n8060), .B2(n8059), .A(n8228), .ZN(n8062) );
  XOR2_X1 U6194 ( .A(n8092), .B(n8060), .Z(n7878) );
  NAND2_X1 U6195 ( .A1(n5768), .A2(n6373), .ZN(n5785) );
  OAI21_X1 U6196 ( .B1(n6373), .B2(n4896), .A(n4895), .ZN(n4897) );
  NAND2_X1 U6197 ( .A1(n4888), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4889) );
  INV_X1 U6198 ( .A(n5739), .ZN(n8939) );
  NAND2_X2 U6199 ( .A1(n5438), .A2(n6376), .ZN(n5446) );
  INV_X1 U6200 ( .A(n8423), .ZN(n8766) );
  AND3_X1 U6201 ( .A1(n6028), .A2(n6027), .A3(n6026), .ZN(n8833) );
  INV_X1 U6202 ( .A(n8833), .ZN(n6029) );
  AND4_X1 U6203 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8705)
         );
  OR2_X1 U6204 ( .A1(n8893), .A2(n8811), .ZN(n4868) );
  INV_X1 U6205 ( .A(n8893), .ZN(n6126) );
  INV_X1 U6206 ( .A(n8662), .ZN(n8905) );
  AND2_X1 U6207 ( .A1(n7784), .A2(n8424), .ZN(n4869) );
  OR2_X1 U6208 ( .A1(n9679), .A2(n9126), .ZN(n4870) );
  OR2_X1 U6209 ( .A1(n9106), .A2(n6226), .ZN(n4871) );
  OR2_X1 U6210 ( .A1(n8285), .A2(n9530), .ZN(n4872) );
  AND2_X1 U6211 ( .A1(n8008), .A2(n8767), .ZN(n4873) );
  OR2_X1 U6212 ( .A1(n9562), .A2(n6240), .ZN(n4875) );
  OR2_X1 U6213 ( .A1(n8285), .A2(n9586), .ZN(n4876) );
  AND2_X1 U6214 ( .A1(n7951), .A2(n7950), .ZN(n4877) );
  AND2_X1 U6215 ( .A1(n8982), .A2(n8981), .ZN(n4878) );
  INV_X1 U6216 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4902) );
  NOR2_X1 U6217 ( .A1(n6198), .A2(n8869), .ZN(n6199) );
  INV_X1 U6218 ( .A(n8908), .ZN(n6019) );
  INV_X1 U6219 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5719) );
  NAND2_X2 U6220 ( .A1(n5740), .A2(n8939), .ZN(n6093) );
  INV_X1 U6221 ( .A(n6093), .ZN(n5805) );
  NAND2_X1 U6222 ( .A1(n5038), .A2(n5035), .ZN(n5036) );
  AND2_X1 U6223 ( .A1(n4933), .A2(n4932), .ZN(n4879) );
  OR2_X1 U6224 ( .A1(n9863), .A2(n10129), .ZN(n4880) );
  OR2_X1 U6225 ( .A1(n5768), .A2(n9760), .ZN(n4881) );
  INV_X1 U6226 ( .A(n9812), .ZN(n5761) );
  AND3_X1 U6227 ( .A1(n5192), .A2(n5287), .A3(n5194), .ZN(n4882) );
  NAND2_X1 U6228 ( .A1(n8112), .A2(n8117), .ZN(n4883) );
  NOR2_X1 U6229 ( .A1(n7530), .A2(n7529), .ZN(n4884) );
  AND2_X1 U6230 ( .A1(n6118), .A2(n8165), .ZN(n4885) );
  NOR2_X1 U6231 ( .A1(n6596), .A2(n6595), .ZN(n9095) );
  INV_X1 U6232 ( .A(n9439), .ZN(n9709) );
  NAND2_X2 U6233 ( .A1(n6957), .A2(n9441), .ZN(n9439) );
  INV_X1 U6234 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5029) );
  INV_X1 U6235 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5973) );
  OR4_X1 U6236 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6169) );
  INV_X1 U6237 ( .A(n9121), .ZN(n6220) );
  INV_X1 U6238 ( .A(n8772), .ZN(n5918) );
  AND2_X1 U6239 ( .A1(n5608), .A2(n5604), .ZN(n6249) );
  INV_X1 U6240 ( .A(n9123), .ZN(n6216) );
  INV_X1 U6241 ( .A(n6308), .ZN(n6302) );
  INV_X1 U6242 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8343) );
  INV_X1 U6243 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5911) );
  OR2_X1 U6244 ( .A1(n6964), .A2(n7971), .ZN(n6565) );
  NOR2_X1 U6245 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  NAND2_X1 U6246 ( .A1(n7965), .A2(n6204), .ZN(n6485) );
  INV_X1 U6247 ( .A(n5312), .ZN(n5068) );
  INV_X1 U6248 ( .A(n7919), .ZN(n7917) );
  INV_X1 U6249 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5251) );
  NOR2_X1 U6250 ( .A1(n7264), .A2(n6216), .ZN(n6217) );
  INV_X1 U6251 ( .A(n9131), .ZN(n6207) );
  INV_X1 U6252 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5047) );
  NOR2_X1 U6253 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5034) );
  INV_X1 U6254 ( .A(n5161), .ZN(n4979) );
  INV_X1 U6255 ( .A(SI_19_), .ZN(n4968) );
  INV_X1 U6256 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5287) );
  INV_X1 U6257 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5861) );
  AND2_X1 U6258 ( .A1(n8359), .A2(n8360), .ZN(n8018) );
  OR2_X1 U6259 ( .A1(n6033), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6035) );
  INV_X1 U6260 ( .A(n7685), .ZN(n7742) );
  INV_X1 U6261 ( .A(n8092), .ZN(n6099) );
  OR2_X1 U6262 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  INV_X1 U6263 ( .A(n7365), .ZN(n8095) );
  NAND2_X1 U6264 ( .A1(n6144), .A2(n6154), .ZN(n6145) );
  NOR2_X1 U6265 ( .A1(n9075), .A2(n8991), .ZN(n8981) );
  OR2_X1 U6266 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  OAI21_X1 U6267 ( .B1(n7971), .B2(n7113), .A(n6485), .ZN(n6486) );
  INV_X1 U6268 ( .A(n5253), .ZN(n5070) );
  NAND2_X1 U6269 ( .A1(n5075), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5133) );
  AND2_X1 U6270 ( .A1(n9220), .A2(n9219), .ZN(n9663) );
  AND2_X1 U6271 ( .A1(n6478), .A2(n6262), .ZN(n6594) );
  NOR2_X1 U6272 ( .A1(n8287), .A2(n8281), .ZN(n6269) );
  NOR2_X1 U6273 ( .A1(n7204), .A2(n6217), .ZN(n6218) );
  AND2_X1 U6274 ( .A1(n6434), .A2(n6594), .ZN(n9070) );
  NAND2_X1 U6275 ( .A1(n4998), .A2(n4997), .ZN(n5119) );
  OR2_X1 U6276 ( .A1(n5272), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5260) );
  AND2_X1 U6277 ( .A1(n5954), .A2(n5953), .ZN(n5998) );
  NAND2_X1 U6278 ( .A1(n8011), .A2(n8853), .ZN(n8012) );
  AND2_X1 U6279 ( .A1(n5976), .A2(n5963), .ZN(n6024) );
  INV_X1 U6280 ( .A(n8409), .ZN(n10131) );
  INV_X1 U6281 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7276) );
  AND2_X1 U6282 ( .A1(n6641), .A2(n6640), .ZN(n8559) );
  NAND2_X1 U6283 ( .A1(n6089), .A2(n6088), .ZN(n6098) );
  INV_X1 U6284 ( .A(n8088), .ZN(n7905) );
  INV_X1 U6285 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U6286 ( .A1(n6163), .A2(n6553), .ZN(n6194) );
  INV_X1 U6287 ( .A(n8143), .ZN(n7749) );
  INV_X1 U6288 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5732) );
  INV_X1 U6289 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6813) );
  OR2_X1 U6290 ( .A1(n5468), .A2(n5072), .ZN(n5202) );
  AND2_X1 U6291 ( .A1(n7945), .A2(n7944), .ZN(n8962) );
  AND2_X1 U6292 ( .A1(n9078), .A2(n9079), .ZN(n7983) );
  OR2_X1 U6293 ( .A1(n8988), .A2(n5180), .ZN(n5095) );
  OR2_X1 U6294 ( .A1(n9258), .A2(n9108), .ZN(n6243) );
  OR2_X1 U6295 ( .A1(n6591), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6289) );
  INV_X1 U6296 ( .A(n6291), .ZN(n8285) );
  INV_X1 U6297 ( .A(n7264), .ZN(n7267) );
  INV_X1 U6298 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5037) );
  AND2_X1 U6299 ( .A1(n4991), .A2(n4990), .ZN(n5140) );
  INV_X1 U6300 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6301 ( .A1(n5187), .A2(n5188), .ZN(n5367) );
  OR2_X1 U6302 ( .A1(n6359), .A2(n6360), .ZN(n10128) );
  INV_X1 U6303 ( .A(n10128), .ZN(n8408) );
  NAND2_X1 U6304 ( .A1(n6356), .A2(n8773), .ZN(n10134) );
  OR2_X1 U6305 ( .A1(n6346), .A2(n7625), .ZN(n6631) );
  AND4_X1 U6306 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n7796)
         );
  INV_X1 U6307 ( .A(n8559), .ZN(n9783) );
  INV_X1 U6308 ( .A(n9804), .ZN(n8773) );
  INV_X1 U6309 ( .A(n8740), .ZN(n8777) );
  NOR2_X1 U6310 ( .A1(n9897), .A2(n6200), .ZN(n6201) );
  AND2_X1 U6311 ( .A1(n9897), .A2(n9877), .ZN(n8835) );
  AND2_X1 U6312 ( .A1(n6191), .A2(n6190), .ZN(n6196) );
  NAND2_X1 U6313 ( .A1(n7573), .A2(n8069), .ZN(n9865) );
  INV_X1 U6314 ( .A(n9865), .ZN(n9877) );
  INV_X1 U6315 ( .A(n9872), .ZN(n9869) );
  XNOR2_X1 U6316 ( .A(n6175), .B(n6174), .ZN(n6369) );
  AND2_X1 U6317 ( .A1(n6159), .A2(n6158), .ZN(n6161) );
  INV_X1 U6318 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5814) );
  AND2_X1 U6319 ( .A1(n6572), .A2(n6571), .ZN(n6625) );
  INV_X1 U6320 ( .A(n9105), .ZN(n9088) );
  AND2_X1 U6321 ( .A1(n5095), .A2(n5094), .ZN(n8978) );
  AND4_X1 U6322 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n7920)
         );
  INV_X1 U6323 ( .A(n9645), .ZN(n9664) );
  AOI21_X1 U6324 ( .B1(n9396), .B2(n6231), .A(n6230), .ZN(n9380) );
  AND2_X1 U6325 ( .A1(n9439), .A2(n9699), .ZN(n9686) );
  NAND2_X1 U6326 ( .A1(n6264), .A2(n6263), .ZN(n9391) );
  NAND2_X1 U6327 ( .A1(n6289), .A2(n9591), .ZN(n6953) );
  INV_X1 U6328 ( .A(n7320), .ZN(n6937) );
  AND2_X1 U6329 ( .A1(n6479), .A2(n9720), .ZN(n9722) );
  INV_X1 U6330 ( .A(n9716), .ZN(n9735) );
  MUX2_X1 U6331 ( .A(n9596), .B(n9592), .S(n6397), .Z(n9719) );
  NAND2_X1 U6332 ( .A1(n4910), .A2(n4909), .ZN(n5395) );
  AND2_X1 U6333 ( .A1(n6376), .A2(P1_U3086), .ZN(n7888) );
  INV_X1 U6334 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10052) );
  INV_X1 U6335 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10100) );
  OR3_X1 U6336 ( .A1(n6343), .A2(n6342), .A3(n6341), .ZN(n8383) );
  AND4_X1 U6337 ( .A1(n7063), .A2(n7062), .A3(n7061), .A4(n7060), .ZN(n8569)
         );
  INV_X1 U6338 ( .A(n8613), .ZN(n8588) );
  INV_X1 U6339 ( .A(n8767), .ZN(n8729) );
  INV_X1 U6340 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10055) );
  OR2_X1 U6341 ( .A1(P2_U3150), .A2(n6639), .ZN(n9768) );
  NAND2_X1 U6342 ( .A1(n6650), .A2(n8251), .ZN(n9778) );
  OR2_X1 U6343 ( .A1(n7139), .A2(n8752), .ZN(n8721) );
  NAND2_X2 U6344 ( .A1(n7139), .A2(n8773), .ZN(n9807) );
  AND2_X1 U6345 ( .A1(n9801), .A2(n7156), .ZN(n8740) );
  INV_X1 U6346 ( .A(n8879), .ZN(n8785) );
  INV_X1 U6347 ( .A(n8835), .ZN(n8869) );
  INV_X1 U6348 ( .A(n9897), .ZN(n9894) );
  INV_X1 U6349 ( .A(n6185), .ZN(n6186) );
  OR2_X1 U6350 ( .A1(n8858), .A2(n8857), .ZN(n8927) );
  AND3_X1 U6351 ( .A1(n9839), .A2(n9838), .A3(n9837), .ZN(n9888) );
  AND2_X1 U6352 ( .A1(n6183), .A2(n6182), .ZN(n9878) );
  AND2_X1 U6353 ( .A1(n6369), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6554) );
  INV_X1 U6354 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7875) );
  INV_X1 U6355 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9927) );
  INV_X1 U6356 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6400) );
  INV_X1 U6357 ( .A(n8941), .ZN(n8937) );
  NAND2_X1 U6358 ( .A1(n8983), .A2(n4878), .ZN(n8996) );
  INV_X1 U6359 ( .A(n9486), .ZN(n9329) );
  INV_X1 U6360 ( .A(n9095), .ZN(n9075) );
  AND2_X1 U6361 ( .A1(n6601), .A2(n9441), .ZN(n9105) );
  INV_X1 U6362 ( .A(n8978), .ZN(n9108) );
  OR2_X1 U6363 ( .A1(n6432), .A2(n6431), .ZN(n9599) );
  INV_X1 U6364 ( .A(n9597), .ZN(n9676) );
  INV_X1 U6365 ( .A(n9686), .ZN(n9247) );
  INV_X1 U6366 ( .A(n9439), .ZN(n9689) );
  NAND2_X1 U6367 ( .A1(n9745), .A2(n9722), .ZN(n9530) );
  INV_X1 U6368 ( .A(n9745), .ZN(n9743) );
  OR2_X1 U6369 ( .A1(n6293), .A2(n6590), .ZN(n7727) );
  NAND2_X1 U6370 ( .A1(n6600), .A2(n6591), .ZN(n9711) );
  INV_X1 U6371 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7623) );
  INV_X1 U6372 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6926) );
  INV_X1 U6373 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U6374 ( .A1(n6373), .A2(P1_U3086), .ZN(n8271) );
  INV_X1 U6375 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10086) );
  INV_X2 U6376 ( .A(n8532), .ZN(P2_U3893) );
  NOR2_X2 U6377 ( .A1(n6605), .A2(n6298), .ZN(P1_U3973) );
  INV_X1 U6378 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6379 ( .A1(n4887), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4888) );
  INV_X1 U6380 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6393) );
  OR2_X1 U6381 ( .A1(n6376), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4892) );
  INV_X1 U6382 ( .A(SI_1_), .ZN(n4893) );
  NAND2_X1 U6383 ( .A1(n5439), .A2(n4893), .ZN(n4898) );
  INV_X1 U6384 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4894) );
  INV_X1 U6385 ( .A(n5439), .ZN(n4899) );
  NAND2_X1 U6386 ( .A1(n4899), .A2(SI_1_), .ZN(n4900) );
  NAND2_X1 U6387 ( .A1(n4901), .A2(n4900), .ZN(n5421) );
  INV_X1 U6388 ( .A(SI_2_), .ZN(n4903) );
  XNOR2_X1 U6389 ( .A(n4904), .B(n4903), .ZN(n5422) );
  NAND2_X1 U6390 ( .A1(n5421), .A2(n5422), .ZN(n4906) );
  NAND2_X1 U6391 ( .A1(n4904), .A2(SI_2_), .ZN(n4905) );
  NAND2_X1 U6392 ( .A1(n4906), .A2(n4905), .ZN(n5379) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6378) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6374) );
  MUX2_X1 U6395 ( .A(n6378), .B(n6374), .S(n6373), .Z(n4907) );
  NAND2_X1 U6396 ( .A1(n5379), .A2(n5378), .ZN(n4910) );
  INV_X1 U6397 ( .A(n4907), .ZN(n4908) );
  NAND2_X1 U6398 ( .A1(n4908), .A2(SI_3_), .ZN(n4909) );
  MUX2_X1 U6399 ( .A(n6390), .B(n6375), .S(n6373), .Z(n4911) );
  XNOR2_X1 U6400 ( .A(n4911), .B(SI_4_), .ZN(n5394) );
  NAND2_X1 U6401 ( .A1(n5395), .A2(n5394), .ZN(n4914) );
  INV_X1 U6402 ( .A(n4911), .ZN(n4912) );
  NAND2_X1 U6403 ( .A1(n4912), .A2(SI_4_), .ZN(n4913) );
  INV_X1 U6404 ( .A(n4915), .ZN(n4916) );
  NAND2_X1 U6405 ( .A1(n4916), .A2(SI_5_), .ZN(n4917) );
  INV_X1 U6406 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6388) );
  INV_X1 U6407 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U6408 ( .A(n4918), .B(SI_6_), .ZN(n5413) );
  INV_X1 U6409 ( .A(n4918), .ZN(n4919) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6384) );
  INV_X1 U6411 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6386) );
  MUX2_X1 U6412 ( .A(n6384), .B(n6386), .S(n6373), .Z(n4920) );
  XNOR2_X1 U6413 ( .A(n4920), .B(SI_7_), .ZN(n5341) );
  INV_X1 U6414 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6415 ( .A1(n4921), .A2(SI_7_), .ZN(n4922) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4923) );
  MUX2_X1 U6417 ( .A(n6400), .B(n4923), .S(n6373), .Z(n4925) );
  INV_X1 U6418 ( .A(SI_8_), .ZN(n4924) );
  NAND2_X1 U6419 ( .A1(n4925), .A2(n4924), .ZN(n4928) );
  INV_X1 U6420 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6421 ( .A1(n4926), .A2(SI_8_), .ZN(n4927) );
  MUX2_X1 U6422 ( .A(n6406), .B(n6408), .S(n6373), .Z(n4930) );
  INV_X1 U6423 ( .A(SI_9_), .ZN(n4929) );
  NAND2_X1 U6424 ( .A1(n4930), .A2(n4929), .ZN(n4933) );
  INV_X1 U6425 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6426 ( .A1(n4931), .A2(SI_9_), .ZN(n4932) );
  INV_X1 U6427 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4935) );
  MUX2_X1 U6428 ( .A(n6410), .B(n4935), .S(n6373), .Z(n4936) );
  XNOR2_X1 U6429 ( .A(n4936), .B(SI_10_), .ZN(n5298) );
  INV_X1 U6430 ( .A(n5298), .ZN(n4939) );
  INV_X1 U6431 ( .A(n4936), .ZN(n4937) );
  NAND2_X1 U6432 ( .A1(n4937), .A2(SI_10_), .ZN(n4938) );
  MUX2_X1 U6433 ( .A(n6414), .B(n6412), .S(n6373), .Z(n4941) );
  INV_X1 U6434 ( .A(SI_11_), .ZN(n4940) );
  NAND2_X1 U6435 ( .A1(n4941), .A2(n4940), .ZN(n4944) );
  INV_X1 U6436 ( .A(n4941), .ZN(n4942) );
  NAND2_X1 U6437 ( .A1(n4942), .A2(SI_11_), .ZN(n4943) );
  NAND2_X1 U6438 ( .A1(n4944), .A2(n4943), .ZN(n5283) );
  MUX2_X1 U6439 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6373), .Z(n4946) );
  INV_X1 U6440 ( .A(SI_12_), .ZN(n4945) );
  XNOR2_X1 U6441 ( .A(n4946), .B(n4945), .ZN(n5270) );
  INV_X1 U6442 ( .A(n5270), .ZN(n4948) );
  NAND2_X1 U6443 ( .A1(n4946), .A2(SI_12_), .ZN(n4947) );
  MUX2_X1 U6444 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6373), .Z(n4949) );
  XNOR2_X1 U6445 ( .A(n4949), .B(SI_13_), .ZN(n5258) );
  NAND2_X1 U6446 ( .A1(n4949), .A2(SI_13_), .ZN(n4950) );
  NAND2_X1 U6447 ( .A1(n4951), .A2(n4950), .ZN(n5247) );
  MUX2_X1 U6448 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6373), .Z(n4953) );
  XNOR2_X1 U6449 ( .A(n4953), .B(SI_14_), .ZN(n5246) );
  INV_X1 U6450 ( .A(n5246), .ZN(n4952) );
  NAND2_X1 U6451 ( .A1(n4953), .A2(SI_14_), .ZN(n4954) );
  MUX2_X1 U6452 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6373), .Z(n5230) );
  NOR2_X1 U6453 ( .A1(n4956), .A2(n4955), .ZN(n4957) );
  MUX2_X1 U6454 ( .A(n6714), .B(n4958), .S(n6373), .Z(n5217) );
  MUX2_X1 U6455 ( .A(n6872), .B(n6874), .S(n6373), .Z(n4961) );
  NAND2_X1 U6456 ( .A1(n4961), .A2(n4960), .ZN(n4964) );
  INV_X1 U6457 ( .A(n4961), .ZN(n4962) );
  NAND2_X1 U6458 ( .A1(n4962), .A2(SI_17_), .ZN(n4963) );
  NAND2_X1 U6459 ( .A1(n4964), .A2(n4963), .ZN(n5455) );
  MUX2_X1 U6460 ( .A(n6924), .B(n6926), .S(n6373), .Z(n4965) );
  XNOR2_X1 U6461 ( .A(n4965), .B(SI_18_), .ZN(n5208) );
  INV_X1 U6462 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6463 ( .A1(n4966), .A2(SI_18_), .ZN(n4967) );
  INV_X1 U6464 ( .A(n5186), .ZN(n4973) );
  MUX2_X1 U6465 ( .A(n7155), .B(n8276), .S(n6373), .Z(n4969) );
  NAND2_X1 U6466 ( .A1(n4969), .A2(n4968), .ZN(n4974) );
  INV_X1 U6467 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U6468 ( .A1(n4970), .A2(SI_19_), .ZN(n4971) );
  NAND2_X1 U6469 ( .A1(n4974), .A2(n4971), .ZN(n5185) );
  INV_X1 U6470 ( .A(n5185), .ZN(n4972) );
  NAND2_X1 U6471 ( .A1(n4973), .A2(n4972), .ZN(n4975) );
  NAND2_X1 U6472 ( .A1(n4975), .A2(n4974), .ZN(n5171) );
  MUX2_X1 U6473 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6373), .Z(n5173) );
  INV_X1 U6474 ( .A(n5173), .ZN(n4976) );
  NAND2_X1 U6475 ( .A1(n5171), .A2(n5172), .ZN(n4977) );
  MUX2_X1 U6476 ( .A(n7492), .B(n7489), .S(n6373), .Z(n5161) );
  NOR2_X1 U6477 ( .A1(n4979), .A2(SI_21_), .ZN(n4981) );
  NAND2_X1 U6478 ( .A1(n4979), .A2(SI_21_), .ZN(n4980) );
  MUX2_X1 U6479 ( .A(n9963), .B(n7576), .S(n6373), .Z(n4983) );
  INV_X1 U6480 ( .A(SI_22_), .ZN(n4982) );
  NAND2_X1 U6481 ( .A1(n4983), .A2(n4982), .ZN(n4986) );
  INV_X1 U6482 ( .A(n4983), .ZN(n4984) );
  NAND2_X1 U6483 ( .A1(n4984), .A2(SI_22_), .ZN(n4985) );
  NAND2_X1 U6484 ( .A1(n4986), .A2(n4985), .ZN(n5153) );
  MUX2_X1 U6485 ( .A(n9927), .B(n7623), .S(n6373), .Z(n4988) );
  INV_X1 U6486 ( .A(SI_23_), .ZN(n4987) );
  NAND2_X1 U6487 ( .A1(n4988), .A2(n4987), .ZN(n4991) );
  INV_X1 U6488 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6489 ( .A1(n4989), .A2(SI_23_), .ZN(n4990) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7808) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7806) );
  MUX2_X1 U6492 ( .A(n7808), .B(n7806), .S(n6373), .Z(n4994) );
  INV_X1 U6493 ( .A(SI_24_), .ZN(n4993) );
  NAND2_X1 U6494 ( .A1(n4994), .A2(n4993), .ZN(n4997) );
  INV_X1 U6495 ( .A(n4994), .ZN(n4995) );
  NAND2_X1 U6496 ( .A1(n4995), .A2(SI_24_), .ZN(n4996) );
  NAND2_X1 U6497 ( .A1(n5128), .A2(n5129), .ZN(n4998) );
  INV_X1 U6498 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9939) );
  INV_X1 U6499 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7865) );
  MUX2_X1 U6500 ( .A(n9939), .B(n7865), .S(n6373), .Z(n5000) );
  INV_X1 U6501 ( .A(SI_25_), .ZN(n4999) );
  NAND2_X1 U6502 ( .A1(n5000), .A2(n4999), .ZN(n5003) );
  INV_X1 U6503 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U6504 ( .A1(n5001), .A2(SI_25_), .ZN(n5002) );
  NAND2_X1 U6505 ( .A1(n5119), .A2(n5120), .ZN(n5004) );
  INV_X1 U6506 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10085) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7869) );
  MUX2_X1 U6508 ( .A(n10085), .B(n7869), .S(n6373), .Z(n5006) );
  INV_X1 U6509 ( .A(SI_26_), .ZN(n5005) );
  NAND2_X1 U6510 ( .A1(n5006), .A2(n5005), .ZN(n5096) );
  INV_X1 U6511 ( .A(n5006), .ZN(n5007) );
  NAND2_X1 U6512 ( .A1(n5007), .A2(SI_26_), .ZN(n5008) );
  INV_X1 U6513 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8051) );
  MUX2_X1 U6514 ( .A(n7875), .B(n8051), .S(n6373), .Z(n5010) );
  INV_X1 U6515 ( .A(SI_27_), .ZN(n5009) );
  NAND2_X1 U6516 ( .A1(n5010), .A2(n5009), .ZN(n5099) );
  INV_X1 U6517 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6518 ( .A1(n5011), .A2(SI_27_), .ZN(n5098) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6373), .Z(n5012) );
  INV_X1 U6520 ( .A(SI_28_), .ZN(n10073) );
  XNOR2_X1 U6521 ( .A(n5012), .B(n10073), .ZN(n5084) );
  NAND2_X1 U6522 ( .A1(n5085), .A2(n5084), .ZN(n5015) );
  INV_X1 U6523 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6524 ( .A1(n5013), .A2(n10073), .ZN(n5014) );
  INV_X1 U6525 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8940) );
  INV_X1 U6526 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7884) );
  MUX2_X1 U6527 ( .A(n8940), .B(n7884), .S(n6373), .Z(n5016) );
  INV_X1 U6528 ( .A(SI_29_), .ZN(n5019) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8272) );
  INV_X1 U6530 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8278) );
  MUX2_X1 U6531 ( .A(n8272), .B(n8278), .S(n6376), .Z(n5021) );
  INV_X1 U6532 ( .A(SI_30_), .ZN(n5020) );
  NAND2_X1 U6533 ( .A1(n5021), .A2(n5020), .ZN(n5024) );
  INV_X1 U6534 ( .A(n5021), .ZN(n5022) );
  NAND2_X1 U6535 ( .A1(n5022), .A2(SI_30_), .ZN(n5023) );
  NAND2_X1 U6536 ( .A1(n5024), .A2(n5023), .ZN(n5056) );
  MUX2_X1 U6537 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6376), .Z(n5025) );
  XNOR2_X1 U6538 ( .A(n5025), .B(SI_31_), .ZN(n5026) );
  MUX2_X1 U6539 ( .A(n5028), .B(n7885), .S(n6373), .Z(n5043) );
  NOR2_X1 U6540 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5031) );
  NOR2_X1 U6541 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5032) );
  NOR2_X2 U6542 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5038) );
  NAND2_X1 U6543 ( .A1(n5037), .A2(n5038), .ZN(n5039) );
  OR2_X2 U6544 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n5039), .ZN(n5040) );
  NAND2_X1 U6545 ( .A1(n5046), .A2(n5041), .ZN(n5044) );
  OAI21_X1 U6546 ( .B1(n5046), .B2(n7886), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n5042) );
  NOR2_X1 U6547 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5045) );
  NAND2_X1 U6548 ( .A1(n5046), .A2(n5045), .ZN(n5051) );
  NAND2_X1 U6549 ( .A1(n5051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6550 ( .A(n5052), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5079) );
  INV_X1 U6551 ( .A(n5079), .ZN(n8270) );
  NAND2_X1 U6552 ( .A1(n5464), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5055) );
  INV_X4 U6554 ( .A(n5373), .ZN(n5469) );
  NAND2_X1 U6555 ( .A1(n5469), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6557 ( .A1(n5463), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5053) );
  NAND3_X1 U6558 ( .A1(n5055), .A2(n5054), .A3(n5053), .ZN(n9238) );
  NAND2_X1 U6559 ( .A1(n8269), .A2(n5457), .ZN(n5059) );
  OR2_X1 U6560 ( .A1(n5446), .A2(n8272), .ZN(n5058) );
  INV_X1 U6561 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U6562 ( .A1(n5469), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6563 ( .A1(n5463), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5060) );
  OAI211_X1 U6564 ( .C1(n5149), .C2(n9462), .A(n5061), .B(n5060), .ZN(n9107)
         );
  INV_X1 U6565 ( .A(n9107), .ZN(n5062) );
  NOR2_X1 U6566 ( .A1(n5642), .A2(n5062), .ZN(n5524) );
  NOR2_X1 U6567 ( .A1(n5706), .A2(n5524), .ZN(n5687) );
  INV_X1 U6568 ( .A(n5687), .ZN(n5483) );
  NOR2_X1 U6569 ( .A1(n9550), .A2(n9107), .ZN(n5523) );
  XNOR2_X1 U6570 ( .A(n5063), .B(SI_29_), .ZN(n7882) );
  NAND2_X1 U6571 ( .A1(n7882), .A2(n5457), .ZN(n5065) );
  OR2_X1 U6572 ( .A1(n5446), .A2(n7884), .ZN(n5064) );
  NAND2_X1 U6573 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5388) );
  INV_X1 U6574 ( .A(n5388), .ZN(n5066) );
  NAND2_X1 U6575 ( .A1(n5066), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5402) );
  INV_X1 U6576 ( .A(n5402), .ZN(n5067) );
  NAND2_X1 U6577 ( .A1(n5067), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6578 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5072) );
  OR2_X2 U6579 ( .A1(n5202), .A2(n10070), .ZN(n5178) );
  INV_X1 U6580 ( .A(n5167), .ZN(n5074) );
  INV_X1 U6581 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8953) );
  INV_X1 U6582 ( .A(n5145), .ZN(n5075) );
  INV_X1 U6583 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9009) );
  OR2_X2 U6584 ( .A1(n5133), .A2(n9009), .ZN(n5124) );
  INV_X1 U6585 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5111) );
  OR2_X2 U6586 ( .A1(n5124), .A2(n5111), .ZN(n5113) );
  INV_X1 U6587 ( .A(n5113), .ZN(n5077) );
  AND2_X1 U6588 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5076) );
  NAND2_X1 U6589 ( .A1(n5077), .A2(n5076), .ZN(n5090) );
  INV_X1 U6590 ( .A(n5090), .ZN(n8282) );
  AND2_X2 U6591 ( .A1(n5079), .A2(n5078), .ZN(n5429) );
  INV_X1 U6592 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6593 ( .A1(n5463), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6594 ( .A1(n5469), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5080) );
  OAI211_X1 U6595 ( .C1(n5149), .C2(n5082), .A(n5081), .B(n5080), .ZN(n5083)
         );
  AOI21_X1 U6596 ( .B1(n8282), .B2(n5362), .A(n5083), .ZN(n8985) );
  OR2_X1 U6597 ( .A1(n6291), .A2(n8985), .ZN(n5639) );
  NAND2_X1 U6598 ( .A1(n6291), .A2(n8985), .ZN(n5638) );
  NAND2_X1 U6599 ( .A1(n8942), .A2(n5457), .ZN(n5087) );
  INV_X1 U6600 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7896) );
  OR2_X1 U6601 ( .A1(n5446), .A2(n7896), .ZN(n5086) );
  INV_X1 U6602 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7999) );
  INV_X1 U6603 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5088) );
  OAI21_X1 U6604 ( .B1(n5113), .B2(n7999), .A(n5088), .ZN(n5089) );
  NAND2_X1 U6605 ( .A1(n5090), .A2(n5089), .ZN(n8988) );
  INV_X1 U6606 ( .A(n5362), .ZN(n5180) );
  INV_X1 U6607 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U6608 ( .A1(n5469), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6609 ( .A1(n5463), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5091) );
  OAI211_X1 U6610 ( .C1(n5149), .C2(n9467), .A(n5092), .B(n5091), .ZN(n5093)
         );
  INV_X1 U6611 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6612 ( .A1(n5633), .A2(n6259), .ZN(n9249) );
  INV_X1 U6613 ( .A(n9249), .ZN(n9251) );
  NAND2_X1 U6614 ( .A1(n5097), .A2(n5096), .ZN(n5101) );
  AND2_X1 U6615 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  NAND2_X1 U6616 ( .A1(n8049), .A2(n5457), .ZN(n5103) );
  OR2_X1 U6617 ( .A1(n5446), .A2(n8051), .ZN(n5102) );
  XNOR2_X1 U6618 ( .A(n5113), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9279) );
  INV_X1 U6619 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U6620 ( .A1(n5463), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6621 ( .A1(n5469), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5104) );
  OAI211_X1 U6622 ( .C1(n5149), .C2(n9472), .A(n5105), .B(n5104), .ZN(n5106)
         );
  AOI21_X1 U6623 ( .B1(n9279), .B2(n5362), .A(n5106), .ZN(n9081) );
  OR2_X1 U6624 ( .A1(n9278), .A2(n9081), .ZN(n5634) );
  NAND2_X1 U6625 ( .A1(n9278), .A2(n9081), .ZN(n6258) );
  XNOR2_X1 U6626 ( .A(n5108), .B(n5107), .ZN(n7868) );
  NAND2_X1 U6627 ( .A1(n7868), .A2(n5457), .ZN(n5110) );
  OR2_X1 U6628 ( .A1(n5446), .A2(n7869), .ZN(n5109) );
  NAND2_X1 U6629 ( .A1(n5124), .A2(n5111), .ZN(n5112) );
  NAND2_X1 U6630 ( .A1(n9294), .A2(n5362), .ZN(n5118) );
  INV_X1 U6631 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U6632 ( .A1(n5469), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6633 ( .A1(n5463), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5114) );
  OAI211_X1 U6634 ( .C1(n5149), .C2(n9477), .A(n5115), .B(n5114), .ZN(n5116)
         );
  INV_X1 U6635 ( .A(n5116), .ZN(n5117) );
  INV_X1 U6636 ( .A(n9109), .ZN(n6240) );
  OR2_X1 U6637 ( .A1(n9293), .A2(n6240), .ZN(n5628) );
  NAND2_X1 U6638 ( .A1(n9293), .A2(n6240), .ZN(n6256) );
  INV_X1 U6639 ( .A(n9286), .ZN(n5480) );
  XNOR2_X1 U6640 ( .A(n5119), .B(n5120), .ZN(n7863) );
  NAND2_X1 U6641 ( .A1(n7863), .A2(n5457), .ZN(n5122) );
  OR2_X1 U6642 ( .A1(n5446), .A2(n7865), .ZN(n5121) );
  INV_X1 U6643 ( .A(n9566), .ZN(n9310) );
  NAND2_X1 U6644 ( .A1(n5133), .A2(n9009), .ZN(n5123) );
  INV_X1 U6645 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U6646 ( .A1(n5463), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6647 ( .A1(n5469), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5125) );
  OAI211_X1 U6648 ( .C1(n5149), .C2(n9482), .A(n5126), .B(n5125), .ZN(n5127)
         );
  AOI21_X1 U6649 ( .B1(n9311), .B2(n5362), .A(n5127), .ZN(n9083) );
  OR2_X1 U6650 ( .A1(n9310), .A2(n9083), .ZN(n5627) );
  NAND2_X1 U6651 ( .A1(n9310), .A2(n9083), .ZN(n6255) );
  NAND2_X1 U6652 ( .A1(n5627), .A2(n6255), .ZN(n9301) );
  XNOR2_X1 U6653 ( .A(n5128), .B(n5129), .ZN(n7805) );
  NAND2_X1 U6654 ( .A1(n7805), .A2(n5457), .ZN(n5131) );
  OR2_X1 U6655 ( .A1(n5446), .A2(n7806), .ZN(n5130) );
  INV_X1 U6656 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U6657 ( .A1(n5145), .A2(n9041), .ZN(n5132) );
  NAND2_X1 U6658 ( .A1(n5133), .A2(n5132), .ZN(n9325) );
  OR2_X1 U6659 ( .A1(n9325), .A2(n5180), .ZN(n5139) );
  INV_X1 U6660 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6661 ( .A1(n5463), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6662 ( .A1(n5469), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5134) );
  OAI211_X1 U6663 ( .C1(n5149), .C2(n5136), .A(n5135), .B(n5134), .ZN(n5137)
         );
  INV_X1 U6664 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6665 ( .A1(n5139), .A2(n5138), .ZN(n9110) );
  INV_X1 U6666 ( .A(n9110), .ZN(n7966) );
  NAND2_X1 U6667 ( .A1(n9486), .A2(n7966), .ZN(n5620) );
  XNOR2_X1 U6668 ( .A(n5141), .B(n5140), .ZN(n7624) );
  NAND2_X1 U6669 ( .A1(n7624), .A2(n5457), .ZN(n5143) );
  OR2_X1 U6670 ( .A1(n5446), .A2(n7623), .ZN(n5142) );
  NAND2_X1 U6671 ( .A1(n5158), .A2(n8953), .ZN(n5144) );
  AND2_X1 U6672 ( .A1(n5145), .A2(n5144), .ZN(n9341) );
  NAND2_X1 U6673 ( .A1(n9341), .A2(n5362), .ZN(n5152) );
  INV_X1 U6674 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6675 ( .A1(n5469), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6676 ( .A1(n5463), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5146) );
  OAI211_X1 U6677 ( .C1(n5149), .C2(n5148), .A(n5147), .B(n5146), .ZN(n5150)
         );
  INV_X1 U6678 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6679 ( .A1(n9491), .A2(n9058), .ZN(n6253) );
  NAND2_X1 U6680 ( .A1(n5618), .A2(n6253), .ZN(n9336) );
  INV_X1 U6681 ( .A(n9336), .ZN(n5478) );
  NAND2_X1 U6682 ( .A1(n7572), .A2(n5457), .ZN(n5156) );
  OR2_X1 U6683 ( .A1(n5446), .A2(n7576), .ZN(n5155) );
  INV_X1 U6684 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9350) );
  INV_X1 U6685 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U6686 ( .A1(n5167), .A2(n9994), .ZN(n5157) );
  NAND2_X1 U6687 ( .A1(n5158), .A2(n5157), .ZN(n9351) );
  OR2_X1 U6688 ( .A1(n9351), .A2(n5180), .ZN(n5160) );
  AOI22_X1 U6689 ( .A1(n5464), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n5463), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5159) );
  OAI211_X1 U6690 ( .C1(n5373), .C2(n9350), .A(n5160), .B(n5159), .ZN(n9112)
         );
  INV_X1 U6691 ( .A(n9112), .ZN(n7956) );
  OR2_X1 U6692 ( .A1(n9349), .A2(n7956), .ZN(n6252) );
  NAND2_X1 U6693 ( .A1(n9349), .A2(n7956), .ZN(n5494) );
  NAND2_X1 U6694 ( .A1(n6252), .A2(n5494), .ZN(n9357) );
  INV_X1 U6695 ( .A(n9357), .ZN(n5477) );
  XNOR2_X1 U6696 ( .A(n5161), .B(SI_21_), .ZN(n5162) );
  XNOR2_X1 U6697 ( .A(n5163), .B(n5162), .ZN(n7488) );
  NAND2_X1 U6698 ( .A1(n7488), .A2(n5457), .ZN(n5165) );
  OR2_X1 U6699 ( .A1(n5446), .A2(n7489), .ZN(n5164) );
  INV_X1 U6700 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U6701 ( .A1(n5178), .A2(n8999), .ZN(n5166) );
  AND2_X1 U6702 ( .A1(n5167), .A2(n5166), .ZN(n9373) );
  NAND2_X1 U6703 ( .A1(n9373), .A2(n5362), .ZN(n5170) );
  AOI22_X1 U6704 ( .A1(n5464), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5469), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6705 ( .A1(n5463), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6706 ( .A1(n9372), .A2(n9057), .ZN(n5608) );
  NAND2_X1 U6707 ( .A1(n9372), .A2(n9057), .ZN(n5609) );
  NAND2_X1 U6708 ( .A1(n5608), .A2(n5609), .ZN(n9365) );
  XNOR2_X1 U6709 ( .A(n5173), .B(n5172), .ZN(n5174) );
  NAND2_X1 U6710 ( .A1(n7364), .A2(n5457), .ZN(n5176) );
  INV_X1 U6711 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7436) );
  OR2_X1 U6712 ( .A1(n5446), .A2(n7436), .ZN(n5175) );
  NAND2_X1 U6713 ( .A1(n5202), .A2(n10070), .ZN(n5177) );
  NAND2_X1 U6714 ( .A1(n5178), .A2(n5177), .ZN(n9383) );
  NAND2_X1 U6715 ( .A1(n5469), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5179) );
  OAI21_X1 U6716 ( .B1(n9383), .B2(n5180), .A(n5179), .ZN(n5184) );
  NAND2_X1 U6717 ( .A1(n5463), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6718 ( .A1(n5464), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6719 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  XNOR2_X1 U6720 ( .A(n9386), .B(n9113), .ZN(n9379) );
  NAND2_X1 U6721 ( .A1(n7154), .A2(n5457), .ZN(n5201) );
  NOR2_X2 U6722 ( .A1(n5367), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6723 ( .A1(n5343), .A2(n5189), .ZN(n5322) );
  NOR2_X1 U6724 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5191) );
  NOR2_X1 U6725 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5190) );
  NAND2_X1 U6726 ( .A1(n5458), .A2(n5194), .ZN(n5195) );
  NAND2_X1 U6727 ( .A1(n5210), .A2(n5196), .ZN(n5197) );
  XNOR2_X2 U6728 ( .A(n5199), .B(n5198), .ZN(n6480) );
  AOI22_X1 U6729 ( .A1(n5460), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5459), .B2(
        n9229), .ZN(n5200) );
  NAND2_X1 U6730 ( .A1(n5464), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5207) );
  INV_X1 U6731 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9071) );
  INV_X1 U6732 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8966) );
  OAI21_X1 U6733 ( .B1(n5468), .B2(n9071), .A(n8966), .ZN(n5203) );
  AND2_X1 U6734 ( .A1(n5203), .A2(n5202), .ZN(n9406) );
  NAND2_X1 U6735 ( .A1(n5362), .A2(n9406), .ZN(n5206) );
  NAND2_X1 U6736 ( .A1(n5469), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6737 ( .A1(n5463), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5204) );
  NAND4_X1 U6738 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n9114)
         );
  INV_X1 U6739 ( .A(n9114), .ZN(n9049) );
  OR2_X1 U6740 ( .A1(n9512), .A2(n9049), .ZN(n5603) );
  NAND2_X1 U6741 ( .A1(n9512), .A2(n9049), .ZN(n5677) );
  NAND2_X1 U6742 ( .A1(n5603), .A2(n5677), .ZN(n9400) );
  XNOR2_X1 U6743 ( .A(n5209), .B(n5208), .ZN(n6923) );
  NAND2_X1 U6744 ( .A1(n6923), .A2(n5457), .ZN(n5212) );
  XNOR2_X1 U6745 ( .A(n5210), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9221) );
  AOI22_X1 U6746 ( .A1(n5460), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5459), .B2(
        n9221), .ZN(n5211) );
  NAND2_X1 U6747 ( .A1(n5464), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6748 ( .A1(n5469), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5215) );
  XNOR2_X1 U6749 ( .A(n5468), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U6750 ( .A1(n5429), .A2(n9421), .ZN(n5214) );
  NAND2_X1 U6751 ( .A1(n5463), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6752 ( .A1(n9420), .A2(n8965), .ZN(n5597) );
  XNOR2_X1 U6753 ( .A(n5217), .B(SI_16_), .ZN(n5218) );
  XNOR2_X1 U6754 ( .A(n5219), .B(n5218), .ZN(n6710) );
  NAND2_X1 U6755 ( .A1(n6710), .A2(n5457), .ZN(n5223) );
  NAND2_X1 U6756 ( .A1(n5220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6757 ( .A(n5221), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7441) );
  AOI22_X1 U6758 ( .A1(n5460), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5459), .B2(
        n7441), .ZN(n5222) );
  NAND2_X1 U6759 ( .A1(n5464), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6760 ( .A1(n5469), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6761 ( .A1(n5241), .A2(n5224), .ZN(n5225) );
  AND2_X1 U6762 ( .A1(n5466), .A2(n5225), .ZN(n9017) );
  NAND2_X1 U6763 ( .A1(n5429), .A2(n9017), .ZN(n5227) );
  NAND2_X1 U6764 ( .A1(n5463), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6765 ( .A1(n9022), .A2(n7920), .ZN(n5590) );
  NAND2_X1 U6766 ( .A1(n9022), .A2(n7920), .ZN(n5671) );
  XNOR2_X1 U6767 ( .A(n5230), .B(SI_15_), .ZN(n5231) );
  XNOR2_X1 U6768 ( .A(n5232), .B(n5231), .ZN(n6662) );
  NAND2_X1 U6769 ( .A1(n6662), .A2(n5457), .ZN(n5239) );
  NOR2_X1 U6770 ( .A1(n5233), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5286) );
  NOR2_X1 U6771 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5234) );
  NAND2_X1 U6772 ( .A1(n5286), .A2(n5234), .ZN(n5272) );
  OAI21_X1 U6773 ( .B1(n5260), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5248) );
  INV_X1 U6774 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6775 ( .A1(n5248), .A2(n5235), .ZN(n5236) );
  NAND2_X1 U6776 ( .A1(n5236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6777 ( .A(n5237), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U6778 ( .A1(n5460), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5459), .B2(
        n9655), .ZN(n5238) );
  NAND2_X1 U6779 ( .A1(n5464), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6780 ( .A1(n5463), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5244) );
  INV_X1 U6781 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U6782 ( .A1(n5253), .A2(n10098), .ZN(n5240) );
  AND2_X1 U6783 ( .A1(n5241), .A2(n5240), .ZN(n9102) );
  NAND2_X1 U6784 ( .A1(n5429), .A2(n9102), .ZN(n5243) );
  NAND2_X1 U6785 ( .A1(n5469), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5242) );
  NAND4_X1 U6786 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n9118)
         );
  INV_X1 U6787 ( .A(n9118), .ZN(n6226) );
  OR2_X1 U6788 ( .A1(n9532), .A2(n6226), .ZN(n5583) );
  NAND2_X1 U6789 ( .A1(n9532), .A2(n6226), .ZN(n5580) );
  NAND2_X1 U6790 ( .A1(n5583), .A2(n5580), .ZN(n7641) );
  XNOR2_X1 U6791 ( .A(n5247), .B(n5246), .ZN(n6621) );
  NAND2_X1 U6792 ( .A1(n6621), .A2(n5457), .ZN(n5250) );
  XNOR2_X1 U6793 ( .A(n5248), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9633) );
  AOI22_X1 U6794 ( .A1(n5460), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5459), .B2(
        n9633), .ZN(n5249) );
  NAND2_X1 U6795 ( .A1(n5464), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6796 ( .A1(n5469), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6797 ( .A1(n5265), .A2(n5251), .ZN(n5252) );
  AND2_X1 U6798 ( .A1(n5253), .A2(n5252), .ZN(n7716) );
  NAND2_X1 U6799 ( .A1(n5362), .A2(n7716), .ZN(n5255) );
  NAND2_X1 U6800 ( .A1(n5463), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5254) );
  NAND4_X1 U6801 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n9119)
         );
  INV_X1 U6802 ( .A(n9119), .ZN(n7536) );
  OR2_X1 U6803 ( .A1(n9538), .A2(n7536), .ZN(n5667) );
  NAND2_X1 U6804 ( .A1(n9538), .A2(n7536), .ZN(n5581) );
  NAND2_X1 U6805 ( .A1(n5667), .A2(n5581), .ZN(n7704) );
  XNOR2_X1 U6806 ( .A(n5259), .B(n5258), .ZN(n6557) );
  NAND2_X1 U6807 ( .A1(n6557), .A2(n5457), .ZN(n5263) );
  NAND2_X1 U6808 ( .A1(n5260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6809 ( .A(n5261), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9624) );
  AOI22_X1 U6810 ( .A1(n5460), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5459), .B2(
        n9624), .ZN(n5262) );
  NAND2_X1 U6811 ( .A1(n5463), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6812 ( .A1(n5464), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6813 ( .A1(n5278), .A2(n7393), .ZN(n5264) );
  AND2_X1 U6814 ( .A1(n5265), .A2(n5264), .ZN(n7660) );
  NAND2_X1 U6815 ( .A1(n5362), .A2(n7660), .ZN(n5267) );
  NAND2_X1 U6816 ( .A1(n5469), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6817 ( .A1(n7729), .A2(n7545), .ZN(n7707) );
  NAND2_X1 U6818 ( .A1(n5666), .A2(n7707), .ZN(n7656) );
  XNOR2_X1 U6819 ( .A(n5271), .B(n5270), .ZN(n6544) );
  NAND2_X1 U6820 ( .A1(n6544), .A2(n5457), .ZN(n5275) );
  NAND2_X1 U6821 ( .A1(n5272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6822 ( .A(n5273), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7126) );
  AOI22_X1 U6823 ( .A1(n5460), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5459), .B2(
        n7126), .ZN(n5274) );
  NAND2_X1 U6824 ( .A1(n5464), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6825 ( .A1(n5463), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5281) );
  INV_X1 U6826 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6827 ( .A1(n5293), .A2(n5276), .ZN(n5277) );
  AND2_X1 U6828 ( .A1(n5278), .A2(n5277), .ZN(n7499) );
  NAND2_X1 U6829 ( .A1(n5429), .A2(n7499), .ZN(n5280) );
  NAND2_X1 U6830 ( .A1(n5469), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5279) );
  NAND4_X1 U6831 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n9121)
         );
  OR2_X1 U6832 ( .A1(n7235), .A2(n6220), .ZN(n7652) );
  NAND2_X1 U6833 ( .A1(n7235), .A2(n6220), .ZN(n5568) );
  NAND2_X1 U6834 ( .A1(n6411), .A2(n5457), .ZN(n5291) );
  OR2_X1 U6835 ( .A1(n5286), .A2(n7886), .ZN(n5300) );
  NAND2_X1 U6836 ( .A1(n5300), .A2(n5287), .ZN(n5288) );
  NAND2_X1 U6837 ( .A1(n5288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6838 ( .A(n5289), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6538) );
  AOI22_X1 U6839 ( .A1(n5460), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5459), .B2(
        n6538), .ZN(n5290) );
  NAND2_X1 U6840 ( .A1(n5464), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6841 ( .A1(n5469), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6842 ( .A1(n5305), .A2(n7314), .ZN(n5292) );
  AND2_X1 U6843 ( .A1(n5293), .A2(n5292), .ZN(n7481) );
  NAND2_X1 U6844 ( .A1(n5362), .A2(n7481), .ZN(n5295) );
  NAND2_X1 U6845 ( .A1(n5463), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5294) );
  NAND4_X1 U6846 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n9122)
         );
  INV_X1 U6847 ( .A(n9122), .ZN(n6219) );
  NAND2_X1 U6848 ( .A1(n7463), .A2(n6219), .ZN(n5567) );
  XNOR2_X1 U6849 ( .A(n5299), .B(n5298), .ZN(n6403) );
  NAND2_X1 U6850 ( .A1(n6403), .A2(n5457), .ZN(n5302) );
  XNOR2_X1 U6851 ( .A(n5300), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6533) );
  AOI22_X1 U6852 ( .A1(n5460), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5459), .B2(
        n6533), .ZN(n5301) );
  NAND2_X1 U6853 ( .A1(n5302), .A2(n5301), .ZN(n7264) );
  NAND2_X1 U6854 ( .A1(n5464), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6855 ( .A1(n5463), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5308) );
  INV_X1 U6856 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6857 ( .A1(n5312), .A2(n5303), .ZN(n5304) );
  AND2_X1 U6858 ( .A1(n5305), .A2(n5304), .ZN(n7208) );
  NAND2_X1 U6859 ( .A1(n5429), .A2(n7208), .ZN(n5307) );
  NAND2_X1 U6860 ( .A1(n5469), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6861 ( .A1(n7264), .A2(n9123), .ZN(n5563) );
  NAND2_X1 U6862 ( .A1(n5567), .A2(n5563), .ZN(n5558) );
  INV_X1 U6863 ( .A(n5558), .ZN(n5453) );
  OR2_X1 U6864 ( .A1(n7463), .A2(n6219), .ZN(n5557) );
  OR2_X1 U6865 ( .A1(n7264), .A2(n9123), .ZN(n5515) );
  AND2_X1 U6866 ( .A1(n5557), .A2(n5515), .ZN(n5663) );
  NAND2_X1 U6867 ( .A1(n5463), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6868 ( .A1(n5464), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6869 ( .A1(n5329), .A2(n5310), .ZN(n5311) );
  AND2_X1 U6870 ( .A1(n5312), .A2(n5311), .ZN(n7252) );
  NAND2_X1 U6871 ( .A1(n5362), .A2(n7252), .ZN(n5314) );
  NAND2_X1 U6872 ( .A1(n5469), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U6873 ( .A(n5317), .B(n4879), .ZN(n6405) );
  NAND2_X1 U6874 ( .A1(n6405), .A2(n5457), .ZN(n5320) );
  NAND2_X1 U6875 ( .A1(n5233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6876 ( .A(n5318), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6467) );
  AOI22_X1 U6877 ( .A1(n5460), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5459), .B2(
        n6467), .ZN(n5319) );
  OR2_X1 U6878 ( .A1(n7192), .A2(n9432), .ZN(n5562) );
  NAND2_X1 U6879 ( .A1(n9432), .A2(n7192), .ZN(n5555) );
  NAND2_X1 U6880 ( .A1(n5562), .A2(n5555), .ZN(n7039) );
  XNOR2_X1 U6881 ( .A(n5321), .B(n4376), .ZN(n6399) );
  OR2_X1 U6882 ( .A1(n6399), .A2(n5442), .ZN(n5326) );
  NAND2_X1 U6883 ( .A1(n5322), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5323) );
  MUX2_X1 U6884 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5323), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5324) );
  AND2_X1 U6885 ( .A1(n5324), .A2(n5233), .ZN(n9201) );
  AOI22_X1 U6886 ( .A1(n5460), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5459), .B2(
        n9201), .ZN(n5325) );
  INV_X1 U6887 ( .A(n9445), .ZN(n7011) );
  NAND2_X1 U6888 ( .A1(n5463), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6889 ( .A1(n5464), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6890 ( .A1(n5336), .A2(n5327), .ZN(n5328) );
  NAND2_X1 U6891 ( .A1(n5329), .A2(n5328), .ZN(n9442) );
  INV_X1 U6892 ( .A(n9442), .ZN(n5330) );
  NAND2_X1 U6893 ( .A1(n5429), .A2(n5330), .ZN(n5332) );
  NAND2_X1 U6894 ( .A1(n5469), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5331) );
  INV_X1 U6895 ( .A(n7041), .ZN(n9125) );
  NAND2_X1 U6896 ( .A1(n7011), .A2(n9125), .ZN(n7004) );
  NAND2_X1 U6897 ( .A1(n5404), .A2(n6813), .ZN(n5335) );
  AND2_X1 U6898 ( .A1(n5336), .A2(n5335), .ZN(n9677) );
  NAND2_X1 U6899 ( .A1(n5362), .A2(n9677), .ZN(n5340) );
  NAND2_X1 U6900 ( .A1(n5464), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6901 ( .A1(n5469), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6902 ( .A1(n5463), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5337) );
  NAND4_X1 U6903 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(n9126)
         );
  XNOR2_X1 U6904 ( .A(n5342), .B(n5341), .ZN(n6385) );
  OR2_X1 U6905 ( .A1(n6385), .A2(n5442), .ZN(n5349) );
  INV_X1 U6906 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U6907 ( .A1(n5344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5410) );
  INV_X1 U6908 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6909 ( .A1(n5410), .A2(n5409), .ZN(n5412) );
  NAND2_X1 U6910 ( .A1(n5412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5346) );
  INV_X1 U6911 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U6912 ( .A(n5346), .B(n5345), .ZN(n9184) );
  OR2_X1 U6913 ( .A1(n6397), .A2(n9184), .ZN(n5348) );
  OR2_X1 U6914 ( .A1(n5446), .A2(n6386), .ZN(n5347) );
  NAND2_X1 U6915 ( .A1(n9126), .A2(n7096), .ZN(n5350) );
  NAND2_X1 U6916 ( .A1(n5429), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6917 ( .A1(n5428), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6918 ( .A1(n5430), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6919 ( .A1(n5431), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5351) );
  INV_X1 U6920 ( .A(SI_0_), .ZN(n5355) );
  NOR2_X1 U6921 ( .A1(n6376), .A2(n5355), .ZN(n5356) );
  XNOR2_X1 U6922 ( .A(n5356), .B(n4894), .ZN(n9592) );
  INV_X1 U6923 ( .A(n9719), .ZN(n7113) );
  NAND2_X1 U6924 ( .A1(n6204), .A2(n7113), .ZN(n5656) );
  INV_X1 U6925 ( .A(n5656), .ZN(n5357) );
  NOR2_X1 U6926 ( .A1(n6204), .A2(n7113), .ZN(n7100) );
  OR2_X1 U6927 ( .A1(n5357), .A2(n7100), .ZN(n9713) );
  NAND2_X1 U6928 ( .A1(n5358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6929 ( .A1(n5464), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6930 ( .A1(n5463), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5365) );
  INV_X1 U6931 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6932 ( .A1(n5388), .A2(n5360), .ZN(n5361) );
  AND2_X1 U6933 ( .A1(n5402), .A2(n5361), .ZN(n7471) );
  NAND2_X1 U6934 ( .A1(n5362), .A2(n7471), .ZN(n5364) );
  NAND2_X1 U6935 ( .A1(n5469), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6936 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5369) );
  INV_X1 U6937 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5368) );
  XNOR2_X1 U6938 ( .A(n5369), .B(n5368), .ZN(n6445) );
  OR2_X1 U6939 ( .A1(n5446), .A2(n6381), .ZN(n5372) );
  NAND2_X1 U6940 ( .A1(n6830), .A2(n6940), .ZN(n5536) );
  INV_X1 U6941 ( .A(n6830), .ZN(n9128) );
  NAND2_X1 U6942 ( .A1(n9128), .A2(n7474), .ZN(n5657) );
  NAND2_X1 U6943 ( .A1(n5536), .A2(n5657), .ZN(n6840) );
  NOR3_X1 U6944 ( .A1(n9713), .A2(n6262), .A3(n6840), .ZN(n5450) );
  NAND2_X1 U6945 ( .A1(n5428), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6946 ( .A1(n5469), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6947 ( .A1(n5431), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5375) );
  INV_X1 U6948 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U6949 ( .A1(n5429), .A2(n6961), .ZN(n5374) );
  OR2_X1 U6950 ( .A1(n5446), .A2(n6374), .ZN(n5386) );
  XNOR2_X1 U6951 ( .A(n5379), .B(n5378), .ZN(n6377) );
  OR2_X1 U6952 ( .A1(n5442), .A2(n6377), .ZN(n5385) );
  OR2_X1 U6953 ( .A1(n5380), .A2(n7886), .ZN(n5424) );
  NAND2_X1 U6954 ( .A1(n5424), .A2(n5381), .ZN(n5423) );
  NAND2_X1 U6955 ( .A1(n5423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5383) );
  INV_X1 U6956 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5382) );
  XNOR2_X1 U6957 ( .A(n5383), .B(n5382), .ZN(n6441) );
  OR2_X1 U6958 ( .A1(n6397), .A2(n6441), .ZN(n5384) );
  XNOR2_X1 U6959 ( .A(n9130), .B(n6964), .ZN(n6864) );
  NAND2_X1 U6960 ( .A1(n5463), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6961 ( .A1(n5464), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5392) );
  INV_X1 U6962 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6963 ( .A1(n6961), .A2(n5387), .ZN(n5389) );
  AND2_X1 U6964 ( .A1(n5389), .A2(n5388), .ZN(n6720) );
  NAND2_X1 U6965 ( .A1(n5429), .A2(n6720), .ZN(n5391) );
  NAND2_X1 U6966 ( .A1(n5469), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U6967 ( .A(n5395), .B(n5394), .ZN(n6389) );
  OR2_X1 U6968 ( .A1(n5442), .A2(n6389), .ZN(n5400) );
  OR2_X1 U6969 ( .A1(n5446), .A2(n6375), .ZN(n5399) );
  OAI21_X1 U6970 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6971 ( .A1(n5424), .A2(n5396), .ZN(n5397) );
  XNOR2_X1 U6972 ( .A(n5397), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6443) );
  OR2_X1 U6973 ( .A1(n6397), .A2(n6443), .ZN(n5398) );
  XNOR2_X1 U6974 ( .A(n9129), .B(n7320), .ZN(n6852) );
  NAND2_X1 U6975 ( .A1(n5463), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6976 ( .A1(n5464), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5407) );
  INV_X1 U6977 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6978 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  AND2_X1 U6979 ( .A1(n5404), .A2(n5403), .ZN(n9688) );
  NAND2_X1 U6980 ( .A1(n5362), .A2(n9688), .ZN(n5406) );
  NAND2_X1 U6981 ( .A1(n5469), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5405) );
  OR2_X1 U6982 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  NAND2_X1 U6983 ( .A1(n5412), .A2(n5411), .ZN(n9170) );
  XNOR2_X1 U6984 ( .A(n5414), .B(n5413), .ZN(n6387) );
  OR2_X1 U6985 ( .A1(n5442), .A2(n6387), .ZN(n5416) );
  OR2_X1 U6986 ( .A1(n5446), .A2(n6382), .ZN(n5415) );
  OAI211_X1 U6987 ( .C1(n6397), .C2(n9170), .A(n5416), .B(n5415), .ZN(n6934)
         );
  NAND2_X1 U6988 ( .A1(n6795), .A2(n6934), .ZN(n5535) );
  NAND2_X1 U6989 ( .A1(n9127), .A2(n9693), .ZN(n6996) );
  NAND2_X1 U6990 ( .A1(n5535), .A2(n6996), .ZN(n6828) );
  NOR3_X1 U6991 ( .A1(n6864), .A2(n6852), .A3(n6828), .ZN(n5449) );
  NAND2_X1 U6992 ( .A1(n5428), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6993 ( .A1(n5429), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6994 ( .A1(n5430), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6995 ( .A1(n5431), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5417) );
  OR2_X1 U6996 ( .A1(n5446), .A2(n4538), .ZN(n5427) );
  XNOR2_X1 U6997 ( .A(n5422), .B(n5421), .ZN(n6391) );
  OR2_X1 U6998 ( .A1(n5442), .A2(n6391), .ZN(n5426) );
  OAI21_X1 U6999 ( .B1(n5424), .B2(n5381), .A(n5423), .ZN(n6436) );
  OR2_X1 U7000 ( .A1(n6397), .A2(n6436), .ZN(n5425) );
  INV_X1 U7001 ( .A(n6881), .ZN(n5503) );
  NAND2_X1 U7002 ( .A1(n5428), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U7003 ( .A1(n5429), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U7004 ( .A1(n5430), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7005 ( .A1(n5431), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5432) );
  NAND4_X2 U7006 ( .A1(n5435), .A2(n5432), .A3(n5433), .A4(n5434), .ZN(n5502)
         );
  INV_X1 U7007 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7008 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9596), .ZN(n5436) );
  XNOR2_X1 U7009 ( .A(n5437), .B(n5436), .ZN(n6438) );
  OR2_X1 U7010 ( .A1(n5438), .A2(n6438), .ZN(n5444) );
  XNOR2_X1 U7011 ( .A(n5439), .B(SI_1_), .ZN(n5440) );
  XNOR2_X1 U7012 ( .A(n5441), .B(n5440), .ZN(n5758) );
  INV_X1 U7013 ( .A(n5758), .ZN(n6392) );
  INV_X1 U7014 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5445) );
  INV_X1 U7015 ( .A(n6205), .ZN(n5501) );
  NAND4_X1 U7016 ( .A1(n5450), .A2(n5449), .A3(n5503), .A4(n5501), .ZN(n5451)
         );
  NAND2_X1 U7017 ( .A1(n7041), .A2(n9445), .ZN(n6214) );
  INV_X1 U7018 ( .A(n9126), .ZN(n6831) );
  INV_X1 U7019 ( .A(n7096), .ZN(n9679) );
  NAND2_X1 U7020 ( .A1(n6831), .A2(n9679), .ZN(n7001) );
  NAND2_X1 U7021 ( .A1(n6214), .A2(n7001), .ZN(n6998) );
  NOR4_X1 U7022 ( .A1(n7039), .A2(n4520), .A3(n5451), .A4(n6998), .ZN(n5452)
         );
  NAND4_X1 U7023 ( .A1(n7495), .A2(n5453), .A3(n5663), .A4(n5452), .ZN(n5454)
         );
  NOR4_X1 U7024 ( .A1(n7641), .A2(n7704), .A3(n7656), .A4(n5454), .ZN(n5474)
         );
  XNOR2_X1 U7025 ( .A(n5456), .B(n5455), .ZN(n6871) );
  NAND2_X1 U7026 ( .A1(n6871), .A2(n5457), .ZN(n5462) );
  XNOR2_X1 U7027 ( .A(n5458), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9218) );
  AOI22_X1 U7028 ( .A1(n5460), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5459), .B2(
        n9218), .ZN(n5461) );
  NAND2_X1 U7029 ( .A1(n5463), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7030 ( .A1(n5464), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5472) );
  INV_X1 U7031 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7032 ( .A1(n5466), .A2(n5465), .ZN(n5467) );
  AND2_X1 U7033 ( .A1(n5468), .A2(n5467), .ZN(n9027) );
  NAND2_X1 U7034 ( .A1(n5362), .A2(n9027), .ZN(n5471) );
  NAND2_X1 U7035 ( .A1(n5469), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5470) );
  NAND4_X1 U7036 ( .A1(n5473), .A2(n5472), .A3(n5471), .A4(n5470), .ZN(n9116)
         );
  INV_X1 U7037 ( .A(n9116), .ZN(n7930) );
  XNOR2_X1 U7038 ( .A(n9521), .B(n7930), .ZN(n5519) );
  NAND4_X1 U7039 ( .A1(n9413), .A2(n4393), .A3(n5474), .A4(n7855), .ZN(n5475)
         );
  NOR4_X1 U7040 ( .A1(n9365), .A2(n9379), .A3(n9400), .A4(n5475), .ZN(n5476)
         );
  NAND4_X1 U7041 ( .A1(n9319), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n5479)
         );
  NOR3_X1 U7042 ( .A1(n5480), .A2(n9301), .A3(n5479), .ZN(n5481) );
  NAND4_X1 U7043 ( .A1(n6260), .A2(n9251), .A3(n9268), .A4(n5481), .ZN(n5482)
         );
  INV_X1 U7044 ( .A(n5648), .ZN(n5533) );
  INV_X1 U7045 ( .A(n5706), .ZN(n5531) );
  INV_X1 U7046 ( .A(n5486), .ZN(n5484) );
  NAND2_X1 U7047 ( .A1(n5484), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7048 ( .A1(n5618), .A2(n6252), .ZN(n5616) );
  NAND2_X1 U7049 ( .A1(n5616), .A2(n6253), .ZN(n5488) );
  NAND2_X1 U7050 ( .A1(n6254), .A2(n5488), .ZN(n5489) );
  NAND2_X1 U7051 ( .A1(n5489), .A2(n5620), .ZN(n5490) );
  AND2_X1 U7052 ( .A1(n5627), .A2(n5490), .ZN(n5497) );
  INV_X1 U7053 ( .A(n5497), .ZN(n5492) );
  OR2_X1 U7054 ( .A1(n9505), .A2(n7947), .ZN(n5604) );
  INV_X1 U7055 ( .A(n6249), .ZN(n5491) );
  OR2_X1 U7056 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  NAND2_X1 U7057 ( .A1(n5634), .A2(n5628), .ZN(n5498) );
  AOI21_X1 U7058 ( .B1(n6256), .B2(n5493), .A(n5498), .ZN(n5500) );
  AND2_X1 U7059 ( .A1(n6253), .A2(n5494), .ZN(n5614) );
  AND2_X1 U7060 ( .A1(n9505), .A2(n7947), .ZN(n5606) );
  NAND2_X1 U7061 ( .A1(n5608), .A2(n5606), .ZN(n5495) );
  AND2_X1 U7062 ( .A1(n5495), .A2(n5609), .ZN(n6250) );
  NAND3_X1 U7063 ( .A1(n5620), .A2(n5614), .A3(n6250), .ZN(n5496) );
  INV_X1 U7064 ( .A(n6255), .ZN(n5630) );
  AOI21_X1 U7065 ( .B1(n5497), .B2(n5496), .A(n5630), .ZN(n5499) );
  OAI21_X1 U7066 ( .B1(n5499), .B2(n5498), .A(n5624), .ZN(n5681) );
  OAI211_X1 U7067 ( .C1(n5500), .C2(n5681), .A(n5639), .B(n5633), .ZN(n5683)
         );
  INV_X1 U7068 ( .A(n6256), .ZN(n9267) );
  INV_X1 U7069 ( .A(n5502), .ZN(n6206) );
  NAND2_X1 U7070 ( .A1(n6206), .A2(n7117), .ZN(n6880) );
  NAND2_X1 U7071 ( .A1(n7103), .A2(n6880), .ZN(n5504) );
  NAND2_X1 U7072 ( .A1(n6207), .A2(n7050), .ZN(n5505) );
  NAND2_X1 U7073 ( .A1(n6883), .A2(n5505), .ZN(n6865) );
  NAND2_X1 U7074 ( .A1(n9130), .A2(n6964), .ZN(n5653) );
  NAND2_X1 U7075 ( .A1(n6865), .A2(n5653), .ZN(n5507) );
  INV_X1 U7076 ( .A(n6964), .ZN(n6863) );
  NAND2_X1 U7077 ( .A1(n6209), .A2(n6863), .ZN(n5506) );
  NAND2_X1 U7078 ( .A1(n5507), .A2(n5506), .ZN(n6853) );
  NAND2_X1 U7079 ( .A1(n9129), .A2(n7320), .ZN(n5655) );
  INV_X1 U7080 ( .A(n9129), .ZN(n6784) );
  NAND2_X1 U7081 ( .A1(n6784), .A2(n6937), .ZN(n5534) );
  INV_X1 U7082 ( .A(n5536), .ZN(n5508) );
  INV_X1 U7083 ( .A(n5555), .ZN(n5509) );
  OR2_X1 U7084 ( .A1(n5509), .A2(n6998), .ZN(n5510) );
  OR2_X2 U7085 ( .A1(n6997), .A2(n5510), .ZN(n5514) );
  NAND2_X1 U7086 ( .A1(n6998), .A2(n7004), .ZN(n5511) );
  NAND2_X1 U7087 ( .A1(n5511), .A2(n5555), .ZN(n5512) );
  NAND2_X1 U7088 ( .A1(n5512), .A2(n5562), .ZN(n5660) );
  NAND3_X1 U7089 ( .A1(n5554), .A2(n5562), .A3(n6996), .ZN(n5513) );
  NAND2_X1 U7090 ( .A1(n5660), .A2(n5513), .ZN(n5662) );
  NAND2_X1 U7091 ( .A1(n5515), .A2(n5563), .ZN(n7206) );
  INV_X1 U7092 ( .A(n7206), .ZN(n7200) );
  NAND2_X1 U7093 ( .A1(n5557), .A2(n5567), .ZN(n7456) );
  INV_X1 U7094 ( .A(n5563), .ZN(n7457) );
  NOR2_X1 U7095 ( .A1(n7456), .A2(n7457), .ZN(n5516) );
  INV_X1 U7096 ( .A(n7652), .ZN(n5569) );
  NOR2_X1 U7097 ( .A1(n7656), .A2(n5569), .ZN(n5517) );
  INV_X1 U7098 ( .A(n7707), .ZN(n5578) );
  NOR2_X1 U7099 ( .A1(n7704), .A2(n5578), .ZN(n5574) );
  NAND2_X1 U7100 ( .A1(n7708), .A2(n5574), .ZN(n7640) );
  INV_X1 U7101 ( .A(n5667), .ZN(n7642) );
  NOR2_X1 U7102 ( .A1(n7641), .A2(n7642), .ZN(n5518) );
  NAND2_X1 U7103 ( .A1(n7643), .A2(n5580), .ZN(n7840) );
  OR2_X1 U7104 ( .A1(n9521), .A2(n7930), .ZN(n5595) );
  NOR3_X1 U7105 ( .A1(n5681), .A2(n9267), .A3(n9389), .ZN(n5521) );
  NOR2_X1 U7106 ( .A1(n5683), .A2(n5521), .ZN(n5528) );
  INV_X1 U7107 ( .A(n5638), .ZN(n5522) );
  NOR2_X1 U7108 ( .A1(n5523), .A2(n5522), .ZN(n5682) );
  INV_X1 U7109 ( .A(n5682), .ZN(n5527) );
  INV_X1 U7110 ( .A(n5524), .ZN(n5526) );
  INV_X1 U7111 ( .A(n9238), .ZN(n5525) );
  OAI22_X1 U7112 ( .A1(n5528), .A2(n5527), .B1(n5526), .B2(n5525), .ZN(n5529)
         );
  OAI211_X1 U7113 ( .C1(n9550), .C2(n9238), .A(n5529), .B(n5711), .ZN(n5530)
         );
  NAND3_X1 U7114 ( .A1(n5531), .A2(n6594), .A3(n5530), .ZN(n5532) );
  NAND2_X1 U7115 ( .A1(n5533), .A2(n5532), .ZN(n5650) );
  NAND4_X1 U7116 ( .A1(n6841), .A2(n6248), .A3(n5657), .A4(n6996), .ZN(n5552)
         );
  AND4_X1 U7117 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5707), .ZN(n5549)
         );
  NAND2_X1 U7118 ( .A1(n6830), .A2(n6248), .ZN(n5542) );
  OAI21_X1 U7119 ( .B1(n5542), .B2(n9127), .A(n6940), .ZN(n5538) );
  OR2_X1 U7120 ( .A1(n6830), .A2(n6248), .ZN(n5539) );
  INV_X1 U7121 ( .A(n6940), .ZN(n7474) );
  OAI21_X1 U7122 ( .B1(n5539), .B2(n6795), .A(n7474), .ZN(n5537) );
  NAND2_X1 U7123 ( .A1(n5538), .A2(n5537), .ZN(n5547) );
  OAI22_X1 U7124 ( .A1(n5539), .A2(n6940), .B1(n6795), .B2(n6248), .ZN(n5540)
         );
  NAND2_X1 U7125 ( .A1(n5540), .A2(n9693), .ZN(n5546) );
  XNOR2_X1 U7126 ( .A(n9126), .B(n7096), .ZN(n7089) );
  INV_X1 U7127 ( .A(n7089), .ZN(n5545) );
  NAND2_X1 U7128 ( .A1(n6795), .A2(n6248), .ZN(n5541) );
  OAI21_X1 U7129 ( .B1(n5542), .B2(n7474), .A(n5541), .ZN(n5543) );
  NAND2_X1 U7130 ( .A1(n5543), .A2(n6934), .ZN(n5544) );
  NAND4_X1 U7131 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n5548)
         );
  AOI21_X1 U7132 ( .B1(n5550), .B2(n5549), .A(n5548), .ZN(n5551) );
  INV_X1 U7133 ( .A(n7004), .ZN(n7037) );
  NAND2_X1 U7134 ( .A1(n5555), .A2(n6214), .ZN(n5553) );
  NAND2_X1 U7135 ( .A1(n5565), .A2(n5562), .ZN(n5556) );
  NAND2_X1 U7136 ( .A1(n5556), .A2(n5555), .ZN(n5561) );
  AND2_X1 U7137 ( .A1(n7652), .A2(n5663), .ZN(n5560) );
  NAND3_X1 U7138 ( .A1(n7652), .A2(n5558), .A3(n5557), .ZN(n5559) );
  NAND2_X1 U7139 ( .A1(n5559), .A2(n5568), .ZN(n5668) );
  AOI21_X1 U7140 ( .B1(n5561), .B2(n5560), .A(n5668), .ZN(n5573) );
  INV_X1 U7141 ( .A(n5562), .ZN(n5564) );
  NAND2_X1 U7142 ( .A1(n5566), .A2(n5663), .ZN(n5571) );
  AND2_X1 U7143 ( .A1(n5568), .A2(n5567), .ZN(n5570) );
  AOI21_X1 U7144 ( .B1(n5571), .B2(n5570), .A(n5569), .ZN(n5572) );
  MUX2_X1 U7145 ( .A(n5573), .B(n5572), .S(n6248), .Z(n5579) );
  INV_X1 U7146 ( .A(n5666), .ZN(n5575) );
  OAI21_X1 U7147 ( .B1(n5579), .B2(n5575), .A(n5574), .ZN(n5577) );
  NAND2_X1 U7148 ( .A1(n5590), .A2(n5583), .ZN(n5670) );
  INV_X1 U7149 ( .A(n5670), .ZN(n5576) );
  NAND3_X1 U7150 ( .A1(n5577), .A2(n5576), .A3(n5667), .ZN(n5589) );
  INV_X1 U7151 ( .A(n7704), .ZN(n7706) );
  OAI211_X1 U7152 ( .C1(n5579), .C2(n5578), .A(n7706), .B(n5666), .ZN(n5587)
         );
  NAND2_X1 U7153 ( .A1(n5671), .A2(n5580), .ZN(n5591) );
  INV_X1 U7154 ( .A(n5581), .ZN(n5582) );
  NOR2_X1 U7155 ( .A1(n5591), .A2(n5582), .ZN(n5673) );
  INV_X1 U7156 ( .A(n5583), .ZN(n5584) );
  NAND2_X1 U7157 ( .A1(n5671), .A2(n5584), .ZN(n5585) );
  NAND2_X1 U7158 ( .A1(n5585), .A2(n5590), .ZN(n5586) );
  AOI21_X1 U7159 ( .B1(n5587), .B2(n5673), .A(n5586), .ZN(n5588) );
  MUX2_X1 U7160 ( .A(n5589), .B(n5588), .S(n6248), .Z(n5593) );
  NAND3_X1 U7161 ( .A1(n5591), .A2(n5590), .A3(n5707), .ZN(n5592) );
  NAND2_X1 U7162 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7163 ( .A1(n5594), .A2(n7855), .ZN(n5599) );
  AND2_X1 U7164 ( .A1(n5600), .A2(n5595), .ZN(n5676) );
  NAND2_X1 U7165 ( .A1(n9521), .A2(n7930), .ZN(n5596) );
  NAND2_X1 U7166 ( .A1(n5597), .A2(n5596), .ZN(n5674) );
  INV_X1 U7167 ( .A(n5674), .ZN(n5598) );
  NAND2_X1 U7168 ( .A1(n5603), .A2(n5600), .ZN(n5678) );
  INV_X1 U7169 ( .A(n5677), .ZN(n5601) );
  OR2_X1 U7170 ( .A1(n5606), .A2(n5601), .ZN(n5602) );
  NAND2_X1 U7171 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  INV_X1 U7172 ( .A(n5606), .ZN(n9364) );
  AND2_X1 U7173 ( .A1(n5609), .A2(n9364), .ZN(n5607) );
  MUX2_X1 U7174 ( .A(n5607), .B(n6249), .S(n5707), .Z(n5612) );
  MUX2_X1 U7175 ( .A(n5609), .B(n5608), .S(n6248), .Z(n5610) );
  INV_X1 U7176 ( .A(n5610), .ZN(n5611) );
  AOI21_X1 U7177 ( .B1(n5613), .B2(n5612), .A(n5611), .ZN(n5615) );
  AND2_X1 U7178 ( .A1(n5616), .A2(n6248), .ZN(n5617) );
  OAI21_X1 U7179 ( .B1(n6253), .B2(n5707), .A(n9319), .ZN(n5619) );
  MUX2_X1 U7180 ( .A(n5620), .B(n6254), .S(n6248), .Z(n5621) );
  NAND2_X1 U7181 ( .A1(n5631), .A2(n6255), .ZN(n5623) );
  AND4_X1 U7182 ( .A1(n5634), .A2(n6248), .A3(n5628), .A4(n5627), .ZN(n5622)
         );
  NAND2_X1 U7183 ( .A1(n5623), .A2(n5622), .ZN(n5626) );
  AND3_X1 U7184 ( .A1(n5628), .A2(n5627), .A3(n5707), .ZN(n5629) );
  OAI21_X1 U7185 ( .B1(n5631), .B2(n5630), .A(n5629), .ZN(n5632) );
  OAI21_X1 U7186 ( .B1(n5635), .B2(n5634), .A(n5633), .ZN(n5636) );
  NAND2_X1 U7187 ( .A1(n5636), .A2(n5707), .ZN(n5637) );
  MUX2_X1 U7188 ( .A(n5639), .B(n5638), .S(n6248), .Z(n5640) );
  NAND2_X1 U7189 ( .A1(n5641), .A2(n5640), .ZN(n5644) );
  NOR2_X1 U7190 ( .A1(n5644), .A2(n9550), .ZN(n5647) );
  INV_X1 U7191 ( .A(n9546), .ZN(n9235) );
  OAI211_X1 U7192 ( .C1(n5642), .C2(n5707), .A(n9235), .B(n9107), .ZN(n5646)
         );
  AOI22_X1 U7193 ( .A1(n5642), .A2(n5707), .B1(n9238), .B2(n9107), .ZN(n5643)
         );
  OAI211_X1 U7194 ( .C1(n5647), .C2(n5644), .A(n5643), .B(n5711), .ZN(n5645)
         );
  OAI21_X1 U7195 ( .B1(n5647), .B2(n5646), .A(n5645), .ZN(n5708) );
  OAI21_X1 U7196 ( .B1(n5708), .B2(n5706), .A(n6478), .ZN(n5649) );
  NAND2_X1 U7197 ( .A1(n4401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  INV_X1 U7198 ( .A(n6997), .ZN(n5661) );
  CLKBUF_X1 U7199 ( .A(n5502), .Z(n9133) );
  OAI21_X1 U7200 ( .B1(n6207), .B2(n7050), .A(n5653), .ZN(n5654) );
  AOI211_X1 U7201 ( .C1(n9724), .C2(n9133), .A(n7490), .B(n5654), .ZN(n5658)
         );
  NAND4_X1 U7202 ( .A1(n5658), .A2(n5657), .A3(n5656), .A4(n5655), .ZN(n5659)
         );
  NAND3_X1 U7203 ( .A1(n5661), .A2(n5660), .A3(n5659), .ZN(n5664) );
  NAND4_X1 U7204 ( .A1(n5664), .A2(n5663), .A3(n7652), .A4(n5662), .ZN(n5665)
         );
  NAND2_X1 U7205 ( .A1(n5665), .A2(n7707), .ZN(n5669) );
  OAI211_X1 U7206 ( .C1(n5669), .C2(n5668), .A(n5667), .B(n5666), .ZN(n5672)
         );
  AOI22_X1 U7207 ( .A1(n5673), .A2(n5672), .B1(n5671), .B2(n5670), .ZN(n5675)
         );
  AOI21_X1 U7208 ( .B1(n5676), .B2(n5675), .A(n5674), .ZN(n5679) );
  OAI211_X1 U7209 ( .C1(n5679), .C2(n5678), .A(n6256), .B(n5677), .ZN(n5680)
         );
  NOR2_X1 U7210 ( .A1(n5681), .A2(n5680), .ZN(n5684) );
  OAI21_X1 U7211 ( .B1(n5684), .B2(n5683), .A(n5682), .ZN(n5686) );
  AOI21_X1 U7212 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5693) );
  INV_X1 U7213 ( .A(n6479), .ZN(n5692) );
  NAND2_X1 U7214 ( .A1(n5688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5690) );
  INV_X1 U7215 ( .A(n7435), .ZN(n6597) );
  NOR3_X1 U7216 ( .A1(n5693), .A2(n6597), .A3(n9699), .ZN(n5691) );
  AOI211_X1 U7217 ( .C1(n5693), .C2(n5692), .A(n7621), .B(n5691), .ZN(n5694)
         );
  NOR2_X1 U7218 ( .A1(n5695), .A2(n5696), .ZN(n6494) );
  XNOR2_X2 U7219 ( .A(n5698), .B(n5697), .ZN(n7870) );
  NAND2_X1 U7220 ( .A1(n5701), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7221 ( .A1(n6270), .A2(n6271), .ZN(n5703) );
  OR2_X4 U7222 ( .A1(n7870), .A2(n5703), .ZN(n6605) );
  NAND2_X1 U7223 ( .A1(n6480), .A2(n6478), .ZN(n6482) );
  NAND2_X1 U7224 ( .A1(n6262), .A2(n7435), .ZN(n6483) );
  OR2_X1 U7225 ( .A1(n6482), .A2(n6483), .ZN(n6246) );
  INV_X1 U7226 ( .A(n6246), .ZN(n5704) );
  NAND3_X1 U7227 ( .A1(n6494), .A2(n6600), .A3(n5704), .ZN(n5705) );
  OAI211_X1 U7228 ( .C1(n6478), .C2(n7621), .A(n5705), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5716) );
  MUX2_X1 U7229 ( .A(n5708), .B(n5707), .S(n5706), .Z(n5709) );
  NOR4_X1 U7230 ( .A1(n7621), .A2(n6478), .A3(n7490), .A4(n7435), .ZN(n5710)
         );
  OAI21_X1 U7231 ( .B1(n5711), .B2(n9699), .A(n5710), .ZN(n5712) );
  INV_X1 U7232 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7233 ( .A1(n5807), .A2(n5806), .ZN(n5820) );
  NAND2_X1 U7234 ( .A1(n5862), .A2(n5861), .ZN(n5871) );
  NAND2_X1 U7235 ( .A1(n5912), .A2(n5911), .ZN(n5926) );
  INV_X1 U7236 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5953) );
  INV_X1 U7237 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5963) );
  INV_X1 U7238 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6023) );
  OR2_X2 U7239 ( .A1(n6035), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7240 ( .A1(n6035), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7241 ( .A1(n6040), .A2(n5717), .ZN(n8636) );
  INV_X1 U7242 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5721) );
  NOR2_X1 U7243 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5725) );
  NOR2_X1 U7244 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5724) );
  NOR2_X1 U7245 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5723) );
  NAND4_X1 U7246 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n5727)
         );
  NOR2_X1 U7247 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5730) );
  NOR2_X1 U7248 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5729) );
  NOR2_X1 U7249 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5728) );
  NAND2_X1 U7250 ( .A1(n5747), .A2(n5736), .ZN(n5731) );
  NOR2_X2 U7251 ( .A1(n5734), .A2(n5731), .ZN(n7890) );
  XNOR2_X2 U7252 ( .A(n5733), .B(n5732), .ZN(n5740) );
  INV_X1 U7253 ( .A(n5740), .ZN(n5738) );
  NAND2_X1 U7254 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5735) );
  XNOR2_X2 U7255 ( .A(n5737), .B(n5736), .ZN(n5739) );
  NAND2_X1 U7256 ( .A1(n8636), .A2(n6070), .ZN(n5746) );
  INV_X1 U7257 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5743) );
  NAND2_X2 U7258 ( .A1(n5739), .A2(n5740), .ZN(n6091) );
  NAND2_X1 U7259 ( .A1(n7059), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5742) );
  INV_X2 U7260 ( .A(n6093), .ZN(n6137) );
  NAND2_X1 U7261 ( .A1(n5805), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5741) );
  OAI211_X1 U7262 ( .C1(n6094), .C2(n5743), .A(n5742), .B(n5741), .ZN(n5744)
         );
  INV_X1 U7263 ( .A(n5744), .ZN(n5745) );
  XNOR2_X1 U7264 ( .A(n5749), .B(n10039), .ZN(n6134) );
  NAND2_X1 U7265 ( .A1(n7624), .A2(n8052), .ZN(n5751) );
  OR2_X1 U7266 ( .A1(n8055), .A2(n9927), .ZN(n5750) );
  NAND2_X1 U7267 ( .A1(n5805), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7268 ( .A1(n4346), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7269 ( .A1(n5778), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7270 ( .A1(n5804), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5752) );
  NAND4_X2 U7271 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n6304)
         );
  NAND2_X1 U7272 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5756) );
  AND2_X1 U7273 ( .A1(n5757), .A2(n4881), .ZN(n5760) );
  OR2_X1 U7274 ( .A1(n8056), .A2(n5758), .ZN(n5759) );
  NAND2_X1 U7275 ( .A1(n5805), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5765) );
  INV_X1 U7276 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6632) );
  OR2_X1 U7277 ( .A1(n6091), .A2(n6632), .ZN(n5764) );
  NAND2_X1 U7278 ( .A1(n5804), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5763) );
  INV_X1 U7279 ( .A(n7159), .ZN(n5766) );
  NAND2_X1 U7280 ( .A1(n6376), .A2(SI_0_), .ZN(n5767) );
  XNOR2_X1 U7281 ( .A(n5767), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U7282 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8946), .S(n5768), .Z(n8872) );
  NAND2_X1 U7283 ( .A1(n5766), .A2(n8872), .ZN(n7158) );
  NAND2_X1 U7284 ( .A1(n7157), .A2(n7158), .ZN(n5770) );
  OR2_X1 U7285 ( .A1(n6304), .A2(n5761), .ZN(n5769) );
  NAND2_X1 U7286 ( .A1(n5778), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7287 ( .A1(n4346), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7288 ( .A1(n5805), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7289 ( .A1(n5804), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5771) );
  NAND4_X2 U7290 ( .A1(n5774), .A2(n5773), .A3(n5772), .A4(n5771), .ZN(n8431)
         );
  OR2_X1 U7291 ( .A1(n8056), .A2(n6391), .ZN(n5777) );
  OR2_X1 U7292 ( .A1(n5785), .A2(n4902), .ZN(n5776) );
  OR2_X1 U7293 ( .A1(n5768), .A2(n6658), .ZN(n5775) );
  AND3_X2 U7294 ( .A1(n5777), .A2(n5776), .A3(n5775), .ZN(n6979) );
  NAND2_X1 U7295 ( .A1(n6979), .A2(n8431), .ZN(n8099) );
  NAND2_X1 U7296 ( .A1(n5778), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7297 ( .A1(n6137), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5781) );
  INV_X1 U7298 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7301) );
  OR2_X1 U7299 ( .A1(n5779), .A2(n7301), .ZN(n5780) );
  NAND4_X4 U7300 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .ZN(n8430)
         );
  NAND2_X1 U7301 ( .A1(n4502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5784) );
  XNOR2_X1 U7302 ( .A(n5784), .B(n5718), .ZN(n6673) );
  OR2_X1 U7303 ( .A1(n8056), .A2(n6377), .ZN(n5787) );
  OR2_X1 U7304 ( .A1(n5785), .A2(n6378), .ZN(n5786) );
  OAI211_X1 U7305 ( .C1(n5768), .C2(n6673), .A(n5787), .B(n5786), .ZN(n6915)
         );
  NAND2_X1 U7306 ( .A1(n8430), .A2(n6915), .ZN(n5790) );
  AND2_X1 U7307 ( .A1(n8105), .A2(n5790), .ZN(n5788) );
  OR2_X1 U7308 ( .A1(n8430), .A2(n6915), .ZN(n5789) );
  INV_X1 U7309 ( .A(n6979), .ZN(n6902) );
  OR2_X1 U7310 ( .A1(n8431), .A2(n6902), .ZN(n6909) );
  AND2_X1 U7311 ( .A1(n5789), .A2(n6909), .ZN(n5792) );
  INV_X1 U7312 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7313 ( .A1(n5804), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7314 ( .A1(n7059), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7315 ( .A1(n6137), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5796) );
  AND2_X1 U7316 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5794) );
  NOR2_X1 U7317 ( .A1(n5807), .A2(n5794), .ZN(n6949) );
  NAND2_X1 U7318 ( .A1(n5799), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5801) );
  INV_X1 U7319 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U7320 ( .A(n5801), .B(n5800), .ZN(n6698) );
  OR2_X1 U7321 ( .A1(n8056), .A2(n6389), .ZN(n5803) );
  OR2_X1 U7322 ( .A1(n8055), .A2(n6390), .ZN(n5802) );
  OAI211_X1 U7323 ( .C1(n5768), .C2(n6698), .A(n5803), .B(n5802), .ZN(n7170)
         );
  NAND2_X1 U7324 ( .A1(n7058), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7325 ( .A1(n7059), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7326 ( .A1(n6137), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7327 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  AND2_X1 U7328 ( .A1(n5820), .A2(n5808), .ZN(n7343) );
  OR2_X1 U7329 ( .A1(n6090), .A2(n7343), .ZN(n5809) );
  NAND4_X1 U7330 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .ZN(n8428)
         );
  OR2_X1 U7331 ( .A1(n5813), .A2(n4505), .ZN(n5815) );
  XNOR2_X1 U7332 ( .A(n5814), .B(n5815), .ZN(n6745) );
  OR2_X1 U7333 ( .A1(n8056), .A2(n6380), .ZN(n5817) );
  OR2_X1 U7334 ( .A1(n8055), .A2(n6379), .ZN(n5816) );
  OAI211_X1 U7335 ( .C1(n5768), .C2(n6745), .A(n5817), .B(n5816), .ZN(n9830)
         );
  NAND2_X1 U7336 ( .A1(n8428), .A2(n9830), .ZN(n5818) );
  NAND2_X1 U7337 ( .A1(n5819), .A2(n5818), .ZN(n7353) );
  NAND2_X1 U7338 ( .A1(n7058), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5825) );
  INV_X1 U7339 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6759) );
  OR2_X1 U7340 ( .A1(n6091), .A2(n6759), .ZN(n5824) );
  NAND2_X1 U7341 ( .A1(n6137), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7342 ( .A1(n5820), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5821) );
  AND2_X1 U7343 ( .A1(n5833), .A2(n5821), .ZN(n7358) );
  OR2_X1 U7344 ( .A1(n6090), .A2(n7358), .ZN(n5822) );
  NAND4_X1 U7345 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(n8427)
         );
  NAND2_X1 U7346 ( .A1(n5826), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5827) );
  MUX2_X1 U7347 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5827), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5828) );
  NAND2_X1 U7348 ( .A1(n5828), .A2(n4385), .ZN(n6764) );
  OR2_X1 U7349 ( .A1(n8055), .A2(n6388), .ZN(n5830) );
  OR2_X1 U7350 ( .A1(n8056), .A2(n6387), .ZN(n5829) );
  OAI211_X1 U7351 ( .C1(n5768), .C2(n6764), .A(n5830), .B(n5829), .ZN(n9836)
         );
  AND2_X1 U7352 ( .A1(n8427), .A2(n9836), .ZN(n5831) );
  OAI22_X1 U7353 ( .A1(n7353), .A2(n5831), .B1(n8427), .B2(n9836), .ZN(n7338)
         );
  NAND2_X1 U7354 ( .A1(n6137), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5838) );
  INV_X1 U7355 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7334) );
  OR2_X1 U7356 ( .A1(n6094), .A2(n7334), .ZN(n5837) );
  INV_X1 U7357 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5832) );
  OR2_X1 U7358 ( .A1(n6091), .A2(n5832), .ZN(n5836) );
  AND2_X1 U7359 ( .A1(n5833), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5834) );
  NOR2_X1 U7360 ( .A1(n5844), .A2(n5834), .ZN(n7376) );
  OR2_X1 U7361 ( .A1(n6090), .A2(n7376), .ZN(n5835) );
  NAND2_X1 U7362 ( .A1(n4385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5839) );
  XNOR2_X1 U7363 ( .A(n5839), .B(n5719), .ZN(n7288) );
  OR2_X1 U7364 ( .A1(n8056), .A2(n6385), .ZN(n5841) );
  OR2_X1 U7365 ( .A1(n8055), .A2(n6384), .ZN(n5840) );
  OAI211_X1 U7366 ( .C1(n5768), .C2(n7288), .A(n5841), .B(n5840), .ZN(n9841)
         );
  NAND2_X1 U7367 ( .A1(n7564), .A2(n9841), .ZN(n8136) );
  INV_X1 U7368 ( .A(n9841), .ZN(n7335) );
  INV_X1 U7369 ( .A(n7564), .ZN(n8426) );
  NAND2_X1 U7370 ( .A1(n7335), .A2(n8426), .ZN(n7560) );
  NAND2_X1 U7371 ( .A1(n8136), .A2(n7560), .ZN(n8132) );
  NAND2_X1 U7372 ( .A1(n7338), .A2(n8132), .ZN(n5843) );
  NAND2_X1 U7373 ( .A1(n7564), .A2(n7335), .ZN(n5842) );
  NAND2_X1 U7374 ( .A1(n5843), .A2(n5842), .ZN(n7563) );
  NAND2_X1 U7375 ( .A1(n7058), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5850) );
  INV_X1 U7376 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7291) );
  OR2_X1 U7377 ( .A1(n6091), .A2(n7291), .ZN(n5849) );
  NOR2_X1 U7378 ( .A1(n5844), .A2(n7276), .ZN(n5845) );
  OR2_X1 U7379 ( .A1(n6090), .A2(n4413), .ZN(n5848) );
  INV_X1 U7380 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5846) );
  OR2_X1 U7381 ( .A1(n6093), .A2(n5846), .ZN(n5847) );
  NAND2_X1 U7382 ( .A1(n5851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7383 ( .A(n5852), .B(n4574), .ZN(n7506) );
  OR2_X1 U7384 ( .A1(n8056), .A2(n6399), .ZN(n5854) );
  OR2_X1 U7385 ( .A1(n8055), .A2(n6400), .ZN(n5853) );
  OAI211_X1 U7386 ( .C1(n5768), .C2(n7506), .A(n5854), .B(n5853), .ZN(n7557)
         );
  NAND2_X1 U7387 ( .A1(n10130), .A2(n7557), .ZN(n8137) );
  NAND2_X1 U7388 ( .A1(n9851), .A2(n10120), .ZN(n8129) );
  AND2_X1 U7389 ( .A1(n8137), .A2(n8129), .ZN(n7562) );
  NAND2_X1 U7390 ( .A1(n10120), .A2(n7557), .ZN(n5855) );
  OR2_X1 U7391 ( .A1(n5856), .A2(n4505), .ZN(n5857) );
  XNOR2_X1 U7392 ( .A(n5857), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7577) );
  AOI22_X1 U7393 ( .A1(n5996), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6371), .B2(
        n7577), .ZN(n5859) );
  NAND2_X1 U7394 ( .A1(n6405), .A2(n8052), .ZN(n5858) );
  NAND2_X1 U7395 ( .A1(n6137), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5868) );
  INV_X1 U7396 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5860) );
  OR2_X1 U7397 ( .A1(n6091), .A2(n5860), .ZN(n5867) );
  OR2_X1 U7398 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  AND2_X1 U7399 ( .A1(n5871), .A2(n5863), .ZN(n10139) );
  OR2_X1 U7400 ( .A1(n6090), .A2(n10139), .ZN(n5866) );
  INV_X1 U7401 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7402 ( .A1(n6094), .A2(n5864), .ZN(n5865) );
  NAND2_X1 U7403 ( .A1(n10135), .A2(n10122), .ZN(n5869) );
  NAND2_X1 U7404 ( .A1(n5870), .A2(n5869), .ZN(n7610) );
  NAND2_X1 U7405 ( .A1(n7058), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5876) );
  INV_X1 U7406 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7589) );
  OR2_X1 U7407 ( .A1(n6091), .A2(n7589), .ZN(n5875) );
  NAND2_X1 U7408 ( .A1(n6137), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7409 ( .A1(n5871), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5872) );
  AND2_X1 U7410 ( .A1(n5888), .A2(n5872), .ZN(n7616) );
  OR2_X1 U7411 ( .A1(n6090), .A2(n7616), .ZN(n5873) );
  NAND4_X1 U7412 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n8425)
         );
  NAND2_X1 U7413 ( .A1(n6403), .A2(n8052), .ZN(n5881) );
  NAND2_X1 U7414 ( .A1(n5877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5878) );
  MUX2_X1 U7415 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5878), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5879) );
  AND2_X1 U7416 ( .A1(n5879), .A2(n5884), .ZN(n7676) );
  AOI22_X1 U7417 ( .A1(n5996), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6371), .B2(
        n7676), .ZN(n5880) );
  NAND2_X1 U7418 ( .A1(n5881), .A2(n5880), .ZN(n9863) );
  OR2_X1 U7419 ( .A1(n8425), .A2(n9863), .ZN(n7608) );
  NAND2_X1 U7420 ( .A1(n7610), .A2(n7608), .ZN(n5882) );
  NAND2_X1 U7421 ( .A1(n9863), .A2(n8425), .ZN(n7607) );
  NAND2_X1 U7422 ( .A1(n5882), .A2(n7607), .ZN(n7629) );
  NAND2_X1 U7423 ( .A1(n6411), .A2(n8052), .ZN(n5887) );
  NAND2_X1 U7424 ( .A1(n5884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  MUX2_X1 U7425 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5883), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5885) );
  NAND2_X1 U7426 ( .A1(n5885), .A2(n4678), .ZN(n7685) );
  AOI22_X1 U7427 ( .A1(n5996), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6371), .B2(
        n7742), .ZN(n5886) );
  NAND2_X1 U7428 ( .A1(n5887), .A2(n5886), .ZN(n7632) );
  NAND2_X1 U7429 ( .A1(n6137), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5893) );
  INV_X1 U7430 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7683) );
  OR2_X1 U7431 ( .A1(n6094), .A2(n7683), .ZN(n5892) );
  INV_X1 U7432 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7682) );
  OR2_X1 U7433 ( .A1(n6091), .A2(n7682), .ZN(n5891) );
  NAND2_X1 U7434 ( .A1(n5888), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5889) );
  AND2_X1 U7435 ( .A1(n5898), .A2(n5889), .ZN(n7760) );
  OR2_X1 U7436 ( .A1(n6090), .A2(n7760), .ZN(n5890) );
  OR2_X1 U7437 ( .A1(n7632), .A2(n7796), .ZN(n8147) );
  NAND2_X1 U7438 ( .A1(n7632), .A2(n7796), .ZN(n8150) );
  NAND2_X1 U7439 ( .A1(n8147), .A2(n8150), .ZN(n8143) );
  NAND2_X1 U7440 ( .A1(n7629), .A2(n8143), .ZN(n7628) );
  INV_X1 U7441 ( .A(n7796), .ZN(n8424) );
  NAND2_X1 U7442 ( .A1(n7632), .A2(n8424), .ZN(n5894) );
  NAND2_X1 U7443 ( .A1(n7628), .A2(n5894), .ZN(n7794) );
  NAND2_X1 U7444 ( .A1(n6544), .A2(n8052), .ZN(n5897) );
  OR2_X1 U7445 ( .A1(n5908), .A2(n4505), .ZN(n5895) );
  XNOR2_X1 U7446 ( .A(n5895), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7696) );
  AOI22_X1 U7447 ( .A1(n5996), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6371), .B2(
        n7696), .ZN(n5896) );
  NAND2_X1 U7448 ( .A1(n5897), .A2(n5896), .ZN(n9876) );
  NAND2_X1 U7449 ( .A1(n7059), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7450 ( .A1(n6137), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7451 ( .A1(n7058), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5901) );
  AND2_X1 U7452 ( .A1(n5898), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5899) );
  NOR2_X1 U7453 ( .A1(n5912), .A2(n5899), .ZN(n7793) );
  OR2_X1 U7454 ( .A1(n6090), .A2(n7793), .ZN(n5900) );
  NAND4_X1 U7455 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n8423)
         );
  OR2_X1 U7456 ( .A1(n9876), .A2(n8423), .ZN(n5904) );
  NAND2_X1 U7457 ( .A1(n7794), .A2(n5904), .ZN(n5906) );
  NAND2_X1 U7458 ( .A1(n9876), .A2(n8423), .ZN(n5905) );
  NAND2_X1 U7459 ( .A1(n5906), .A2(n5905), .ZN(n8764) );
  INV_X1 U7460 ( .A(n8764), .ZN(n5919) );
  NAND2_X1 U7461 ( .A1(n6557), .A2(n8052), .ZN(n5910) );
  OR2_X1 U7462 ( .A1(n5949), .A2(n4505), .ZN(n5921) );
  XNOR2_X1 U7463 ( .A(n5921), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7812) );
  AOI22_X1 U7464 ( .A1(n5996), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6371), .B2(
        n7812), .ZN(n5909) );
  NAND2_X1 U7465 ( .A1(n5910), .A2(n5909), .ZN(n8864) );
  NAND2_X1 U7466 ( .A1(n6137), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5917) );
  INV_X1 U7467 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8775) );
  OR2_X1 U7468 ( .A1(n6094), .A2(n8775), .ZN(n5916) );
  INV_X1 U7469 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8867) );
  OR2_X1 U7470 ( .A1(n6091), .A2(n8867), .ZN(n5915) );
  OR2_X1 U7471 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  AND2_X1 U7472 ( .A1(n5913), .A2(n5926), .ZN(n8774) );
  OR2_X1 U7473 ( .A1(n6090), .A2(n8774), .ZN(n5914) );
  OR2_X1 U7474 ( .A1(n8864), .A2(n8746), .ZN(n8160) );
  NAND2_X1 U7475 ( .A1(n8864), .A2(n8746), .ZN(n8159) );
  INV_X1 U7476 ( .A(n8746), .ZN(n8422) );
  OR2_X1 U7477 ( .A1(n8864), .A2(n8422), .ZN(n5920) );
  NAND2_X1 U7478 ( .A1(n6621), .A2(n8052), .ZN(n5925) );
  NAND2_X1 U7479 ( .A1(n5921), .A2(n5947), .ZN(n5922) );
  NAND2_X1 U7480 ( .A1(n5922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7481 ( .A1(n5923), .A2(n5946), .ZN(n5933) );
  INV_X1 U7482 ( .A(n8454), .ZN(n7824) );
  AOI22_X1 U7483 ( .A1(n5996), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7824), .B2(
        n6371), .ZN(n5924) );
  NAND2_X1 U7484 ( .A1(n5925), .A2(n5924), .ZN(n8750) );
  NAND2_X1 U7485 ( .A1(n6137), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5931) );
  INV_X1 U7486 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8862) );
  OR2_X1 U7487 ( .A1(n6091), .A2(n8862), .ZN(n5930) );
  INV_X1 U7488 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7823) );
  OR2_X1 U7489 ( .A1(n6094), .A2(n7823), .ZN(n5929) );
  NAND2_X1 U7490 ( .A1(n5926), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5927) );
  AND2_X1 U7491 ( .A1(n4368), .A2(n5927), .ZN(n8751) );
  OR2_X1 U7492 ( .A1(n6090), .A2(n8751), .ZN(n5928) );
  OR2_X1 U7493 ( .A1(n8750), .A2(n8767), .ZN(n8165) );
  NAND2_X1 U7494 ( .A1(n8750), .A2(n8767), .ZN(n8164) );
  NAND2_X1 U7495 ( .A1(n8750), .A2(n8729), .ZN(n5932) );
  NAND2_X1 U7496 ( .A1(n8748), .A2(n5932), .ZN(n8725) );
  NAND2_X1 U7497 ( .A1(n6662), .A2(n8052), .ZN(n5936) );
  NAND2_X1 U7498 ( .A1(n5933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7499 ( .A(n5934), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8477) );
  AOI22_X1 U7500 ( .A1(n6371), .A2(n8477), .B1(n5996), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7501 ( .A1(n5936), .A2(n5935), .ZN(n8854) );
  NAND2_X1 U7502 ( .A1(n6137), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5942) );
  INV_X1 U7503 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8735) );
  OR2_X1 U7504 ( .A1(n6094), .A2(n8735), .ZN(n5941) );
  INV_X1 U7505 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5937) );
  OR2_X1 U7506 ( .A1(n6091), .A2(n5937), .ZN(n5940) );
  AND2_X1 U7507 ( .A1(n4368), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5938) );
  NOR2_X1 U7508 ( .A1(n5954), .A2(n5938), .ZN(n8734) );
  OR2_X1 U7509 ( .A1(n6090), .A2(n8734), .ZN(n5939) );
  OR2_X1 U7510 ( .A1(n8854), .A2(n8745), .ZN(n8168) );
  NAND2_X1 U7511 ( .A1(n8854), .A2(n8745), .ZN(n8169) );
  NAND2_X1 U7512 ( .A1(n8168), .A2(n8169), .ZN(n8163) );
  NAND2_X1 U7513 ( .A1(n8725), .A2(n8163), .ZN(n5944) );
  INV_X1 U7514 ( .A(n8745), .ZN(n8421) );
  NAND2_X1 U7515 ( .A1(n8854), .A2(n8421), .ZN(n5943) );
  NAND2_X1 U7516 ( .A1(n5944), .A2(n5943), .ZN(n7897) );
  NAND2_X1 U7517 ( .A1(n6710), .A2(n8052), .ZN(n5952) );
  INV_X1 U7518 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5945) );
  AND3_X1 U7519 ( .A1(n5947), .A2(n5946), .A3(n5945), .ZN(n5948) );
  NAND2_X1 U7520 ( .A1(n5970), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7521 ( .A(n5950), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8502) );
  AOI22_X1 U7522 ( .A1(n5996), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6371), .B2(
        n8502), .ZN(n5951) );
  NAND2_X1 U7523 ( .A1(n5952), .A2(n5951), .ZN(n8332) );
  NAND2_X1 U7524 ( .A1(n6137), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5960) );
  INV_X1 U7525 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8479) );
  OR2_X1 U7526 ( .A1(n6094), .A2(n8479), .ZN(n5959) );
  INV_X1 U7527 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8851) );
  OR2_X1 U7528 ( .A1(n6091), .A2(n8851), .ZN(n5958) );
  NOR2_X1 U7529 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  OR2_X1 U7530 ( .A1(n5998), .A2(n5955), .ZN(n8719) );
  INV_X1 U7531 ( .A(n8719), .ZN(n5956) );
  OR2_X1 U7532 ( .A1(n6090), .A2(n5956), .ZN(n5957) );
  OR2_X1 U7533 ( .A1(n8332), .A2(n8705), .ZN(n8175) );
  NAND2_X1 U7534 ( .A1(n8332), .A2(n8705), .ZN(n8187) );
  NAND2_X1 U7535 ( .A1(n8175), .A2(n8187), .ZN(n8717) );
  NAND2_X1 U7536 ( .A1(n7364), .A2(n8052), .ZN(n5962) );
  INV_X1 U7537 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7366) );
  OR2_X1 U7538 ( .A1(n8055), .A2(n7366), .ZN(n5961) );
  NOR2_X1 U7539 ( .A1(n5976), .A2(n5963), .ZN(n5964) );
  OR2_X1 U7540 ( .A1(n6024), .A2(n5964), .ZN(n8365) );
  NAND2_X1 U7541 ( .A1(n8365), .A2(n6070), .ZN(n5969) );
  NAND2_X1 U7542 ( .A1(n7058), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5966) );
  INV_X1 U7543 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10083) );
  OR2_X1 U7544 ( .A1(n6091), .A2(n10083), .ZN(n5965) );
  AND2_X1 U7545 ( .A1(n5966), .A2(n5965), .ZN(n5968) );
  NAND2_X1 U7546 ( .A1(n6137), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7547 ( .A1(n8908), .A2(n8656), .ZN(n8651) );
  NAND2_X1 U7548 ( .A1(n8196), .A2(n8651), .ZN(n8088) );
  NAND2_X1 U7549 ( .A1(n7154), .A2(n8052), .ZN(n5975) );
  NAND2_X1 U7550 ( .A1(n5993), .A2(n5971), .ZN(n5972) );
  AOI22_X1 U7551 ( .A1(n6299), .A2(n6371), .B1(n5996), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5974) );
  AND2_X1 U7552 ( .A1(n5988), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5977) );
  OR2_X1 U7553 ( .A1(n5977), .A2(n5976), .ZN(n8678) );
  NAND2_X1 U7554 ( .A1(n8678), .A2(n6070), .ZN(n5982) );
  NAND2_X1 U7555 ( .A1(n6137), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5981) );
  INV_X1 U7556 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7557 ( .A1(n6094), .A2(n5978), .ZN(n5980) );
  INV_X1 U7558 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8839) );
  OR2_X1 U7559 ( .A1(n6091), .A2(n8839), .ZN(n5979) );
  INV_X1 U7560 ( .A(n8689), .ZN(n8419) );
  NAND2_X1 U7561 ( .A1(n5983), .A2(n8419), .ZN(n6014) );
  NAND2_X1 U7562 ( .A1(n5983), .A2(n8689), .ZN(n8192) );
  NAND2_X1 U7563 ( .A1(n6923), .A2(n8052), .ZN(n5986) );
  XNOR2_X1 U7564 ( .A(n5984), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8541) );
  AOI22_X1 U7565 ( .A1(n5996), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8541), .B2(
        n6371), .ZN(n5985) );
  NAND2_X1 U7566 ( .A1(n7058), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7567 ( .A1(n7059), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7568 ( .A1(n6000), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7569 ( .A1(n5988), .A2(n5987), .ZN(n8698) );
  NAND2_X1 U7570 ( .A1(n6070), .A2(n8698), .ZN(n5990) );
  NAND2_X1 U7571 ( .A1(n6137), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5989) );
  NAND4_X1 U7572 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n8674)
         );
  OR2_X1 U7573 ( .A1(n8385), .A2(n8674), .ZN(n6008) );
  INV_X1 U7574 ( .A(n6008), .ZN(n6007) );
  NAND2_X1 U7575 ( .A1(n8385), .A2(n8674), .ZN(n6005) );
  INV_X1 U7576 ( .A(n5993), .ZN(n5994) );
  NAND2_X1 U7577 ( .A1(n5994), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5995) );
  XNOR2_X1 U7578 ( .A(n5995), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8524) );
  AOI22_X1 U7579 ( .A1(n5996), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6371), .B2(
        n8524), .ZN(n5997) );
  NAND2_X1 U7580 ( .A1(n6137), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6004) );
  INV_X1 U7581 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8710) );
  OR2_X1 U7582 ( .A1(n6094), .A2(n8710), .ZN(n6003) );
  INV_X1 U7583 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8847) );
  OR2_X1 U7584 ( .A1(n6091), .A2(n8847), .ZN(n6002) );
  OR2_X1 U7585 ( .A1(n5998), .A2(n8343), .ZN(n5999) );
  AND2_X1 U7586 ( .A1(n6000), .A2(n5999), .ZN(n8709) );
  OR2_X1 U7587 ( .A1(n6090), .A2(n8709), .ZN(n6001) );
  INV_X1 U7588 ( .A(n8716), .ZN(n8420) );
  NAND2_X1 U7589 ( .A1(n8708), .A2(n8420), .ZN(n8685) );
  AND2_X1 U7590 ( .A1(n6005), .A2(n8685), .ZN(n6006) );
  OR2_X1 U7591 ( .A1(n6007), .A2(n6006), .ZN(n6013) );
  INV_X1 U7592 ( .A(n6013), .ZN(n6010) );
  NAND2_X1 U7593 ( .A1(n8708), .A2(n8716), .ZN(n8692) );
  AND2_X1 U7594 ( .A1(n8707), .A2(n6008), .ZN(n6009) );
  OR2_X1 U7595 ( .A1(n6010), .A2(n6009), .ZN(n8667) );
  NAND2_X1 U7596 ( .A1(n7897), .A2(n6011), .ZN(n6018) );
  INV_X1 U7597 ( .A(n6012), .ZN(n6016) );
  INV_X1 U7598 ( .A(n8705), .ZN(n8853) );
  NAND2_X1 U7599 ( .A1(n8332), .A2(n8853), .ZN(n8683) );
  AND2_X1 U7600 ( .A1(n8683), .A2(n6013), .ZN(n8666) );
  AND2_X1 U7601 ( .A1(n8666), .A2(n6014), .ZN(n7898) );
  AND2_X1 U7602 ( .A1(n7898), .A2(n8088), .ZN(n6015) );
  NAND2_X1 U7603 ( .A1(n6018), .A2(n6017), .ZN(n7901) );
  NAND2_X1 U7604 ( .A1(n6019), .A2(n8656), .ZN(n6020) );
  NAND2_X1 U7605 ( .A1(n7901), .A2(n6020), .ZN(n8655) );
  NAND2_X1 U7606 ( .A1(n7488), .A2(n8052), .ZN(n6022) );
  OR2_X1 U7607 ( .A1(n8055), .A2(n7492), .ZN(n6021) );
  OR2_X1 U7608 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  NAND2_X1 U7609 ( .A1(n6033), .A2(n6025), .ZN(n8658) );
  NAND2_X1 U7610 ( .A1(n8658), .A2(n6070), .ZN(n6028) );
  AOI22_X1 U7611 ( .A1(n7058), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n7059), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7612 ( .A1(n6137), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7613 ( .A1(n8662), .A2(n8833), .ZN(n8181) );
  NAND2_X1 U7614 ( .A1(n8179), .A2(n8181), .ZN(n8654) );
  OR2_X1 U7615 ( .A1(n8055), .A2(n9963), .ZN(n6031) );
  INV_X1 U7616 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U7617 ( .A1(n6033), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7618 ( .A1(n6035), .A2(n6034), .ZN(n8646) );
  NAND2_X1 U7619 ( .A1(n8646), .A2(n6070), .ZN(n6037) );
  AOI22_X1 U7620 ( .A1(n7058), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n7059), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U7621 ( .C1(n6093), .C2(n8899), .A(n6037), .B(n6036), .ZN(n8418)
         );
  NAND2_X1 U7622 ( .A1(n7805), .A2(n8052), .ZN(n6039) );
  OR2_X1 U7623 ( .A1(n8055), .A2(n7808), .ZN(n6038) );
  AND2_X1 U7624 ( .A1(n6040), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6041) );
  NOR2_X2 U7625 ( .A1(n6040), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6049) );
  OR2_X1 U7626 ( .A1(n6041), .A2(n6049), .ZN(n8625) );
  INV_X1 U7627 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7628 ( .A1(n7059), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7629 ( .A1(n6137), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6042) );
  OAI211_X1 U7630 ( .C1(n6094), .C2(n6044), .A(n6043), .B(n6042), .ZN(n6045)
         );
  INV_X1 U7631 ( .A(n8811), .ZN(n8416) );
  NAND2_X1 U7632 ( .A1(n7863), .A2(n8052), .ZN(n6048) );
  OR2_X1 U7633 ( .A1(n8055), .A2(n9939), .ZN(n6047) );
  INV_X1 U7634 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U7635 ( .A1(n6049), .A2(n8327), .ZN(n6057) );
  OR2_X1 U7636 ( .A1(n6049), .A2(n8327), .ZN(n6050) );
  NAND2_X1 U7637 ( .A1(n6057), .A2(n6050), .ZN(n8615) );
  INV_X1 U7638 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7639 ( .A1(n6137), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7640 ( .A1(n7059), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7641 ( .C1(n6094), .C2(n6053), .A(n6052), .B(n6051), .ZN(n6054)
         );
  OR2_X1 U7642 ( .A1(n8614), .A2(n8623), .ZN(n6127) );
  NAND2_X1 U7643 ( .A1(n8614), .A2(n8623), .ZN(n8212) );
  NAND2_X1 U7644 ( .A1(n6127), .A2(n8212), .ZN(n8616) );
  NAND2_X1 U7645 ( .A1(n7868), .A2(n8052), .ZN(n6056) );
  OR2_X1 U7646 ( .A1(n8055), .A2(n10085), .ZN(n6055) );
  NAND2_X1 U7647 ( .A1(n6057), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7648 ( .A1(n6068), .A2(n6058), .ZN(n8602) );
  NAND2_X1 U7649 ( .A1(n8602), .A2(n6070), .ZN(n6064) );
  INV_X1 U7650 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7651 ( .A1(n5805), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7652 ( .A1(n7059), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7653 ( .C1(n6094), .C2(n6061), .A(n6060), .B(n6059), .ZN(n6062)
         );
  INV_X1 U7654 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7655 ( .A1(n8404), .A2(n8613), .ZN(n6065) );
  NAND2_X1 U7656 ( .A1(n8049), .A2(n8052), .ZN(n6067) );
  OR2_X1 U7657 ( .A1(n8055), .A2(n7875), .ZN(n6066) );
  NAND2_X1 U7658 ( .A1(n6068), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7659 ( .A1(n6069), .A2(n4369), .ZN(n8590) );
  NAND2_X1 U7660 ( .A1(n8590), .A2(n6070), .ZN(n6076) );
  INV_X1 U7661 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7662 ( .A1(n7059), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7663 ( .A1(n6137), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6071) );
  OAI211_X1 U7664 ( .C1(n6073), .C2(n6094), .A(n6072), .B(n6071), .ZN(n6074)
         );
  INV_X1 U7665 ( .A(n6074), .ZN(n6075) );
  NAND2_X1 U7666 ( .A1(n8794), .A2(n8798), .ZN(n6077) );
  NAND2_X1 U7667 ( .A1(n8942), .A2(n8052), .ZN(n6079) );
  INV_X1 U7668 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8945) );
  OR2_X1 U7669 ( .A1(n8055), .A2(n8945), .ZN(n6078) );
  NAND2_X1 U7670 ( .A1(n7058), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6085) );
  INV_X1 U7671 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6080) );
  OR2_X1 U7672 ( .A1(n6091), .A2(n6080), .ZN(n6084) );
  NOR2_X1 U7673 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n4369), .ZN(n8571) );
  AND2_X1 U7674 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n4369), .ZN(n6081) );
  INV_X1 U7675 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10059) );
  OR2_X1 U7676 ( .A1(n6093), .A2(n10059), .ZN(n6082) );
  NAND2_X1 U7677 ( .A1(n8236), .A2(n8592), .ZN(n6086) );
  NAND2_X1 U7678 ( .A1(n8576), .A2(n6086), .ZN(n6087) );
  INV_X2 U7679 ( .A(n8592), .ZN(n8793) );
  NAND2_X1 U7680 ( .A1(n7882), .A2(n8052), .ZN(n6089) );
  OR2_X1 U7681 ( .A1(n8055), .A2(n8940), .ZN(n6088) );
  INV_X1 U7682 ( .A(n4348), .ZN(n7877) );
  OR2_X1 U7683 ( .A1(n6090), .A2(n7877), .ZN(n7063) );
  OR2_X1 U7684 ( .A1(n6091), .A2(n6200), .ZN(n6097) );
  INV_X1 U7685 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7686 ( .A1(n6093), .A2(n6092), .ZN(n6096) );
  OR2_X1 U7687 ( .A1(n6094), .A2(n10069), .ZN(n6095) );
  NAND2_X1 U7688 ( .A1(n6098), .A2(n8581), .ZN(n8058) );
  NAND2_X1 U7689 ( .A1(n8241), .A2(n8058), .ZN(n8092) );
  NAND2_X1 U7690 ( .A1(n6299), .A2(n8254), .ZN(n6109) );
  INV_X1 U7691 ( .A(n6102), .ZN(n6103) );
  NAND2_X1 U7692 ( .A1(n6103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6104) );
  INV_X1 U7693 ( .A(n6100), .ZN(n6106) );
  NAND2_X1 U7694 ( .A1(n6106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6108) );
  INV_X1 U7695 ( .A(n8105), .ZN(n6981) );
  NAND2_X1 U7696 ( .A1(n6969), .A2(n8104), .ZN(n6913) );
  INV_X1 U7697 ( .A(n7170), .ZN(n9825) );
  NAND2_X1 U7698 ( .A1(n9825), .A2(n8429), .ZN(n8118) );
  INV_X1 U7699 ( .A(n8430), .ZN(n6983) );
  NAND2_X1 U7700 ( .A1(n6983), .A2(n6915), .ZN(n8117) );
  INV_X1 U7701 ( .A(n6915), .ZN(n7299) );
  NAND2_X1 U7702 ( .A1(n7299), .A2(n8430), .ZN(n8111) );
  AND2_X1 U7703 ( .A1(n8118), .A2(n6908), .ZN(n6110) );
  NAND2_X1 U7704 ( .A1(n7146), .A2(n7170), .ZN(n8112) );
  NAND2_X1 U7705 ( .A1(n8118), .A2(n4883), .ZN(n6111) );
  INV_X1 U7706 ( .A(n9830), .ZN(n7344) );
  NAND2_X1 U7707 ( .A1(n7344), .A2(n8428), .ZN(n8119) );
  NAND2_X1 U7708 ( .A1(n7242), .A2(n9830), .ZN(n8122) );
  INV_X1 U7709 ( .A(n8427), .ZN(n7373) );
  AND2_X1 U7710 ( .A1(n7373), .A2(n9836), .ZN(n8115) );
  INV_X1 U7711 ( .A(n9836), .ZN(n7359) );
  NAND2_X1 U7712 ( .A1(n7359), .A2(n8427), .ZN(n8125) );
  OAI21_X1 U7713 ( .B1(n7361), .B2(n8115), .A(n8125), .ZN(n7330) );
  INV_X1 U7714 ( .A(n8132), .ZN(n8076) );
  NAND2_X1 U7715 ( .A1(n7330), .A2(n8076), .ZN(n7331) );
  AND2_X1 U7716 ( .A1(n7560), .A2(n8129), .ZN(n8135) );
  NAND2_X1 U7717 ( .A1(n7331), .A2(n8135), .ZN(n6112) );
  NAND2_X1 U7718 ( .A1(n6112), .A2(n8137), .ZN(n9793) );
  NAND2_X1 U7719 ( .A1(n6332), .A2(n10122), .ZN(n8134) );
  NAND2_X1 U7720 ( .A1(n7611), .A2(n10135), .ZN(n8138) );
  NAND2_X1 U7721 ( .A1(n8134), .A2(n8138), .ZN(n9795) );
  NAND2_X1 U7722 ( .A1(n9863), .A2(n10129), .ZN(n8149) );
  NAND2_X1 U7723 ( .A1(n6113), .A2(n8149), .ZN(n7627) );
  NAND2_X1 U7724 ( .A1(n7627), .A2(n7749), .ZN(n6114) );
  NAND2_X1 U7725 ( .A1(n6114), .A2(n8150), .ZN(n7798) );
  XNOR2_X1 U7726 ( .A(n9876), .B(n8766), .ZN(n8157) );
  INV_X1 U7727 ( .A(n8159), .ZN(n6116) );
  OR2_X1 U7728 ( .A1(n8157), .A2(n6116), .ZN(n8755) );
  INV_X1 U7729 ( .A(n8164), .ZN(n6117) );
  OR2_X1 U7730 ( .A1(n8755), .A2(n6117), .ZN(n6119) );
  OR2_X1 U7731 ( .A1(n9876), .A2(n8766), .ZN(n8769) );
  AND2_X1 U7732 ( .A1(n8769), .A2(n8160), .ZN(n6115) );
  OR2_X1 U7733 ( .A1(n6116), .A2(n6115), .ZN(n8756) );
  OR2_X1 U7734 ( .A1(n6117), .A2(n8756), .ZN(n6118) );
  OAI21_X1 U7735 ( .B1(n7798), .B2(n6119), .A(n4885), .ZN(n8733) );
  INV_X1 U7736 ( .A(n8188), .ZN(n8691) );
  INV_X1 U7737 ( .A(n8189), .ZN(n6121) );
  OR2_X1 U7738 ( .A1(n8691), .A2(n6121), .ZN(n6120) );
  NAND2_X1 U7739 ( .A1(n8385), .A2(n8706), .ZN(n8193) );
  NAND2_X1 U7740 ( .A1(n8189), .A2(n8193), .ZN(n8697) );
  INV_X1 U7741 ( .A(n8697), .ZN(n8086) );
  AND2_X1 U7742 ( .A1(n8086), .A2(n8692), .ZN(n8693) );
  OR2_X1 U7743 ( .A1(n6121), .A2(n8693), .ZN(n6122) );
  INV_X1 U7744 ( .A(n8181), .ZN(n6125) );
  INV_X1 U7745 ( .A(n8651), .ZN(n6124) );
  NOR2_X1 U7746 ( .A1(n6125), .A2(n6124), .ZN(n8200) );
  INV_X1 U7747 ( .A(n8179), .ZN(n8198) );
  INV_X1 U7748 ( .A(n8418), .ZN(n8824) );
  OR2_X1 U7749 ( .A1(n8817), .A2(n8824), .ZN(n8185) );
  NAND2_X1 U7750 ( .A1(n6126), .A2(n8811), .ZN(n8205) );
  NAND2_X1 U7751 ( .A1(n8639), .A2(n8818), .ZN(n8067) );
  NAND2_X1 U7752 ( .A1(n8205), .A2(n8067), .ZN(n8208) );
  INV_X1 U7753 ( .A(n6127), .ZN(n8214) );
  NAND2_X1 U7754 ( .A1(n8794), .A2(n8604), .ZN(n8065) );
  AOI21_X1 U7755 ( .B1(n8593), .B2(n8065), .A(n8222), .ZN(n8583) );
  NOR2_X1 U7756 ( .A1(n8236), .A2(n8793), .ZN(n6128) );
  OAI22_X1 U7757 ( .A1(n8583), .A2(n6128), .B1(n8592), .B2(n8787), .ZN(n8060)
         );
  NAND2_X1 U7758 ( .A1(n7573), .A2(n8095), .ZN(n6129) );
  AND2_X1 U7759 ( .A1(n9865), .A2(n6129), .ZN(n6130) );
  AND2_X1 U7760 ( .A1(n8558), .A2(n6130), .ZN(n6132) );
  NOR2_X1 U7761 ( .A1(n8227), .A2(n8095), .ZN(n6131) );
  NAND2_X1 U7762 ( .A1(n8558), .A2(n6131), .ZN(n6176) );
  NAND2_X1 U7763 ( .A1(n6132), .A2(n6176), .ZN(n7615) );
  INV_X1 U7764 ( .A(n6133), .ZN(n8251) );
  NAND2_X1 U7765 ( .A1(n8251), .A2(n8549), .ZN(n6135) );
  NAND2_X1 U7766 ( .A1(n5768), .A2(n6135), .ZN(n6141) );
  AND2_X1 U7767 ( .A1(n5768), .A2(P2_B_REG_SCAN_IN), .ZN(n6136) );
  NOR2_X1 U7768 ( .A1(n9813), .A2(n6136), .ZN(n8568) );
  NAND2_X1 U7769 ( .A1(n7058), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7770 ( .A1(n7059), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7771 ( .A1(n6137), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6138) );
  NAND4_X1 U7772 ( .A1(n7063), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n8415)
         );
  INV_X1 U7773 ( .A(n6141), .ZN(n6360) );
  AOI22_X1 U7774 ( .A1(n8568), .A2(n8415), .B1(n8793), .B2(n8728), .ZN(n6142)
         );
  OAI21_X1 U7775 ( .B1(n7878), .B2(n7615), .A(n6142), .ZN(n6143) );
  XNOR2_X1 U7776 ( .A(n7810), .B(P2_B_REG_SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7777 ( .A1(n7864), .A2(n6151), .ZN(n6160) );
  NAND4_X1 U7778 ( .A1(n6154), .A2(n6153), .A3(n6174), .A4(n6152), .ZN(n6155)
         );
  OAI21_X1 U7779 ( .B1(n6156), .B2(n6155), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6157) );
  MUX2_X1 U7780 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6157), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6159) );
  NAND2_X1 U7781 ( .A1(n7864), .A2(n7872), .ZN(n6550) );
  NAND2_X1 U7782 ( .A1(n7810), .A2(n7872), .ZN(n6553) );
  NOR4_X1 U7783 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6172) );
  NOR4_X1 U7784 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6167) );
  NOR4_X1 U7785 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6166) );
  NOR4_X1 U7786 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6165) );
  NOR4_X1 U7787 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7788 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n6168)
         );
  NOR4_X1 U7789 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6169), .A4(n6168), .ZN(n6171) );
  NOR4_X1 U7790 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6170) );
  AND3_X1 U7791 ( .A1(n6172), .A2(n6171), .A3(n6170), .ZN(n6173) );
  INV_X1 U7792 ( .A(n6176), .ZN(n7140) );
  NAND2_X1 U7793 ( .A1(n6974), .A2(n7140), .ZN(n6357) );
  AND3_X1 U7794 ( .A1(n8254), .A2(n8095), .A3(n8069), .ZN(n6177) );
  NAND2_X1 U7795 ( .A1(n6299), .A2(n6177), .ZN(n6338) );
  INV_X1 U7796 ( .A(n6338), .ZN(n6339) );
  NAND2_X1 U7797 ( .A1(n6974), .A2(n6339), .ZN(n6178) );
  NAND2_X1 U7798 ( .A1(n6357), .A2(n6178), .ZN(n6179) );
  NAND2_X1 U7799 ( .A1(n6353), .A2(n6179), .ZN(n6183) );
  NAND2_X1 U7800 ( .A1(n6195), .A2(n6194), .ZN(n6191) );
  NAND2_X1 U7801 ( .A1(n6989), .A2(n9877), .ZN(n8752) );
  NOR2_X1 U7802 ( .A1(n9877), .A2(n8246), .ZN(n6340) );
  NAND2_X1 U7803 ( .A1(n6338), .A2(n6340), .ZN(n6181) );
  NAND2_X1 U7804 ( .A1(n8752), .A2(n6181), .ZN(n6345) );
  NAND3_X1 U7805 ( .A1(n6358), .A2(n6974), .A3(n6345), .ZN(n6182) );
  OR2_X1 U7806 ( .A1(n9880), .A2(n6092), .ZN(n6184) );
  NAND2_X1 U7807 ( .A1(n6187), .A2(n6186), .ZN(P2_U3456) );
  NAND2_X1 U7808 ( .A1(n8558), .A2(n7365), .ZN(n6189) );
  NAND2_X1 U7809 ( .A1(n6189), .A2(n8246), .ZN(n6972) );
  AND4_X1 U7810 ( .A1(n6973), .A2(n6974), .A3(n6354), .A4(n6972), .ZN(n6190)
         );
  NAND3_X1 U7811 ( .A1(n8558), .A2(n8095), .A3(n8254), .ZN(n6192) );
  NAND2_X1 U7812 ( .A1(n6192), .A2(n8227), .ZN(n6193) );
  MUX2_X1 U7813 ( .A(n6195), .B(n6194), .S(n6193), .Z(n6971) );
  NAND2_X1 U7814 ( .A1(n6197), .A2(n9897), .ZN(n6203) );
  INV_X1 U7815 ( .A(n6098), .ZN(n6198) );
  NAND2_X1 U7816 ( .A1(n6203), .A2(n6202), .ZN(P2_U3488) );
  NAND2_X1 U7817 ( .A1(n6204), .A2(n9719), .ZN(n7108) );
  NAND2_X1 U7818 ( .A1(n6876), .A2(n6881), .ZN(n6875) );
  NAND2_X1 U7819 ( .A1(n6859), .A2(n6210), .ZN(n6849) );
  NAND2_X1 U7820 ( .A1(n6849), .A2(n6852), .ZN(n6848) );
  NAND2_X1 U7821 ( .A1(n7320), .A2(n6784), .ZN(n6211) );
  NAND2_X1 U7822 ( .A1(n6848), .A2(n6211), .ZN(n6838) );
  NAND2_X1 U7823 ( .A1(n6838), .A2(n6840), .ZN(n6837) );
  NAND2_X1 U7824 ( .A1(n6830), .A2(n7474), .ZN(n6212) );
  NAND2_X1 U7825 ( .A1(n6837), .A2(n6212), .ZN(n6826) );
  NAND2_X1 U7826 ( .A1(n6826), .A2(n6828), .ZN(n6825) );
  NAND2_X1 U7827 ( .A1(n6795), .A2(n9693), .ZN(n6213) );
  NAND2_X1 U7828 ( .A1(n6825), .A2(n6213), .ZN(n7082) );
  NAND2_X1 U7829 ( .A1(n7082), .A2(n7089), .ZN(n7081) );
  NAND2_X1 U7830 ( .A1(n7081), .A2(n4870), .ZN(n6994) );
  NAND2_X1 U7831 ( .A1(n7004), .A2(n6214), .ZN(n6999) );
  NAND2_X1 U7832 ( .A1(n6994), .A2(n6999), .ZN(n6993) );
  NAND2_X1 U7833 ( .A1(n7011), .A2(n7041), .ZN(n6215) );
  INV_X1 U7834 ( .A(n7192), .ZN(n9124) );
  NAND2_X1 U7835 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  INV_X1 U7836 ( .A(n7545), .ZN(n9120) );
  AOI21_X1 U7837 ( .B1(n7651), .B2(n7656), .A(n6223), .ZN(n7705) );
  NAND2_X1 U7838 ( .A1(n9538), .A2(n9119), .ZN(n6224) );
  AOI22_X1 U7839 ( .A1(n7705), .A2(n6224), .B1(n7536), .B2(n7719), .ZN(n7637)
         );
  INV_X1 U7840 ( .A(n7920), .ZN(n9117) );
  INV_X1 U7841 ( .A(n9521), .ZN(n7931) );
  NAND2_X1 U7842 ( .A1(n9581), .A2(n8965), .ZN(n6229) );
  NAND2_X1 U7843 ( .A1(n9512), .A2(n9114), .ZN(n6231) );
  NOR2_X1 U7844 ( .A1(n9512), .A2(n9114), .ZN(n6230) );
  NAND2_X1 U7845 ( .A1(n9386), .A2(n7947), .ZN(n6232) );
  NAND2_X1 U7846 ( .A1(n9380), .A2(n6232), .ZN(n6234) );
  NAND2_X1 U7847 ( .A1(n9505), .A2(n9113), .ZN(n6233) );
  NAND2_X1 U7848 ( .A1(n6234), .A2(n6233), .ZN(n9363) );
  NOR2_X1 U7849 ( .A1(n9575), .A2(n9057), .ZN(n6236) );
  NAND2_X1 U7850 ( .A1(n9575), .A2(n9057), .ZN(n6235) );
  NOR2_X1 U7851 ( .A1(n9344), .A2(n9058), .ZN(n6237) );
  NOR2_X1 U7852 ( .A1(n9566), .A2(n9083), .ZN(n6239) );
  NAND2_X1 U7853 ( .A1(n9566), .A2(n9083), .ZN(n6238) );
  OAI21_X1 U7854 ( .B1(n9300), .B2(n6239), .A(n6238), .ZN(n9285) );
  NOR2_X1 U7855 ( .A1(n9293), .A2(n9109), .ZN(n6241) );
  NAND2_X1 U7856 ( .A1(n9558), .A2(n9081), .ZN(n6242) );
  OAI21_X1 U7857 ( .B1(n9265), .B2(n9268), .A(n6242), .ZN(n9250) );
  NAND2_X1 U7858 ( .A1(n9250), .A2(n9249), .ZN(n9248) );
  NAND2_X1 U7859 ( .A1(n9248), .A2(n6243), .ZN(n6244) );
  INV_X1 U7860 ( .A(n9720), .ZN(n6245) );
  AND2_X1 U7861 ( .A1(n6246), .A2(n6245), .ZN(n9707) );
  NAND2_X1 U7862 ( .A1(n6479), .A2(n6482), .ZN(n6247) );
  AND2_X1 U7863 ( .A1(n9707), .A2(n6247), .ZN(n9446) );
  NAND2_X1 U7864 ( .A1(n6251), .A2(n6250), .ZN(n9356) );
  OR2_X2 U7865 ( .A1(n9356), .A2(n9357), .ZN(n9354) );
  OR2_X2 U7866 ( .A1(n9335), .A2(n9336), .ZN(n9333) );
  NAND2_X1 U7867 ( .A1(n9304), .A2(n6255), .ZN(n9287) );
  NAND2_X1 U7868 ( .A1(n9269), .A2(n6256), .ZN(n6257) );
  INV_X1 U7869 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U7870 ( .A1(n9229), .A2(n6478), .ZN(n6264) );
  NAND2_X1 U7871 ( .A1(n6262), .A2(n6597), .ZN(n6263) );
  NAND2_X1 U7872 ( .A1(n6265), .A2(n9391), .ZN(n6268) );
  INV_X1 U7873 ( .A(n5695), .ZN(n6434) );
  NAND2_X1 U7874 ( .A1(n5695), .A2(n6594), .ZN(n9080) );
  INV_X1 U7875 ( .A(n5696), .ZN(n9594) );
  AND2_X1 U7876 ( .A1(n9594), .A2(P1_B_REG_SCAN_IN), .ZN(n6266) );
  NOR2_X1 U7877 ( .A1(n9080), .A2(n6266), .ZN(n9237) );
  AOI22_X1 U7878 ( .A1(n9108), .A2(n9070), .B1(n9237), .B2(n9107), .ZN(n6267)
         );
  NAND2_X1 U7879 ( .A1(n6268), .A2(n6267), .ZN(n8287) );
  NAND2_X1 U7880 ( .A1(n6860), .A2(n6964), .ZN(n6861) );
  AND2_X1 U7881 ( .A1(n6839), .A2(n9693), .ZN(n7083) );
  NAND2_X1 U7882 ( .A1(n7452), .A2(n4772), .ZN(n7453) );
  OR2_X2 U7883 ( .A1(n7853), .A2(n9521), .ZN(n9419) );
  INV_X1 U7884 ( .A(n9512), .ZN(n9409) );
  AND2_X2 U7885 ( .A1(n9323), .A2(n9566), .ZN(n9308) );
  INV_X2 U7886 ( .A(n9242), .ZN(n9418) );
  AOI211_X1 U7887 ( .C1(n6291), .C2(n9256), .A(n9418), .B(n9243), .ZN(n8281)
         );
  OAI21_X1 U7888 ( .B1(n8289), .B2(n9716), .A(n6269), .ZN(n6294) );
  NAND2_X1 U7889 ( .A1(n7867), .A2(P1_B_REG_SCAN_IN), .ZN(n6272) );
  MUX2_X1 U7890 ( .A(P1_B_REG_SCAN_IN), .B(n6272), .S(n7807), .Z(n6274) );
  INV_X1 U7891 ( .A(n7870), .ZN(n6273) );
  NOR2_X1 U7892 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n6278) );
  NOR4_X1 U7893 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6277) );
  NOR4_X1 U7894 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6276) );
  NOR4_X1 U7895 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6275) );
  NAND4_X1 U7896 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n6284)
         );
  NOR4_X1 U7897 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6282) );
  NOR4_X1 U7898 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6281) );
  NOR4_X1 U7899 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6280) );
  NOR4_X1 U7900 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6279) );
  NAND4_X1 U7901 ( .A1(n6282), .A2(n6281), .A3(n6280), .A4(n6279), .ZN(n6283)
         );
  NOR2_X1 U7902 ( .A1(n6284), .A2(n6283), .ZN(n6592) );
  NAND2_X1 U7903 ( .A1(n6600), .A2(n6592), .ZN(n6285) );
  NAND2_X1 U7904 ( .A1(n9711), .A2(n6285), .ZN(n6286) );
  NAND2_X1 U7905 ( .A1(n6479), .A2(n6594), .ZN(n6606) );
  NAND2_X1 U7906 ( .A1(n6286), .A2(n6606), .ZN(n6956) );
  OR2_X1 U7907 ( .A1(n6591), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7908 ( .A1(n7870), .A2(n7867), .ZN(n9590) );
  NAND2_X1 U7909 ( .A1(n6287), .A2(n9590), .ZN(n6589) );
  NAND2_X1 U7910 ( .A1(n9229), .A2(n9242), .ZN(n6603) );
  NAND2_X1 U7911 ( .A1(n6589), .A2(n6603), .ZN(n6288) );
  NAND2_X1 U7912 ( .A1(n7870), .A2(n7807), .ZN(n9591) );
  INV_X1 U7913 ( .A(n6953), .ZN(n6590) );
  MUX2_X1 U7914 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n6294), .S(n9738), .Z(n6290)
         );
  INV_X1 U7915 ( .A(n6290), .ZN(n6292) );
  NAND2_X1 U7916 ( .A1(n6292), .A2(n4876), .ZN(P1_U3519) );
  MUX2_X1 U7917 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n6294), .S(n9745), .Z(n6295)
         );
  INV_X1 U7918 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7919 ( .A1(n6296), .A2(n4872), .ZN(P1_U3551) );
  INV_X1 U7920 ( .A(n6297), .ZN(n6298) );
  INV_X1 U7921 ( .A(n6369), .ZN(n7625) );
  NAND2_X1 U7922 ( .A1(n6299), .A2(n8069), .ZN(n6301) );
  NAND2_X2 U7923 ( .A1(n6301), .A2(n6300), .ZN(n6308) );
  INV_X1 U7924 ( .A(n8872), .ZN(n6927) );
  NAND2_X1 U7925 ( .A1(n6308), .A2(n6927), .ZN(n6303) );
  NAND2_X1 U7926 ( .A1(n8070), .A2(n6303), .ZN(n6894) );
  NAND2_X1 U7927 ( .A1(n6894), .A2(n6895), .ZN(n6307) );
  NAND2_X1 U7928 ( .A1(n6305), .A2(n6984), .ZN(n6306) );
  NAND2_X1 U7929 ( .A1(n6307), .A2(n6306), .ZN(n6900) );
  XNOR2_X1 U7930 ( .A(n6308), .B(n6979), .ZN(n6309) );
  XNOR2_X1 U7931 ( .A(n6309), .B(n8431), .ZN(n6901) );
  NAND2_X1 U7932 ( .A1(n6900), .A2(n6901), .ZN(n6311) );
  INV_X1 U7933 ( .A(n8431), .ZN(n9814) );
  NAND2_X1 U7934 ( .A1(n6309), .A2(n9814), .ZN(n6310) );
  NAND2_X1 U7935 ( .A1(n6311), .A2(n6310), .ZN(n6819) );
  INV_X1 U7936 ( .A(n6819), .ZN(n6313) );
  XNOR2_X1 U7937 ( .A(n6308), .B(n6915), .ZN(n6314) );
  XNOR2_X1 U7938 ( .A(n6314), .B(n8430), .ZN(n6820) );
  INV_X1 U7939 ( .A(n6820), .ZN(n6312) );
  NAND2_X1 U7940 ( .A1(n6314), .A2(n8430), .ZN(n6315) );
  NAND2_X1 U7941 ( .A1(n6821), .A2(n6315), .ZN(n6945) );
  INV_X1 U7942 ( .A(n6945), .ZN(n6317) );
  XNOR2_X1 U7943 ( .A(n6318), .B(n8429), .ZN(n6946) );
  INV_X1 U7944 ( .A(n6946), .ZN(n6316) );
  NAND2_X1 U7945 ( .A1(n6317), .A2(n6316), .ZN(n6943) );
  INV_X1 U7946 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U7947 ( .A1(n6319), .A2(n7146), .ZN(n6320) );
  NAND2_X1 U7948 ( .A1(n6943), .A2(n6320), .ZN(n7149) );
  XNOR2_X1 U7949 ( .A(n8261), .B(n9830), .ZN(n6321) );
  XNOR2_X1 U7950 ( .A(n6321), .B(n7242), .ZN(n7150) );
  NAND2_X1 U7951 ( .A1(n7149), .A2(n7150), .ZN(n6324) );
  INV_X1 U7952 ( .A(n6321), .ZN(n6322) );
  NAND2_X1 U7953 ( .A1(n6322), .A2(n7242), .ZN(n6323) );
  NAND2_X1 U7954 ( .A1(n6324), .A2(n6323), .ZN(n7238) );
  XNOR2_X1 U7955 ( .A(n8261), .B(n9836), .ZN(n6327) );
  XNOR2_X1 U7956 ( .A(n6327), .B(n8427), .ZN(n7239) );
  XNOR2_X1 U7957 ( .A(n8261), .B(n9841), .ZN(n6326) );
  INV_X1 U7958 ( .A(n6326), .ZN(n6325) );
  AND2_X1 U7959 ( .A1(n6325), .A2(n7564), .ZN(n6329) );
  OR2_X1 U7960 ( .A1(n7239), .A2(n6329), .ZN(n6331) );
  XNOR2_X1 U7961 ( .A(n6326), .B(n8426), .ZN(n7372) );
  INV_X1 U7962 ( .A(n7372), .ZN(n6328) );
  NAND2_X1 U7963 ( .A1(n6327), .A2(n8427), .ZN(n7367) );
  AND2_X1 U7964 ( .A1(n6328), .A2(n7367), .ZN(n7368) );
  OR2_X1 U7965 ( .A1(n6329), .A2(n7368), .ZN(n6330) );
  OAI21_X1 U7966 ( .B1(n7238), .B2(n6331), .A(n6330), .ZN(n7553) );
  XNOR2_X1 U7967 ( .A(n6332), .B(n8261), .ZN(n10123) );
  XNOR2_X1 U7968 ( .A(n8261), .B(n7557), .ZN(n10119) );
  INV_X1 U7969 ( .A(n10119), .ZN(n6333) );
  AOI22_X1 U7970 ( .A1(n7611), .A2(n10123), .B1(n6333), .B2(n10130), .ZN(n6337) );
  AOI21_X1 U7971 ( .B1(n10119), .B2(n10120), .A(n10122), .ZN(n6335) );
  NAND3_X1 U7972 ( .A1(n10119), .A2(n10120), .A3(n10122), .ZN(n6334) );
  OAI21_X1 U7973 ( .B1(n6335), .B2(n10123), .A(n6334), .ZN(n6336) );
  XNOR2_X1 U7974 ( .A(n7750), .B(n10129), .ZN(n7753) );
  XNOR2_X1 U7975 ( .A(n9863), .B(n8261), .ZN(n7752) );
  XOR2_X1 U7976 ( .A(n7753), .B(n7752), .Z(n6344) );
  OR2_X1 U7977 ( .A1(n6358), .A2(n6338), .ZN(n6348) );
  INV_X1 U7978 ( .A(n6348), .ZN(n6343) );
  AOI21_X1 U7979 ( .B1(n6353), .B2(n6340), .A(n6339), .ZN(n6342) );
  INV_X1 U7980 ( .A(n6974), .ZN(n6341) );
  NOR2_X1 U7981 ( .A1(n6344), .A2(n8383), .ZN(n6368) );
  INV_X1 U7982 ( .A(n6345), .ZN(n6349) );
  AND3_X1 U7983 ( .A1(n6346), .A2(n6369), .A3(n6972), .ZN(n6347) );
  OAI211_X1 U7984 ( .C1(n6353), .C2(n6349), .A(n6348), .B(n6347), .ZN(n6350)
         );
  NAND2_X1 U7985 ( .A1(n6350), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6352) );
  OR2_X1 U7986 ( .A1(n6358), .A2(n6357), .ZN(n6351) );
  NOR2_X1 U7987 ( .A1(n10138), .A2(n7616), .ZN(n6367) );
  INV_X1 U7988 ( .A(n8752), .ZN(n8768) );
  NAND3_X1 U7989 ( .A1(n6353), .A2(n6974), .A3(n8768), .ZN(n6356) );
  AND2_X1 U7990 ( .A1(n10134), .A2(n9863), .ZN(n6366) );
  INV_X1 U7991 ( .A(n6357), .ZN(n8252) );
  AND2_X1 U7992 ( .A1(n6358), .A2(n8252), .ZN(n6361) );
  INV_X1 U7993 ( .A(n6361), .ZN(n6359) );
  NAND2_X1 U7994 ( .A1(n8409), .A2(n10122), .ZN(n6364) );
  INV_X1 U7995 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6362) );
  NOR2_X1 U7996 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6362), .ZN(n7600) );
  INV_X1 U7997 ( .A(n7600), .ZN(n6363) );
  OAI211_X1 U7998 ( .C1(n7796), .C2(n10128), .A(n6364), .B(n6363), .ZN(n6365)
         );
  OR4_X1 U7999 ( .A1(n6368), .A2(n6367), .A3(n6366), .A4(n6365), .ZN(P2_U3157)
         );
  NAND2_X1 U8000 ( .A1(n6369), .A2(n8246), .ZN(n6370) );
  NAND2_X1 U8001 ( .A1(n6631), .A2(n6370), .ZN(n6654) );
  OAI21_X1 U8002 ( .B1(n6654), .B2(n6371), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X2 U8003 ( .A(n7888), .ZN(n8273) );
  OAI222_X1 U8004 ( .A1(P1_U3086), .A2(n6436), .B1(n8271), .B2(n6391), .C1(
        n4538), .C2(n8273), .ZN(P1_U3353) );
  OAI222_X1 U8005 ( .A1(P1_U3086), .A2(n6441), .B1(n8271), .B2(n6377), .C1(
        n6374), .C2(n8273), .ZN(P1_U3352) );
  OAI222_X1 U8006 ( .A1(n6375), .A2(n8273), .B1(P1_U3086), .B2(n6443), .C1(
        n8271), .C2(n6389), .ZN(P1_U3351) );
  NOR2_X1 U8007 ( .A1(n6376), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7893) );
  INV_X2 U8008 ( .A(n7893), .ZN(n8277) );
  NAND2_X1 U8009 ( .A1(n6376), .A2(P2_U3151), .ZN(n8280) );
  OAI222_X1 U8010 ( .A1(n8277), .A2(n6378), .B1(n8280), .B2(n6377), .C1(
        P2_U3151), .C2(n6673), .ZN(P2_U3292) );
  INV_X1 U8011 ( .A(n8271), .ZN(n7620) );
  INV_X1 U8012 ( .A(n7620), .ZN(n8275) );
  OAI222_X1 U8013 ( .A1(n8275), .A2(n6392), .B1(n8273), .B2(n5445), .C1(
        P1_U3086), .C2(n6438), .ZN(P1_U3354) );
  OAI222_X1 U8014 ( .A1(n8277), .A2(n6379), .B1(n8280), .B2(n6380), .C1(
        P2_U3151), .C2(n6745), .ZN(P2_U3290) );
  OAI222_X1 U8015 ( .A1(n8273), .A2(n6381), .B1(n8271), .B2(n6380), .C1(
        P1_U3086), .C2(n6445), .ZN(P1_U3350) );
  OAI222_X1 U8016 ( .A1(n8273), .A2(n6382), .B1(n8271), .B2(n6387), .C1(
        P1_U3086), .C2(n9170), .ZN(P1_U3349) );
  NAND2_X1 U8017 ( .A1(n6204), .A2(P1_U3973), .ZN(n6383) );
  OAI21_X1 U8018 ( .B1(P1_U3973), .B2(n4896), .A(n6383), .ZN(P1_U3554) );
  OAI222_X1 U8019 ( .A1(n8277), .A2(n6384), .B1(n8280), .B2(n6385), .C1(
        P2_U3151), .C2(n7288), .ZN(P2_U3288) );
  OAI222_X1 U8020 ( .A1(n8273), .A2(n6386), .B1(n8271), .B2(n6385), .C1(
        P1_U3086), .C2(n9184), .ZN(P1_U3348) );
  INV_X1 U8021 ( .A(n8280), .ZN(n8941) );
  OAI222_X1 U8022 ( .A1(n8277), .A2(n6388), .B1(n8937), .B2(n6387), .C1(
        P2_U3151), .C2(n6764), .ZN(P2_U3289) );
  OAI222_X1 U8023 ( .A1(n8277), .A2(n6390), .B1(n8937), .B2(n6389), .C1(
        P2_U3151), .C2(n6698), .ZN(P2_U3291) );
  OAI222_X1 U8024 ( .A1(n8277), .A2(n4902), .B1(n8937), .B2(n6391), .C1(
        P2_U3151), .C2(n6658), .ZN(P2_U3293) );
  OAI222_X1 U8025 ( .A1(P2_U3151), .A2(n4590), .B1(n8277), .B2(n6393), .C1(
        n8937), .C2(n6392), .ZN(P2_U3294) );
  AOI22_X1 U8026 ( .A1(n9201), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7888), .ZN(n6394) );
  OAI21_X1 U8027 ( .B1(n6399), .B2(n8271), .A(n6394), .ZN(P1_U3347) );
  INV_X1 U8028 ( .A(n7621), .ZN(n6609) );
  NOR2_X1 U8029 ( .A1(n6600), .A2(n6609), .ZN(n6431) );
  INV_X1 U8030 ( .A(n6431), .ZN(n6398) );
  NAND2_X1 U8031 ( .A1(n6594), .A2(n6395), .ZN(n6396) );
  NAND2_X1 U8032 ( .A1(n6397), .A2(n6396), .ZN(n6432) );
  AND2_X1 U8033 ( .A1(n6398), .A2(n6432), .ZN(n9597) );
  NOR2_X1 U8034 ( .A1(n9597), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8035 ( .A1(n8277), .A2(n6400), .B1(n8937), .B2(n6399), .C1(
        P2_U3151), .C2(n7506), .ZN(P2_U3287) );
  INV_X1 U8036 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8037 ( .A1(n9238), .A2(P1_U3973), .ZN(n6401) );
  OAI21_X1 U8038 ( .B1(P1_U3973), .B2(n6402), .A(n6401), .ZN(P1_U3585) );
  INV_X1 U8039 ( .A(n6403), .ZN(n6409) );
  AOI22_X1 U8040 ( .A1(n6533), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7888), .ZN(n6404) );
  OAI21_X1 U8041 ( .B1(n6409), .B2(n8271), .A(n6404), .ZN(P1_U3345) );
  INV_X1 U8042 ( .A(n6405), .ZN(n6407) );
  OAI222_X1 U8043 ( .A1(n8277), .A2(n6406), .B1(n8937), .B2(n6407), .C1(n4690), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8044 ( .A(n6467), .ZN(n6460) );
  OAI222_X1 U8045 ( .A1(n8273), .A2(n6408), .B1(n8275), .B2(n6407), .C1(n6460), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8046 ( .A(n7676), .ZN(n7667) );
  OAI222_X1 U8047 ( .A1(n8277), .A2(n6410), .B1(n8280), .B2(n6409), .C1(n7667), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8048 ( .A(n6411), .ZN(n6413) );
  INV_X1 U8049 ( .A(n6538), .ZN(n9611) );
  OAI222_X1 U8050 ( .A1(n8273), .A2(n6412), .B1(n8271), .B2(n6413), .C1(
        P1_U3086), .C2(n9611), .ZN(P1_U3344) );
  OAI222_X1 U8051 ( .A1(n8277), .A2(n6414), .B1(n8280), .B2(n6413), .C1(
        P2_U3151), .C2(n7685), .ZN(P2_U3284) );
  INV_X1 U8052 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6415) );
  MUX2_X1 U8053 ( .A(n6415), .B(P1_REG1_REG_9__SCAN_IN), .S(n6467), .Z(n6430)
         );
  INV_X1 U8054 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6416) );
  MUX2_X1 U8055 ( .A(n6416), .B(P1_REG1_REG_2__SCAN_IN), .S(n6436), .Z(n6513)
         );
  INV_X1 U8056 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9741) );
  MUX2_X1 U8057 ( .A(n9741), .B(P1_REG1_REG_1__SCAN_IN), .S(n6438), .Z(n9136)
         );
  AND2_X1 U8058 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n9596), .ZN(n9135) );
  NAND2_X1 U8059 ( .A1(n9136), .A2(n9135), .ZN(n9134) );
  INV_X1 U8060 ( .A(n6438), .ZN(n9137) );
  NAND2_X1 U8061 ( .A1(n9137), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8062 ( .A1(n9134), .A2(n6417), .ZN(n6512) );
  NAND2_X1 U8063 ( .A1(n6513), .A2(n6512), .ZN(n6511) );
  INV_X1 U8064 ( .A(n6436), .ZN(n6514) );
  NAND2_X1 U8065 ( .A1(n6514), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8066 ( .A1(n6511), .A2(n6418), .ZN(n9149) );
  XNOR2_X1 U8067 ( .A(n6441), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U8068 ( .A1(n9149), .A2(n9150), .ZN(n9148) );
  INV_X1 U8069 ( .A(n6441), .ZN(n9147) );
  NAND2_X1 U8070 ( .A1(n9147), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8071 ( .A1(n9148), .A2(n6419), .ZN(n6499) );
  INV_X1 U8072 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6420) );
  MUX2_X1 U8073 ( .A(n6420), .B(P1_REG1_REG_4__SCAN_IN), .S(n6443), .Z(n6500)
         );
  NAND2_X1 U8074 ( .A1(n6499), .A2(n6500), .ZN(n6498) );
  INV_X1 U8075 ( .A(n6443), .ZN(n6502) );
  NAND2_X1 U8076 ( .A1(n6502), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U8077 ( .A1(n6498), .A2(n6421), .ZN(n9162) );
  INV_X1 U8078 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9929) );
  MUX2_X1 U8079 ( .A(n9929), .B(P1_REG1_REG_5__SCAN_IN), .S(n6445), .Z(n9163)
         );
  NAND2_X1 U8080 ( .A1(n9162), .A2(n9163), .ZN(n9161) );
  INV_X1 U8081 ( .A(n6445), .ZN(n9160) );
  NAND2_X1 U8082 ( .A1(n9160), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U8083 ( .A1(n9161), .A2(n6422), .ZN(n9176) );
  INV_X1 U8084 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6423) );
  MUX2_X1 U8085 ( .A(n6423), .B(P1_REG1_REG_6__SCAN_IN), .S(n9170), .Z(n9177)
         );
  NAND2_X1 U8086 ( .A1(n9176), .A2(n9177), .ZN(n9175) );
  OR2_X1 U8087 ( .A1(n9170), .A2(n6423), .ZN(n6424) );
  NAND2_X1 U8088 ( .A1(n9175), .A2(n6424), .ZN(n9193) );
  INV_X1 U8089 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9952) );
  MUX2_X1 U8090 ( .A(n9952), .B(P1_REG1_REG_7__SCAN_IN), .S(n9184), .Z(n9194)
         );
  NAND2_X1 U8091 ( .A1(n9193), .A2(n9194), .ZN(n9192) );
  OR2_X1 U8092 ( .A1(n9184), .A2(n9952), .ZN(n6425) );
  NAND2_X1 U8093 ( .A1(n9192), .A2(n6425), .ZN(n9206) );
  INV_X1 U8094 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U8095 ( .A(n9201), .B(n6426), .ZN(n9207) );
  NAND2_X1 U8096 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  NAND2_X1 U8097 ( .A1(n9201), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8098 ( .A1(n9205), .A2(n6427), .ZN(n6429) );
  OR2_X1 U8099 ( .A1(n6429), .A2(n6430), .ZN(n6469) );
  INV_X1 U8100 ( .A(n6469), .ZN(n6428) );
  AOI21_X1 U8101 ( .B1(n6430), .B2(n6429), .A(n6428), .ZN(n6458) );
  INV_X1 U8102 ( .A(n9599), .ZN(n6433) );
  NAND2_X1 U8103 ( .A1(n6433), .A2(n5696), .ZN(n9645) );
  NOR2_X2 U8104 ( .A1(n9599), .A2(n6434), .ZN(n9656) );
  INV_X1 U8105 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8106 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7255) );
  OAI21_X1 U8107 ( .B1(n9676), .B2(n6435), .A(n7255), .ZN(n6456) );
  INV_X1 U8108 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6437) );
  MUX2_X1 U8109 ( .A(n6437), .B(P1_REG2_REG_2__SCAN_IN), .S(n6436), .Z(n6517)
         );
  INV_X1 U8110 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7115) );
  MUX2_X1 U8111 ( .A(n7115), .B(P1_REG2_REG_1__SCAN_IN), .S(n6438), .Z(n9140)
         );
  AND2_X1 U8112 ( .A1(n9596), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U8113 ( .A1(n9140), .A2(n9139), .ZN(n9138) );
  NAND2_X1 U8114 ( .A1(n9137), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8115 ( .A1(n9138), .A2(n6439), .ZN(n6516) );
  NAND2_X1 U8116 ( .A1(n6517), .A2(n6516), .ZN(n6515) );
  NAND2_X1 U8117 ( .A1(n6514), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8118 ( .A1(n6515), .A2(n6440), .ZN(n9152) );
  XNOR2_X1 U8119 ( .A(n6441), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U8120 ( .A1(n9152), .A2(n9153), .ZN(n9151) );
  NAND2_X1 U8121 ( .A1(n9147), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8122 ( .A1(n9151), .A2(n6442), .ZN(n6504) );
  INV_X1 U8123 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7322) );
  MUX2_X1 U8124 ( .A(n7322), .B(P1_REG2_REG_4__SCAN_IN), .S(n6443), .Z(n6505)
         );
  NAND2_X1 U8125 ( .A1(n6504), .A2(n6505), .ZN(n6503) );
  NAND2_X1 U8126 ( .A1(n6502), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8127 ( .A1(n6503), .A2(n6444), .ZN(n9165) );
  XNOR2_X1 U8128 ( .A(n6445), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U8129 ( .A1(n9165), .A2(n9166), .ZN(n9164) );
  NAND2_X1 U8130 ( .A1(n9160), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8131 ( .A1(n9164), .A2(n6446), .ZN(n9179) );
  INV_X1 U8132 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U8133 ( .A(n10097), .B(P1_REG2_REG_6__SCAN_IN), .S(n9170), .Z(n9180)
         );
  NAND2_X1 U8134 ( .A1(n9179), .A2(n9180), .ZN(n9178) );
  OR2_X1 U8135 ( .A1(n9170), .A2(n10097), .ZN(n6447) );
  NAND2_X1 U8136 ( .A1(n9178), .A2(n6447), .ZN(n9190) );
  XNOR2_X1 U8137 ( .A(n9184), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U8138 ( .A1(n9190), .A2(n9191), .ZN(n9189) );
  INV_X1 U8139 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8140 ( .A1(n9184), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U8141 ( .A1(n9189), .A2(n6449), .ZN(n9203) );
  INV_X1 U8142 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9443) );
  XNOR2_X1 U8143 ( .A(n9201), .B(n9443), .ZN(n9204) );
  NAND2_X1 U8144 ( .A1(n9203), .A2(n9204), .ZN(n9202) );
  NAND2_X1 U8145 ( .A1(n9201), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8146 ( .A1(n9202), .A2(n6450), .ZN(n6452) );
  XNOR2_X1 U8147 ( .A(n6467), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6451) );
  OR2_X1 U8148 ( .A1(n6452), .A2(n6451), .ZN(n6462) );
  NAND2_X1 U8149 ( .A1(n6452), .A2(n6451), .ZN(n6454) );
  INV_X1 U8150 ( .A(n6494), .ZN(n6453) );
  NOR2_X2 U8151 ( .A1(n9599), .A2(n6453), .ZN(n9660) );
  INV_X1 U8152 ( .A(n9660), .ZN(n9649) );
  AOI21_X1 U8153 ( .B1(n6462), .B2(n6454), .A(n9649), .ZN(n6455) );
  AOI211_X1 U8154 ( .C1(n9656), .C2(n6467), .A(n6456), .B(n6455), .ZN(n6457)
         );
  OAI21_X1 U8155 ( .B1(n6458), .B2(n9645), .A(n6457), .ZN(P1_U3252) );
  NAND2_X1 U8156 ( .A1(n9132), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6459) );
  OAI21_X1 U8157 ( .B1(n9057), .B2(n9132), .A(n6459), .ZN(P1_U3575) );
  XNOR2_X1 U8158 ( .A(n6533), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6465) );
  INV_X1 U8159 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U8160 ( .A1(n6460), .A2(n9430), .ZN(n6461) );
  NAND2_X1 U8161 ( .A1(n6462), .A2(n6461), .ZN(n6464) );
  OR2_X1 U8162 ( .A1(n6464), .A2(n6465), .ZN(n6535) );
  INV_X1 U8163 ( .A(n6535), .ZN(n6463) );
  AOI211_X1 U8164 ( .C1(n6465), .C2(n6464), .A(n9649), .B(n6463), .ZN(n6477)
         );
  INV_X1 U8165 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6466) );
  MUX2_X1 U8166 ( .A(n6466), .B(P1_REG1_REG_10__SCAN_IN), .S(n6533), .Z(n6472)
         );
  OR2_X1 U8167 ( .A1(n6467), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8168 ( .A1(n6469), .A2(n6468), .ZN(n6471) );
  OR2_X1 U8169 ( .A1(n6471), .A2(n6472), .ZN(n6525) );
  INV_X1 U8170 ( .A(n6525), .ZN(n6470) );
  AOI211_X1 U8171 ( .C1(n6472), .C2(n6471), .A(n9645), .B(n6470), .ZN(n6476)
         );
  INV_X1 U8172 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U8173 ( .A1(n9656), .A2(n6533), .ZN(n6474) );
  NAND2_X1 U8174 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n6473) );
  OAI211_X1 U8175 ( .C1(n7413), .C2(n9676), .A(n6474), .B(n6473), .ZN(n6475)
         );
  OR3_X1 U8176 ( .A1(n6477), .A2(n6476), .A3(n6475), .ZN(P1_U3253) );
  NAND3_X4 U8177 ( .A1(n6481), .A2(n6605), .A3(n7049), .ZN(n8977) );
  NAND3_X4 U8178 ( .A1(n6482), .A2(n6605), .A3(n6483), .ZN(n7975) );
  INV_X1 U8179 ( .A(n6483), .ZN(n6484) );
  AND2_X2 U8180 ( .A1(n6605), .A2(n6484), .ZN(n7965) );
  INV_X1 U8181 ( .A(n6605), .ZN(n6488) );
  NAND2_X1 U8182 ( .A1(n6488), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8183 ( .A1(n6204), .A2(n7977), .ZN(n6490) );
  AOI22_X1 U8184 ( .A1(n9719), .A2(n7965), .B1(n9596), .B2(n6488), .ZN(n6489)
         );
  NAND2_X1 U8185 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  NAND2_X1 U8186 ( .A1(n6492), .A2(n6491), .ZN(n6572) );
  OAI21_X1 U8187 ( .B1(n6492), .B2(n6491), .A(n6572), .ZN(n6719) );
  NOR2_X1 U8188 ( .A1(n5695), .A2(n9594), .ZN(n6497) );
  INV_X1 U8189 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U8190 ( .A1(n5696), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6493) );
  NOR2_X1 U8191 ( .A1(n5695), .A2(n6493), .ZN(n9593) );
  NAND2_X1 U8192 ( .A1(n6494), .A2(n9139), .ZN(n6495) );
  OAI211_X1 U8193 ( .C1(n9593), .C2(n9596), .A(n6495), .B(P1_U3973), .ZN(n6496) );
  AOI21_X1 U8194 ( .B1(n6719), .B2(n6497), .A(n6496), .ZN(n6523) );
  OAI211_X1 U8195 ( .C1(n6500), .C2(n6499), .A(n9664), .B(n6498), .ZN(n6509)
         );
  NAND2_X1 U8196 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6740) );
  INV_X1 U8197 ( .A(n6740), .ZN(n6501) );
  AOI21_X1 U8198 ( .B1(n9597), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6501), .ZN(
        n6508) );
  NAND2_X1 U8199 ( .A1(n9656), .A2(n6502), .ZN(n6507) );
  OAI211_X1 U8200 ( .C1(n6505), .C2(n6504), .A(n9660), .B(n6503), .ZN(n6506)
         );
  NAND4_X1 U8201 ( .A1(n6509), .A2(n6508), .A3(n6507), .A4(n6506), .ZN(n6510)
         );
  OR2_X1 U8202 ( .A1(n6523), .A2(n6510), .ZN(P1_U3247) );
  OAI211_X1 U8203 ( .C1(n6513), .C2(n6512), .A(n9664), .B(n6511), .ZN(n6521)
         );
  AOI22_X1 U8204 ( .A1(n9597), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6520) );
  NAND2_X1 U8205 ( .A1(n9656), .A2(n6514), .ZN(n6519) );
  OAI211_X1 U8206 ( .C1(n6517), .C2(n6516), .A(n9660), .B(n6515), .ZN(n6518)
         );
  NAND4_X1 U8207 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n6522)
         );
  OR2_X1 U8208 ( .A1(n6523), .A2(n6522), .ZN(P1_U3245) );
  NAND2_X1 U8209 ( .A1(n6533), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8210 ( .A1(n6525), .A2(n6524), .ZN(n9602) );
  INV_X1 U8211 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6526) );
  MUX2_X1 U8212 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6526), .S(n6538), .Z(n9601)
         );
  AND2_X1 U8213 ( .A1(n9602), .A2(n9601), .ZN(n9604) );
  AOI21_X1 U8214 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6538), .A(n9604), .ZN(
        n6528) );
  INV_X1 U8215 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10067) );
  INV_X1 U8216 ( .A(n7126), .ZN(n6545) );
  AOI22_X1 U8217 ( .A1(n7126), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n10067), .B2(
        n6545), .ZN(n6527) );
  NAND2_X1 U8218 ( .A1(n6528), .A2(n6527), .ZN(n7121) );
  OAI21_X1 U8219 ( .B1(n6528), .B2(n6527), .A(n7121), .ZN(n6531) );
  INV_X1 U8220 ( .A(n9656), .ZN(n9671) );
  NAND2_X1 U8221 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7232) );
  NAND2_X1 U8222 ( .A1(n9597), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6529) );
  OAI211_X1 U8223 ( .C1(n9671), .C2(n6545), .A(n7232), .B(n6529), .ZN(n6530)
         );
  AOI21_X1 U8224 ( .B1(n6531), .B2(n9664), .A(n6530), .ZN(n6543) );
  NOR2_X1 U8225 ( .A1(n7126), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6532) );
  AOI21_X1 U8226 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7126), .A(n6532), .ZN(
        n6540) );
  NAND2_X1 U8227 ( .A1(n6533), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8228 ( .A1(n6535), .A2(n6534), .ZN(n9606) );
  OR2_X1 U8229 ( .A1(n6538), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8230 ( .A1(n6538), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6536) );
  AND2_X1 U8231 ( .A1(n6537), .A2(n6536), .ZN(n9605) );
  AND2_X1 U8232 ( .A1(n9606), .A2(n9605), .ZN(n9608) );
  AOI21_X1 U8233 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6538), .A(n9608), .ZN(
        n6539) );
  NAND2_X1 U8234 ( .A1(n6540), .A2(n6539), .ZN(n7125) );
  OAI21_X1 U8235 ( .B1(n6540), .B2(n6539), .A(n7125), .ZN(n6541) );
  NAND2_X1 U8236 ( .A1(n6541), .A2(n9660), .ZN(n6542) );
  NAND2_X1 U8237 ( .A1(n6543), .A2(n6542), .ZN(P1_U3255) );
  INV_X1 U8238 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6546) );
  INV_X1 U8239 ( .A(n6544), .ZN(n6547) );
  OAI222_X1 U8240 ( .A1(n8273), .A2(n6546), .B1(n8271), .B2(n6547), .C1(n6545), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8241 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6548) );
  INV_X1 U8242 ( .A(n7696), .ZN(n7764) );
  OAI222_X1 U8243 ( .A1(n8277), .A2(n6548), .B1(n8280), .B2(n6547), .C1(n7764), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8244 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6552) );
  INV_X1 U8245 ( .A(n6550), .ZN(n6551) );
  AOI22_X1 U8246 ( .A1(n6561), .A2(n6552), .B1(n6551), .B2(n6554), .ZN(
        P2_U3377) );
  INV_X1 U8247 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6556) );
  INV_X1 U8248 ( .A(n6553), .ZN(n6555) );
  AOI22_X1 U8249 ( .A1(n6561), .A2(n6556), .B1(n6555), .B2(n6554), .ZN(
        P2_U3376) );
  INV_X1 U8250 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10104) );
  INV_X1 U8251 ( .A(n6557), .ZN(n6559) );
  INV_X1 U8252 ( .A(n9624), .ZN(n6558) );
  OAI222_X1 U8253 ( .A1(n8273), .A2(n10104), .B1(n8275), .B2(n6559), .C1(
        P1_U3086), .C2(n6558), .ZN(P1_U3342) );
  INV_X1 U8254 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6560) );
  INV_X1 U8255 ( .A(n7812), .ZN(n7818) );
  OAI222_X1 U8256 ( .A1(n8277), .A2(n6560), .B1(n8280), .B2(n6559), .C1(
        P2_U3151), .C2(n7818), .ZN(P2_U3282) );
  AND2_X1 U8257 ( .A1(n6561), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8258 ( .A1(n6561), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8259 ( .A1(n6561), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8260 ( .A1(n6561), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8261 ( .A1(n6561), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8262 ( .A1(n6561), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8263 ( .A1(n6561), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8264 ( .A1(n6561), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8265 ( .A1(n6561), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8266 ( .A1(n6561), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8267 ( .A1(n6561), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8268 ( .A1(n6561), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8269 ( .A1(n6561), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8270 ( .A1(n6561), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8271 ( .A1(n6561), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8272 ( .A1(n6561), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8273 ( .A1(n6561), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8274 ( .A1(n6561), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8275 ( .A1(n6561), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8276 ( .A1(n6561), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8277 ( .A1(n6561), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8278 ( .A1(n6561), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8279 ( .A1(n6561), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8280 ( .A1(n6561), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8281 ( .A1(n6561), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8282 ( .A1(n6561), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8283 ( .A1(n6561), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  INV_X1 U8284 ( .A(n6561), .ZN(n6564) );
  INV_X1 U8285 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6562) );
  NOR2_X1 U8286 ( .A1(n6564), .A2(n6562), .ZN(P2_U3237) );
  INV_X1 U8287 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10089) );
  NOR2_X1 U8288 ( .A1(n6564), .A2(n10089), .ZN(P2_U3258) );
  INV_X1 U8289 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U8290 ( .A1(n6564), .A2(n6563), .ZN(P2_U3250) );
  NAND2_X1 U8291 ( .A1(n9130), .A2(n7965), .ZN(n6566) );
  NAND2_X1 U8292 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  XNOR2_X1 U8293 ( .A(n6567), .B(n8973), .ZN(n6723) );
  NAND2_X1 U8294 ( .A1(n9130), .A2(n7977), .ZN(n6569) );
  OR2_X1 U8295 ( .A1(n6964), .A2(n7984), .ZN(n6568) );
  NAND2_X1 U8296 ( .A1(n6569), .A2(n6568), .ZN(n6721) );
  XNOR2_X1 U8297 ( .A(n6723), .B(n6721), .ZN(n6728) );
  NAND2_X1 U8298 ( .A1(n6570), .A2(n8973), .ZN(n6571) );
  NAND2_X1 U8299 ( .A1(n9133), .A2(n7965), .ZN(n6573) );
  XNOR2_X1 U8300 ( .A(n6574), .B(n8973), .ZN(n6579) );
  NAND2_X1 U8301 ( .A1(n9133), .A2(n7977), .ZN(n6576) );
  OR2_X1 U8302 ( .A1(n9724), .A2(n7984), .ZN(n6575) );
  NAND2_X1 U8303 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  XNOR2_X1 U8304 ( .A(n6579), .B(n6577), .ZN(n6624) );
  INV_X1 U8305 ( .A(n6577), .ZN(n6578) );
  NAND2_X1 U8306 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  NAND2_X1 U8307 ( .A1(n9131), .A2(n8975), .ZN(n6581) );
  NAND2_X1 U8308 ( .A1(n9131), .A2(n7977), .ZN(n6584) );
  OR2_X1 U8309 ( .A1(n6582), .A2(n7984), .ZN(n6583) );
  NAND2_X1 U8310 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U8311 ( .A1(n6615), .A2(n6614), .ZN(n6726) );
  INV_X1 U8312 ( .A(n6585), .ZN(n6586) );
  NAND2_X1 U8313 ( .A1(n6587), .A2(n6586), .ZN(n6724) );
  NAND2_X1 U8314 ( .A1(n6726), .A2(n6724), .ZN(n6588) );
  XOR2_X1 U8315 ( .A(n6728), .B(n6588), .Z(n6613) );
  INV_X1 U8316 ( .A(n6589), .ZN(n6954) );
  OAI211_X1 U8317 ( .C1(n6592), .C2(n6591), .A(n6590), .B(n6954), .ZN(n6604)
         );
  INV_X1 U8318 ( .A(n6600), .ZN(n6593) );
  OR2_X1 U8319 ( .A1(n6604), .A2(n6593), .ZN(n6596) );
  OR2_X1 U8320 ( .A1(n9722), .A2(n6594), .ZN(n6595) );
  AOI22_X1 U8321 ( .A1(n9069), .A2(n9129), .B1(n9131), .B2(n9070), .ZN(n6866)
         );
  INV_X1 U8322 ( .A(n6866), .ZN(n6602) );
  NOR2_X2 U8323 ( .A1(n6596), .A2(n6479), .ZN(n9059) );
  INV_X1 U8324 ( .A(n6596), .ZN(n6598) );
  AND2_X1 U8325 ( .A1(n9720), .A2(n6597), .ZN(n9700) );
  NAND2_X1 U8326 ( .A1(n6598), .A2(n9700), .ZN(n6601) );
  INV_X1 U8327 ( .A(n6603), .ZN(n6599) );
  AOI22_X1 U8328 ( .A1(n6602), .A2(n9059), .B1(n6863), .B2(n9088), .ZN(n6612)
         );
  NAND2_X1 U8329 ( .A1(n6604), .A2(n6603), .ZN(n6608) );
  AND2_X1 U8330 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  NAND2_X1 U8331 ( .A1(n6608), .A2(n6607), .ZN(n6610) );
  AOI21_X2 U8332 ( .B1(n6610), .B2(P1_STATE_REG_SCAN_IN), .A(n6609), .ZN(n9061) );
  MUX2_X1 U8333 ( .A(P1_STATE_REG_SCAN_IN), .B(n9061), .S(n6961), .Z(n6611) );
  OAI211_X1 U8334 ( .C1(n6613), .C2(n9075), .A(n6612), .B(n6611), .ZN(P1_U3218) );
  XOR2_X1 U8335 ( .A(n6615), .B(n6614), .Z(n6620) );
  NAND2_X1 U8336 ( .A1(n9133), .A2(n9070), .ZN(n6617) );
  NAND2_X1 U8337 ( .A1(n9130), .A2(n9069), .ZN(n6616) );
  NAND2_X1 U8338 ( .A1(n6617), .A2(n6616), .ZN(n6884) );
  AOI22_X1 U8339 ( .A1(n9088), .A2(n7050), .B1(n6884), .B2(n9059), .ZN(n6619)
         );
  NAND2_X1 U8340 ( .A1(n9061), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8341 ( .A1(n6717), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6618) );
  OAI211_X1 U8342 ( .C1(n6620), .C2(n9075), .A(n6619), .B(n6618), .ZN(P1_U3237) );
  INV_X1 U8343 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6622) );
  INV_X1 U8344 ( .A(n6621), .ZN(n6623) );
  INV_X1 U8345 ( .A(n9633), .ZN(n7127) );
  OAI222_X1 U8346 ( .A1(n8273), .A2(n6622), .B1(n8275), .B2(n6623), .C1(
        P1_U3086), .C2(n7127), .ZN(P1_U3341) );
  INV_X1 U8347 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10058) );
  OAI222_X1 U8348 ( .A1(n8277), .A2(n10058), .B1(n8280), .B2(n6623), .C1(
        P2_U3151), .C2(n8454), .ZN(P2_U3281) );
  XOR2_X1 U8349 ( .A(n6625), .B(n6624), .Z(n6630) );
  NAND2_X1 U8350 ( .A1(n6204), .A2(n9070), .ZN(n6627) );
  NAND2_X1 U8351 ( .A1(n9131), .A2(n9069), .ZN(n6626) );
  NAND2_X1 U8352 ( .A1(n6627), .A2(n6626), .ZN(n7105) );
  AOI22_X1 U8353 ( .A1(n9088), .A2(n7117), .B1(n7105), .B2(n9059), .ZN(n6629)
         );
  NAND2_X1 U8354 ( .A1(n6717), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6628) );
  OAI211_X1 U8355 ( .C1(n6630), .C2(n9075), .A(n6629), .B(n6628), .ZN(P1_U3222) );
  INV_X1 U8356 ( .A(n6631), .ZN(n6639) );
  NOR2_X2 U8357 ( .A1(n8532), .A2(n8251), .ZN(n9788) );
  INV_X1 U8358 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7143) );
  MUX2_X1 U8359 ( .A(n7143), .B(n6632), .S(n8478), .Z(n9746) );
  AND2_X1 U8360 ( .A1(n9746), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9762) );
  INV_X1 U8361 ( .A(n6633), .ZN(n6634) );
  MUX2_X1 U8362 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8478), .Z(n6635) );
  INV_X1 U8363 ( .A(n6658), .ZN(n9784) );
  XNOR2_X1 U8364 ( .A(n6635), .B(n9784), .ZN(n9786) );
  AOI22_X1 U8365 ( .A1(n9785), .A2(n9786), .B1(n6635), .B2(n6658), .ZN(n6637)
         );
  MUX2_X1 U8366 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8478), .Z(n6666) );
  XOR2_X1 U8367 ( .A(n6673), .B(n6666), .Z(n6636) );
  NAND2_X1 U8368 ( .A1(n6637), .A2(n6636), .ZN(n6671) );
  OAI21_X1 U8369 ( .B1(n6637), .B2(n6636), .A(n6671), .ZN(n6653) );
  NAND2_X1 U8370 ( .A1(n8549), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7873) );
  NOR2_X1 U8371 ( .A1(n6654), .A2(n7873), .ZN(n6650) );
  NAND2_X1 U8372 ( .A1(n6650), .A2(n6133), .ZN(n6641) );
  OR2_X1 U8373 ( .A1(n6133), .A2(P2_U3151), .ZN(n8943) );
  INV_X1 U8374 ( .A(n8943), .ZN(n6638) );
  NAND2_X1 U8375 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  INV_X1 U8376 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6642) );
  INV_X1 U8377 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8378 ( .A1(n6655), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U8379 ( .A1(n9760), .A2(n6643), .ZN(n6644) );
  NAND2_X1 U8380 ( .A1(n6644), .A2(n6645), .ZN(n9753) );
  INV_X1 U8381 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9754) );
  OR2_X1 U8382 ( .A1(n9753), .A2(n9754), .ZN(n9751) );
  NAND2_X1 U8383 ( .A1(n9751), .A2(n6645), .ZN(n9774) );
  NAND2_X1 U8384 ( .A1(n6658), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8385 ( .A1(n9773), .A2(n6646), .ZN(n6647) );
  INV_X1 U8386 ( .A(n6682), .ZN(n6648) );
  AOI21_X1 U8387 ( .B1(n7301), .B2(n6649), .A(n6648), .ZN(n6651) );
  OAI22_X1 U8388 ( .A1(n8559), .A2(n6673), .B1(n6651), .B2(n9778), .ZN(n6652)
         );
  AOI21_X1 U8389 ( .B1(n9788), .B2(n6653), .A(n6652), .ZN(n6661) );
  NOR2_X1 U8390 ( .A1(n6654), .A2(n8943), .ZN(n9748) );
  NAND2_X1 U8391 ( .A1(n9748), .A2(n8478), .ZN(n9779) );
  INV_X1 U8392 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U8393 ( .A1(n6655), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6656) );
  AOI21_X1 U8394 ( .B1(n9755), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6657), .ZN(
        n9772) );
  INV_X1 U8395 ( .A(n6673), .ZN(n6667) );
  XNOR2_X1 U8396 ( .A(n6672), .B(n6667), .ZN(n6674) );
  XNOR2_X1 U8397 ( .A(n6674), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6659) );
  AND2_X1 U8398 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6818) );
  AOI21_X1 U8399 ( .B1(n8542), .B2(n6659), .A(n6818), .ZN(n6660) );
  OAI211_X1 U8400 ( .C1(n10055), .C2(n9768), .A(n6661), .B(n6660), .ZN(
        P2_U3185) );
  INV_X1 U8401 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6663) );
  INV_X1 U8402 ( .A(n6662), .ZN(n6664) );
  INV_X1 U8403 ( .A(n9655), .ZN(n7128) );
  OAI222_X1 U8404 ( .A1(n8273), .A2(n6663), .B1(n8275), .B2(n6664), .C1(
        P1_U3086), .C2(n7128), .ZN(P1_U3340) );
  INV_X1 U8405 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6665) );
  INV_X1 U8406 ( .A(n8477), .ZN(n8489) );
  OAI222_X1 U8407 ( .A1(n8277), .A2(n6665), .B1(n8280), .B2(n6664), .C1(
        P2_U3151), .C2(n8489), .ZN(P2_U3280) );
  INV_X1 U8408 ( .A(n6666), .ZN(n6668) );
  NAND2_X1 U8409 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  MUX2_X1 U8410 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8478), .Z(n6691) );
  XOR2_X1 U8411 ( .A(n6698), .B(n6691), .Z(n6669) );
  AOI21_X1 U8412 ( .B1(n6671), .B2(n6670), .A(n6669), .ZN(n6690) );
  NAND3_X1 U8413 ( .A1(n6671), .A2(n6670), .A3(n6669), .ZN(n6692) );
  NAND2_X1 U8414 ( .A1(n6692), .A2(n9788), .ZN(n6689) );
  INV_X1 U8415 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9885) );
  MUX2_X1 U8416 ( .A(n9885), .B(P2_REG1_REG_4__SCAN_IN), .S(n6698), .Z(n6676)
         );
  AOI22_X1 U8417 ( .A1(n6674), .A2(P2_REG1_REG_3__SCAN_IN), .B1(n6673), .B2(
        n6672), .ZN(n6675) );
  NOR2_X1 U8418 ( .A1(n6675), .A2(n6676), .ZN(n6695) );
  AOI21_X1 U8419 ( .B1(n6676), .B2(n6675), .A(n6695), .ZN(n6677) );
  OAI22_X1 U8420 ( .A1(n8559), .A2(n6698), .B1(n6677), .B2(n9779), .ZN(n6687)
         );
  INV_X1 U8421 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7168) );
  XNOR2_X1 U8422 ( .A(n6698), .B(n7168), .ZN(n6679) );
  NAND2_X1 U8423 ( .A1(n6678), .A2(n6679), .ZN(n6700) );
  INV_X1 U8424 ( .A(n6679), .ZN(n6681) );
  NAND3_X1 U8425 ( .A1(n6682), .A2(n6681), .A3(n6680), .ZN(n6683) );
  AOI21_X1 U8426 ( .B1(n6700), .B2(n6683), .A(n9778), .ZN(n6686) );
  INV_X1 U8427 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U8428 ( .A1(n9768), .A2(n6684), .ZN(n6685) );
  AND2_X1 U8429 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6948) );
  NOR4_X1 U8430 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6948), .ZN(n6688)
         );
  OAI21_X1 U8431 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(P2_U3186) );
  INV_X1 U8432 ( .A(n6698), .ZN(n6694) );
  INV_X1 U8433 ( .A(n6691), .ZN(n6693) );
  OAI21_X1 U8434 ( .B1(n6694), .B2(n6693), .A(n6692), .ZN(n6748) );
  MUX2_X1 U8435 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8478), .Z(n6746) );
  XNOR2_X1 U8436 ( .A(n6746), .B(n4486), .ZN(n6747) );
  XNOR2_X1 U8437 ( .A(n6748), .B(n6747), .ZN(n6708) );
  INV_X1 U8438 ( .A(n9768), .ZN(n8555) );
  AOI21_X1 U8439 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6698), .A(n6695), .ZN(
        n6756) );
  XNOR2_X1 U8440 ( .A(n6756), .B(n4486), .ZN(n6758) );
  XNOR2_X1 U8441 ( .A(n6758), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6697) );
  AND2_X1 U8442 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7148) );
  INV_X1 U8443 ( .A(n7148), .ZN(n6696) );
  OAI21_X1 U8444 ( .B1(n9779), .B2(n6697), .A(n6696), .ZN(n6706) );
  INV_X1 U8445 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8446 ( .A1(n6698), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6699) );
  INV_X1 U8447 ( .A(n8444), .ZN(n6702) );
  OAI22_X1 U8448 ( .A1(n8559), .A2(n6745), .B1(n6704), .B2(n9778), .ZN(n6705)
         );
  AOI211_X1 U8449 ( .C1(n8555), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6706), .B(
        n6705), .ZN(n6707) );
  OAI21_X1 U8450 ( .B1(n8534), .B2(n6708), .A(n6707), .ZN(P2_U3187) );
  NAND2_X1 U8451 ( .A1(n9132), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8452 ( .B1(n9083), .B2(n9132), .A(n6709), .ZN(P1_U3579) );
  INV_X1 U8453 ( .A(n6710), .ZN(n6713) );
  AOI22_X1 U8454 ( .A1(n7441), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7888), .ZN(n6711) );
  OAI21_X1 U8455 ( .B1(n6713), .B2(n8275), .A(n6711), .ZN(P1_U3339) );
  NAND2_X1 U8456 ( .A1(P2_U3893), .A2(n5766), .ZN(n6712) );
  OAI21_X1 U8457 ( .B1(P2_U3893), .B2(n4894), .A(n6712), .ZN(P2_U3491) );
  OAI222_X1 U8458 ( .A1(n8277), .A2(n6714), .B1(n8280), .B2(n6713), .C1(n8499), 
        .C2(P2_U3151), .ZN(P2_U3279) );
  NAND2_X1 U8459 ( .A1(n9132), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6715) );
  OAI21_X1 U8460 ( .B1(n8985), .B2(n9132), .A(n6715), .ZN(P1_U3583) );
  NAND2_X1 U8461 ( .A1(n9133), .A2(n9069), .ZN(n9712) );
  OAI22_X1 U8462 ( .A1(n9098), .A2(n9712), .B1(n9105), .B2(n7113), .ZN(n6716)
         );
  AOI21_X1 U8463 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6717), .A(n6716), .ZN(
        n6718) );
  OAI21_X1 U8464 ( .B1(n6719), .B2(n9075), .A(n6718), .ZN(P1_U3232) );
  INV_X1 U8465 ( .A(n6720), .ZN(n7321) );
  INV_X1 U8466 ( .A(n6721), .ZN(n6722) );
  NAND2_X1 U8467 ( .A1(n6723), .A2(n6722), .ZN(n6727) );
  AND2_X1 U8468 ( .A1(n6724), .A2(n6727), .ZN(n6725) );
  NAND2_X1 U8469 ( .A1(n6726), .A2(n6725), .ZN(n6731) );
  INV_X1 U8470 ( .A(n6727), .ZN(n6729) );
  NAND2_X1 U8471 ( .A1(n9129), .A2(n8975), .ZN(n6733) );
  OR2_X1 U8472 ( .A1(n7320), .A2(n7971), .ZN(n6732) );
  NAND2_X1 U8473 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  XNOR2_X1 U8474 ( .A(n6734), .B(n7975), .ZN(n6779) );
  NAND2_X1 U8475 ( .A1(n9129), .A2(n7977), .ZN(n6736) );
  OR2_X1 U8476 ( .A1(n7320), .A2(n7984), .ZN(n6735) );
  NAND2_X1 U8477 ( .A1(n6736), .A2(n6735), .ZN(n6778) );
  XNOR2_X1 U8478 ( .A(n6779), .B(n6778), .ZN(n6737) );
  AOI21_X1 U8479 ( .B1(n6738), .B2(n6737), .A(n9075), .ZN(n6739) );
  NAND2_X1 U8480 ( .A1(n6739), .A2(n6781), .ZN(n6743) );
  AOI22_X1 U8481 ( .A1(n9128), .A2(n9069), .B1(n9070), .B2(n9130), .ZN(n6854)
         );
  OAI21_X1 U8482 ( .B1(n6854), .B2(n9098), .A(n6740), .ZN(n6741) );
  AOI21_X1 U8483 ( .B1(n6937), .B2(n9088), .A(n6741), .ZN(n6742) );
  OAI211_X1 U8484 ( .C1(n9061), .C2(n7321), .A(n6743), .B(n6742), .ZN(P1_U3230) );
  NAND2_X1 U8485 ( .A1(n9132), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6744) );
  OAI21_X1 U8486 ( .B1(n9081), .B2(n9132), .A(n6744), .ZN(P1_U3581) );
  AOI22_X1 U8487 ( .A1(n6748), .A2(n6747), .B1(n6746), .B2(n6745), .ZN(n8434)
         );
  MUX2_X1 U8488 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8478), .Z(n6749) );
  NOR2_X1 U8489 ( .A1(n6749), .A2(n6764), .ZN(n6750) );
  AOI21_X1 U8490 ( .B1(n6749), .B2(n6764), .A(n6750), .ZN(n8433) );
  NAND2_X1 U8491 ( .A1(n8434), .A2(n8433), .ZN(n8432) );
  INV_X1 U8492 ( .A(n6750), .ZN(n6751) );
  NAND2_X1 U8493 ( .A1(n8432), .A2(n6751), .ZN(n6754) );
  MUX2_X1 U8494 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8478), .Z(n6752) );
  NOR2_X1 U8495 ( .A1(n6752), .A2(n7288), .ZN(n7280) );
  AOI21_X1 U8496 ( .B1(n6752), .B2(n7288), .A(n7280), .ZN(n6753) );
  AND2_X1 U8497 ( .A1(n6754), .A2(n6753), .ZN(n7279) );
  NOR2_X1 U8498 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  OAI21_X1 U8499 ( .B1(n7279), .B2(n6755), .A(n9788), .ZN(n6775) );
  INV_X1 U8500 ( .A(n6764), .ZN(n8440) );
  INV_X1 U8501 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6757) );
  OAI22_X1 U8502 ( .A1(n6758), .A2(n6757), .B1(n4486), .B2(n6756), .ZN(n8437)
         );
  MUX2_X1 U8503 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6759), .S(n6764), .Z(n8438)
         );
  NAND2_X1 U8504 ( .A1(n8437), .A2(n8438), .ZN(n8436) );
  OAI21_X1 U8505 ( .B1(n6760), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7289), .ZN(
        n6773) );
  INV_X1 U8506 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U8507 ( .A1(n9768), .A2(n6761), .ZN(n6772) );
  AND2_X1 U8508 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7375) );
  INV_X1 U8509 ( .A(n7375), .ZN(n6770) );
  INV_X1 U8510 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6762) );
  MUX2_X1 U8511 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6762), .S(n6764), .Z(n8441)
         );
  NAND2_X1 U8512 ( .A1(n6763), .A2(n8441), .ZN(n8446) );
  NAND2_X1 U8513 ( .A1(n6764), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8514 ( .A1(n8446), .A2(n6765), .ZN(n6766) );
  AOI21_X1 U8515 ( .B1(n6767), .B2(n7334), .A(n7273), .ZN(n6768) );
  OR2_X1 U8516 ( .A1(n9778), .A2(n6768), .ZN(n6769) );
  OAI211_X1 U8517 ( .C1(n8559), .C2(n7288), .A(n6770), .B(n6769), .ZN(n6771)
         );
  AOI211_X1 U8518 ( .C1(n8542), .C2(n6773), .A(n6772), .B(n6771), .ZN(n6774)
         );
  NAND2_X1 U8519 ( .A1(n6775), .A2(n6774), .ZN(P2_U3189) );
  OR2_X1 U8520 ( .A1(n6830), .A2(n8977), .ZN(n6777) );
  NAND2_X1 U8521 ( .A1(n6940), .A2(n8975), .ZN(n6776) );
  NAND2_X1 U8522 ( .A1(n6777), .A2(n6776), .ZN(n6801) );
  NAND2_X1 U8523 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  OAI22_X1 U8524 ( .A1(n6830), .A2(n7984), .B1(n7474), .B2(n7971), .ZN(n6782)
         );
  XNOR2_X1 U8525 ( .A(n6782), .B(n7975), .ZN(n6802) );
  XNOR2_X1 U8526 ( .A(n6809), .B(n6802), .ZN(n6783) );
  NOR2_X1 U8527 ( .A1(n6783), .A2(n6801), .ZN(n7067) );
  AOI21_X1 U8528 ( .B1(n6801), .B2(n6783), .A(n7067), .ZN(n6788) );
  INV_X1 U8529 ( .A(n9070), .ZN(n9082) );
  OAI22_X1 U8530 ( .A1(n6784), .A2(n9082), .B1(n6795), .B2(n9080), .ZN(n6842)
         );
  AOI22_X1 U8531 ( .A1(n6842), .A2(n9059), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6785) );
  OAI21_X1 U8532 ( .B1(n7474), .B2(n9105), .A(n6785), .ZN(n6786) );
  AOI21_X1 U8533 ( .B1(n7471), .B2(n9101), .A(n6786), .ZN(n6787) );
  OAI21_X1 U8534 ( .B1(n6788), .B2(n9075), .A(n6787), .ZN(P1_U3227) );
  NAND2_X1 U8535 ( .A1(n9126), .A2(n8975), .ZN(n6790) );
  OR2_X1 U8536 ( .A1(n7096), .A2(n7971), .ZN(n6789) );
  NAND2_X1 U8537 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  XNOR2_X1 U8538 ( .A(n6791), .B(n8973), .ZN(n7017) );
  NAND2_X1 U8539 ( .A1(n9126), .A2(n7977), .ZN(n6793) );
  OR2_X1 U8540 ( .A1(n7096), .A2(n7984), .ZN(n6792) );
  NAND2_X1 U8541 ( .A1(n6793), .A2(n6792), .ZN(n7015) );
  XNOR2_X1 U8542 ( .A(n7017), .B(n7015), .ZN(n6811) );
  OAI22_X1 U8543 ( .A1(n6795), .A2(n7984), .B1(n9693), .B2(n7971), .ZN(n6794)
         );
  XNOR2_X1 U8544 ( .A(n6794), .B(n7975), .ZN(n7066) );
  INV_X1 U8545 ( .A(n7066), .ZN(n6798) );
  OR2_X1 U8546 ( .A1(n6795), .A2(n8977), .ZN(n6797) );
  NAND2_X1 U8547 ( .A1(n6934), .A2(n8975), .ZN(n6796) );
  NAND2_X1 U8548 ( .A1(n6797), .A2(n6796), .ZN(n7065) );
  INV_X1 U8549 ( .A(n7065), .ZN(n6806) );
  NAND2_X1 U8550 ( .A1(n6798), .A2(n6806), .ZN(n7072) );
  INV_X1 U8551 ( .A(n6802), .ZN(n7069) );
  INV_X1 U8552 ( .A(n6801), .ZN(n6799) );
  NAND2_X1 U8553 ( .A1(n7069), .A2(n6799), .ZN(n6800) );
  AND2_X1 U8554 ( .A1(n7072), .A2(n6800), .ZN(n6808) );
  NAND2_X1 U8555 ( .A1(n6802), .A2(n6801), .ZN(n6805) );
  NAND2_X1 U8556 ( .A1(n6805), .A2(n6806), .ZN(n6803) );
  NAND2_X1 U8557 ( .A1(n6803), .A2(n7066), .ZN(n6804) );
  OAI21_X1 U8558 ( .B1(n6806), .B2(n6805), .A(n6804), .ZN(n6807) );
  OAI21_X1 U8559 ( .B1(n6811), .B2(n6810), .A(n7019), .ZN(n6812) );
  NAND2_X1 U8560 ( .A1(n6812), .A2(n9095), .ZN(n6816) );
  AOI22_X1 U8561 ( .A1(n9070), .A2(n9127), .B1(n9125), .B2(n9069), .ZN(n7090)
         );
  OAI22_X1 U8562 ( .A1(n7090), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6813), .ZN(n6814) );
  AOI21_X1 U8563 ( .B1(n9677), .B2(n9101), .A(n6814), .ZN(n6815) );
  OAI211_X1 U8564 ( .C1(n7096), .C2(n9105), .A(n6816), .B(n6815), .ZN(P1_U3213) );
  OAI22_X1 U8565 ( .A1(n10131), .A2(n9814), .B1(n7146), .B2(n10128), .ZN(n6817) );
  AOI211_X1 U8566 ( .C1(n6915), .C2(n10134), .A(n6818), .B(n6817), .ZN(n6824)
         );
  AOI21_X1 U8567 ( .B1(n6820), .B2(n6819), .A(n8383), .ZN(n6822) );
  NAND2_X1 U8568 ( .A1(n6822), .A2(n6821), .ZN(n6823) );
  OAI211_X1 U8569 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n10138), .A(n6824), .B(
        n6823), .ZN(P2_U3158) );
  OAI21_X1 U8570 ( .B1(n6826), .B2(n6828), .A(n6825), .ZN(n9696) );
  INV_X1 U8571 ( .A(n6839), .ZN(n6827) );
  AOI211_X1 U8572 ( .C1(n6934), .C2(n6827), .A(n9418), .B(n7083), .ZN(n9687)
         );
  XNOR2_X1 U8573 ( .A(n6829), .B(n6828), .ZN(n6832) );
  OAI22_X1 U8574 ( .A1(n6831), .A2(n9080), .B1(n6830), .B2(n9082), .ZN(n7076)
         );
  AOI21_X1 U8575 ( .B1(n6832), .B2(n9391), .A(n7076), .ZN(n9698) );
  INV_X1 U8576 ( .A(n9698), .ZN(n6833) );
  AOI211_X1 U8577 ( .C1(n9735), .C2(n9696), .A(n9687), .B(n6833), .ZN(n6936)
         );
  INV_X1 U8578 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6834) );
  OAI22_X1 U8579 ( .A1(n9586), .A2(n9693), .B1(n9738), .B2(n6834), .ZN(n6835)
         );
  INV_X1 U8580 ( .A(n6835), .ZN(n6836) );
  OAI21_X1 U8581 ( .B1(n6936), .B2(n7727), .A(n6836), .ZN(P1_U3471) );
  OAI21_X1 U8582 ( .B1(n6838), .B2(n6840), .A(n6837), .ZN(n7476) );
  AOI211_X1 U8583 ( .C1(n6940), .C2(n6850), .A(n9418), .B(n6839), .ZN(n7470)
         );
  XNOR2_X1 U8584 ( .A(n6841), .B(n6840), .ZN(n6844) );
  INV_X1 U8585 ( .A(n6842), .ZN(n6843) );
  OAI21_X1 U8586 ( .B1(n6844), .B2(n9715), .A(n6843), .ZN(n7469) );
  AOI211_X1 U8587 ( .C1(n9735), .C2(n7476), .A(n7470), .B(n7469), .ZN(n6942)
         );
  INV_X1 U8588 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6845) );
  OAI22_X1 U8589 ( .A1(n9586), .A2(n7474), .B1(n9738), .B2(n6845), .ZN(n6846)
         );
  INV_X1 U8590 ( .A(n6846), .ZN(n6847) );
  OAI21_X1 U8591 ( .B1(n6942), .B2(n7727), .A(n6847), .ZN(P1_U3468) );
  OAI21_X1 U8592 ( .B1(n6849), .B2(n6852), .A(n6848), .ZN(n7319) );
  INV_X1 U8593 ( .A(n6850), .ZN(n6851) );
  AOI211_X1 U8594 ( .C1(n6937), .C2(n6861), .A(n9418), .B(n6851), .ZN(n7325)
         );
  XNOR2_X1 U8595 ( .A(n6853), .B(n6852), .ZN(n6855) );
  OAI21_X1 U8596 ( .B1(n6855), .B2(n9715), .A(n6854), .ZN(n7326) );
  AOI211_X1 U8597 ( .C1(n9735), .C2(n7319), .A(n7325), .B(n7326), .ZN(n6939)
         );
  INV_X1 U8598 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6856) );
  OAI22_X1 U8599 ( .A1(n9586), .A2(n7320), .B1(n9738), .B2(n6856), .ZN(n6857)
         );
  INV_X1 U8600 ( .A(n6857), .ZN(n6858) );
  OAI21_X1 U8601 ( .B1(n6939), .B2(n7727), .A(n6858), .ZN(P1_U3465) );
  INV_X1 U8602 ( .A(n6860), .ZN(n6878) );
  INV_X1 U8603 ( .A(n6861), .ZN(n6862) );
  AOI211_X1 U8604 ( .C1(n6863), .C2(n6878), .A(n9418), .B(n6862), .ZN(n6960)
         );
  XNOR2_X1 U8605 ( .A(n6865), .B(n6864), .ZN(n6867) );
  OAI21_X1 U8606 ( .B1(n6867), .B2(n9715), .A(n6866), .ZN(n6958) );
  AOI211_X1 U8607 ( .C1(n9735), .C2(n6966), .A(n6960), .B(n6958), .ZN(n6893)
         );
  INV_X1 U8608 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6868) );
  OAI22_X1 U8609 ( .A1(n9586), .A2(n6964), .B1(n9738), .B2(n6868), .ZN(n6869)
         );
  INV_X1 U8610 ( .A(n6869), .ZN(n6870) );
  OAI21_X1 U8611 ( .B1(n6893), .B2(n7727), .A(n6870), .ZN(P1_U3462) );
  INV_X1 U8612 ( .A(n6871), .ZN(n6873) );
  INV_X1 U8613 ( .A(n8524), .ZN(n8538) );
  OAI222_X1 U8614 ( .A1(n8277), .A2(n6872), .B1(n8280), .B2(n6873), .C1(
        P2_U3151), .C2(n8538), .ZN(P2_U3278) );
  INV_X1 U8615 ( .A(n9218), .ZN(n9211) );
  OAI222_X1 U8616 ( .A1(n8273), .A2(n6874), .B1(n8275), .B2(n6873), .C1(
        P1_U3086), .C2(n9211), .ZN(P1_U3338) );
  OR2_X1 U8617 ( .A1(n6876), .A2(n6881), .ZN(n6877) );
  NAND2_X1 U8618 ( .A1(n6875), .A2(n6877), .ZN(n7056) );
  INV_X1 U8619 ( .A(n7112), .ZN(n6879) );
  OAI211_X1 U8620 ( .C1(n6582), .C2(n6879), .A(n6878), .B(n9242), .ZN(n7052)
         );
  INV_X1 U8621 ( .A(n7052), .ZN(n6888) );
  NAND3_X1 U8622 ( .A1(n7103), .A2(n6881), .A3(n6880), .ZN(n6882) );
  NAND2_X1 U8623 ( .A1(n6883), .A2(n6882), .ZN(n6885) );
  AOI21_X1 U8624 ( .B1(n6885), .B2(n9391), .A(n6884), .ZN(n6887) );
  NAND2_X1 U8625 ( .A1(n7056), .A2(n9446), .ZN(n6886) );
  NAND2_X1 U8626 ( .A1(n6887), .A2(n6886), .ZN(n7053) );
  AOI211_X1 U8627 ( .C1(n9726), .C2(n7056), .A(n6888), .B(n7053), .ZN(n6933)
         );
  INV_X1 U8628 ( .A(n9586), .ZN(n7725) );
  AOI22_X1 U8629 ( .A1(n7725), .A2(n7050), .B1(n7727), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n6889) );
  OAI21_X1 U8630 ( .B1(n6933), .B2(n7727), .A(n6889), .ZN(P1_U3459) );
  INV_X1 U8631 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6890) );
  OAI22_X1 U8632 ( .A1(n9530), .A2(n6964), .B1(n9745), .B2(n6890), .ZN(n6891)
         );
  INV_X1 U8633 ( .A(n6891), .ZN(n6892) );
  OAI21_X1 U8634 ( .B1(n6893), .B2(n9743), .A(n6892), .ZN(P1_U3525) );
  XOR2_X1 U8635 ( .A(n6895), .B(n6894), .Z(n6899) );
  NOR2_X1 U8636 ( .A1(n8400), .A2(P2_U3151), .ZN(n6931) );
  INV_X1 U8637 ( .A(n6931), .ZN(n6905) );
  AOI22_X1 U8638 ( .A1(n8408), .A2(n8431), .B1(n5761), .B2(n10134), .ZN(n6896)
         );
  OAI21_X1 U8639 ( .B1(n7159), .B2(n10131), .A(n6896), .ZN(n6897) );
  AOI21_X1 U8640 ( .B1(n6905), .B2(P2_REG3_REG_1__SCAN_IN), .A(n6897), .ZN(
        n6898) );
  OAI21_X1 U8641 ( .B1(n6899), .B2(n8383), .A(n6898), .ZN(P2_U3162) );
  XOR2_X1 U8642 ( .A(n6900), .B(n6901), .Z(n6907) );
  AOI22_X1 U8643 ( .A1(n8408), .A2(n8430), .B1(n6902), .B2(n10134), .ZN(n6903)
         );
  OAI21_X1 U8644 ( .B1(n6984), .B2(n10131), .A(n6903), .ZN(n6904) );
  AOI21_X1 U8645 ( .B1(n6905), .B2(P2_REG3_REG_2__SCAN_IN), .A(n6904), .ZN(
        n6906) );
  OAI21_X1 U8646 ( .B1(n8383), .B2(n6907), .A(n6906), .ZN(P2_U3177) );
  INV_X1 U8647 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8648 ( .A1(n6982), .A2(n8105), .ZN(n6910) );
  NAND2_X1 U8649 ( .A1(n6910), .A2(n6909), .ZN(n6911) );
  XOR2_X1 U8650 ( .A(n6908), .B(n6911), .Z(n6912) );
  AOI22_X1 U8651 ( .A1(n6912), .A2(n8726), .B1(n8728), .B2(n8431), .ZN(n7302)
         );
  NAND2_X1 U8652 ( .A1(n6913), .A2(n6908), .ZN(n7165) );
  OAI21_X1 U8653 ( .B1(n6913), .B2(n6908), .A(n7165), .ZN(n7298) );
  AOI22_X1 U8654 ( .A1(n7298), .A2(n9869), .B1(n9842), .B2(n8429), .ZN(n6914)
         );
  NAND2_X1 U8655 ( .A1(n7302), .A2(n6914), .ZN(n6921) );
  NAND2_X1 U8656 ( .A1(n6921), .A2(n9897), .ZN(n6917) );
  NAND2_X1 U8657 ( .A1(n8835), .A2(n6915), .ZN(n6916) );
  OAI211_X1 U8658 ( .C1(n9897), .C2(n6918), .A(n6917), .B(n6916), .ZN(P2_U3462) );
  INV_X1 U8659 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6919) );
  OAI22_X1 U8660 ( .A1(n7299), .A2(n8935), .B1(n9880), .B2(n6919), .ZN(n6920)
         );
  AOI21_X1 U8661 ( .B1(n9880), .B2(n6921), .A(n6920), .ZN(n6922) );
  INV_X1 U8662 ( .A(n6922), .ZN(P2_U3399) );
  INV_X1 U8663 ( .A(n8541), .ZN(n8560) );
  INV_X1 U8664 ( .A(n6923), .ZN(n6925) );
  OAI222_X1 U8665 ( .A1(P2_U3151), .A2(n8560), .B1(n8280), .B2(n6925), .C1(
        n6924), .C2(n8277), .ZN(P2_U3277) );
  INV_X1 U8666 ( .A(n9221), .ZN(n9670) );
  OAI222_X1 U8667 ( .A1(n8273), .A2(n6926), .B1(n8275), .B2(n6925), .C1(n9670), 
        .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U8668 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8669 ( .A1(n6927), .A2(n5766), .ZN(n8072) );
  NAND2_X1 U8670 ( .A1(n8070), .A2(n8072), .ZN(n8870) );
  OAI22_X1 U8671 ( .A1(n8403), .A2(n6927), .B1(n10128), .B2(n6984), .ZN(n6928)
         );
  AOI21_X1 U8672 ( .B1(n10126), .B2(n8870), .A(n6928), .ZN(n6929) );
  OAI21_X1 U8673 ( .B1(n6931), .B2(n6930), .A(n6929), .ZN(P2_U3172) );
  AOI22_X1 U8674 ( .A1(n7728), .A2(n7050), .B1(n9743), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6932) );
  OAI21_X1 U8675 ( .B1(n6933), .B2(n9743), .A(n6932), .ZN(P1_U3524) );
  AOI22_X1 U8676 ( .A1(n7728), .A2(n6934), .B1(n9743), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6935) );
  OAI21_X1 U8677 ( .B1(n6936), .B2(n9743), .A(n6935), .ZN(P1_U3528) );
  AOI22_X1 U8678 ( .A1(n7728), .A2(n6937), .B1(n9743), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U8679 ( .B1(n6939), .B2(n9743), .A(n6938), .ZN(P1_U3526) );
  AOI22_X1 U8680 ( .A1(n7728), .A2(n6940), .B1(n9743), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6941) );
  OAI21_X1 U8681 ( .B1(n6942), .B2(n9743), .A(n6941), .ZN(P1_U3527) );
  INV_X1 U8682 ( .A(n6943), .ZN(n6944) );
  AOI21_X1 U8683 ( .B1(n6946), .B2(n6945), .A(n6944), .ZN(n6952) );
  OAI22_X1 U8684 ( .A1(n10131), .A2(n6983), .B1(n7242), .B2(n10128), .ZN(n6947) );
  AOI211_X1 U8685 ( .C1(n7170), .C2(n10134), .A(n6948), .B(n6947), .ZN(n6951)
         );
  INV_X1 U8686 ( .A(n6949), .ZN(n7169) );
  NAND2_X1 U8687 ( .A1(n8400), .A2(n7169), .ZN(n6950) );
  OAI211_X1 U8688 ( .C1(n6952), .C2(n8383), .A(n6951), .B(n6950), .ZN(P2_U3170) );
  NAND2_X1 U8689 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  INV_X1 U8690 ( .A(n6958), .ZN(n6968) );
  INV_X1 U8691 ( .A(n7049), .ZN(n6959) );
  OAI21_X2 U8692 ( .B1(n9446), .B2(n6959), .A(n9439), .ZN(n9426) );
  INV_X1 U8693 ( .A(n9426), .ZN(n9695) );
  NAND2_X2 U8694 ( .A1(n9439), .A2(n9700), .ZN(n9692) );
  NAND2_X1 U8695 ( .A1(n6960), .A2(n9686), .ZN(n6963) );
  INV_X2 U8696 ( .A(n9441), .ZN(n9703) );
  AOI22_X1 U8697 ( .A1(n9689), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9703), .B2(
        n6961), .ZN(n6962) );
  OAI211_X1 U8698 ( .C1(n6964), .C2(n9692), .A(n6963), .B(n6962), .ZN(n6965)
         );
  AOI21_X1 U8699 ( .B1(n9695), .B2(n6966), .A(n6965), .ZN(n6967) );
  OAI21_X1 U8700 ( .B1(n9709), .B2(n6968), .A(n6967), .ZN(P1_U3290) );
  OAI21_X1 U8701 ( .B1(n6970), .B2(n6981), .A(n6969), .ZN(n9821) );
  INV_X1 U8702 ( .A(n9821), .ZN(n6992) );
  INV_X1 U8703 ( .A(n6971), .ZN(n6977) );
  NOR2_X1 U8704 ( .A1(n6989), .A2(n8069), .ZN(n6978) );
  NAND2_X1 U8705 ( .A1(n9807), .A2(n6978), .ZN(n9801) );
  NOR2_X1 U8706 ( .A1(n6979), .A2(n9865), .ZN(n9820) );
  INV_X1 U8707 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U8708 ( .A1(n8773), .A2(n6980), .ZN(n6988) );
  XNOR2_X1 U8709 ( .A(n6982), .B(n6981), .ZN(n6987) );
  INV_X1 U8710 ( .A(n7615), .ZN(n9848) );
  OAI22_X1 U8711 ( .A1(n6984), .A2(n9794), .B1(n6983), .B2(n9813), .ZN(n6985)
         );
  AOI21_X1 U8712 ( .B1(n9821), .B2(n9848), .A(n6985), .ZN(n6986) );
  OAI21_X1 U8713 ( .B1(n9797), .B2(n6987), .A(n6986), .ZN(n9819) );
  AOI211_X1 U8714 ( .C1(n9820), .C2(n6989), .A(n6988), .B(n9819), .ZN(n6990)
         );
  MUX2_X1 U8715 ( .A(n6642), .B(n6990), .S(n9807), .Z(n6991) );
  OAI21_X1 U8716 ( .B1(n6992), .B2(n9801), .A(n6991), .ZN(P2_U3231) );
  OAI21_X1 U8717 ( .B1(n6994), .B2(n6999), .A(n6993), .ZN(n9448) );
  AOI21_X1 U8718 ( .B1(n7084), .B2(n9445), .A(n9418), .ZN(n6995) );
  AND2_X1 U8719 ( .A1(n6995), .A2(n7032), .ZN(n9451) );
  NAND2_X1 U8720 ( .A1(n6997), .A2(n6996), .ZN(n7088) );
  NOR2_X1 U8721 ( .A1(n7088), .A2(n7089), .ZN(n7087) );
  NOR2_X1 U8722 ( .A1(n7087), .A2(n6998), .ZN(n7038) );
  INV_X1 U8723 ( .A(n7087), .ZN(n7002) );
  INV_X1 U8724 ( .A(n6999), .ZN(n7000) );
  AOI21_X1 U8725 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7003) );
  AOI211_X1 U8726 ( .C1(n7038), .C2(n7004), .A(n9715), .B(n7003), .ZN(n7007)
         );
  OR2_X1 U8727 ( .A1(n7192), .A2(n9080), .ZN(n7006) );
  NAND2_X1 U8728 ( .A1(n9126), .A2(n9070), .ZN(n7005) );
  NAND2_X1 U8729 ( .A1(n7006), .A2(n7005), .ZN(n7025) );
  OR2_X1 U8730 ( .A1(n7007), .A2(n7025), .ZN(n9440) );
  AOI211_X1 U8731 ( .C1(n9735), .C2(n9448), .A(n9451), .B(n9440), .ZN(n7014)
         );
  INV_X1 U8732 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7008) );
  OAI22_X1 U8733 ( .A1(n7011), .A2(n9586), .B1(n9738), .B2(n7008), .ZN(n7009)
         );
  INV_X1 U8734 ( .A(n7009), .ZN(n7010) );
  OAI21_X1 U8735 ( .B1(n7014), .B2(n7727), .A(n7010), .ZN(P1_U3477) );
  OAI22_X1 U8736 ( .A1(n7011), .A2(n9530), .B1(n9745), .B2(n6426), .ZN(n7012)
         );
  INV_X1 U8737 ( .A(n7012), .ZN(n7013) );
  OAI21_X1 U8738 ( .B1(n7014), .B2(n9743), .A(n7013), .ZN(P1_U3530) );
  INV_X1 U8739 ( .A(n7015), .ZN(n7016) );
  NAND2_X1 U8740 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  NAND2_X1 U8741 ( .A1(n9445), .A2(n8970), .ZN(n7020) );
  OAI21_X1 U8742 ( .B1(n7041), .B2(n7984), .A(n7020), .ZN(n7021) );
  XNOR2_X1 U8743 ( .A(n7187), .B(n7247), .ZN(n7024) );
  OR2_X1 U8744 ( .A1(n7041), .A2(n8977), .ZN(n7023) );
  NAND2_X1 U8745 ( .A1(n9445), .A2(n8975), .ZN(n7022) );
  NAND2_X1 U8746 ( .A1(n7023), .A2(n7022), .ZN(n7180) );
  NOR2_X1 U8747 ( .A1(n7024), .A2(n7180), .ZN(n7246) );
  AOI21_X1 U8748 ( .B1(n7024), .B2(n7180), .A(n7246), .ZN(n7029) );
  AOI22_X1 U8749 ( .A1(n7025), .A2(n9059), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7026) );
  OAI21_X1 U8750 ( .B1(n9061), .B2(n9442), .A(n7026), .ZN(n7027) );
  AOI21_X1 U8751 ( .B1(n9445), .B2(n9088), .A(n7027), .ZN(n7028) );
  OAI21_X1 U8752 ( .B1(n7029), .B2(n9075), .A(n7028), .ZN(P1_U3221) );
  OAI21_X1 U8753 ( .B1(n7031), .B2(n7039), .A(n7030), .ZN(n9433) );
  NAND2_X1 U8754 ( .A1(n7032), .A2(n9432), .ZN(n7033) );
  NAND2_X1 U8755 ( .A1(n7033), .A2(n9242), .ZN(n7034) );
  OR2_X1 U8756 ( .A1(n7034), .A2(n7207), .ZN(n7036) );
  NOR2_X1 U8757 ( .A1(n9123), .A2(n9080), .ZN(n7253) );
  INV_X1 U8758 ( .A(n7253), .ZN(n7035) );
  NAND2_X1 U8759 ( .A1(n7036), .A2(n7035), .ZN(n9434) );
  NOR2_X1 U8760 ( .A1(n7038), .A2(n7037), .ZN(n7040) );
  XNOR2_X1 U8761 ( .A(n7040), .B(n7039), .ZN(n7043) );
  NOR2_X1 U8762 ( .A1(n7041), .A2(n9082), .ZN(n7254) );
  INV_X1 U8763 ( .A(n7254), .ZN(n7042) );
  OAI21_X1 U8764 ( .B1(n7043), .B2(n9715), .A(n7042), .ZN(n9428) );
  AOI211_X1 U8765 ( .C1(n9735), .C2(n9433), .A(n9434), .B(n9428), .ZN(n7048)
         );
  AOI22_X1 U8766 ( .A1(n7728), .A2(n9432), .B1(n9743), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7044) );
  OAI21_X1 U8767 ( .B1(n7048), .B2(n9743), .A(n7044), .ZN(P1_U3531) );
  INV_X1 U8768 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7045) );
  NOR2_X1 U8769 ( .A1(n9738), .A2(n7045), .ZN(n7046) );
  AOI21_X1 U8770 ( .B1(n7725), .B2(n9432), .A(n7046), .ZN(n7047) );
  OAI21_X1 U8771 ( .B1(n7048), .B2(n7727), .A(n7047), .ZN(P1_U3480) );
  NOR2_X1 U8772 ( .A1(n9689), .A2(n7049), .ZN(n9681) );
  INV_X1 U8773 ( .A(n9692), .ZN(n9678) );
  AOI22_X1 U8774 ( .A1(n9678), .A2(n7050), .B1(n9703), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7051) );
  OAI21_X1 U8775 ( .B1(n7052), .B2(n9247), .A(n7051), .ZN(n7055) );
  MUX2_X1 U8776 ( .A(n7053), .B(P1_REG2_REG_2__SCAN_IN), .S(n9689), .Z(n7054)
         );
  AOI211_X1 U8777 ( .C1(n9681), .C2(n7056), .A(n7055), .B(n7054), .ZN(n7057)
         );
  INV_X1 U8778 ( .A(n7057), .ZN(P1_U3291) );
  NAND2_X1 U8779 ( .A1(n7058), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U8780 ( .A1(n7059), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8781 ( .A1(n6137), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7060) );
  NAND2_X1 U8782 ( .A1(n8532), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7064) );
  OAI21_X1 U8783 ( .B1(n8532), .B2(n8569), .A(n7064), .ZN(P2_U3522) );
  NAND2_X1 U8784 ( .A1(n7066), .A2(n7065), .ZN(n7070) );
  INV_X1 U8785 ( .A(n7070), .ZN(n7075) );
  INV_X1 U8786 ( .A(n6809), .ZN(n7068) );
  AOI21_X1 U8787 ( .B1(n7069), .B2(n7068), .A(n7067), .ZN(n7074) );
  AOI21_X1 U8788 ( .B1(n7072), .B2(n7070), .A(n7074), .ZN(n7071) );
  AOI21_X1 U8789 ( .B1(n7074), .B2(n7072), .A(n7071), .ZN(n7073) );
  AOI21_X1 U8790 ( .B1(n7075), .B2(n7074), .A(n7073), .ZN(n7080) );
  AOI22_X1 U8791 ( .A1(n7076), .A2(n9059), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7077) );
  OAI21_X1 U8792 ( .B1(n9693), .B2(n9105), .A(n7077), .ZN(n7078) );
  AOI21_X1 U8793 ( .B1(n9688), .B2(n9101), .A(n7078), .ZN(n7079) );
  OAI21_X1 U8794 ( .B1(n7080), .B2(n9075), .A(n7079), .ZN(P1_U3239) );
  OAI21_X1 U8795 ( .B1(n7082), .B2(n7089), .A(n7081), .ZN(n9682) );
  INV_X1 U8796 ( .A(n7083), .ZN(n7086) );
  INV_X1 U8797 ( .A(n7084), .ZN(n7085) );
  AOI211_X1 U8798 ( .C1(n9679), .C2(n7086), .A(n9418), .B(n7085), .ZN(n9680)
         );
  AOI21_X1 U8799 ( .B1(n7089), .B2(n7088), .A(n7087), .ZN(n7091) );
  OAI21_X1 U8800 ( .B1(n7091), .B2(n9715), .A(n7090), .ZN(n7092) );
  AOI21_X1 U8801 ( .B1(n9446), .B2(n9682), .A(n7092), .ZN(n9685) );
  INV_X1 U8802 ( .A(n9685), .ZN(n7093) );
  AOI211_X1 U8803 ( .C1(n9726), .C2(n9682), .A(n9680), .B(n7093), .ZN(n7099)
         );
  AOI22_X1 U8804 ( .A1(n7728), .A2(n9679), .B1(n9743), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7094) );
  OAI21_X1 U8805 ( .B1(n7099), .B2(n9743), .A(n7094), .ZN(P1_U3529) );
  INV_X1 U8806 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7095) );
  OAI22_X1 U8807 ( .A1(n9586), .A2(n7096), .B1(n9738), .B2(n7095), .ZN(n7097)
         );
  INV_X1 U8808 ( .A(n7097), .ZN(n7098) );
  OAI21_X1 U8809 ( .B1(n7099), .B2(n7727), .A(n7098), .ZN(P1_U3474) );
  INV_X1 U8810 ( .A(n7100), .ZN(n7102) );
  NAND2_X1 U8811 ( .A1(n7102), .A2(n7109), .ZN(n7104) );
  NAND2_X1 U8812 ( .A1(n7104), .A2(n7103), .ZN(n7106) );
  AOI21_X1 U8813 ( .B1(n7106), .B2(n9391), .A(n7105), .ZN(n7111) );
  OAI21_X1 U8814 ( .B1(n7109), .B2(n7108), .A(n7107), .ZN(n9727) );
  NAND2_X1 U8815 ( .A1(n9727), .A2(n9446), .ZN(n7110) );
  AND2_X1 U8816 ( .A1(n7111), .A2(n7110), .ZN(n9729) );
  OAI211_X1 U8817 ( .C1(n7113), .C2(n9724), .A(n9242), .B(n7112), .ZN(n9723)
         );
  INV_X1 U8818 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7114) );
  OAI22_X1 U8819 ( .A1(n9439), .A2(n7115), .B1(n7114), .B2(n9441), .ZN(n7116)
         );
  AOI21_X1 U8820 ( .B1(n9678), .B2(n7117), .A(n7116), .ZN(n7118) );
  OAI21_X1 U8821 ( .B1(n9723), .B2(n9247), .A(n7118), .ZN(n7119) );
  AOI21_X1 U8822 ( .B1(n9727), .B2(n9681), .A(n7119), .ZN(n7120) );
  OAI21_X1 U8823 ( .B1(n9729), .B2(n9709), .A(n7120), .ZN(P1_U3292) );
  XNOR2_X1 U8824 ( .A(n9624), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9617) );
  OAI21_X1 U8825 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7126), .A(n7121), .ZN(
        n9618) );
  NOR2_X1 U8826 ( .A1(n9617), .A2(n9618), .ZN(n9616) );
  AOI21_X1 U8827 ( .B1(n9624), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9616), .ZN(
        n9628) );
  XNOR2_X1 U8828 ( .A(n9633), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9629) );
  NOR2_X1 U8829 ( .A1(n9628), .A2(n9629), .ZN(n9630) );
  AOI21_X1 U8830 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9633), .A(n9630), .ZN(
        n7122) );
  NOR2_X1 U8831 ( .A1(n7122), .A2(n7128), .ZN(n7123) );
  INV_X1 U8832 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9647) );
  XNOR2_X1 U8833 ( .A(n7128), .B(n7122), .ZN(n9648) );
  NOR2_X1 U8834 ( .A1(n9647), .A2(n9648), .ZN(n9646) );
  NOR2_X1 U8835 ( .A1(n7123), .A2(n9646), .ZN(n7437) );
  XNOR2_X1 U8836 ( .A(n7441), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7438) );
  XNOR2_X1 U8837 ( .A(n7437), .B(n7438), .ZN(n7138) );
  NAND2_X1 U8838 ( .A1(n9624), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7124) );
  OAI21_X1 U8839 ( .B1(n9624), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7124), .ZN(
        n9620) );
  OAI21_X1 U8840 ( .B1(n7126), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7125), .ZN(
        n9621) );
  NOR2_X1 U8841 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  AOI21_X1 U8842 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9624), .A(n9619), .ZN(
        n9635) );
  INV_X1 U8843 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U8844 ( .A1(n9633), .A2(n10082), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7127), .ZN(n9636) );
  NOR2_X1 U8845 ( .A1(n9635), .A2(n9636), .ZN(n9634) );
  AOI21_X1 U8846 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9633), .A(n9634), .ZN(
        n7129) );
  NOR2_X1 U8847 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  INV_X1 U8848 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9651) );
  XOR2_X1 U8849 ( .A(n9655), .B(n7129), .Z(n9652) );
  NOR2_X1 U8850 ( .A1(n9651), .A2(n9652), .ZN(n9650) );
  NOR2_X1 U8851 ( .A1(n7130), .A2(n9650), .ZN(n7132) );
  XNOR2_X1 U8852 ( .A(n7441), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n7131) );
  AOI21_X1 U8853 ( .B1(n7132), .B2(n7131), .A(n9649), .ZN(n7136) );
  OR2_X1 U8854 ( .A1(n7132), .A2(n7131), .ZN(n7443) );
  INV_X1 U8855 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U8856 ( .A1(n9656), .A2(n7441), .ZN(n7133) );
  NAND2_X1 U8857 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9018) );
  OAI211_X1 U8858 ( .C1(n9676), .C2(n7134), .A(n7133), .B(n9018), .ZN(n7135)
         );
  AOI21_X1 U8859 ( .B1(n7136), .B2(n7443), .A(n7135), .ZN(n7137) );
  OAI21_X1 U8860 ( .B1(n7138), .B2(n9645), .A(n7137), .ZN(P1_U3259) );
  NAND2_X1 U8861 ( .A1(n9807), .A2(n9842), .ZN(n8660) );
  INV_X1 U8862 ( .A(n8660), .ZN(n8737) );
  AOI22_X1 U8863 ( .A1(n8737), .A2(n6304), .B1(n8872), .B2(n9802), .ZN(n7145)
         );
  NOR2_X1 U8864 ( .A1(n7140), .A2(n9877), .ZN(n7141) );
  AOI22_X1 U8865 ( .A1(n9804), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n7141), .B2(
        n8870), .ZN(n7142) );
  MUX2_X1 U8866 ( .A(n7143), .B(n7142), .S(n9807), .Z(n7144) );
  NAND2_X1 U8867 ( .A1(n7145), .A2(n7144), .ZN(P2_U3233) );
  OAI22_X1 U8868 ( .A1(n10131), .A2(n7146), .B1(n7373), .B2(n10128), .ZN(n7147) );
  AOI211_X1 U8869 ( .C1(n9830), .C2(n10134), .A(n7148), .B(n7147), .ZN(n7153)
         );
  XNOR2_X1 U8870 ( .A(n7149), .B(n7150), .ZN(n7151) );
  NAND2_X1 U8871 ( .A1(n7151), .A2(n10126), .ZN(n7152) );
  OAI211_X1 U8872 ( .C1(n7343), .C2(n10138), .A(n7153), .B(n7152), .ZN(
        P2_U3167) );
  INV_X1 U8873 ( .A(n7154), .ZN(n8274) );
  OAI222_X1 U8874 ( .A1(n8277), .A2(n7155), .B1(n8937), .B2(n8274), .C1(
        P2_U3151), .C2(n8558), .ZN(P2_U3276) );
  NAND2_X1 U8875 ( .A1(n9807), .A2(n9848), .ZN(n7156) );
  XOR2_X1 U8876 ( .A(n8070), .B(n7157), .Z(n9811) );
  XOR2_X1 U8877 ( .A(n7158), .B(n7157), .Z(n7160) );
  OAI22_X1 U8878 ( .A1(n7160), .A2(n9797), .B1(n7159), .B2(n9794), .ZN(n9815)
         );
  NAND2_X1 U8879 ( .A1(n9807), .A2(n9815), .ZN(n7161) );
  OAI21_X1 U8880 ( .B1(n9807), .B2(n9754), .A(n7161), .ZN(n7163) );
  INV_X1 U8881 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9766) );
  OAI22_X1 U8882 ( .A1(n8721), .A2(n9812), .B1(n9766), .B2(n8773), .ZN(n7162)
         );
  AOI211_X1 U8883 ( .C1(n8737), .C2(n8431), .A(n7163), .B(n7162), .ZN(n7164)
         );
  OAI21_X1 U8884 ( .B1(n8740), .B2(n9811), .A(n7164), .ZN(P2_U3232) );
  NAND2_X1 U8885 ( .A1(n7165), .A2(n8117), .ZN(n7166) );
  XOR2_X1 U8886 ( .A(n8109), .B(n7166), .Z(n9823) );
  XNOR2_X1 U8887 ( .A(n4432), .B(n8109), .ZN(n7167) );
  AOI222_X1 U8888 ( .A1(n8726), .A2(n7167), .B1(n8430), .B2(n8728), .C1(n8428), 
        .C2(n9842), .ZN(n9824) );
  MUX2_X1 U8889 ( .A(n7168), .B(n9824), .S(n9807), .Z(n7172) );
  AOI22_X1 U8890 ( .A1(n9802), .A2(n7170), .B1(n9804), .B2(n7169), .ZN(n7171)
         );
  OAI211_X1 U8891 ( .C1(n8740), .C2(n9823), .A(n7172), .B(n7171), .ZN(P2_U3229) );
  NOR2_X1 U8892 ( .A1(n9123), .A2(n8977), .ZN(n7173) );
  AOI21_X1 U8893 ( .B1(n7264), .B2(n7965), .A(n7173), .ZN(n7217) );
  NAND2_X1 U8894 ( .A1(n9432), .A2(n8970), .ZN(n7175) );
  OR2_X1 U8895 ( .A1(n7192), .A2(n7984), .ZN(n7174) );
  NAND2_X1 U8896 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  XNOR2_X1 U8897 ( .A(n7176), .B(n7975), .ZN(n7249) );
  NAND2_X1 U8898 ( .A1(n9432), .A2(n8975), .ZN(n7178) );
  OR2_X1 U8899 ( .A1(n7192), .A2(n8977), .ZN(n7177) );
  NAND2_X1 U8900 ( .A1(n7178), .A2(n7177), .ZN(n7182) );
  NAND2_X1 U8901 ( .A1(n7247), .A2(n4446), .ZN(n7179) );
  OAI21_X1 U8902 ( .B1(n7249), .B2(n7182), .A(n7179), .ZN(n7186) );
  INV_X1 U8903 ( .A(n7182), .ZN(n7248) );
  NAND2_X1 U8904 ( .A1(n7181), .A2(n7248), .ZN(n7184) );
  INV_X1 U8905 ( .A(n7181), .ZN(n7183) );
  AOI22_X1 U8906 ( .A1(n7249), .A2(n7184), .B1(n7183), .B2(n7182), .ZN(n7185)
         );
  NAND2_X1 U8907 ( .A1(n7264), .A2(n8970), .ZN(n7189) );
  OR2_X1 U8908 ( .A1(n9123), .A2(n7984), .ZN(n7188) );
  NAND2_X1 U8909 ( .A1(n7189), .A2(n7188), .ZN(n7190) );
  XNOR2_X1 U8910 ( .A(n7190), .B(n8973), .ZN(n7221) );
  XNOR2_X1 U8911 ( .A(n7225), .B(n7221), .ZN(n7191) );
  NAND2_X1 U8912 ( .A1(n7191), .A2(n7217), .ZN(n7306) );
  OAI21_X1 U8913 ( .B1(n7217), .B2(n7191), .A(n7306), .ZN(n7198) );
  OR2_X1 U8914 ( .A1(n7192), .A2(n9082), .ZN(n7194) );
  NAND2_X1 U8915 ( .A1(n9122), .A2(n9069), .ZN(n7193) );
  NAND2_X1 U8916 ( .A1(n7194), .A2(n7193), .ZN(n7201) );
  AOI22_X1 U8917 ( .A1(n7201), .A2(n9059), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7196) );
  NAND2_X1 U8918 ( .A1(n9101), .A2(n7208), .ZN(n7195) );
  OAI211_X1 U8919 ( .C1(n7267), .C2(n9105), .A(n7196), .B(n7195), .ZN(n7197)
         );
  AOI21_X1 U8920 ( .B1(n7198), .B2(n9095), .A(n7197), .ZN(n7199) );
  INV_X1 U8921 ( .A(n7199), .ZN(P1_U3217) );
  OAI21_X1 U8922 ( .B1(n4435), .B2(n7200), .A(n7455), .ZN(n7202) );
  AOI21_X1 U8923 ( .B1(n7202), .B2(n9391), .A(n7201), .ZN(n7260) );
  INV_X1 U8924 ( .A(n7204), .ZN(n7205) );
  OAI21_X1 U8925 ( .B1(n7203), .B2(n7206), .A(n7205), .ZN(n7263) );
  NAND2_X1 U8926 ( .A1(n7263), .A2(n9695), .ZN(n7212) );
  AOI211_X1 U8927 ( .C1(n7264), .C2(n4701), .A(n9418), .B(n7452), .ZN(n7262)
         );
  AOI22_X1 U8928 ( .A1(n9689), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7208), .B2(
        n9703), .ZN(n7209) );
  OAI21_X1 U8929 ( .B1(n7267), .B2(n9692), .A(n7209), .ZN(n7210) );
  AOI21_X1 U8930 ( .B1(n7262), .B2(n9686), .A(n7210), .ZN(n7211) );
  OAI211_X1 U8931 ( .C1(n9709), .C2(n7260), .A(n7212), .B(n7211), .ZN(P1_U3283) );
  NAND2_X1 U8932 ( .A1(n7463), .A2(n8970), .ZN(n7214) );
  NAND2_X1 U8933 ( .A1(n9122), .A2(n8975), .ZN(n7213) );
  NAND2_X1 U8934 ( .A1(n7214), .A2(n7213), .ZN(n7215) );
  XNOR2_X1 U8935 ( .A(n7215), .B(n8973), .ZN(n7309) );
  NAND2_X1 U8936 ( .A1(n9122), .A2(n7977), .ZN(n7216) );
  OAI22_X1 U8937 ( .A1(n7309), .A2(n7308), .B1(n7217), .B2(n7221), .ZN(n7224)
         );
  INV_X1 U8938 ( .A(n7221), .ZN(n7307) );
  INV_X1 U8939 ( .A(n7217), .ZN(n7218) );
  OAI21_X1 U8940 ( .B1(n7307), .B2(n7218), .A(n7219), .ZN(n7222) );
  NOR2_X1 U8941 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  AOI22_X1 U8942 ( .A1(n7222), .A2(n7309), .B1(n7221), .B2(n7220), .ZN(n7223)
         );
  NAND2_X1 U8943 ( .A1(n7235), .A2(n8970), .ZN(n7227) );
  NAND2_X1 U8944 ( .A1(n9121), .A2(n8975), .ZN(n7226) );
  NAND2_X1 U8945 ( .A1(n7227), .A2(n7226), .ZN(n7228) );
  XNOR2_X1 U8946 ( .A(n7228), .B(n7975), .ZN(n7387) );
  AND2_X1 U8947 ( .A1(n9121), .A2(n7977), .ZN(n7229) );
  AOI21_X1 U8948 ( .B1(n7235), .B2(n7965), .A(n7229), .ZN(n7388) );
  XNOR2_X1 U8949 ( .A(n7387), .B(n7388), .ZN(n7385) );
  XOR2_X1 U8950 ( .A(n7386), .B(n7385), .Z(n7237) );
  OR2_X1 U8951 ( .A1(n7545), .A2(n9080), .ZN(n7231) );
  NAND2_X1 U8952 ( .A1(n9122), .A2(n9070), .ZN(n7230) );
  AND2_X1 U8953 ( .A1(n7231), .A2(n7230), .ZN(n7496) );
  NAND2_X1 U8954 ( .A1(n9101), .A2(n7499), .ZN(n7233) );
  OAI211_X1 U8955 ( .C1(n7496), .C2(n9098), .A(n7233), .B(n7232), .ZN(n7234)
         );
  AOI21_X1 U8956 ( .B1(n7235), .B2(n9088), .A(n7234), .ZN(n7236) );
  OAI21_X1 U8957 ( .B1(n7237), .B2(n9075), .A(n7236), .ZN(P1_U3224) );
  AOI21_X1 U8958 ( .B1(n7238), .B2(n7239), .A(n8383), .ZN(n7240) );
  OR2_X1 U8959 ( .A1(n7238), .A2(n7239), .ZN(n7369) );
  NAND2_X1 U8960 ( .A1(n7240), .A2(n7369), .ZN(n7245) );
  INV_X1 U8961 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7241) );
  NOR2_X1 U8962 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7241), .ZN(n8448) );
  OAI22_X1 U8963 ( .A1(n10131), .A2(n7242), .B1(n7564), .B2(n10128), .ZN(n7243) );
  AOI211_X1 U8964 ( .C1(n9836), .C2(n10134), .A(n8448), .B(n7243), .ZN(n7244)
         );
  OAI211_X1 U8965 ( .C1(n7358), .C2(n10138), .A(n7245), .B(n7244), .ZN(
        P2_U3179) );
  AOI21_X1 U8966 ( .B1(n7247), .B2(n7187), .A(n7246), .ZN(n7251) );
  XNOR2_X1 U8967 ( .A(n7249), .B(n7248), .ZN(n7250) );
  XNOR2_X1 U8968 ( .A(n7251), .B(n7250), .ZN(n7259) );
  INV_X1 U8969 ( .A(n7252), .ZN(n9429) );
  OAI21_X1 U8970 ( .B1(n7254), .B2(n7253), .A(n9059), .ZN(n7256) );
  OAI211_X1 U8971 ( .C1(n9061), .C2(n9429), .A(n7256), .B(n7255), .ZN(n7257)
         );
  AOI21_X1 U8972 ( .B1(n9432), .B2(n9088), .A(n7257), .ZN(n7258) );
  OAI21_X1 U8973 ( .B1(n7259), .B2(n9075), .A(n7258), .ZN(P1_U3231) );
  INV_X1 U8974 ( .A(n7260), .ZN(n7261) );
  AOI211_X1 U8975 ( .C1(n7263), .C2(n9735), .A(n7262), .B(n7261), .ZN(n7270)
         );
  AOI22_X1 U8976 ( .A1(n7264), .A2(n7728), .B1(n9743), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7265) );
  OAI21_X1 U8977 ( .B1(n7270), .B2(n9743), .A(n7265), .ZN(P1_U3532) );
  INV_X1 U8978 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7266) );
  OAI22_X1 U8979 ( .A1(n7267), .A2(n9586), .B1(n9738), .B2(n7266), .ZN(n7268)
         );
  INV_X1 U8980 ( .A(n7268), .ZN(n7269) );
  OAI21_X1 U8981 ( .B1(n7270), .B2(n7727), .A(n7269), .ZN(P1_U3483) );
  INV_X1 U8982 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7297) );
  INV_X1 U8983 ( .A(n9778), .ZN(n7286) );
  INV_X1 U8984 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7271) );
  MUX2_X1 U8985 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7271), .S(n7506), .Z(n7275)
         );
  INV_X1 U8986 ( .A(n7272), .ZN(n7274) );
  NAND2_X1 U8987 ( .A1(n7275), .A2(n4371), .ZN(n7505) );
  OAI21_X1 U8988 ( .B1(n7275), .B2(n4371), .A(n7505), .ZN(n7285) );
  NOR2_X1 U8989 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7276), .ZN(n7556) );
  MUX2_X1 U8990 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8478), .Z(n7277) );
  NOR2_X1 U8991 ( .A1(n7277), .A2(n7506), .ZN(n7513) );
  AOI21_X1 U8992 ( .B1(n7277), .B2(n7506), .A(n7513), .ZN(n7278) );
  INV_X1 U8993 ( .A(n7278), .ZN(n7282) );
  AOI21_X1 U8994 ( .B1(n7282), .B2(n7281), .A(n7512), .ZN(n7283) );
  NOR2_X1 U8995 ( .A1(n8534), .A2(n7283), .ZN(n7284) );
  AOI211_X1 U8996 ( .C1(n7286), .C2(n7285), .A(n7556), .B(n7284), .ZN(n7296)
         );
  INV_X1 U8997 ( .A(n7506), .ZN(n7509) );
  NAND2_X1 U8998 ( .A1(n7288), .A2(n7287), .ZN(n7290) );
  MUX2_X1 U8999 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7291), .S(n7506), .Z(n7292)
         );
  NAND2_X1 U9000 ( .A1(n7292), .A2(n7293), .ZN(n7508) );
  OAI21_X1 U9001 ( .B1(n7293), .B2(n7292), .A(n7508), .ZN(n7294) );
  AOI22_X1 U9002 ( .A1(n9783), .A2(n7509), .B1(n8542), .B2(n7294), .ZN(n7295)
         );
  OAI211_X1 U9003 ( .C1(n9768), .C2(n7297), .A(n7296), .B(n7295), .ZN(P2_U3190) );
  INV_X1 U9004 ( .A(n7298), .ZN(n7305) );
  OAI22_X1 U9005 ( .A1(n8721), .A2(n7299), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8773), .ZN(n7300) );
  AOI21_X1 U9006 ( .B1(n8737), .B2(n8429), .A(n7300), .ZN(n7304) );
  MUX2_X1 U9007 ( .A(n7302), .B(n7301), .S(n9808), .Z(n7303) );
  OAI211_X1 U9008 ( .C1(n8740), .C2(n7305), .A(n7304), .B(n7303), .ZN(P2_U3230) );
  OAI21_X1 U9009 ( .B1(n7307), .B2(n7225), .A(n7306), .ZN(n7311) );
  XNOR2_X1 U9010 ( .A(n7309), .B(n7308), .ZN(n7310) );
  XNOR2_X1 U9011 ( .A(n7311), .B(n7310), .ZN(n7318) );
  OR2_X1 U9012 ( .A1(n9123), .A2(n9082), .ZN(n7313) );
  NAND2_X1 U9013 ( .A1(n9121), .A2(n9069), .ZN(n7312) );
  AND2_X1 U9014 ( .A1(n7313), .A2(n7312), .ZN(n7461) );
  OAI22_X1 U9015 ( .A1(n7461), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7314), .ZN(n7316) );
  NOR2_X1 U9016 ( .A1(n4772), .A2(n9105), .ZN(n7315) );
  AOI211_X1 U9017 ( .C1(n7481), .C2(n9101), .A(n7316), .B(n7315), .ZN(n7317)
         );
  OAI21_X1 U9018 ( .B1(n7318), .B2(n9075), .A(n7317), .ZN(P1_U3236) );
  INV_X1 U9019 ( .A(n7319), .ZN(n7329) );
  NOR2_X1 U9020 ( .A1(n9692), .A2(n7320), .ZN(n7324) );
  OAI22_X1 U9021 ( .A1(n9439), .A2(n7322), .B1(n7321), .B2(n9441), .ZN(n7323)
         );
  AOI211_X1 U9022 ( .C1(n7325), .C2(n9450), .A(n7324), .B(n7323), .ZN(n7328)
         );
  NAND2_X1 U9023 ( .A1(n7326), .A2(n9439), .ZN(n7327) );
  OAI211_X1 U9024 ( .C1(n7329), .C2(n9426), .A(n7328), .B(n7327), .ZN(P1_U3289) );
  INV_X1 U9025 ( .A(n7330), .ZN(n7333) );
  INV_X1 U9026 ( .A(n7331), .ZN(n7332) );
  AOI21_X1 U9027 ( .B1(n7333), .B2(n8132), .A(n7332), .ZN(n9847) );
  INV_X1 U9028 ( .A(n9847), .ZN(n9844) );
  NOR2_X1 U9029 ( .A1(n9807), .A2(n7334), .ZN(n7337) );
  OAI22_X1 U9030 ( .A1(n8721), .A2(n7335), .B1(n7376), .B2(n8773), .ZN(n7336)
         );
  AOI211_X1 U9031 ( .C1(n8737), .C2(n10120), .A(n7337), .B(n7336), .ZN(n7341)
         );
  XNOR2_X1 U9032 ( .A(n7338), .B(n8076), .ZN(n7339) );
  OAI22_X1 U9033 ( .A1(n7339), .A2(n9797), .B1(n7373), .B2(n9794), .ZN(n9845)
         );
  NAND2_X1 U9034 ( .A1(n9845), .A2(n9807), .ZN(n7340) );
  OAI211_X1 U9035 ( .C1(n9844), .C2(n8740), .A(n7341), .B(n7340), .ZN(P2_U3226) );
  XNOR2_X1 U9036 ( .A(n8428), .B(n9830), .ZN(n8074) );
  XNOR2_X1 U9037 ( .A(n7342), .B(n8074), .ZN(n9829) );
  OAI22_X1 U9038 ( .A1(n8721), .A2(n7344), .B1(n7343), .B2(n8773), .ZN(n7351)
         );
  INV_X1 U9039 ( .A(n8074), .ZN(n7345) );
  XNOR2_X1 U9040 ( .A(n7346), .B(n7345), .ZN(n7347) );
  NAND2_X1 U9041 ( .A1(n7347), .A2(n8726), .ZN(n7349) );
  AOI22_X1 U9042 ( .A1(n8728), .A2(n8429), .B1(n8427), .B2(n9842), .ZN(n7348)
         );
  NAND2_X1 U9043 ( .A1(n7349), .A2(n7348), .ZN(n9833) );
  MUX2_X1 U9044 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9833), .S(n9807), .Z(n7350)
         );
  AOI211_X1 U9045 ( .C1(n8777), .C2(n9829), .A(n7351), .B(n7350), .ZN(n7352)
         );
  INV_X1 U9046 ( .A(n7352), .ZN(P2_U3228) );
  INV_X1 U9047 ( .A(n8125), .ZN(n7354) );
  NOR2_X1 U9048 ( .A1(n8115), .A2(n7354), .ZN(n8075) );
  XNOR2_X1 U9049 ( .A(n7353), .B(n8075), .ZN(n7357) );
  NAND2_X1 U9050 ( .A1(n8428), .A2(n8728), .ZN(n7355) );
  OAI21_X1 U9051 ( .B1(n7564), .B2(n9813), .A(n7355), .ZN(n7356) );
  AOI21_X1 U9052 ( .B1(n7357), .B2(n8726), .A(n7356), .ZN(n9839) );
  OAI22_X1 U9053 ( .A1(n8721), .A2(n7359), .B1(n7358), .B2(n8773), .ZN(n7360)
         );
  AOI21_X1 U9054 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9808), .A(n7360), .ZN(
        n7363) );
  XNOR2_X1 U9055 ( .A(n7361), .B(n8075), .ZN(n9835) );
  NAND2_X1 U9056 ( .A1(n9835), .A2(n8777), .ZN(n7362) );
  OAI211_X1 U9057 ( .C1(n9839), .C2(n9808), .A(n7363), .B(n7362), .ZN(P2_U3227) );
  INV_X1 U9058 ( .A(n7364), .ZN(n7434) );
  OAI222_X1 U9059 ( .A1(n8277), .A2(n7366), .B1(n8937), .B2(n7434), .C1(n7365), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  NAND2_X1 U9060 ( .A1(n7369), .A2(n7367), .ZN(n7371) );
  AND2_X1 U9061 ( .A1(n7369), .A2(n7368), .ZN(n7370) );
  AOI21_X1 U9062 ( .B1(n7372), .B2(n7371), .A(n7370), .ZN(n7380) );
  OAI22_X1 U9063 ( .A1(n10131), .A2(n7373), .B1(n10130), .B2(n10128), .ZN(
        n7374) );
  AOI211_X1 U9064 ( .C1(n9841), .C2(n10134), .A(n7375), .B(n7374), .ZN(n7379)
         );
  INV_X1 U9065 ( .A(n7376), .ZN(n7377) );
  NAND2_X1 U9066 ( .A1(n8400), .A2(n7377), .ZN(n7378) );
  OAI211_X1 U9067 ( .C1(n7380), .C2(n8383), .A(n7379), .B(n7378), .ZN(P2_U3153) );
  NAND2_X1 U9068 ( .A1(n7729), .A2(n8970), .ZN(n7382) );
  OR2_X1 U9069 ( .A1(n7545), .A2(n7984), .ZN(n7381) );
  NAND2_X1 U9070 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  XNOR2_X1 U9071 ( .A(n7383), .B(n7975), .ZN(n7524) );
  NOR2_X1 U9072 ( .A1(n7545), .A2(n8977), .ZN(n7384) );
  AOI21_X1 U9073 ( .B1(n7729), .B2(n7965), .A(n7384), .ZN(n7525) );
  XNOR2_X1 U9074 ( .A(n7524), .B(n7525), .ZN(n7529) );
  INV_X1 U9075 ( .A(n7387), .ZN(n7389) );
  NAND2_X1 U9076 ( .A1(n7389), .A2(n7388), .ZN(n7527) );
  NAND2_X1 U9077 ( .A1(n7532), .A2(n7527), .ZN(n7390) );
  XOR2_X1 U9078 ( .A(n7529), .B(n7390), .Z(n7397) );
  NAND2_X1 U9079 ( .A1(n9119), .A2(n9069), .ZN(n7392) );
  NAND2_X1 U9080 ( .A1(n9121), .A2(n9070), .ZN(n7391) );
  AND2_X1 U9081 ( .A1(n7392), .A2(n7391), .ZN(n7657) );
  OAI22_X1 U9082 ( .A1(n7657), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7393), .ZN(n7395) );
  INV_X1 U9083 ( .A(n7729), .ZN(n7663) );
  NOR2_X1 U9084 ( .A1(n7663), .A2(n9105), .ZN(n7394) );
  AOI211_X1 U9085 ( .C1(n7660), .C2(n9101), .A(n7395), .B(n7394), .ZN(n7396)
         );
  OAI21_X1 U9086 ( .B1(n7397), .B2(n9075), .A(n7396), .ZN(P1_U3234) );
  NOR2_X1 U9087 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7429) );
  NOR2_X1 U9088 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7426) );
  NOR2_X1 U9089 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7424) );
  NOR2_X1 U9090 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7422) );
  NOR2_X1 U9091 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7420) );
  INV_X1 U9092 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7699) );
  NOR2_X1 U9093 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7417) );
  NOR2_X1 U9094 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7415) );
  NOR2_X1 U9095 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7412) );
  NOR2_X1 U9096 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7410) );
  NOR2_X1 U9097 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7408) );
  NOR2_X1 U9098 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7406) );
  NOR2_X1 U9099 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7404) );
  NOR2_X1 U9100 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7402) );
  AOI22_X1 U9101 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n10055), .B2(n10052), .ZN(n10155) );
  NAND2_X1 U9102 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7399) );
  AOI21_X1 U9103 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9902) );
  INV_X1 U9104 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U9105 ( .A1(n10086), .A2(n9904), .ZN(n9903) );
  AOI21_X1 U9106 ( .B1(n9903), .B2(P1_ADDR_REG_1__SCAN_IN), .A(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n9898) );
  NOR2_X1 U9107 ( .A1(n9902), .A2(n9898), .ZN(n10153) );
  XOR2_X1 U9108 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10152) );
  NAND2_X1 U9109 ( .A1(n10153), .A2(n10152), .ZN(n7398) );
  NAND2_X1 U9110 ( .A1(n7399), .A2(n7398), .ZN(n10154) );
  NAND2_X1 U9111 ( .A1(n10155), .A2(n10154), .ZN(n7400) );
  OAI21_X1 U9112 ( .B1(n10055), .B2(n10052), .A(n7400), .ZN(n10157) );
  XNOR2_X1 U9113 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10156) );
  NOR2_X1 U9114 ( .A1(n10157), .A2(n10156), .ZN(n7401) );
  NOR2_X1 U9115 ( .A1(n7402), .A2(n7401), .ZN(n10145) );
  XNOR2_X1 U9116 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10144) );
  NOR2_X1 U9117 ( .A1(n10145), .A2(n10144), .ZN(n7403) );
  NOR2_X1 U9118 ( .A1(n7404), .A2(n7403), .ZN(n10143) );
  XNOR2_X1 U9119 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10142) );
  NOR2_X1 U9120 ( .A1(n10143), .A2(n10142), .ZN(n7405) );
  NOR2_X1 U9121 ( .A1(n7406), .A2(n7405), .ZN(n10149) );
  XNOR2_X1 U9122 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10148) );
  NOR2_X1 U9123 ( .A1(n10149), .A2(n10148), .ZN(n7407) );
  NOR2_X1 U9124 ( .A1(n7408), .A2(n7407), .ZN(n10151) );
  XNOR2_X1 U9125 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10150) );
  NOR2_X1 U9126 ( .A1(n10151), .A2(n10150), .ZN(n7409) );
  NOR2_X1 U9127 ( .A1(n7410), .A2(n7409), .ZN(n10147) );
  INV_X1 U9128 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7519) );
  AOI22_X1 U9129 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6435), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7519), .ZN(n10146) );
  NOR2_X1 U9130 ( .A1(n10147), .A2(n10146), .ZN(n7411) );
  NOR2_X1 U9131 ( .A1(n7412), .A2(n7411), .ZN(n9923) );
  INV_X1 U9132 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7602) );
  AOI22_X1 U9133 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7413), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7602), .ZN(n9922) );
  NOR2_X1 U9134 ( .A1(n9923), .A2(n9922), .ZN(n7414) );
  NOR2_X1 U9135 ( .A1(n7415), .A2(n7414), .ZN(n9921) );
  INV_X1 U9136 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9615) );
  INV_X1 U9137 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7744) );
  AOI22_X1 U9138 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9615), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7744), .ZN(n9920) );
  NOR2_X1 U9139 ( .A1(n9921), .A2(n9920), .ZN(n7416) );
  NOR2_X1 U9140 ( .A1(n7417), .A2(n7416), .ZN(n9919) );
  AOI22_X1 U9141 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n7699), .B1(
        P2_ADDR_REG_12__SCAN_IN), .B2(n10100), .ZN(n9918) );
  NOR2_X1 U9142 ( .A1(n9919), .A2(n9918), .ZN(n7418) );
  AOI21_X1 U9143 ( .B1(n10100), .B2(n7699), .A(n7418), .ZN(n9917) );
  INV_X1 U9144 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9627) );
  INV_X1 U9145 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7779) );
  AOI22_X1 U9146 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9627), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n7779), .ZN(n9916) );
  NOR2_X1 U9147 ( .A1(n9917), .A2(n9916), .ZN(n7419) );
  NOR2_X1 U9148 ( .A1(n7420), .A2(n7419), .ZN(n9915) );
  XNOR2_X1 U9149 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9914) );
  NOR2_X1 U9150 ( .A1(n9915), .A2(n9914), .ZN(n7421) );
  NOR2_X1 U9151 ( .A1(n7422), .A2(n7421), .ZN(n9913) );
  INV_X1 U9152 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9659) );
  INV_X1 U9153 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8460) );
  AOI22_X1 U9154 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9659), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8460), .ZN(n9912) );
  NOR2_X1 U9155 ( .A1(n9913), .A2(n9912), .ZN(n7423) );
  NOR2_X1 U9156 ( .A1(n7424), .A2(n7423), .ZN(n9911) );
  INV_X1 U9157 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8483) );
  AOI22_X1 U9158 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7134), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8483), .ZN(n9910) );
  NOR2_X1 U9159 ( .A1(n9911), .A2(n9910), .ZN(n7425) );
  NOR2_X1 U9160 ( .A1(n7426), .A2(n7425), .ZN(n9909) );
  INV_X1 U9161 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7427) );
  INV_X1 U9162 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U9163 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7427), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9991), .ZN(n9908) );
  NOR2_X1 U9164 ( .A1(n9909), .A2(n9908), .ZN(n7428) );
  NOR2_X1 U9165 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  AND2_X1 U9166 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7430), .ZN(n9905) );
  NOR2_X1 U9167 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9905), .ZN(n7431) );
  NOR2_X1 U9168 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7430), .ZN(n9906) );
  NOR2_X1 U9169 ( .A1(n7431), .A2(n9906), .ZN(n7433) );
  XNOR2_X1 U9170 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7432) );
  XNOR2_X1 U9171 ( .A(n7433), .B(n7432), .ZN(ADD_1068_U4) );
  OAI222_X1 U9172 ( .A1(n8273), .A2(n7436), .B1(P1_U3086), .B2(n7435), .C1(
        n8271), .C2(n7434), .ZN(P1_U3335) );
  XOR2_X1 U9173 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9218), .Z(n9213) );
  INV_X1 U9174 ( .A(n7437), .ZN(n7439) );
  OAI22_X1 U9175 ( .A1(n7439), .A2(n7438), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n7441), .ZN(n9214) );
  XOR2_X1 U9176 ( .A(n9213), .B(n9214), .Z(n7450) );
  INV_X1 U9177 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7440) );
  XNOR2_X1 U9178 ( .A(n9218), .B(n7440), .ZN(n7445) );
  NAND2_X1 U9179 ( .A1(n7441), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7442) );
  AND2_X1 U9180 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  NAND2_X1 U9181 ( .A1(n7444), .A2(n7445), .ZN(n9220) );
  OAI21_X1 U9182 ( .B1(n7445), .B2(n7444), .A(n9220), .ZN(n7448) );
  NAND2_X1 U9183 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U9184 ( .A1(n9597), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n7446) );
  OAI211_X1 U9185 ( .C1(n9671), .C2(n9211), .A(n9029), .B(n7446), .ZN(n7447)
         );
  AOI21_X1 U9186 ( .B1(n7448), .B2(n9660), .A(n7447), .ZN(n7449) );
  OAI21_X1 U9187 ( .B1(n9645), .B2(n7450), .A(n7449), .ZN(P1_U3260) );
  XNOR2_X1 U9188 ( .A(n7451), .B(n7456), .ZN(n7479) );
  INV_X1 U9189 ( .A(n7452), .ZN(n7454) );
  INV_X1 U9190 ( .A(n7453), .ZN(n7498) );
  AOI211_X1 U9191 ( .C1(n7463), .C2(n7454), .A(n9418), .B(n7498), .ZN(n7480)
         );
  INV_X1 U9192 ( .A(n7455), .ZN(n7458) );
  OAI21_X1 U9193 ( .B1(n7458), .B2(n7457), .A(n7456), .ZN(n7460) );
  NAND3_X1 U9194 ( .A1(n7460), .A2(n7459), .A3(n9391), .ZN(n7462) );
  NAND2_X1 U9195 ( .A1(n7462), .A2(n7461), .ZN(n7485) );
  AOI211_X1 U9196 ( .C1(n7479), .C2(n9735), .A(n7480), .B(n7485), .ZN(n7468)
         );
  AOI22_X1 U9197 ( .A1(n7463), .A2(n7728), .B1(n9743), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7464) );
  OAI21_X1 U9198 ( .B1(n7468), .B2(n9743), .A(n7464), .ZN(P1_U3533) );
  INV_X1 U9199 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7465) );
  OAI22_X1 U9200 ( .A1(n4772), .A2(n9586), .B1(n9738), .B2(n7465), .ZN(n7466)
         );
  INV_X1 U9201 ( .A(n7466), .ZN(n7467) );
  OAI21_X1 U9202 ( .B1(n7468), .B2(n7727), .A(n7467), .ZN(P1_U3486) );
  INV_X1 U9203 ( .A(n7469), .ZN(n7478) );
  NAND2_X1 U9204 ( .A1(n7470), .A2(n9450), .ZN(n7473) );
  AOI22_X1 U9205 ( .A1(n9709), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7471), .B2(
        n9703), .ZN(n7472) );
  OAI211_X1 U9206 ( .C1(n7474), .C2(n9692), .A(n7473), .B(n7472), .ZN(n7475)
         );
  AOI21_X1 U9207 ( .B1(n7476), .B2(n9695), .A(n7475), .ZN(n7477) );
  OAI21_X1 U9208 ( .B1(n7478), .B2(n9689), .A(n7477), .ZN(P1_U3288) );
  INV_X1 U9209 ( .A(n7479), .ZN(n7487) );
  NAND2_X1 U9210 ( .A1(n7480), .A2(n9450), .ZN(n7483) );
  AOI22_X1 U9211 ( .A1(n9709), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7481), .B2(
        n9703), .ZN(n7482) );
  OAI211_X1 U9212 ( .C1(n4772), .C2(n9692), .A(n7483), .B(n7482), .ZN(n7484)
         );
  AOI21_X1 U9213 ( .B1(n9439), .B2(n7485), .A(n7484), .ZN(n7486) );
  OAI21_X1 U9214 ( .B1(n7487), .B2(n9426), .A(n7486), .ZN(P1_U3282) );
  INV_X1 U9215 ( .A(n7488), .ZN(n7491) );
  OAI222_X1 U9216 ( .A1(P1_U3086), .A2(n7490), .B1(n8275), .B2(n7491), .C1(
        n7489), .C2(n8273), .ZN(P1_U3334) );
  OAI222_X1 U9217 ( .A1(n8277), .A2(n7492), .B1(n8937), .B2(n7491), .C1(n8069), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  XNOR2_X1 U9218 ( .A(n7493), .B(n7495), .ZN(n9736) );
  INV_X1 U9219 ( .A(n9736), .ZN(n7504) );
  OAI211_X1 U9220 ( .C1(n7495), .C2(n7494), .A(n7653), .B(n9391), .ZN(n7497)
         );
  NAND2_X1 U9221 ( .A1(n7497), .A2(n7496), .ZN(n9734) );
  OAI211_X1 U9222 ( .C1(n7498), .C2(n6221), .A(n9242), .B(n7659), .ZN(n9731)
         );
  NOR2_X1 U9223 ( .A1(n9731), .A2(n9247), .ZN(n7502) );
  AOI22_X1 U9224 ( .A1(n9709), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7499), .B2(
        n9703), .ZN(n7500) );
  OAI21_X1 U9225 ( .B1(n6221), .B2(n9692), .A(n7500), .ZN(n7501) );
  AOI211_X1 U9226 ( .C1(n9734), .C2(n9439), .A(n7502), .B(n7501), .ZN(n7503)
         );
  OAI21_X1 U9227 ( .B1(n7504), .B2(n9426), .A(n7503), .ZN(P1_U3281) );
  AOI21_X1 U9228 ( .B1(n5864), .B2(n7507), .A(n7578), .ZN(n7523) );
  OAI21_X1 U9229 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7510), .A(n7584), .ZN(
        n7521) );
  MUX2_X1 U9230 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8478), .Z(n7511) );
  NOR2_X1 U9231 ( .A1(n7511), .A2(n4690), .ZN(n7588) );
  AOI21_X1 U9232 ( .B1(n7511), .B2(n4690), .A(n7588), .ZN(n7515) );
  OAI21_X1 U9233 ( .B1(n7515), .B2(n7514), .A(n7596), .ZN(n7517) );
  AND2_X1 U9234 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U9235 ( .A1(n8559), .A2(n4690), .ZN(n7516) );
  AOI211_X1 U9236 ( .C1(n9788), .C2(n7517), .A(n10133), .B(n7516), .ZN(n7518)
         );
  OAI21_X1 U9237 ( .B1(n7519), .B2(n9768), .A(n7518), .ZN(n7520) );
  AOI21_X1 U9238 ( .B1(n8542), .B2(n7521), .A(n7520), .ZN(n7522) );
  OAI21_X1 U9239 ( .B1(n7523), .B2(n9778), .A(n7522), .ZN(P2_U3191) );
  INV_X1 U9240 ( .A(n7524), .ZN(n7526) );
  NAND2_X1 U9241 ( .A1(n7526), .A2(n7525), .ZN(n7528) );
  AND2_X1 U9242 ( .A1(n7527), .A2(n7528), .ZN(n7531) );
  INV_X1 U9243 ( .A(n7528), .ZN(n7530) );
  NAND2_X1 U9244 ( .A1(n9538), .A2(n8970), .ZN(n7534) );
  NAND2_X1 U9245 ( .A1(n9119), .A2(n8975), .ZN(n7533) );
  NAND2_X1 U9246 ( .A1(n7534), .A2(n7533), .ZN(n7535) );
  XNOR2_X1 U9247 ( .A(n7535), .B(n8973), .ZN(n7537) );
  NAND2_X1 U9248 ( .A1(n7538), .A2(n7537), .ZN(n7544) );
  OAI22_X1 U9249 ( .A1(n7719), .A2(n7984), .B1(n7536), .B2(n8977), .ZN(n7542)
         );
  OR2_X2 U9250 ( .A1(n7538), .A2(n7537), .ZN(n7540) );
  INV_X1 U9251 ( .A(n7539), .ZN(n7541) );
  NAND2_X1 U9252 ( .A1(n7541), .A2(n7540), .ZN(n7543) );
  AOI22_X1 U9253 ( .A1(n4613), .A2(n7544), .B1(n7543), .B2(n7542), .ZN(n7552)
         );
  INV_X1 U9254 ( .A(n7716), .ZN(n7549) );
  OR2_X1 U9255 ( .A1(n7545), .A2(n9082), .ZN(n7547) );
  NAND2_X1 U9256 ( .A1(n9118), .A2(n9069), .ZN(n7546) );
  NAND2_X1 U9257 ( .A1(n7547), .A2(n7546), .ZN(n7711) );
  AOI22_X1 U9258 ( .A1(n7711), .A2(n9059), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n7548) );
  OAI21_X1 U9259 ( .B1(n9061), .B2(n7549), .A(n7548), .ZN(n7550) );
  AOI21_X1 U9260 ( .B1(n9538), .B2(n9088), .A(n7550), .ZN(n7551) );
  OAI21_X1 U9261 ( .B1(n7552), .B2(n9075), .A(n7551), .ZN(P1_U3215) );
  XNOR2_X1 U9262 ( .A(n7553), .B(n10119), .ZN(n10121) );
  XNOR2_X1 U9263 ( .A(n10121), .B(n10120), .ZN(n7554) );
  NAND2_X1 U9264 ( .A1(n7554), .A2(n10126), .ZN(n7559) );
  OAI22_X1 U9265 ( .A1(n10131), .A2(n7564), .B1(n7611), .B2(n10128), .ZN(n7555) );
  AOI211_X1 U9266 ( .C1(n7557), .C2(n10134), .A(n7556), .B(n7555), .ZN(n7558)
         );
  OAI211_X1 U9267 ( .C1(n4413), .C2(n10138), .A(n7559), .B(n7558), .ZN(
        P2_U3161) );
  NAND2_X1 U9268 ( .A1(n7331), .A2(n7560), .ZN(n7561) );
  INV_X1 U9269 ( .A(n7562), .ZN(n8078) );
  XNOR2_X1 U9270 ( .A(n7561), .B(n8078), .ZN(n9853) );
  INV_X1 U9271 ( .A(n9853), .ZN(n7571) );
  OAI22_X1 U9272 ( .A1(n8721), .A2(n9851), .B1(n4413), .B2(n8773), .ZN(n7569)
         );
  AOI21_X1 U9273 ( .B1(n7563), .B2(n7562), .A(n9797), .ZN(n7567) );
  OAI22_X1 U9274 ( .A1(n7611), .A2(n9813), .B1(n7564), .B2(n9794), .ZN(n7565)
         );
  AOI21_X1 U9275 ( .B1(n7567), .B2(n7566), .A(n7565), .ZN(n9850) );
  NOR2_X1 U9276 ( .A1(n9850), .A2(n9808), .ZN(n7568) );
  AOI211_X1 U9277 ( .C1(n9808), .C2(P2_REG2_REG_8__SCAN_IN), .A(n7569), .B(
        n7568), .ZN(n7570) );
  OAI21_X1 U9278 ( .B1(n8740), .B2(n7571), .A(n7570), .ZN(P2_U3225) );
  INV_X1 U9279 ( .A(n7572), .ZN(n7575) );
  OAI222_X1 U9280 ( .A1(n8277), .A2(n9963), .B1(n8937), .B2(n7575), .C1(
        P2_U3151), .C2(n7573), .ZN(P2_U3273) );
  OAI222_X1 U9281 ( .A1(n8273), .A2(n7576), .B1(n8275), .B2(n7575), .C1(
        P1_U3086), .C2(n7574), .ZN(P1_U3333) );
  NOR2_X1 U9282 ( .A1(n7577), .A2(n4411), .ZN(n7579) );
  INV_X1 U9283 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7590) );
  MUX2_X1 U9284 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7590), .S(n7676), .Z(n7581)
         );
  INV_X1 U9285 ( .A(n7669), .ZN(n7580) );
  AOI21_X1 U9286 ( .B1(n7582), .B2(n7581), .A(n7580), .ZN(n7606) );
  NAND2_X1 U9287 ( .A1(n4690), .A2(n7583), .ZN(n7585) );
  MUX2_X1 U9288 ( .A(n7589), .B(P2_REG1_REG_10__SCAN_IN), .S(n7676), .Z(n7586)
         );
  NAND2_X1 U9289 ( .A1(n7587), .A2(n7586), .ZN(n7675) );
  OAI21_X1 U9290 ( .B1(n7587), .B2(n7586), .A(n7675), .ZN(n7604) );
  INV_X1 U9291 ( .A(n7588), .ZN(n7595) );
  MUX2_X1 U9292 ( .A(n7590), .B(n7589), .S(n8478), .Z(n7591) );
  NAND2_X1 U9293 ( .A1(n7591), .A2(n7676), .ZN(n7681) );
  INV_X1 U9294 ( .A(n7591), .ZN(n7592) );
  NAND2_X1 U9295 ( .A1(n7592), .A2(n7667), .ZN(n7593) );
  NAND2_X1 U9296 ( .A1(n7681), .A2(n7593), .ZN(n7594) );
  AOI21_X1 U9297 ( .B1(n7596), .B2(n7595), .A(n7594), .ZN(n7738) );
  INV_X1 U9298 ( .A(n7738), .ZN(n7598) );
  NAND3_X1 U9299 ( .A1(n7596), .A2(n7595), .A3(n7594), .ZN(n7597) );
  AOI21_X1 U9300 ( .B1(n7598), .B2(n7597), .A(n8534), .ZN(n7599) );
  AOI211_X1 U9301 ( .C1(n7676), .C2(n9783), .A(n7600), .B(n7599), .ZN(n7601)
         );
  OAI21_X1 U9302 ( .B1(n7602), .B2(n9768), .A(n7601), .ZN(n7603) );
  AOI21_X1 U9303 ( .B1(n8542), .B2(n7604), .A(n7603), .ZN(n7605) );
  OAI21_X1 U9304 ( .B1(n7606), .B2(n9778), .A(n7605), .ZN(P2_U3192) );
  NAND2_X1 U9305 ( .A1(n7608), .A2(n7607), .ZN(n8080) );
  XNOR2_X1 U9306 ( .A(n7609), .B(n8080), .ZN(n9860) );
  XNOR2_X1 U9307 ( .A(n7610), .B(n8080), .ZN(n7613) );
  OAI22_X1 U9308 ( .A1(n7611), .A2(n9794), .B1(n7796), .B2(n9813), .ZN(n7612)
         );
  AOI21_X1 U9309 ( .B1(n7613), .B2(n8726), .A(n7612), .ZN(n7614) );
  OAI21_X1 U9310 ( .B1(n7615), .B2(n9860), .A(n7614), .ZN(n9861) );
  NAND2_X1 U9311 ( .A1(n9861), .A2(n9807), .ZN(n7619) );
  OAI22_X1 U9312 ( .A1(n9807), .A2(n7590), .B1(n7616), .B2(n8773), .ZN(n7617)
         );
  AOI21_X1 U9313 ( .B1(n9802), .B2(n9863), .A(n7617), .ZN(n7618) );
  OAI211_X1 U9314 ( .C1(n9860), .C2(n9801), .A(n7619), .B(n7618), .ZN(P2_U3223) );
  NAND2_X1 U9315 ( .A1(n7624), .A2(n7620), .ZN(n7622) );
  OAI211_X1 U9316 ( .C1(n7623), .C2(n8273), .A(n7622), .B(n7621), .ZN(P1_U3332) );
  NAND2_X1 U9317 ( .A1(n7624), .A2(n8941), .ZN(n7626) );
  NAND2_X1 U9318 ( .A1(n7625), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8256) );
  OAI211_X1 U9319 ( .C1(n9927), .C2(n8277), .A(n7626), .B(n8256), .ZN(P2_U3272) );
  XNOR2_X1 U9320 ( .A(n7627), .B(n7749), .ZN(n9870) );
  INV_X1 U9321 ( .A(n9870), .ZN(n7636) );
  OAI211_X1 U9322 ( .C1(n7629), .C2(n8143), .A(n7628), .B(n8726), .ZN(n7631)
         );
  AOI22_X1 U9323 ( .A1(n8728), .A2(n8425), .B1(n8423), .B2(n9842), .ZN(n7630)
         );
  NAND2_X1 U9324 ( .A1(n7631), .A2(n7630), .ZN(n9867) );
  INV_X1 U9325 ( .A(n7632), .ZN(n9866) );
  NOR2_X1 U9326 ( .A1(n8721), .A2(n9866), .ZN(n7634) );
  OAI22_X1 U9327 ( .A1(n9807), .A2(n7683), .B1(n7760), .B2(n8773), .ZN(n7633)
         );
  AOI211_X1 U9328 ( .C1(n9867), .C2(n9807), .A(n7634), .B(n7633), .ZN(n7635)
         );
  OAI21_X1 U9329 ( .B1(n8740), .B2(n7636), .A(n7635), .ZN(P2_U3222) );
  XNOR2_X1 U9330 ( .A(n7637), .B(n7641), .ZN(n9535) );
  INV_X1 U9331 ( .A(n7714), .ZN(n7638) );
  AOI211_X1 U9332 ( .C1(n9532), .C2(n7638), .A(n9418), .B(n4708), .ZN(n9531)
         );
  AOI22_X1 U9333 ( .A1(n9709), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9102), .B2(
        n9703), .ZN(n7639) );
  OAI21_X1 U9334 ( .B1(n9106), .B2(n9692), .A(n7639), .ZN(n7649) );
  INV_X1 U9335 ( .A(n7640), .ZN(n7710) );
  OAI21_X1 U9336 ( .B1(n7710), .B2(n7642), .A(n7641), .ZN(n7644) );
  AOI21_X1 U9337 ( .B1(n7644), .B2(n7643), .A(n9715), .ZN(n7647) );
  OR2_X1 U9338 ( .A1(n7920), .A2(n9080), .ZN(n7646) );
  NAND2_X1 U9339 ( .A1(n9119), .A2(n9070), .ZN(n7645) );
  NAND2_X1 U9340 ( .A1(n7646), .A2(n7645), .ZN(n9097) );
  NOR2_X1 U9341 ( .A1(n7647), .A2(n9097), .ZN(n9534) );
  NOR2_X1 U9342 ( .A1(n9534), .A2(n9689), .ZN(n7648) );
  AOI211_X1 U9343 ( .C1(n9531), .C2(n9686), .A(n7649), .B(n7648), .ZN(n7650)
         );
  OAI21_X1 U9344 ( .B1(n9535), .B2(n9426), .A(n7650), .ZN(P1_U3278) );
  XOR2_X1 U9345 ( .A(n7656), .B(n7651), .Z(n7724) );
  INV_X1 U9346 ( .A(n7724), .ZN(n7666) );
  NAND2_X1 U9347 ( .A1(n7653), .A2(n7652), .ZN(n7655) );
  INV_X1 U9348 ( .A(n7708), .ZN(n7654) );
  AOI21_X1 U9349 ( .B1(n7656), .B2(n7655), .A(n7654), .ZN(n7658) );
  OAI21_X1 U9350 ( .B1(n7658), .B2(n9715), .A(n7657), .ZN(n7722) );
  AOI211_X1 U9351 ( .C1(n7729), .C2(n7659), .A(n9418), .B(n7713), .ZN(n7723)
         );
  NAND2_X1 U9352 ( .A1(n7723), .A2(n9450), .ZN(n7662) );
  AOI22_X1 U9353 ( .A1(n9709), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7660), .B2(
        n9703), .ZN(n7661) );
  OAI211_X1 U9354 ( .C1(n7663), .C2(n9692), .A(n7662), .B(n7661), .ZN(n7664)
         );
  AOI21_X1 U9355 ( .B1(n7722), .B2(n9439), .A(n7664), .ZN(n7665) );
  OAI21_X1 U9356 ( .B1(n7666), .B2(n9426), .A(n7665), .ZN(P1_U3280) );
  NAND2_X1 U9357 ( .A1(n7667), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7668) );
  NAND2_X1 U9358 ( .A1(n7764), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7761) );
  INV_X1 U9359 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9360 ( .A1(n7696), .A2(n7688), .ZN(n7671) );
  NAND2_X1 U9361 ( .A1(n7761), .A2(n7671), .ZN(n7673) );
  INV_X1 U9362 ( .A(n7762), .ZN(n7672) );
  AOI21_X1 U9363 ( .B1(n7674), .B2(n7673), .A(n7672), .ZN(n7703) );
  OAI21_X1 U9364 ( .B1(n7676), .B2(n7589), .A(n7675), .ZN(n7677) );
  NAND2_X1 U9365 ( .A1(n7685), .A2(n7677), .ZN(n7678) );
  XNOR2_X1 U9366 ( .A(n7677), .B(n7742), .ZN(n7735) );
  NAND2_X1 U9367 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7735), .ZN(n7734) );
  MUX2_X1 U9368 ( .A(n9895), .B(P2_REG1_REG_12__SCAN_IN), .S(n7696), .Z(n7679)
         );
  OAI21_X1 U9369 ( .B1(n7680), .B2(n7679), .A(n7765), .ZN(n7701) );
  INV_X1 U9370 ( .A(n7681), .ZN(n7737) );
  MUX2_X1 U9371 ( .A(n7683), .B(n7682), .S(n8478), .Z(n7684) );
  NAND2_X1 U9372 ( .A1(n7684), .A2(n7742), .ZN(n7693) );
  INV_X1 U9373 ( .A(n7684), .ZN(n7686) );
  NAND2_X1 U9374 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  AND2_X1 U9375 ( .A1(n7693), .A2(n7687), .ZN(n7736) );
  OAI21_X1 U9376 ( .B1(n7738), .B2(n7737), .A(n7736), .ZN(n7740) );
  MUX2_X1 U9377 ( .A(n7688), .B(n9895), .S(n8478), .Z(n7689) );
  NAND2_X1 U9378 ( .A1(n7689), .A2(n7696), .ZN(n7768) );
  INV_X1 U9379 ( .A(n7689), .ZN(n7690) );
  NAND2_X1 U9380 ( .A1(n7690), .A2(n7764), .ZN(n7691) );
  NAND2_X1 U9381 ( .A1(n7768), .A2(n7691), .ZN(n7692) );
  AOI21_X1 U9382 ( .B1(n7740), .B2(n7693), .A(n7692), .ZN(n7774) );
  AND3_X1 U9383 ( .A1(n7740), .A2(n7693), .A3(n7692), .ZN(n7694) );
  OAI21_X1 U9384 ( .B1(n7774), .B2(n7694), .A(n9788), .ZN(n7698) );
  INV_X1 U9385 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7695) );
  NOR2_X1 U9386 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7695), .ZN(n7787) );
  AOI21_X1 U9387 ( .B1(n9783), .B2(n7696), .A(n7787), .ZN(n7697) );
  OAI211_X1 U9388 ( .C1(n7699), .C2(n9768), .A(n7698), .B(n7697), .ZN(n7700)
         );
  AOI21_X1 U9389 ( .B1(n7701), .B2(n8542), .A(n7700), .ZN(n7702) );
  OAI21_X1 U9390 ( .B1(n7703), .B2(n9778), .A(n7702), .ZN(P2_U3194) );
  XNOR2_X1 U9391 ( .A(n7705), .B(n7704), .ZN(n9536) );
  AOI21_X1 U9392 ( .B1(n7708), .B2(n7707), .A(n7706), .ZN(n7709) );
  NOR3_X1 U9393 ( .A1(n7710), .A2(n7709), .A3(n9715), .ZN(n7712) );
  AOI211_X1 U9394 ( .C1(n9536), .C2(n9446), .A(n7712), .B(n7711), .ZN(n9540)
         );
  INV_X1 U9395 ( .A(n7713), .ZN(n7715) );
  AOI211_X1 U9396 ( .C1(n9538), .C2(n7715), .A(n9418), .B(n7714), .ZN(n9537)
         );
  NAND2_X1 U9397 ( .A1(n9537), .A2(n9450), .ZN(n7718) );
  AOI22_X1 U9398 ( .A1(n9709), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7716), .B2(
        n9703), .ZN(n7717) );
  OAI211_X1 U9399 ( .C1(n7719), .C2(n9692), .A(n7718), .B(n7717), .ZN(n7720)
         );
  AOI21_X1 U9400 ( .B1(n9536), .B2(n9681), .A(n7720), .ZN(n7721) );
  OAI21_X1 U9401 ( .B1(n9540), .B2(n9709), .A(n7721), .ZN(P1_U3279) );
  AOI211_X1 U9402 ( .C1(n7724), .C2(n9735), .A(n7723), .B(n7722), .ZN(n7731)
         );
  AOI22_X1 U9403 ( .A1(n7729), .A2(n7725), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n7727), .ZN(n7726) );
  OAI21_X1 U9404 ( .B1(n7731), .B2(n7727), .A(n7726), .ZN(P1_U3492) );
  AOI22_X1 U9405 ( .A1(n7729), .A2(n7728), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9743), .ZN(n7730) );
  OAI21_X1 U9406 ( .B1(n7731), .B2(n9743), .A(n7730), .ZN(P1_U3535) );
  AOI21_X1 U9407 ( .B1(n7683), .B2(n7733), .A(n7732), .ZN(n7748) );
  OAI21_X1 U9408 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7735), .A(n7734), .ZN(
        n7746) );
  AND2_X1 U9409 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7757) );
  OR3_X1 U9410 ( .A1(n7738), .A2(n7737), .A3(n7736), .ZN(n7739) );
  AOI21_X1 U9411 ( .B1(n7740), .B2(n7739), .A(n8534), .ZN(n7741) );
  AOI211_X1 U9412 ( .C1(n7742), .C2(n9783), .A(n7757), .B(n7741), .ZN(n7743)
         );
  OAI21_X1 U9413 ( .B1(n7744), .B2(n9768), .A(n7743), .ZN(n7745) );
  AOI21_X1 U9414 ( .B1(n7746), .B2(n8542), .A(n7745), .ZN(n7747) );
  OAI21_X1 U9415 ( .B1(n7748), .B2(n9778), .A(n7747), .ZN(P2_U3193) );
  XNOR2_X1 U9416 ( .A(n7749), .B(n8261), .ZN(n7784) );
  INV_X1 U9417 ( .A(n7750), .ZN(n7751) );
  OAI22_X1 U9418 ( .A1(n7753), .A2(n7752), .B1(n8425), .B2(n7751), .ZN(n7754)
         );
  NOR2_X1 U9419 ( .A1(n7754), .A2(n7784), .ZN(n7785) );
  AOI211_X1 U9420 ( .C1(n7784), .C2(n7754), .A(n8383), .B(n7785), .ZN(n7755)
         );
  INV_X1 U9421 ( .A(n7755), .ZN(n7759) );
  OAI22_X1 U9422 ( .A1(n10131), .A2(n10129), .B1(n9866), .B2(n8403), .ZN(n7756) );
  AOI211_X1 U9423 ( .C1(n8408), .C2(n8423), .A(n7757), .B(n7756), .ZN(n7758)
         );
  OAI211_X1 U9424 ( .C1(n7760), .C2(n10138), .A(n7759), .B(n7758), .ZN(
        P2_U3176) );
  AOI21_X1 U9425 ( .B1(n8775), .B2(n7763), .A(n7813), .ZN(n7783) );
  NAND2_X1 U9426 ( .A1(n7764), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U9427 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7767), .ZN(n7819) );
  OAI21_X1 U9428 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7767), .A(n7819), .ZN(
        n7781) );
  INV_X1 U9429 ( .A(n7768), .ZN(n7773) );
  MUX2_X1 U9430 ( .A(n8775), .B(n8867), .S(n8478), .Z(n7769) );
  NAND2_X1 U9431 ( .A1(n7769), .A2(n7812), .ZN(n7829) );
  INV_X1 U9432 ( .A(n7769), .ZN(n7770) );
  NAND2_X1 U9433 ( .A1(n7770), .A2(n7818), .ZN(n7771) );
  AND2_X1 U9434 ( .A1(n7829), .A2(n7771), .ZN(n7772) );
  INV_X1 U9435 ( .A(n7830), .ZN(n7776) );
  NOR3_X1 U9436 ( .A1(n7774), .A2(n7773), .A3(n7772), .ZN(n7775) );
  OAI21_X1 U9437 ( .B1(n7776), .B2(n7775), .A(n9788), .ZN(n7778) );
  AND2_X1 U9438 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8371) );
  AOI21_X1 U9439 ( .B1(n9783), .B2(n7812), .A(n8371), .ZN(n7777) );
  OAI211_X1 U9440 ( .C1(n7779), .C2(n9768), .A(n7778), .B(n7777), .ZN(n7780)
         );
  AOI21_X1 U9441 ( .B1(n7781), .B2(n8542), .A(n7780), .ZN(n7782) );
  OAI21_X1 U9442 ( .B1(n7783), .B2(n9778), .A(n7782), .ZN(P2_U3195) );
  NOR2_X1 U9443 ( .A1(n7785), .A2(n4869), .ZN(n8005) );
  XNOR2_X1 U9444 ( .A(n9876), .B(n8261), .ZN(n8004) );
  XNOR2_X1 U9445 ( .A(n8004), .B(n8423), .ZN(n7786) );
  XNOR2_X1 U9446 ( .A(n8005), .B(n7786), .ZN(n7792) );
  AOI21_X1 U9447 ( .B1(n8408), .B2(n8422), .A(n7787), .ZN(n7789) );
  NAND2_X1 U9448 ( .A1(n8409), .A2(n8424), .ZN(n7788) );
  OAI211_X1 U9449 ( .C1(n10138), .C2(n7793), .A(n7789), .B(n7788), .ZN(n7790)
         );
  AOI21_X1 U9450 ( .B1(n9876), .B2(n10134), .A(n7790), .ZN(n7791) );
  OAI21_X1 U9451 ( .B1(n7792), .B2(n8383), .A(n7791), .ZN(P2_U3164) );
  INV_X1 U9452 ( .A(n7793), .ZN(n7797) );
  XNOR2_X1 U9453 ( .A(n7794), .B(n8157), .ZN(n7795) );
  OAI222_X1 U9454 ( .A1(n9813), .A2(n8746), .B1(n9794), .B2(n7796), .C1(n9797), 
        .C2(n7795), .ZN(n9874) );
  AOI21_X1 U9455 ( .B1(n9804), .B2(n7797), .A(n9874), .ZN(n7804) );
  INV_X1 U9456 ( .A(n7798), .ZN(n7799) );
  INV_X1 U9457 ( .A(n8157), .ZN(n8081) );
  OR2_X1 U9458 ( .A1(n7798), .A2(n8157), .ZN(n8770) );
  OAI21_X1 U9459 ( .B1(n7799), .B2(n8081), .A(n8770), .ZN(n9873) );
  INV_X1 U9460 ( .A(n9873), .ZN(n7802) );
  INV_X1 U9461 ( .A(n9876), .ZN(n7800) );
  OAI22_X1 U9462 ( .A1(n7800), .A2(n8721), .B1(n9807), .B2(n7688), .ZN(n7801)
         );
  AOI21_X1 U9463 ( .B1(n7802), .B2(n8777), .A(n7801), .ZN(n7803) );
  OAI21_X1 U9464 ( .B1(n7804), .B2(n9808), .A(n7803), .ZN(P2_U3221) );
  INV_X1 U9465 ( .A(n7805), .ZN(n7809) );
  OAI222_X1 U9466 ( .A1(n7807), .A2(P1_U3086), .B1(n8275), .B2(n7809), .C1(
        n7806), .C2(n8273), .ZN(P1_U3331) );
  OAI222_X1 U9467 ( .A1(P2_U3151), .A2(n7810), .B1(n8937), .B2(n7809), .C1(
        n7808), .C2(n8277), .ZN(P2_U3271) );
  NOR2_X1 U9468 ( .A1(n7812), .A2(n7811), .ZN(n7814) );
  NAND2_X1 U9469 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8454), .ZN(n7815) );
  OAI21_X1 U9470 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8454), .A(n7815), .ZN(
        n7816) );
  AOI21_X1 U9471 ( .B1(n4430), .B2(n7816), .A(n8452), .ZN(n7837) );
  NAND2_X1 U9472 ( .A1(n7818), .A2(n7817), .ZN(n7820) );
  XNOR2_X1 U9473 ( .A(n8454), .B(n8862), .ZN(n7821) );
  OAI21_X1 U9474 ( .B1(n7822), .B2(n7821), .A(n8455), .ZN(n7835) );
  MUX2_X1 U9475 ( .A(n7823), .B(n8862), .S(n8478), .Z(n7825) );
  NAND2_X1 U9476 ( .A1(n7824), .A2(n7825), .ZN(n8458) );
  INV_X1 U9477 ( .A(n7825), .ZN(n7826) );
  NAND2_X1 U9478 ( .A1(n7826), .A2(n8454), .ZN(n7827) );
  NAND2_X1 U9479 ( .A1(n8458), .A2(n7827), .ZN(n7828) );
  NAND3_X1 U9480 ( .A1(n7830), .A2(n7829), .A3(n7828), .ZN(n7831) );
  AOI21_X1 U9481 ( .B1(n4420), .B2(n7831), .A(n8534), .ZN(n7834) );
  NAND2_X1 U9482 ( .A1(n8555), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7832) );
  NAND2_X1 U9483 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8292) );
  OAI211_X1 U9484 ( .C1(n8559), .C2(n8454), .A(n7832), .B(n8292), .ZN(n7833)
         );
  AOI211_X1 U9485 ( .C1(n7835), .C2(n8542), .A(n7834), .B(n7833), .ZN(n7836)
         );
  OAI21_X1 U9486 ( .B1(n7837), .B2(n9778), .A(n7836), .ZN(P2_U3196) );
  XNOR2_X1 U9487 ( .A(n7838), .B(n4393), .ZN(n9527) );
  INV_X1 U9488 ( .A(n9527), .ZN(n7850) );
  OAI21_X1 U9489 ( .B1(n4393), .B2(n7840), .A(n7839), .ZN(n7841) );
  NAND2_X1 U9490 ( .A1(n7841), .A2(n9391), .ZN(n7844) );
  NAND2_X1 U9491 ( .A1(n9118), .A2(n9070), .ZN(n7843) );
  NAND2_X1 U9492 ( .A1(n9116), .A2(n9069), .ZN(n7842) );
  AND2_X1 U9493 ( .A1(n7843), .A2(n7842), .ZN(n9020) );
  NAND2_X1 U9494 ( .A1(n7844), .A2(n9020), .ZN(n9525) );
  INV_X1 U9495 ( .A(n9022), .ZN(n9587) );
  AOI211_X1 U9496 ( .C1(n9022), .C2(n7845), .A(n9418), .B(n4707), .ZN(n9526)
         );
  NAND2_X1 U9497 ( .A1(n9526), .A2(n9450), .ZN(n7847) );
  AOI22_X1 U9498 ( .A1(n9709), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9017), .B2(
        n9703), .ZN(n7846) );
  OAI211_X1 U9499 ( .C1(n9587), .C2(n9692), .A(n7847), .B(n7846), .ZN(n7848)
         );
  AOI21_X1 U9500 ( .B1(n9439), .B2(n9525), .A(n7848), .ZN(n7849) );
  OAI21_X1 U9501 ( .B1(n7850), .B2(n9426), .A(n7849), .ZN(P1_U3277) );
  XNOR2_X1 U9502 ( .A(n7851), .B(n7855), .ZN(n9524) );
  INV_X1 U9503 ( .A(n9419), .ZN(n7852) );
  AOI211_X1 U9504 ( .C1(n9521), .C2(n7853), .A(n9418), .B(n7852), .ZN(n9520)
         );
  AOI22_X1 U9505 ( .A1(n9709), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9027), .B2(
        n9703), .ZN(n7854) );
  OAI21_X1 U9506 ( .B1(n7931), .B2(n9692), .A(n7854), .ZN(n7861) );
  XNOR2_X1 U9507 ( .A(n7856), .B(n7855), .ZN(n7859) );
  OR2_X1 U9508 ( .A1(n7920), .A2(n9082), .ZN(n7858) );
  OR2_X1 U9509 ( .A1(n8965), .A2(n9080), .ZN(n7857) );
  NAND2_X1 U9510 ( .A1(n7858), .A2(n7857), .ZN(n9028) );
  AOI21_X1 U9511 ( .B1(n7859), .B2(n9391), .A(n9028), .ZN(n9523) );
  NOR2_X1 U9512 ( .A1(n9523), .A2(n9689), .ZN(n7860) );
  AOI211_X1 U9513 ( .C1(n9520), .C2(n9450), .A(n7861), .B(n7860), .ZN(n7862)
         );
  OAI21_X1 U9514 ( .B1(n9524), .B2(n9426), .A(n7862), .ZN(P1_U3276) );
  INV_X1 U9515 ( .A(n7863), .ZN(n7866) );
  OAI222_X1 U9516 ( .A1(P2_U3151), .A2(n7864), .B1(n8937), .B2(n7866), .C1(
        n9939), .C2(n8277), .ZN(P2_U3270) );
  OAI222_X1 U9517 ( .A1(n7867), .A2(P1_U3086), .B1(n8275), .B2(n7866), .C1(
        n7865), .C2(n8273), .ZN(P1_U3330) );
  INV_X1 U9518 ( .A(n7868), .ZN(n7871) );
  OAI222_X1 U9519 ( .A1(n7870), .A2(P1_U3086), .B1(n8275), .B2(n7871), .C1(
        n7869), .C2(n8273), .ZN(P1_U3329) );
  OAI222_X1 U9520 ( .A1(P2_U3151), .A2(n7872), .B1(n8937), .B2(n7871), .C1(
        n10085), .C2(n8277), .ZN(P2_U3269) );
  NAND2_X1 U9521 ( .A1(n8049), .A2(n8941), .ZN(n7874) );
  OAI211_X1 U9522 ( .C1(n8277), .C2(n7875), .A(n7874), .B(n7873), .ZN(P2_U3268) );
  OAI22_X1 U9523 ( .A1(n9807), .A2(n10069), .B1(n7877), .B2(n8773), .ZN(n7880)
         );
  NOR2_X1 U9524 ( .A1(n7878), .A2(n9801), .ZN(n7879) );
  AOI211_X1 U9525 ( .C1(n9802), .C2(n6098), .A(n7880), .B(n7879), .ZN(n7881)
         );
  OAI21_X1 U9526 ( .B1(n7876), .B2(n9808), .A(n7881), .ZN(P2_U3204) );
  INV_X1 U9527 ( .A(n7882), .ZN(n8938) );
  OAI222_X1 U9528 ( .A1(n8273), .A2(n7884), .B1(P1_U3086), .B2(n7883), .C1(
        n8271), .C2(n8938), .ZN(P1_U3326) );
  NOR4_X1 U9529 ( .A1(n5051), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7886), .A4(
        P1_U3086), .ZN(n7887) );
  AOI21_X1 U9530 ( .B1(n7888), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n7887), .ZN(
        n7889) );
  OAI21_X1 U9531 ( .B1(n7885), .B2(n8271), .A(n7889), .ZN(P1_U3324) );
  INV_X1 U9532 ( .A(n7890), .ZN(n7891) );
  NOR4_X1 U9533 ( .A1(n7891), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4505), .A4(
        P2_U3151), .ZN(n7892) );
  AOI21_X1 U9534 ( .B1(n7893), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n7892), .ZN(
        n7894) );
  OAI21_X1 U9535 ( .B1(n7885), .B2(n8937), .A(n7894), .ZN(P2_U3264) );
  INV_X1 U9536 ( .A(n8942), .ZN(n7895) );
  OAI222_X1 U9537 ( .A1(n8273), .A2(n7896), .B1(P1_U3086), .B2(n5695), .C1(
        n8271), .C2(n7895), .ZN(P1_U3327) );
  NAND2_X1 U9538 ( .A1(n7897), .A2(n8717), .ZN(n8684) );
  NAND2_X1 U9539 ( .A1(n8684), .A2(n7898), .ZN(n7900) );
  NAND2_X1 U9540 ( .A1(n7900), .A2(n7899), .ZN(n7902) );
  OAI21_X1 U9541 ( .B1(n7902), .B2(n8088), .A(n7901), .ZN(n7904) );
  NOR2_X1 U9542 ( .A1(n8689), .A2(n9794), .ZN(n7903) );
  AOI21_X1 U9543 ( .B1(n7904), .B2(n8726), .A(n7903), .ZN(n8832) );
  XNOR2_X1 U9544 ( .A(n7906), .B(n7905), .ZN(n8830) );
  NAND2_X1 U9545 ( .A1(n8908), .A2(n9802), .ZN(n7908) );
  AOI22_X1 U9546 ( .A1(n9808), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9804), .B2(
        n8365), .ZN(n7907) );
  OAI211_X1 U9547 ( .C1(n8833), .C2(n8660), .A(n7908), .B(n7907), .ZN(n7909)
         );
  AOI21_X1 U9548 ( .B1(n8830), .B2(n8777), .A(n7909), .ZN(n7910) );
  OAI21_X1 U9549 ( .B1(n8832), .B2(n9808), .A(n7910), .ZN(P2_U3213) );
  NAND2_X1 U9550 ( .A1(n9349), .A2(n8970), .ZN(n7912) );
  NAND2_X1 U9551 ( .A1(n9112), .A2(n8975), .ZN(n7911) );
  NAND2_X1 U9552 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  XNOR2_X1 U9553 ( .A(n7913), .B(n7975), .ZN(n7958) );
  NAND2_X1 U9554 ( .A1(n9532), .A2(n8970), .ZN(n7915) );
  NAND2_X1 U9555 ( .A1(n9118), .A2(n8975), .ZN(n7914) );
  NAND2_X1 U9556 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  XNOR2_X1 U9557 ( .A(n7916), .B(n7975), .ZN(n7919) );
  AOI22_X1 U9558 ( .A1(n9532), .A2(n7965), .B1(n7977), .B2(n9118), .ZN(n9094)
         );
  NAND2_X1 U9559 ( .A1(n9022), .A2(n8970), .ZN(n7922) );
  OR2_X1 U9560 ( .A1(n7920), .A2(n7984), .ZN(n7921) );
  NAND2_X1 U9561 ( .A1(n7922), .A2(n7921), .ZN(n7923) );
  XNOR2_X1 U9562 ( .A(n7923), .B(n7975), .ZN(n7924) );
  AOI22_X1 U9563 ( .A1(n9022), .A2(n7965), .B1(n7977), .B2(n9117), .ZN(n7925)
         );
  XNOR2_X1 U9564 ( .A(n7924), .B(n7925), .ZN(n9016) );
  INV_X1 U9565 ( .A(n7924), .ZN(n7926) );
  NAND2_X1 U9566 ( .A1(n9521), .A2(n8970), .ZN(n7928) );
  NAND2_X1 U9567 ( .A1(n9116), .A2(n8975), .ZN(n7927) );
  NAND2_X1 U9568 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  XNOR2_X1 U9569 ( .A(n7929), .B(n7975), .ZN(n7933) );
  OAI22_X1 U9570 ( .A1(n7931), .A2(n7984), .B1(n7930), .B2(n8977), .ZN(n7932)
         );
  XNOR2_X1 U9571 ( .A(n7933), .B(n7932), .ZN(n9026) );
  OAI22_X1 U9572 ( .A1(n9581), .A2(n7971), .B1(n8965), .B2(n7984), .ZN(n7934)
         );
  XNOR2_X1 U9573 ( .A(n7934), .B(n7975), .ZN(n9067) );
  OR2_X1 U9574 ( .A1(n9581), .A2(n7984), .ZN(n7936) );
  OR2_X1 U9575 ( .A1(n8965), .A2(n8977), .ZN(n7935) );
  NAND2_X1 U9576 ( .A1(n7936), .A2(n7935), .ZN(n9066) );
  NOR2_X1 U9577 ( .A1(n9067), .A2(n9066), .ZN(n7939) );
  INV_X1 U9578 ( .A(n9067), .ZN(n7938) );
  INV_X1 U9579 ( .A(n9066), .ZN(n7937) );
  NAND2_X1 U9580 ( .A1(n9512), .A2(n8970), .ZN(n7941) );
  NAND2_X1 U9581 ( .A1(n9114), .A2(n8975), .ZN(n7940) );
  NAND2_X1 U9582 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  XNOR2_X1 U9583 ( .A(n7942), .B(n8973), .ZN(n7945) );
  AND2_X1 U9584 ( .A1(n9114), .A2(n7977), .ZN(n7943) );
  AOI21_X1 U9585 ( .B1(n9512), .B2(n7965), .A(n7943), .ZN(n7944) );
  NOR2_X1 U9586 ( .A1(n7945), .A2(n7944), .ZN(n8960) );
  OAI22_X1 U9587 ( .A1(n9386), .A2(n7971), .B1(n7947), .B2(n7984), .ZN(n7946)
         );
  XNOR2_X1 U9588 ( .A(n7946), .B(n7975), .ZN(n7948) );
  OAI22_X1 U9589 ( .A1(n9386), .A2(n7984), .B1(n7947), .B2(n8977), .ZN(n7949)
         );
  XNOR2_X1 U9590 ( .A(n7948), .B(n7949), .ZN(n9047) );
  INV_X1 U9591 ( .A(n7948), .ZN(n7951) );
  INV_X1 U9592 ( .A(n7949), .ZN(n7950) );
  OAI22_X1 U9593 ( .A1(n9575), .A2(n7971), .B1(n9057), .B2(n7984), .ZN(n7952)
         );
  XNOR2_X1 U9594 ( .A(n7952), .B(n7975), .ZN(n7954) );
  OAI22_X1 U9595 ( .A1(n9575), .A2(n7984), .B1(n9057), .B2(n8977), .ZN(n7953)
         );
  XNOR2_X1 U9596 ( .A(n7954), .B(n7953), .ZN(n8997) );
  OR2_X1 U9597 ( .A1(n7954), .A2(n7953), .ZN(n7955) );
  OAI22_X1 U9598 ( .A1(n9571), .A2(n7984), .B1(n7956), .B2(n8977), .ZN(n9055)
         );
  OAI22_X1 U9599 ( .A1(n9344), .A2(n7971), .B1(n9058), .B2(n7984), .ZN(n7961)
         );
  XOR2_X1 U9600 ( .A(n7975), .B(n7961), .Z(n7963) );
  INV_X1 U9601 ( .A(n9058), .ZN(n9111) );
  AOI22_X1 U9602 ( .A1(n9491), .A2(n7965), .B1(n7977), .B2(n9111), .ZN(n7962)
         );
  NOR2_X1 U9603 ( .A1(n7963), .A2(n7962), .ZN(n8950) );
  NAND2_X1 U9604 ( .A1(n7963), .A2(n7962), .ZN(n8948) );
  AOI22_X1 U9605 ( .A1(n9486), .A2(n8970), .B1(n7965), .B2(n9110), .ZN(n7964)
         );
  XOR2_X1 U9606 ( .A(n7975), .B(n7964), .Z(n7968) );
  OAI22_X1 U9607 ( .A1(n9329), .A2(n7984), .B1(n7966), .B2(n8977), .ZN(n7967)
         );
  NOR2_X1 U9608 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  AOI21_X1 U9609 ( .B1(n7968), .B2(n7967), .A(n7969), .ZN(n9037) );
  NAND2_X1 U9610 ( .A1(n9036), .A2(n9037), .ZN(n9035) );
  INV_X1 U9611 ( .A(n7969), .ZN(n7970) );
  OAI22_X1 U9612 ( .A1(n9566), .A2(n7984), .B1(n9083), .B2(n8977), .ZN(n7980)
         );
  OAI22_X1 U9613 ( .A1(n9566), .A2(n7971), .B1(n9083), .B2(n7984), .ZN(n7972)
         );
  XNOR2_X1 U9614 ( .A(n7972), .B(n7975), .ZN(n7979) );
  XOR2_X1 U9615 ( .A(n7980), .B(n7979), .Z(n9006) );
  NAND2_X1 U9616 ( .A1(n9293), .A2(n8970), .ZN(n7974) );
  NAND2_X1 U9617 ( .A1(n9109), .A2(n8975), .ZN(n7973) );
  NAND2_X1 U9618 ( .A1(n7974), .A2(n7973), .ZN(n7976) );
  XNOR2_X1 U9619 ( .A(n7976), .B(n7975), .ZN(n7995) );
  AND2_X1 U9620 ( .A1(n9109), .A2(n7977), .ZN(n7978) );
  AOI21_X1 U9621 ( .B1(n9293), .B2(n7965), .A(n7978), .ZN(n7993) );
  XNOR2_X1 U9622 ( .A(n7995), .B(n7993), .ZN(n9078) );
  INV_X1 U9623 ( .A(n7979), .ZN(n7982) );
  INV_X1 U9624 ( .A(n7980), .ZN(n7981) );
  NAND2_X1 U9625 ( .A1(n7982), .A2(n7981), .ZN(n9079) );
  NAND2_X1 U9626 ( .A1(n9278), .A2(n8970), .ZN(n7986) );
  OR2_X1 U9627 ( .A1(n9081), .A2(n7984), .ZN(n7985) );
  NAND2_X1 U9628 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  XNOR2_X1 U9629 ( .A(n7987), .B(n8973), .ZN(n7990) );
  INV_X1 U9630 ( .A(n7990), .ZN(n7992) );
  NOR2_X1 U9631 ( .A1(n9081), .A2(n8977), .ZN(n7988) );
  AOI21_X1 U9632 ( .B1(n9278), .B2(n7965), .A(n7988), .ZN(n7989) );
  INV_X1 U9633 ( .A(n7989), .ZN(n7991) );
  AOI21_X1 U9634 ( .B1(n7992), .B2(n7991), .A(n8991), .ZN(n7996) );
  INV_X1 U9635 ( .A(n7993), .ZN(n7994) );
  NAND2_X1 U9636 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  AND2_X1 U9637 ( .A1(n9109), .A2(n9070), .ZN(n7998) );
  AOI21_X1 U9638 ( .B1(n9108), .B2(n9069), .A(n7998), .ZN(n9273) );
  INV_X1 U9639 ( .A(n9273), .ZN(n8002) );
  INV_X1 U9640 ( .A(n9279), .ZN(n8000) );
  OAI22_X1 U9641 ( .A1(n8000), .A2(n9061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7999), .ZN(n8001) );
  AOI21_X1 U9642 ( .B1(n8002), .B2(n9059), .A(n8001), .ZN(n8003) );
  XNOR2_X1 U9643 ( .A(n8864), .B(n6302), .ZN(n8006) );
  NOR2_X1 U9644 ( .A1(n8006), .A2(n8746), .ZN(n8368) );
  XNOR2_X1 U9645 ( .A(n8750), .B(n8261), .ZN(n8007) );
  XNOR2_X1 U9646 ( .A(n8007), .B(n8767), .ZN(n8291) );
  INV_X1 U9647 ( .A(n8007), .ZN(n8008) );
  XNOR2_X1 U9648 ( .A(n8854), .B(n8261), .ZN(n8009) );
  XNOR2_X1 U9649 ( .A(n8009), .B(n8745), .ZN(n8406) );
  NAND2_X1 U9650 ( .A1(n8407), .A2(n8406), .ZN(n8405) );
  INV_X1 U9651 ( .A(n8009), .ZN(n8010) );
  NAND2_X1 U9652 ( .A1(n8405), .A2(n4874), .ZN(n8335) );
  XNOR2_X1 U9653 ( .A(n8332), .B(n8261), .ZN(n8011) );
  XNOR2_X1 U9654 ( .A(n8011), .B(n8705), .ZN(n8334) );
  NAND2_X1 U9655 ( .A1(n8335), .A2(n8334), .ZN(n8333) );
  XNOR2_X1 U9656 ( .A(n8708), .B(n6302), .ZN(n8340) );
  INV_X1 U9657 ( .A(n8340), .ZN(n8013) );
  XNOR2_X1 U9658 ( .A(n8385), .B(n8261), .ZN(n8014) );
  XNOR2_X1 U9659 ( .A(n8014), .B(n8706), .ZN(n8388) );
  XNOR2_X1 U9660 ( .A(n5983), .B(n8261), .ZN(n8017) );
  XNOR2_X1 U9661 ( .A(n8017), .B(n8689), .ZN(n8308) );
  INV_X1 U9662 ( .A(n8014), .ZN(n8015) );
  NAND2_X1 U9663 ( .A1(n8015), .A2(n8706), .ZN(n8306) );
  XNOR2_X1 U9664 ( .A(n8908), .B(n8261), .ZN(n8016) );
  NOR2_X1 U9665 ( .A1(n8016), .A2(n8675), .ZN(n8019) );
  AOI21_X1 U9666 ( .B1(n8675), .B2(n8016), .A(n8019), .ZN(n8359) );
  NAND2_X1 U9667 ( .A1(n8017), .A2(n8419), .ZN(n8360) );
  NAND2_X1 U9668 ( .A1(n8307), .A2(n8018), .ZN(n8358) );
  INV_X1 U9669 ( .A(n8019), .ZN(n8315) );
  XNOR2_X1 U9670 ( .A(n8662), .B(n6302), .ZN(n8020) );
  NAND2_X1 U9671 ( .A1(n8020), .A2(n8833), .ZN(n8023) );
  INV_X1 U9672 ( .A(n8020), .ZN(n8021) );
  NAND2_X1 U9673 ( .A1(n8021), .A2(n6029), .ZN(n8022) );
  NAND2_X1 U9674 ( .A1(n8023), .A2(n8022), .ZN(n8314) );
  INV_X1 U9675 ( .A(n8023), .ZN(n8024) );
  XNOR2_X1 U9676 ( .A(n8817), .B(n8261), .ZN(n8025) );
  XNOR2_X1 U9677 ( .A(n8025), .B(n8418), .ZN(n8377) );
  INV_X1 U9678 ( .A(n8025), .ZN(n8026) );
  XNOR2_X1 U9679 ( .A(n8639), .B(n8261), .ZN(n8031) );
  NAND2_X1 U9680 ( .A1(n8030), .A2(n8031), .ZN(n8298) );
  XNOR2_X1 U9681 ( .A(n8893), .B(n8261), .ZN(n8027) );
  NAND2_X1 U9682 ( .A1(n8027), .A2(n8811), .ZN(n8322) );
  INV_X1 U9683 ( .A(n8027), .ZN(n8028) );
  NAND2_X1 U9684 ( .A1(n8028), .A2(n8416), .ZN(n8029) );
  AND2_X1 U9685 ( .A1(n8322), .A2(n8029), .ZN(n8350) );
  INV_X1 U9686 ( .A(n8031), .ZN(n8032) );
  NAND2_X1 U9687 ( .A1(n4666), .A2(n8032), .ZN(n8299) );
  NAND2_X1 U9688 ( .A1(n8299), .A2(n8417), .ZN(n8351) );
  NAND2_X1 U9689 ( .A1(n8033), .A2(n8351), .ZN(n8349) );
  XNOR2_X1 U9690 ( .A(n8614), .B(n8261), .ZN(n8037) );
  INV_X1 U9691 ( .A(n8037), .ZN(n8034) );
  NAND2_X1 U9692 ( .A1(n8034), .A2(n8623), .ZN(n8036) );
  AND2_X1 U9693 ( .A1(n8322), .A2(n8036), .ZN(n8035) );
  NAND2_X1 U9694 ( .A1(n8349), .A2(n8035), .ZN(n8040) );
  INV_X1 U9695 ( .A(n8036), .ZN(n8038) );
  XNOR2_X1 U9696 ( .A(n8037), .B(n8623), .ZN(n8325) );
  OR2_X1 U9697 ( .A1(n8038), .A2(n8325), .ZN(n8039) );
  XNOR2_X1 U9698 ( .A(n8404), .B(n8261), .ZN(n8394) );
  XNOR2_X1 U9699 ( .A(n8794), .B(n6302), .ZN(n8041) );
  NOR2_X1 U9700 ( .A1(n8041), .A2(n8604), .ZN(n8258) );
  AOI21_X1 U9701 ( .B1(n8041), .B2(n8604), .A(n8258), .ZN(n8042) );
  OAI211_X1 U9702 ( .C1(n8043), .C2(n8042), .A(n8260), .B(n10126), .ZN(n8047)
         );
  AOI22_X1 U9703 ( .A1(n8409), .A2(n8588), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8044) );
  OAI21_X1 U9704 ( .B1(n8592), .B2(n10128), .A(n8044), .ZN(n8045) );
  AOI21_X1 U9705 ( .B1(n8590), .B2(n8400), .A(n8045), .ZN(n8046) );
  OAI211_X1 U9706 ( .C1(n8048), .C2(n8403), .A(n8047), .B(n8046), .ZN(P2_U3154) );
  INV_X1 U9707 ( .A(n8049), .ZN(n8050) );
  OAI222_X1 U9708 ( .A1(n8273), .A2(n8051), .B1(P1_U3086), .B2(n5696), .C1(
        n8271), .C2(n8050), .ZN(P1_U3328) );
  NAND2_X1 U9709 ( .A1(n8269), .A2(n8052), .ZN(n8054) );
  OR2_X1 U9710 ( .A1(n8055), .A2(n8278), .ZN(n8053) );
  NAND2_X1 U9711 ( .A1(n8054), .A2(n8053), .ZN(n8879) );
  AND2_X1 U9712 ( .A1(n8785), .A2(n8415), .ZN(n8245) );
  OAI22_X1 U9713 ( .A1(n7885), .A2(n8056), .B1(n8055), .B2(n6402), .ZN(n8780)
         );
  INV_X1 U9714 ( .A(n8241), .ZN(n8059) );
  INV_X1 U9715 ( .A(n8415), .ZN(n8057) );
  NAND2_X1 U9716 ( .A1(n8879), .A2(n8057), .ZN(n8243) );
  AND2_X1 U9717 ( .A1(n8243), .A2(n8058), .ZN(n8228) );
  NAND2_X1 U9718 ( .A1(n8780), .A2(n8569), .ZN(n8064) );
  INV_X1 U9719 ( .A(n8780), .ZN(n8878) );
  NAND2_X1 U9720 ( .A1(n8785), .A2(n8569), .ZN(n8061) );
  AOI22_X1 U9721 ( .A1(n8062), .A2(n8064), .B1(n8878), .B2(n8061), .ZN(n8063)
         );
  INV_X1 U9722 ( .A(n8064), .ZN(n8233) );
  NOR2_X1 U9723 ( .A1(n8780), .A2(n8569), .ZN(n8247) );
  XNOR2_X2 U9724 ( .A(n8236), .B(n8793), .ZN(n8582) );
  INV_X1 U9725 ( .A(n8065), .ZN(n8223) );
  INV_X1 U9726 ( .A(n8219), .ZN(n8066) );
  INV_X1 U9727 ( .A(n8616), .ZN(n8610) );
  INV_X1 U9728 ( .A(n8067), .ZN(n8626) );
  INV_X1 U9729 ( .A(n8707), .ZN(n8172) );
  INV_X1 U9730 ( .A(n8743), .ZN(n8758) );
  INV_X1 U9731 ( .A(n8068), .ZN(n8101) );
  NOR2_X1 U9732 ( .A1(n8105), .A2(n8101), .ZN(n8097) );
  NAND2_X1 U9733 ( .A1(n8070), .A2(n8069), .ZN(n8102) );
  NAND2_X1 U9734 ( .A1(n8072), .A2(n8071), .ZN(n8098) );
  NOR2_X1 U9735 ( .A1(n8102), .A2(n8098), .ZN(n8073) );
  AND4_X1 U9736 ( .A1(n8097), .A2(n8109), .A3(n8073), .A4(n6908), .ZN(n8077)
         );
  NAND4_X1 U9737 ( .A1(n8077), .A2(n8076), .A3(n8075), .A4(n8074), .ZN(n8079)
         );
  NOR4_X1 U9738 ( .A1(n8079), .A2(n8143), .A3(n9795), .A4(n8078), .ZN(n8082)
         );
  NAND4_X1 U9739 ( .A1(n8772), .A2(n8082), .A3(n8081), .A4(n8080), .ZN(n8083)
         );
  OR3_X1 U9740 ( .A1(n8758), .A2(n8083), .A3(n8163), .ZN(n8084) );
  NOR2_X1 U9741 ( .A1(n8717), .A2(n8084), .ZN(n8085) );
  NAND4_X1 U9742 ( .A1(n8668), .A2(n8172), .A3(n8086), .A4(n8085), .ZN(n8087)
         );
  OR3_X1 U9743 ( .A1(n8654), .A2(n8088), .A3(n8087), .ZN(n8089) );
  NOR3_X1 U9744 ( .A1(n8634), .A2(n8643), .A3(n8089), .ZN(n8090) );
  NAND4_X1 U9745 ( .A1(n8598), .A2(n8610), .A3(n8629), .A4(n8090), .ZN(n8091)
         );
  INV_X1 U9746 ( .A(n8245), .ZN(n8239) );
  NAND2_X1 U9747 ( .A1(n8239), .A2(n8243), .ZN(n8093) );
  INV_X1 U9748 ( .A(n8097), .ZN(n8100) );
  INV_X1 U9749 ( .A(n8098), .ZN(n8103) );
  OAI211_X1 U9750 ( .C1(n8100), .C2(n8103), .A(n8111), .B(n8099), .ZN(n8108)
         );
  AOI21_X1 U9751 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8106) );
  OAI211_X1 U9752 ( .C1(n8106), .C2(n8105), .A(n8104), .B(n8117), .ZN(n8107)
         );
  NAND2_X1 U9753 ( .A1(n8110), .A2(n8109), .ZN(n8121) );
  INV_X1 U9754 ( .A(n8111), .ZN(n8113) );
  OAI211_X1 U9755 ( .C1(n8121), .C2(n8113), .A(n8122), .B(n8112), .ZN(n8114)
         );
  NAND3_X1 U9756 ( .A1(n8114), .A2(n8125), .A3(n8119), .ZN(n8116) );
  INV_X1 U9757 ( .A(n8115), .ZN(n8123) );
  NAND2_X1 U9758 ( .A1(n8116), .A2(n8123), .ZN(n8128) );
  INV_X1 U9759 ( .A(n8117), .ZN(n8120) );
  OAI211_X1 U9760 ( .C1(n8121), .C2(n8120), .A(n8119), .B(n8118), .ZN(n8124)
         );
  NAND3_X1 U9761 ( .A1(n8124), .A2(n8123), .A3(n8122), .ZN(n8126) );
  NAND2_X1 U9762 ( .A1(n8126), .A2(n8125), .ZN(n8127) );
  MUX2_X1 U9763 ( .A(n8128), .B(n8127), .S(n8246), .Z(n8133) );
  NAND2_X1 U9764 ( .A1(n8134), .A2(n8129), .ZN(n8131) );
  NAND2_X1 U9765 ( .A1(n8137), .A2(n8138), .ZN(n8130) );
  OAI211_X1 U9766 ( .C1(n8140), .C2(n8135), .A(n4880), .B(n8134), .ZN(n8142)
         );
  AND2_X1 U9767 ( .A1(n8137), .A2(n8136), .ZN(n8139) );
  OAI211_X1 U9768 ( .C1(n8140), .C2(n8139), .A(n8138), .B(n8149), .ZN(n8141)
         );
  MUX2_X1 U9769 ( .A(n8142), .B(n8141), .S(n8246), .Z(n8144) );
  NOR3_X1 U9770 ( .A1(n8145), .A2(n8144), .A3(n8143), .ZN(n8154) );
  INV_X1 U9771 ( .A(n8150), .ZN(n8146) );
  OAI21_X1 U9772 ( .B1(n8146), .B2(n4880), .A(n8147), .ZN(n8152) );
  INV_X1 U9773 ( .A(n8147), .ZN(n8148) );
  AOI21_X1 U9774 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8151) );
  MUX2_X1 U9775 ( .A(n8152), .B(n8151), .S(n8227), .Z(n8153) );
  NOR2_X1 U9776 ( .A1(n8154), .A2(n8153), .ZN(n8158) );
  NAND2_X1 U9777 ( .A1(n9876), .A2(n8766), .ZN(n8155) );
  MUX2_X1 U9778 ( .A(n8769), .B(n8155), .S(n8227), .Z(n8156) );
  OAI211_X1 U9779 ( .C1(n8158), .C2(n8157), .A(n8772), .B(n8156), .ZN(n8162)
         );
  MUX2_X1 U9780 ( .A(n8160), .B(n8159), .S(n8246), .Z(n8161) );
  MUX2_X1 U9781 ( .A(n8165), .B(n8164), .S(n8227), .Z(n8166) );
  NAND2_X1 U9782 ( .A1(n8167), .A2(n8175), .ZN(n8174) );
  INV_X1 U9783 ( .A(n8168), .ZN(n8171) );
  NAND2_X1 U9784 ( .A1(n8187), .A2(n8169), .ZN(n8170) );
  MUX2_X1 U9785 ( .A(n8171), .B(n8170), .S(n8246), .Z(n8173) );
  INV_X1 U9786 ( .A(n8175), .ZN(n8176) );
  OAI211_X1 U9787 ( .C1(n8191), .C2(n8176), .A(n8692), .B(n8193), .ZN(n8177)
         );
  NAND3_X1 U9788 ( .A1(n8177), .A2(n8189), .A3(n8195), .ZN(n8178) );
  NAND3_X1 U9789 ( .A1(n8178), .A2(n8651), .A3(n8192), .ZN(n8180) );
  NAND3_X1 U9790 ( .A1(n8180), .A2(n8179), .A3(n8196), .ZN(n8183) );
  NAND3_X1 U9791 ( .A1(n8183), .A2(n8182), .A3(n8181), .ZN(n8186) );
  INV_X1 U9792 ( .A(n8184), .ZN(n8204) );
  AND3_X1 U9793 ( .A1(n8186), .A2(n8204), .A3(n8185), .ZN(n8203) );
  INV_X1 U9794 ( .A(n8187), .ZN(n8190) );
  OAI211_X1 U9795 ( .C1(n8191), .C2(n8190), .A(n8189), .B(n8188), .ZN(n8194)
         );
  NAND3_X1 U9796 ( .A1(n8194), .A2(n8193), .A3(n8192), .ZN(n8197) );
  NAND3_X1 U9797 ( .A1(n8197), .A2(n8196), .A3(n8195), .ZN(n8199) );
  AOI211_X1 U9798 ( .C1(n8824), .C2(n8817), .A(n8626), .B(n8201), .ZN(n8202)
         );
  NAND2_X1 U9799 ( .A1(n8204), .A2(n8207), .ZN(n8206) );
  OAI21_X1 U9800 ( .B1(n8209), .B2(n8206), .A(n8205), .ZN(n8211) );
  OAI21_X1 U9801 ( .B1(n8209), .B2(n8208), .A(n8207), .ZN(n8210) );
  MUX2_X1 U9802 ( .A(n8211), .B(n8210), .S(n8246), .Z(n8216) );
  INV_X1 U9803 ( .A(n8212), .ZN(n8213) );
  MUX2_X1 U9804 ( .A(n8214), .B(n8213), .S(n8227), .Z(n8215) );
  INV_X1 U9805 ( .A(n8217), .ZN(n8218) );
  MUX2_X1 U9806 ( .A(n8219), .B(n8218), .S(n8227), .Z(n8220) );
  MUX2_X1 U9807 ( .A(n8223), .B(n8222), .S(n8246), .Z(n8224) );
  NAND2_X1 U9808 ( .A1(n6098), .A2(n8246), .ZN(n8226) );
  INV_X1 U9809 ( .A(n8581), .ZN(n8786) );
  AOI22_X1 U9810 ( .A1(n8241), .A2(n8226), .B1(n8246), .B2(n8786), .ZN(n8230)
         );
  MUX2_X1 U9811 ( .A(n8592), .B(n8236), .S(n8227), .Z(n8231) );
  INV_X1 U9812 ( .A(n8228), .ZN(n8229) );
  NOR3_X1 U9813 ( .A1(n8238), .A2(n8246), .A3(n8229), .ZN(n8235) );
  AOI21_X1 U9814 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8237) );
  NAND2_X1 U9815 ( .A1(n8237), .A2(n8592), .ZN(n8234) );
  AOI21_X1 U9816 ( .B1(n8235), .B2(n8234), .A(n8233), .ZN(n8249) );
  NAND2_X1 U9817 ( .A1(n8237), .A2(n8236), .ZN(n8242) );
  INV_X1 U9818 ( .A(n8238), .ZN(n8240) );
  NAND4_X1 U9819 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n8244)
         );
  OAI211_X1 U9820 ( .C1(n8246), .C2(n8245), .A(n8244), .B(n8243), .ZN(n8248)
         );
  NAND3_X1 U9821 ( .A1(n8252), .A2(n8251), .A3(n8478), .ZN(n8253) );
  OAI211_X1 U9822 ( .C1(n8254), .C2(n8256), .A(n8253), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8255) );
  OAI21_X1 U9823 ( .B1(n8257), .B2(n8256), .A(n8255), .ZN(P2_U3296) );
  INV_X1 U9824 ( .A(n8258), .ZN(n8259) );
  XNOR2_X1 U9825 ( .A(n8582), .B(n8261), .ZN(n8262) );
  XNOR2_X1 U9826 ( .A(n8263), .B(n8262), .ZN(n8268) );
  NOR2_X1 U9827 ( .A1(n10138), .A2(n8578), .ZN(n8266) );
  AOI22_X1 U9828 ( .A1(n8409), .A2(n8798), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8264) );
  OAI21_X1 U9829 ( .B1(n8581), .B2(n10128), .A(n8264), .ZN(n8265) );
  AOI211_X1 U9830 ( .C1(n8787), .C2(n10134), .A(n8266), .B(n8265), .ZN(n8267)
         );
  OAI21_X1 U9831 ( .B1(n8268), .B2(n8383), .A(n8267), .ZN(P2_U3160) );
  INV_X1 U9832 ( .A(n8269), .ZN(n8279) );
  OAI222_X1 U9833 ( .A1(n8273), .A2(n8272), .B1(n8271), .B2(n8279), .C1(n8270), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U9834 ( .A1(n8273), .A2(n8276), .B1(n8275), .B2(n8274), .C1(
        P1_U3086), .C2(n9699), .ZN(P1_U3336) );
  OAI222_X1 U9835 ( .A1(P2_U3151), .A2(n5740), .B1(n8280), .B2(n8279), .C1(
        n8278), .C2(n8277), .ZN(P2_U3265) );
  NAND2_X1 U9836 ( .A1(n8281), .A2(n9686), .ZN(n8284) );
  AOI22_X1 U9837 ( .A1(n8282), .A2(n9703), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9709), .ZN(n8283) );
  OAI211_X1 U9838 ( .C1(n8285), .C2(n9692), .A(n8284), .B(n8283), .ZN(n8286)
         );
  AOI21_X1 U9839 ( .B1(n8287), .B2(n9439), .A(n8286), .ZN(n8288) );
  OAI21_X1 U9840 ( .B1(n8289), .B2(n9426), .A(n8288), .ZN(P1_U3356) );
  XOR2_X1 U9841 ( .A(n8291), .B(n8290), .Z(n8297) );
  NAND2_X1 U9842 ( .A1(n8409), .A2(n8422), .ZN(n8293) );
  OAI211_X1 U9843 ( .C1(n8745), .C2(n10128), .A(n8293), .B(n8292), .ZN(n8295)
         );
  NOR2_X1 U9844 ( .A1(n10138), .A2(n8751), .ZN(n8294) );
  AOI211_X1 U9845 ( .C1(n8750), .C2(n10134), .A(n8295), .B(n8294), .ZN(n8296)
         );
  OAI21_X1 U9846 ( .B1(n8297), .B2(n8383), .A(n8296), .ZN(P2_U3155) );
  NAND2_X1 U9847 ( .A1(n8298), .A2(n8299), .ZN(n8300) );
  XNOR2_X1 U9848 ( .A(n8300), .B(n8818), .ZN(n8305) );
  NAND2_X1 U9849 ( .A1(n8400), .A2(n8636), .ZN(n8302) );
  AOI22_X1 U9850 ( .A1(n8408), .A2(n8416), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8301) );
  OAI211_X1 U9851 ( .C1(n8824), .C2(n10131), .A(n8302), .B(n8301), .ZN(n8303)
         );
  AOI21_X1 U9852 ( .B1(n8639), .B2(n10134), .A(n8303), .ZN(n8304) );
  OAI21_X1 U9853 ( .B1(n8305), .B2(n8383), .A(n8304), .ZN(P2_U3156) );
  AND2_X1 U9854 ( .A1(n8386), .A2(n8306), .ZN(n8309) );
  OAI211_X1 U9855 ( .C1(n8309), .C2(n8308), .A(n10126), .B(n8307), .ZN(n8313)
         );
  NAND2_X1 U9856 ( .A1(n8409), .A2(n8674), .ZN(n8310) );
  NAND2_X1 U9857 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U9858 ( .C1(n8656), .C2(n10128), .A(n8310), .B(n8556), .ZN(n8311)
         );
  AOI21_X1 U9859 ( .B1(n8400), .B2(n8678), .A(n8311), .ZN(n8312) );
  OAI211_X1 U9860 ( .C1(n8914), .C2(n8403), .A(n8313), .B(n8312), .ZN(P2_U3159) );
  AND3_X1 U9861 ( .A1(n8358), .A2(n8315), .A3(n8314), .ZN(n8316) );
  OAI21_X1 U9862 ( .B1(n8317), .B2(n8316), .A(n10126), .ZN(n8321) );
  AOI22_X1 U9863 ( .A1(n8408), .A2(n8418), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8318) );
  OAI21_X1 U9864 ( .B1(n8656), .B2(n10131), .A(n8318), .ZN(n8319) );
  AOI21_X1 U9865 ( .B1(n8658), .B2(n8400), .A(n8319), .ZN(n8320) );
  OAI211_X1 U9866 ( .C1(n8905), .C2(n8403), .A(n8321), .B(n8320), .ZN(P2_U3163) );
  NAND2_X1 U9867 ( .A1(n8349), .A2(n8322), .ZN(n8324) );
  NAND2_X1 U9868 ( .A1(n8324), .A2(n8325), .ZN(n8323) );
  OAI21_X1 U9869 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(n8326) );
  NAND2_X1 U9870 ( .A1(n8326), .A2(n10126), .ZN(n8331) );
  OAI22_X1 U9871 ( .A1(n10128), .A2(n8613), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8327), .ZN(n8329) );
  NOR2_X1 U9872 ( .A1(n10131), .A2(n8811), .ZN(n8328) );
  AOI211_X1 U9873 ( .C1(n8615), .C2(n8400), .A(n8329), .B(n8328), .ZN(n8330)
         );
  OAI211_X1 U9874 ( .C1(n8889), .C2(n8403), .A(n8331), .B(n8330), .ZN(P2_U3165) );
  INV_X1 U9875 ( .A(n8332), .ZN(n8926) );
  OAI211_X1 U9876 ( .C1(n8335), .C2(n8334), .A(n8333), .B(n10126), .ZN(n8339)
         );
  NAND2_X1 U9877 ( .A1(n8409), .A2(n8421), .ZN(n8336) );
  NAND2_X1 U9878 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8484) );
  OAI211_X1 U9879 ( .C1(n8716), .C2(n10128), .A(n8336), .B(n8484), .ZN(n8337)
         );
  AOI21_X1 U9880 ( .B1(n8400), .B2(n8719), .A(n8337), .ZN(n8338) );
  OAI211_X1 U9881 ( .C1(n8926), .C2(n8403), .A(n8339), .B(n8338), .ZN(P2_U3166) );
  XNOR2_X1 U9882 ( .A(n8340), .B(n8420), .ZN(n8341) );
  XNOR2_X1 U9883 ( .A(n8342), .B(n8341), .ZN(n8348) );
  NOR2_X1 U9884 ( .A1(n8343), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8509) );
  NOR2_X1 U9885 ( .A1(n10128), .A2(n8706), .ZN(n8344) );
  AOI211_X1 U9886 ( .C1(n8409), .C2(n8853), .A(n8509), .B(n8344), .ZN(n8345)
         );
  OAI21_X1 U9887 ( .B1(n8709), .B2(n10138), .A(n8345), .ZN(n8346) );
  AOI21_X1 U9888 ( .B1(n8708), .B2(n10134), .A(n8346), .ZN(n8347) );
  OAI21_X1 U9889 ( .B1(n8348), .B2(n8383), .A(n8347), .ZN(P2_U3168) );
  INV_X1 U9890 ( .A(n8349), .ZN(n8353) );
  AOI21_X1 U9891 ( .B1(n8298), .B2(n8351), .A(n8350), .ZN(n8352) );
  OAI21_X1 U9892 ( .B1(n8353), .B2(n8352), .A(n10126), .ZN(n8357) );
  INV_X1 U9893 ( .A(n8623), .ZN(n8600) );
  AOI22_X1 U9894 ( .A1(n8408), .A2(n8600), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8354) );
  OAI21_X1 U9895 ( .B1(n8818), .B2(n10131), .A(n8354), .ZN(n8355) );
  AOI21_X1 U9896 ( .B1(n8625), .B2(n8400), .A(n8355), .ZN(n8356) );
  OAI211_X1 U9897 ( .C1(n8893), .C2(n8403), .A(n8357), .B(n8356), .ZN(P2_U3169) );
  INV_X1 U9898 ( .A(n8358), .ZN(n8362) );
  AOI21_X1 U9899 ( .B1(n8307), .B2(n8360), .A(n8359), .ZN(n8361) );
  OAI21_X1 U9900 ( .B1(n8362), .B2(n8361), .A(n10126), .ZN(n8367) );
  AOI22_X1 U9901 ( .A1(n8408), .A2(n6029), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8363) );
  OAI21_X1 U9902 ( .B1(n8689), .B2(n10131), .A(n8363), .ZN(n8364) );
  AOI21_X1 U9903 ( .B1(n8365), .B2(n8400), .A(n8364), .ZN(n8366) );
  OAI211_X1 U9904 ( .C1(n6019), .C2(n8403), .A(n8367), .B(n8366), .ZN(P2_U3173) );
  NOR2_X1 U9905 ( .A1(n8368), .A2(n4433), .ZN(n8369) );
  XNOR2_X1 U9906 ( .A(n8370), .B(n8369), .ZN(n8376) );
  AOI21_X1 U9907 ( .B1(n8408), .B2(n8729), .A(n8371), .ZN(n8373) );
  NAND2_X1 U9908 ( .A1(n8409), .A2(n8423), .ZN(n8372) );
  OAI211_X1 U9909 ( .C1(n10138), .C2(n8774), .A(n8373), .B(n8372), .ZN(n8374)
         );
  AOI21_X1 U9910 ( .B1(n8864), .B2(n10134), .A(n8374), .ZN(n8375) );
  OAI21_X1 U9911 ( .B1(n8376), .B2(n8383), .A(n8375), .ZN(P2_U3174) );
  AOI21_X1 U9912 ( .B1(n8378), .B2(n8377), .A(n4389), .ZN(n8384) );
  NAND2_X1 U9913 ( .A1(n8400), .A2(n8646), .ZN(n8380) );
  AOI22_X1 U9914 ( .A1(n8408), .A2(n8417), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8379) );
  OAI211_X1 U9915 ( .C1(n8833), .C2(n10131), .A(n8380), .B(n8379), .ZN(n8381)
         );
  AOI21_X1 U9916 ( .B1(n8817), .B2(n10134), .A(n8381), .ZN(n8382) );
  OAI21_X1 U9917 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(P2_U3175) );
  OAI21_X1 U9918 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8389) );
  NAND2_X1 U9919 ( .A1(n8389), .A2(n10126), .ZN(n8393) );
  AND2_X1 U9920 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8536) );
  AOI21_X1 U9921 ( .B1(n8408), .B2(n8419), .A(n8536), .ZN(n8390) );
  OAI21_X1 U9922 ( .B1(n10131), .B2(n8716), .A(n8390), .ZN(n8391) );
  AOI21_X1 U9923 ( .B1(n8698), .B2(n8400), .A(n8391), .ZN(n8392) );
  OAI211_X1 U9924 ( .C1(n8918), .C2(n8403), .A(n8393), .B(n8392), .ZN(P2_U3178) );
  XNOR2_X1 U9925 ( .A(n8394), .B(n8613), .ZN(n8395) );
  XNOR2_X1 U9926 ( .A(n8396), .B(n8395), .ZN(n8397) );
  NAND2_X1 U9927 ( .A1(n8397), .A2(n10126), .ZN(n8402) );
  NOR2_X1 U9928 ( .A1(n8604), .A2(n10128), .ZN(n8399) );
  INV_X1 U9929 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10088) );
  OAI22_X1 U9930 ( .A1(n10131), .A2(n8623), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10088), .ZN(n8398) );
  AOI211_X1 U9931 ( .C1(n8602), .C2(n8400), .A(n8399), .B(n8398), .ZN(n8401)
         );
  OAI211_X1 U9932 ( .C1(n8404), .C2(n8403), .A(n8402), .B(n8401), .ZN(P2_U3180) );
  OAI211_X1 U9933 ( .C1(n8407), .C2(n8406), .A(n8405), .B(n10126), .ZN(n8414)
         );
  AND2_X1 U9934 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8462) );
  AOI21_X1 U9935 ( .B1(n8408), .B2(n8853), .A(n8462), .ZN(n8411) );
  NAND2_X1 U9936 ( .A1(n8409), .A2(n8729), .ZN(n8410) );
  OAI211_X1 U9937 ( .C1(n10138), .C2(n8734), .A(n8411), .B(n8410), .ZN(n8412)
         );
  AOI21_X1 U9938 ( .B1(n8854), .B2(n10134), .A(n8412), .ZN(n8413) );
  NAND2_X1 U9939 ( .A1(n8414), .A2(n8413), .ZN(P2_U3181) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8415), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8786), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8793), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8798), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8588), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8600), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8416), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8417), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8418), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n6029), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8675), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8419), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9952 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8674), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9953 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8420), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8853), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8421), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8729), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9957 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8422), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9958 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8423), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8424), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8425), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9961 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n10122), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9962 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n10120), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8426), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9964 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8427), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8428), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8429), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9967 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8430), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8431), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6304), .S(P2_U3893), .Z(
        P2_U3492) );
  OAI21_X1 U9970 ( .B1(n8434), .B2(n8433), .A(n8432), .ZN(n8435) );
  NAND2_X1 U9971 ( .A1(n8435), .A2(n9788), .ZN(n8451) );
  OAI21_X1 U9972 ( .B1(n8438), .B2(n8437), .A(n8436), .ZN(n8439) );
  AOI22_X1 U9973 ( .A1(n9783), .A2(n8440), .B1(n8542), .B2(n8439), .ZN(n8450)
         );
  INV_X1 U9974 ( .A(n8441), .ZN(n8443) );
  NAND3_X1 U9975 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8445) );
  AOI21_X1 U9976 ( .B1(n8446), .B2(n8445), .A(n9778), .ZN(n8447) );
  AOI211_X1 U9977 ( .C1(n8555), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n8448), .B(
        n8447), .ZN(n8449) );
  NAND3_X1 U9978 ( .A1(n8451), .A2(n8450), .A3(n8449), .ZN(P2_U3188) );
  AOI21_X1 U9979 ( .B1(n8735), .B2(n8453), .A(n8470), .ZN(n8468) );
  NAND2_X1 U9980 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8454), .ZN(n8456) );
  NAND2_X1 U9981 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8457), .ZN(n8490) );
  OAI21_X1 U9982 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8457), .A(n8490), .ZN(
        n8466) );
  MUX2_X1 U9983 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8478), .Z(n8474) );
  XNOR2_X1 U9984 ( .A(n8489), .B(n8474), .ZN(n8459) );
  AOI21_X1 U9985 ( .B1(n4421), .B2(n8459), .A(n8475), .ZN(n8464) );
  NOR2_X1 U9986 ( .A1(n9768), .A2(n8460), .ZN(n8461) );
  AOI211_X1 U9987 ( .C1(n8477), .C2(n9783), .A(n8462), .B(n8461), .ZN(n8463)
         );
  OAI21_X1 U9988 ( .B1(n8464), .B2(n8534), .A(n8463), .ZN(n8465) );
  AOI21_X1 U9989 ( .B1(n8466), .B2(n8542), .A(n8465), .ZN(n8467) );
  OAI21_X1 U9990 ( .B1(n8468), .B2(n9778), .A(n8467), .ZN(P2_U3197) );
  NOR2_X1 U9991 ( .A1(n8477), .A2(n8469), .ZN(n8471) );
  NAND2_X1 U9992 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8499), .ZN(n8472) );
  OAI21_X1 U9993 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8499), .A(n8472), .ZN(
        n8473) );
  AOI21_X1 U9994 ( .B1(n4383), .B2(n8473), .A(n8498), .ZN(n8497) );
  INV_X1 U9995 ( .A(n8474), .ZN(n8476) );
  AOI21_X1 U9996 ( .B1(n8477), .B2(n8476), .A(n8475), .ZN(n8505) );
  MUX2_X1 U9997 ( .A(n8479), .B(n8851), .S(n8478), .Z(n8480) );
  NOR2_X1 U9998 ( .A1(n8480), .A2(n8502), .ZN(n8506) );
  INV_X1 U9999 ( .A(n8506), .ZN(n8481) );
  NAND2_X1 U10000 ( .A1(n8480), .A2(n8502), .ZN(n8504) );
  NAND2_X1 U10001 ( .A1(n8481), .A2(n8504), .ZN(n8482) );
  XNOR2_X1 U10002 ( .A(n8505), .B(n8482), .ZN(n8487) );
  NOR2_X1 U10003 ( .A1(n9768), .A2(n8483), .ZN(n8486) );
  OAI21_X1 U10004 ( .B1(n8559), .B2(n8499), .A(n8484), .ZN(n8485) );
  AOI211_X1 U10005 ( .C1(n8487), .C2(n9788), .A(n8486), .B(n8485), .ZN(n8496)
         );
  AOI22_X1 U10006 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8499), .B1(n8502), .B2(
        n8851), .ZN(n8493) );
  NAND2_X1 U10007 ( .A1(n8489), .A2(n8488), .ZN(n8491) );
  NAND2_X1 U10008 ( .A1(n8491), .A2(n8490), .ZN(n8492) );
  OAI21_X1 U10009 ( .B1(n8493), .B2(n8492), .A(n8501), .ZN(n8494) );
  NAND2_X1 U10010 ( .A1(n8494), .A2(n8542), .ZN(n8495) );
  OAI211_X1 U10011 ( .C1(n8497), .C2(n9778), .A(n8496), .B(n8495), .ZN(
        P2_U3198) );
  AOI21_X1 U10012 ( .B1(n8710), .B2(n8500), .A(n8518), .ZN(n8516) );
  OAI21_X1 U10013 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8503), .A(n8539), .ZN(
        n8514) );
  MUX2_X1 U10014 ( .A(n8710), .B(n8847), .S(n8478), .Z(n8525) );
  XNOR2_X1 U10015 ( .A(n8538), .B(n8525), .ZN(n8508) );
  OAI21_X1 U10016 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8507) );
  OAI21_X1 U10017 ( .B1(n8508), .B2(n8507), .A(n8523), .ZN(n8510) );
  AOI21_X1 U10018 ( .B1(n9788), .B2(n8510), .A(n8509), .ZN(n8512) );
  NAND2_X1 U10019 ( .A1(n8555), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8511) );
  OAI211_X1 U10020 ( .C1(n8559), .C2(n8538), .A(n8512), .B(n8511), .ZN(n8513)
         );
  AOI21_X1 U10021 ( .B1(n8514), .B2(n8542), .A(n8513), .ZN(n8515) );
  OAI21_X1 U10022 ( .B1(n8516), .B2(n9778), .A(n8515), .ZN(P2_U3199) );
  NOR2_X1 U10023 ( .A1(n8524), .A2(n8517), .ZN(n8519) );
  INV_X1 U10024 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8520) );
  MUX2_X1 U10025 ( .A(n8520), .B(P2_REG2_REG_18__SCAN_IN), .S(n8541), .Z(n8521) );
  INV_X1 U10026 ( .A(n8521), .ZN(n8522) );
  AOI21_X1 U10027 ( .B1(n4384), .B2(n8522), .A(n8547), .ZN(n8546) );
  MUX2_X1 U10028 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8478), .Z(n8527) );
  AND2_X1 U10029 ( .A1(n8526), .A2(n8527), .ZN(n8552) );
  INV_X1 U10030 ( .A(n8527), .ZN(n8528) );
  NAND2_X1 U10031 ( .A1(n8529), .A2(n8528), .ZN(n8551) );
  INV_X1 U10032 ( .A(n8551), .ZN(n8530) );
  INV_X1 U10033 ( .A(n8533), .ZN(n8531) );
  OAI21_X1 U10034 ( .B1(n8532), .B2(n8531), .A(n8559), .ZN(n8535) );
  NAND2_X1 U10035 ( .A1(n8538), .A2(n8537), .ZN(n8540) );
  NAND2_X1 U10036 ( .A1(n8540), .A2(n8539), .ZN(n8562) );
  XNOR2_X1 U10037 ( .A(n8541), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8561) );
  XNOR2_X1 U10038 ( .A(n8562), .B(n8561), .ZN(n8543) );
  NAND2_X1 U10039 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  OAI211_X1 U10040 ( .C1(n8546), .C2(n9778), .A(n8545), .B(n8544), .ZN(
        P2_U3200) );
  AOI21_X1 U10041 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8560), .A(n8547), .ZN(
        n8548) );
  MUX2_X1 U10042 ( .A(n5978), .B(P2_REG2_REG_19__SCAN_IN), .S(n6299), .Z(n8550) );
  XNOR2_X1 U10043 ( .A(n8548), .B(n8550), .ZN(n8567) );
  XNOR2_X1 U10044 ( .A(n6299), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8563) );
  MUX2_X1 U10045 ( .A(n8563), .B(n8550), .S(n8549), .Z(n8554) );
  OAI21_X1 U10046 ( .B1(n8552), .B2(n8560), .A(n8551), .ZN(n8553) );
  XNOR2_X1 U10047 ( .A(n8554), .B(n8553), .ZN(n8566) );
  NAND2_X1 U10048 ( .A1(n8555), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8557) );
  OAI211_X1 U10049 ( .C1(n8559), .C2(n8558), .A(n8557), .B(n8556), .ZN(n8565)
         );
  AOI22_X1 U10050 ( .A1(n8562), .A2(n8561), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8560), .ZN(n8564) );
  NAND2_X1 U10051 ( .A1(n9808), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8573) );
  INV_X1 U10052 ( .A(n8568), .ZN(n8570) );
  NOR2_X1 U10053 ( .A1(n8570), .A2(n8569), .ZN(n8876) );
  AND2_X1 U10054 ( .A1(n4348), .A2(n9804), .ZN(n8572) );
  OAI21_X1 U10055 ( .B1(n8876), .B2(n8572), .A(n9807), .ZN(n8574) );
  OAI211_X1 U10056 ( .C1(n8878), .C2(n8721), .A(n8573), .B(n8574), .ZN(
        P2_U3202) );
  NAND2_X1 U10057 ( .A1(n9808), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8575) );
  OAI211_X1 U10058 ( .C1(n8785), .C2(n8721), .A(n8575), .B(n8574), .ZN(
        P2_U3203) );
  INV_X1 U10059 ( .A(n8576), .ZN(n8577) );
  INV_X1 U10060 ( .A(n8578), .ZN(n8579) );
  AOI22_X1 U10061 ( .A1(n9808), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9804), .B2(
        n8579), .ZN(n8580) );
  OAI21_X1 U10062 ( .B1(n8581), .B2(n8660), .A(n8580), .ZN(n8585) );
  XNOR2_X1 U10063 ( .A(n8583), .B(n8582), .ZN(n8789) );
  NOR2_X1 U10064 ( .A1(n8789), .A2(n8740), .ZN(n8584) );
  AOI211_X1 U10065 ( .C1(n9802), .C2(n8787), .A(n8585), .B(n8584), .ZN(n8586)
         );
  OAI21_X1 U10066 ( .B1(n8792), .B2(n9808), .A(n8586), .ZN(P2_U3205) );
  XNOR2_X1 U10067 ( .A(n8587), .B(n8594), .ZN(n8589) );
  AOI22_X1 U10068 ( .A1(n8589), .A2(n8726), .B1(n8728), .B2(n8588), .ZN(n8796)
         );
  AOI22_X1 U10069 ( .A1(n9808), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n9804), .B2(
        n8590), .ZN(n8591) );
  OAI21_X1 U10070 ( .B1(n8592), .B2(n8660), .A(n8591), .ZN(n8596) );
  XOR2_X1 U10071 ( .A(n8594), .B(n8593), .Z(n8797) );
  NOR2_X1 U10072 ( .A1(n8797), .A2(n8740), .ZN(n8595) );
  AOI211_X1 U10073 ( .C1(n9802), .C2(n8794), .A(n8596), .B(n8595), .ZN(n8597)
         );
  OAI21_X1 U10074 ( .B1(n8796), .B2(n9808), .A(n8597), .ZN(P2_U3206) );
  XNOR2_X1 U10075 ( .A(n8599), .B(n8598), .ZN(n8601) );
  AOI22_X1 U10076 ( .A1(n8601), .A2(n8726), .B1(n8728), .B2(n8600), .ZN(n8801)
         );
  AOI22_X1 U10077 ( .A1(n9808), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9804), .B2(
        n8602), .ZN(n8603) );
  OAI21_X1 U10078 ( .B1(n8604), .B2(n8660), .A(n8603), .ZN(n8608) );
  XNOR2_X1 U10079 ( .A(n8606), .B(n8605), .ZN(n8802) );
  NOR2_X1 U10080 ( .A1(n8802), .A2(n8740), .ZN(n8607) );
  AOI211_X1 U10081 ( .C1(n9802), .C2(n8799), .A(n8608), .B(n8607), .ZN(n8609)
         );
  OAI21_X1 U10082 ( .B1(n8801), .B2(n9808), .A(n8609), .ZN(P2_U3207) );
  XNOR2_X1 U10083 ( .A(n8611), .B(n8610), .ZN(n8612) );
  OAI222_X1 U10084 ( .A1(n9813), .A2(n8613), .B1(n9794), .B2(n8811), .C1(n9797), .C2(n8612), .ZN(n8803) );
  AOI21_X1 U10085 ( .B1(n8768), .B2(n8614), .A(n8803), .ZN(n8620) );
  AOI22_X1 U10086 ( .A1(n9808), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9804), .B2(
        n8615), .ZN(n8619) );
  XNOR2_X1 U10087 ( .A(n8617), .B(n8616), .ZN(n8804) );
  NAND2_X1 U10088 ( .A1(n8804), .A2(n8777), .ZN(n8618) );
  OAI211_X1 U10089 ( .C1(n8620), .C2(n9808), .A(n8619), .B(n8618), .ZN(
        P2_U3208) );
  NOR2_X1 U10090 ( .A1(n8893), .A2(n8752), .ZN(n8624) );
  XNOR2_X1 U10091 ( .A(n8621), .B(n8629), .ZN(n8622) );
  OAI222_X1 U10092 ( .A1(n9794), .A2(n8818), .B1(n9813), .B2(n8623), .C1(n8622), .C2(n9797), .ZN(n8807) );
  AOI211_X1 U10093 ( .C1(n9804), .C2(n8625), .A(n8624), .B(n8807), .ZN(n8631)
         );
  NOR2_X1 U10094 ( .A1(n8627), .A2(n8626), .ZN(n8628) );
  XOR2_X1 U10095 ( .A(n8629), .B(n8628), .Z(n8808) );
  AOI22_X1 U10096 ( .A1(n8808), .A2(n8777), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9808), .ZN(n8630) );
  OAI21_X1 U10097 ( .B1(n8631), .B2(n9808), .A(n8630), .ZN(P2_U3209) );
  XOR2_X1 U10098 ( .A(n8634), .B(n8632), .Z(n8812) );
  XOR2_X1 U10099 ( .A(n8634), .B(n8633), .Z(n8635) );
  OAI22_X1 U10100 ( .A1(n8635), .A2(n9797), .B1(n8824), .B2(n9794), .ZN(n8814)
         );
  NAND2_X1 U10101 ( .A1(n8814), .A2(n9807), .ZN(n8641) );
  AOI22_X1 U10102 ( .A1(n9808), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9804), .B2(
        n8636), .ZN(n8637) );
  OAI21_X1 U10103 ( .B1(n8811), .B2(n8660), .A(n8637), .ZN(n8638) );
  AOI21_X1 U10104 ( .B1(n8639), .B2(n9802), .A(n8638), .ZN(n8640) );
  OAI211_X1 U10105 ( .C1(n8740), .C2(n8812), .A(n8641), .B(n8640), .ZN(
        P2_U3210) );
  XNOR2_X1 U10106 ( .A(n8642), .B(n8643), .ZN(n8819) );
  XNOR2_X1 U10107 ( .A(n8644), .B(n8643), .ZN(n8645) );
  OAI22_X1 U10108 ( .A1(n8645), .A2(n9797), .B1(n8833), .B2(n9794), .ZN(n8821)
         );
  NAND2_X1 U10109 ( .A1(n8821), .A2(n9807), .ZN(n8650) );
  AOI22_X1 U10110 ( .A1(n9808), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9804), .B2(
        n8646), .ZN(n8647) );
  OAI21_X1 U10111 ( .B1(n8818), .B2(n8660), .A(n8647), .ZN(n8648) );
  AOI21_X1 U10112 ( .B1(n8817), .B2(n9802), .A(n8648), .ZN(n8649) );
  OAI211_X1 U10113 ( .C1(n8740), .C2(n8819), .A(n8650), .B(n8649), .ZN(
        P2_U3211) );
  NAND2_X1 U10114 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  XNOR2_X1 U10115 ( .A(n8653), .B(n8654), .ZN(n8825) );
  XOR2_X1 U10116 ( .A(n8655), .B(n8654), .Z(n8657) );
  OAI22_X1 U10117 ( .A1(n8657), .A2(n9797), .B1(n8656), .B2(n9794), .ZN(n8827)
         );
  NAND2_X1 U10118 ( .A1(n8827), .A2(n9807), .ZN(n8664) );
  AOI22_X1 U10119 ( .A1(n9808), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9804), .B2(
        n8658), .ZN(n8659) );
  OAI21_X1 U10120 ( .B1(n8824), .B2(n8660), .A(n8659), .ZN(n8661) );
  AOI21_X1 U10121 ( .B1(n8662), .B2(n9802), .A(n8661), .ZN(n8663) );
  OAI211_X1 U10122 ( .C1(n8740), .C2(n8825), .A(n8664), .B(n8663), .ZN(
        P2_U3212) );
  XOR2_X1 U10123 ( .A(n8668), .B(n8665), .Z(n8838) );
  INV_X1 U10124 ( .A(n8838), .ZN(n8682) );
  NAND2_X1 U10125 ( .A1(n8684), .A2(n8666), .ZN(n8670) );
  AND2_X1 U10126 ( .A1(n8670), .A2(n8667), .ZN(n8673) );
  INV_X1 U10127 ( .A(n8668), .ZN(n8672) );
  NAND2_X1 U10128 ( .A1(n8670), .A2(n8669), .ZN(n8671) );
  OAI211_X1 U10129 ( .C1(n8673), .C2(n8672), .A(n8726), .B(n8671), .ZN(n8677)
         );
  AOI22_X1 U10130 ( .A1(n8675), .A2(n9842), .B1(n8728), .B2(n8674), .ZN(n8676)
         );
  NAND2_X1 U10131 ( .A1(n8677), .A2(n8676), .ZN(n8837) );
  AOI22_X1 U10132 ( .A1(n9808), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9804), .B2(
        n8678), .ZN(n8679) );
  OAI21_X1 U10133 ( .B1(n8914), .B2(n8721), .A(n8679), .ZN(n8680) );
  AOI21_X1 U10134 ( .B1(n8837), .B2(n9807), .A(n8680), .ZN(n8681) );
  OAI21_X1 U10135 ( .B1(n8740), .B2(n8682), .A(n8681), .ZN(P2_U3214) );
  NAND2_X1 U10136 ( .A1(n8684), .A2(n8683), .ZN(n8703) );
  NAND2_X1 U10137 ( .A1(n8703), .A2(n8707), .ZN(n8686) );
  NAND2_X1 U10138 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  XNOR2_X1 U10139 ( .A(n8687), .B(n8697), .ZN(n8688) );
  OAI222_X1 U10140 ( .A1(n9794), .A2(n8716), .B1(n9813), .B2(n8689), .C1(n8688), .C2(n9797), .ZN(n8841) );
  INV_X1 U10141 ( .A(n8841), .ZN(n8702) );
  OR2_X1 U10142 ( .A1(n8690), .A2(n8691), .ZN(n8694) );
  NAND2_X1 U10143 ( .A1(n8694), .A2(n8692), .ZN(n8696) );
  AND2_X1 U10144 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  AOI21_X1 U10145 ( .B1(n8697), .B2(n8696), .A(n8695), .ZN(n8842) );
  AOI22_X1 U10146 ( .A1(n9808), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9804), .B2(
        n8698), .ZN(n8699) );
  OAI21_X1 U10147 ( .B1(n8918), .B2(n8721), .A(n8699), .ZN(n8700) );
  AOI21_X1 U10148 ( .B1(n8842), .B2(n8777), .A(n8700), .ZN(n8701) );
  OAI21_X1 U10149 ( .B1(n8702), .B2(n9808), .A(n8701), .ZN(P2_U3215) );
  XNOR2_X1 U10150 ( .A(n8703), .B(n8707), .ZN(n8704) );
  OAI222_X1 U10151 ( .A1(n9813), .A2(n8706), .B1(n9794), .B2(n8705), .C1(n8704), .C2(n9797), .ZN(n8845) );
  INV_X1 U10152 ( .A(n8845), .ZN(n8714) );
  XNOR2_X1 U10153 ( .A(n8690), .B(n8707), .ZN(n8846) );
  INV_X1 U10154 ( .A(n8708), .ZN(n8922) );
  NOR2_X1 U10155 ( .A1(n8922), .A2(n8721), .ZN(n8712) );
  OAI22_X1 U10156 ( .A1(n9807), .A2(n8710), .B1(n8709), .B2(n8773), .ZN(n8711)
         );
  AOI211_X1 U10157 ( .C1(n8846), .C2(n8777), .A(n8712), .B(n8711), .ZN(n8713)
         );
  OAI21_X1 U10158 ( .B1(n8714), .B2(n9808), .A(n8713), .ZN(P2_U3216) );
  XNOR2_X1 U10159 ( .A(n7897), .B(n8717), .ZN(n8715) );
  OAI222_X1 U10160 ( .A1(n9794), .A2(n8745), .B1(n9813), .B2(n8716), .C1(n8715), .C2(n9797), .ZN(n8849) );
  INV_X1 U10161 ( .A(n8849), .ZN(n8724) );
  XNOR2_X1 U10162 ( .A(n8718), .B(n8717), .ZN(n8850) );
  AOI22_X1 U10163 ( .A1(n9808), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9804), .B2(
        n8719), .ZN(n8720) );
  OAI21_X1 U10164 ( .B1(n8926), .B2(n8721), .A(n8720), .ZN(n8722) );
  AOI21_X1 U10165 ( .B1(n8850), .B2(n8777), .A(n8722), .ZN(n8723) );
  OAI21_X1 U10166 ( .B1(n8724), .B2(n9808), .A(n8723), .ZN(P2_U3217) );
  XNOR2_X1 U10167 ( .A(n8725), .B(n8732), .ZN(n8727) );
  NAND2_X1 U10168 ( .A1(n8727), .A2(n8726), .ZN(n8731) );
  NAND2_X1 U10169 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U10170 ( .A1(n8731), .A2(n8730), .ZN(n8858) );
  XNOR2_X1 U10171 ( .A(n8733), .B(n8732), .ZN(n8856) );
  OAI22_X1 U10172 ( .A1(n9807), .A2(n8735), .B1(n8734), .B2(n8773), .ZN(n8736)
         );
  AOI21_X1 U10173 ( .B1(n8737), .B2(n8853), .A(n8736), .ZN(n8739) );
  NAND2_X1 U10174 ( .A1(n8854), .A2(n9802), .ZN(n8738) );
  OAI211_X1 U10175 ( .C1(n8856), .C2(n8740), .A(n8739), .B(n8738), .ZN(n8741)
         );
  AOI21_X1 U10176 ( .B1(n8858), .B2(n9807), .A(n8741), .ZN(n8742) );
  INV_X1 U10177 ( .A(n8742), .ZN(P2_U3218) );
  AOI21_X1 U10178 ( .B1(n8744), .B2(n8743), .A(n9797), .ZN(n8749) );
  OAI22_X1 U10179 ( .A1(n8746), .A2(n9794), .B1(n8745), .B2(n9813), .ZN(n8747)
         );
  AOI21_X1 U10180 ( .B1(n8749), .B2(n8748), .A(n8747), .ZN(n8861) );
  INV_X1 U10181 ( .A(n8861), .ZN(n8754) );
  INV_X1 U10182 ( .A(n8750), .ZN(n8931) );
  OAI22_X1 U10183 ( .A1(n8931), .A2(n8752), .B1(n8751), .B2(n8773), .ZN(n8753)
         );
  OAI21_X1 U10184 ( .B1(n8754), .B2(n8753), .A(n9807), .ZN(n8761) );
  OR2_X1 U10185 ( .A1(n7798), .A2(n8755), .ZN(n8757) );
  NAND2_X1 U10186 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  XNOR2_X1 U10187 ( .A(n8759), .B(n8758), .ZN(n8859) );
  AOI22_X1 U10188 ( .A1(n8859), .A2(n8777), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9808), .ZN(n8760) );
  NAND2_X1 U10189 ( .A1(n8761), .A2(n8760), .ZN(P2_U3219) );
  INV_X1 U10190 ( .A(n8762), .ZN(n8763) );
  AOI21_X1 U10191 ( .B1(n8772), .B2(n8764), .A(n8763), .ZN(n8765) );
  OAI222_X1 U10192 ( .A1(n9813), .A2(n8767), .B1(n9794), .B2(n8766), .C1(n9797), .C2(n8765), .ZN(n8865) );
  AOI21_X1 U10193 ( .B1(n8768), .B2(n8864), .A(n8865), .ZN(n8779) );
  NAND2_X1 U10194 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  XOR2_X1 U10195 ( .A(n8772), .B(n8771), .Z(n8866) );
  OAI22_X1 U10196 ( .A1(n9807), .A2(n8775), .B1(n8774), .B2(n8773), .ZN(n8776)
         );
  AOI21_X1 U10197 ( .B1(n8866), .B2(n8777), .A(n8776), .ZN(n8778) );
  OAI21_X1 U10198 ( .B1(n8779), .B2(n9808), .A(n8778), .ZN(P2_U3220) );
  INV_X1 U10199 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U10200 ( .A1(n8780), .A2(n8835), .ZN(n8781) );
  NAND2_X1 U10201 ( .A1(n9897), .A2(n8876), .ZN(n8783) );
  OAI211_X1 U10202 ( .C1(n9897), .C2(n8782), .A(n8781), .B(n8783), .ZN(
        P2_U3490) );
  NAND2_X1 U10203 ( .A1(n9894), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8784) );
  OAI211_X1 U10204 ( .C1(n8785), .C2(n8869), .A(n8784), .B(n8783), .ZN(
        P2_U3489) );
  AOI22_X1 U10205 ( .A1(n8787), .A2(n9877), .B1(n9842), .B2(n8786), .ZN(n8788)
         );
  OAI21_X1 U10206 ( .B1(n8789), .B2(n9872), .A(n8788), .ZN(n8790) );
  INV_X1 U10207 ( .A(n8790), .ZN(n8791) );
  AOI22_X1 U10208 ( .A1(n8794), .A2(n9877), .B1(n9842), .B2(n8793), .ZN(n8795)
         );
  OAI211_X1 U10209 ( .C1(n9872), .C2(n8797), .A(n8796), .B(n8795), .ZN(n8884)
         );
  MUX2_X1 U10210 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8884), .S(n9897), .Z(
        P2_U3486) );
  AOI22_X1 U10211 ( .A1(n8799), .A2(n9877), .B1(n9842), .B2(n8798), .ZN(n8800)
         );
  OAI211_X1 U10212 ( .C1(n9872), .C2(n8802), .A(n8801), .B(n8800), .ZN(n8885)
         );
  MUX2_X1 U10213 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8885), .S(n9897), .Z(
        P2_U3485) );
  INV_X1 U10214 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8805) );
  AOI21_X1 U10215 ( .B1(n9869), .B2(n8804), .A(n8803), .ZN(n8886) );
  MUX2_X1 U10216 ( .A(n8805), .B(n8886), .S(n9897), .Z(n8806) );
  OAI21_X1 U10217 ( .B1(n8889), .B2(n8869), .A(n8806), .ZN(P2_U3484) );
  INV_X1 U10218 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8809) );
  AOI21_X1 U10219 ( .B1(n8808), .B2(n9869), .A(n8807), .ZN(n8890) );
  MUX2_X1 U10220 ( .A(n8809), .B(n8890), .S(n9897), .Z(n8810) );
  OAI21_X1 U10221 ( .B1(n8893), .B2(n8869), .A(n8810), .ZN(P2_U3483) );
  INV_X1 U10222 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8815) );
  OAI22_X1 U10223 ( .A1(n8812), .A2(n9872), .B1(n8811), .B2(n9813), .ZN(n8813)
         );
  NOR2_X1 U10224 ( .A1(n8814), .A2(n8813), .ZN(n8894) );
  MUX2_X1 U10225 ( .A(n8815), .B(n8894), .S(n9897), .Z(n8816) );
  OAI21_X1 U10226 ( .B1(n8897), .B2(n8869), .A(n8816), .ZN(P2_U3482) );
  INV_X1 U10227 ( .A(n8817), .ZN(n8901) );
  INV_X1 U10228 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8822) );
  OAI22_X1 U10229 ( .A1(n8819), .A2(n9872), .B1(n8818), .B2(n9813), .ZN(n8820)
         );
  NOR2_X1 U10230 ( .A1(n8821), .A2(n8820), .ZN(n8898) );
  MUX2_X1 U10231 ( .A(n8822), .B(n8898), .S(n9897), .Z(n8823) );
  OAI21_X1 U10232 ( .B1(n8901), .B2(n8869), .A(n8823), .ZN(P2_U3481) );
  INV_X1 U10233 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8828) );
  OAI22_X1 U10234 ( .A1(n8825), .A2(n9872), .B1(n8824), .B2(n9813), .ZN(n8826)
         );
  NOR2_X1 U10235 ( .A1(n8827), .A2(n8826), .ZN(n8902) );
  MUX2_X1 U10236 ( .A(n8828), .B(n8902), .S(n9897), .Z(n8829) );
  OAI21_X1 U10237 ( .B1(n8905), .B2(n8869), .A(n8829), .ZN(P2_U3480) );
  NAND2_X1 U10238 ( .A1(n8830), .A2(n9869), .ZN(n8831) );
  OAI211_X1 U10239 ( .C1(n8833), .C2(n9813), .A(n8832), .B(n8831), .ZN(n8906)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8906), .S(n9897), .Z(n8834) );
  AOI21_X1 U10241 ( .B1(n8835), .B2(n8908), .A(n8834), .ZN(n8836) );
  INV_X1 U10242 ( .A(n8836), .ZN(P2_U3479) );
  AOI21_X1 U10243 ( .B1(n9869), .B2(n8838), .A(n8837), .ZN(n8911) );
  MUX2_X1 U10244 ( .A(n8839), .B(n8911), .S(n9897), .Z(n8840) );
  OAI21_X1 U10245 ( .B1(n8914), .B2(n8869), .A(n8840), .ZN(P2_U3478) );
  INV_X1 U10246 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8843) );
  AOI21_X1 U10247 ( .B1(n8842), .B2(n9869), .A(n8841), .ZN(n8915) );
  MUX2_X1 U10248 ( .A(n8843), .B(n8915), .S(n9897), .Z(n8844) );
  OAI21_X1 U10249 ( .B1(n8918), .B2(n8869), .A(n8844), .ZN(P2_U3477) );
  AOI21_X1 U10250 ( .B1(n9869), .B2(n8846), .A(n8845), .ZN(n8919) );
  MUX2_X1 U10251 ( .A(n8847), .B(n8919), .S(n9897), .Z(n8848) );
  OAI21_X1 U10252 ( .B1(n8922), .B2(n8869), .A(n8848), .ZN(P2_U3476) );
  AOI21_X1 U10253 ( .B1(n9869), .B2(n8850), .A(n8849), .ZN(n8923) );
  MUX2_X1 U10254 ( .A(n8851), .B(n8923), .S(n9897), .Z(n8852) );
  OAI21_X1 U10255 ( .B1(n8926), .B2(n8869), .A(n8852), .ZN(P2_U3475) );
  AOI22_X1 U10256 ( .A1(n8854), .A2(n9877), .B1(n9842), .B2(n8853), .ZN(n8855)
         );
  OAI21_X1 U10257 ( .B1(n8856), .B2(n9872), .A(n8855), .ZN(n8857) );
  MUX2_X1 U10258 ( .A(n8927), .B(P2_REG1_REG_15__SCAN_IN), .S(n9894), .Z(
        P2_U3474) );
  NAND2_X1 U10259 ( .A1(n8859), .A2(n9869), .ZN(n8860) );
  AND2_X1 U10260 ( .A1(n8861), .A2(n8860), .ZN(n8928) );
  MUX2_X1 U10261 ( .A(n8862), .B(n8928), .S(n9897), .Z(n8863) );
  OAI21_X1 U10262 ( .B1(n8931), .B2(n8869), .A(n8863), .ZN(P2_U3473) );
  INV_X1 U10263 ( .A(n8864), .ZN(n8936) );
  AOI21_X1 U10264 ( .B1(n9869), .B2(n8866), .A(n8865), .ZN(n8932) );
  MUX2_X1 U10265 ( .A(n8867), .B(n8932), .S(n9897), .Z(n8868) );
  OAI21_X1 U10266 ( .B1(n8936), .B2(n8869), .A(n8868), .ZN(P2_U3472) );
  NAND2_X1 U10267 ( .A1(n9872), .A2(n9797), .ZN(n8871) );
  NAND2_X1 U10268 ( .A1(n8871), .A2(n8870), .ZN(n8874) );
  AOI22_X1 U10269 ( .A1(n6304), .A2(n9842), .B1(n8872), .B2(n9877), .ZN(n8873)
         );
  AND2_X1 U10270 ( .A1(n8874), .A2(n8873), .ZN(n9810) );
  INV_X1 U10271 ( .A(n9810), .ZN(n8875) );
  MUX2_X1 U10272 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8875), .S(n9897), .Z(
        P2_U3459) );
  NAND2_X1 U10273 ( .A1(n9878), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U10274 ( .A1(n9880), .A2(n8876), .ZN(n8880) );
  OAI211_X1 U10275 ( .C1(n8878), .C2(n8935), .A(n8877), .B(n8880), .ZN(
        P2_U3458) );
  INV_X1 U10276 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8882) );
  INV_X1 U10277 ( .A(n8935), .ZN(n8909) );
  NAND2_X1 U10278 ( .A1(n8879), .A2(n8909), .ZN(n8881) );
  OAI211_X1 U10279 ( .C1(n8882), .C2(n9880), .A(n8881), .B(n8880), .ZN(
        P2_U3457) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8883), .S(n9880), .Z(
        P2_U3455) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8884), .S(n9880), .Z(
        P2_U3454) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8885), .S(n9880), .Z(
        P2_U3453) );
  INV_X1 U10283 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8887) );
  MUX2_X1 U10284 ( .A(n8887), .B(n8886), .S(n9880), .Z(n8888) );
  OAI21_X1 U10285 ( .B1(n8889), .B2(n8935), .A(n8888), .ZN(P2_U3452) );
  INV_X1 U10286 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8891) );
  MUX2_X1 U10287 ( .A(n8891), .B(n8890), .S(n9880), .Z(n8892) );
  OAI21_X1 U10288 ( .B1(n8893), .B2(n8935), .A(n8892), .ZN(P2_U3451) );
  INV_X1 U10289 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10290 ( .A(n8895), .B(n8894), .S(n9880), .Z(n8896) );
  OAI21_X1 U10291 ( .B1(n8897), .B2(n8935), .A(n8896), .ZN(P2_U3450) );
  MUX2_X1 U10292 ( .A(n8899), .B(n8898), .S(n9880), .Z(n8900) );
  OAI21_X1 U10293 ( .B1(n8901), .B2(n8935), .A(n8900), .ZN(P2_U3449) );
  INV_X1 U10294 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8903) );
  MUX2_X1 U10295 ( .A(n8903), .B(n8902), .S(n9880), .Z(n8904) );
  OAI21_X1 U10296 ( .B1(n8905), .B2(n8935), .A(n8904), .ZN(P2_U3448) );
  MUX2_X1 U10297 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8906), .S(n9880), .Z(n8907) );
  AOI21_X1 U10298 ( .B1(n8909), .B2(n8908), .A(n8907), .ZN(n8910) );
  INV_X1 U10299 ( .A(n8910), .ZN(P2_U3447) );
  INV_X1 U10300 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8912) );
  MUX2_X1 U10301 ( .A(n8912), .B(n8911), .S(n9880), .Z(n8913) );
  OAI21_X1 U10302 ( .B1(n8914), .B2(n8935), .A(n8913), .ZN(P2_U3446) );
  INV_X1 U10303 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8916) );
  MUX2_X1 U10304 ( .A(n8916), .B(n8915), .S(n9880), .Z(n8917) );
  OAI21_X1 U10305 ( .B1(n8918), .B2(n8935), .A(n8917), .ZN(P2_U3444) );
  INV_X1 U10306 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U10307 ( .A(n8920), .B(n8919), .S(n9880), .Z(n8921) );
  OAI21_X1 U10308 ( .B1(n8922), .B2(n8935), .A(n8921), .ZN(P2_U3441) );
  INV_X1 U10309 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8924) );
  MUX2_X1 U10310 ( .A(n8924), .B(n8923), .S(n9880), .Z(n8925) );
  OAI21_X1 U10311 ( .B1(n8926), .B2(n8935), .A(n8925), .ZN(P2_U3438) );
  MUX2_X1 U10312 ( .A(n8927), .B(P2_REG0_REG_15__SCAN_IN), .S(n9878), .Z(
        P2_U3435) );
  INV_X1 U10313 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8929) );
  MUX2_X1 U10314 ( .A(n8929), .B(n8928), .S(n9880), .Z(n8930) );
  OAI21_X1 U10315 ( .B1(n8931), .B2(n8935), .A(n8930), .ZN(P2_U3432) );
  INV_X1 U10316 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8933) );
  MUX2_X1 U10317 ( .A(n8933), .B(n8932), .S(n9880), .Z(n8934) );
  OAI21_X1 U10318 ( .B1(n8936), .B2(n8935), .A(n8934), .ZN(P2_U3429) );
  OAI222_X1 U10319 ( .A1(n8277), .A2(n8940), .B1(P2_U3151), .B2(n8939), .C1(
        n8938), .C2(n8937), .ZN(P2_U3266) );
  NAND2_X1 U10320 ( .A1(n8942), .A2(n8941), .ZN(n8944) );
  OAI211_X1 U10321 ( .C1(n8277), .C2(n8945), .A(n8944), .B(n8943), .ZN(
        P2_U3267) );
  MUX2_X1 U10322 ( .A(n8946), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10323 ( .A(n8948), .ZN(n8949) );
  NOR2_X1 U10324 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  XNOR2_X1 U10325 ( .A(n8947), .B(n8951), .ZN(n8957) );
  AND2_X1 U10326 ( .A1(n9112), .A2(n9070), .ZN(n8952) );
  AOI21_X1 U10327 ( .B1(n9110), .B2(n9069), .A(n8952), .ZN(n9337) );
  OAI22_X1 U10328 ( .A1(n9337), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8953), .ZN(n8955) );
  NOR2_X1 U10329 ( .A1(n9344), .A2(n9105), .ZN(n8954) );
  AOI211_X1 U10330 ( .C1(n9341), .C2(n9101), .A(n8955), .B(n8954), .ZN(n8956)
         );
  OAI21_X1 U10331 ( .B1(n8957), .B2(n9075), .A(n8956), .ZN(P1_U3216) );
  INV_X1 U10332 ( .A(n8958), .ZN(n8963) );
  OAI21_X1 U10333 ( .B1(n8960), .B2(n8962), .A(n8959), .ZN(n8961) );
  OAI21_X1 U10334 ( .B1(n8963), .B2(n8962), .A(n8961), .ZN(n8964) );
  NAND2_X1 U10335 ( .A1(n8964), .A2(n9095), .ZN(n8969) );
  INV_X1 U10336 ( .A(n8965), .ZN(n9115) );
  AOI22_X1 U10337 ( .A1(n9113), .A2(n9069), .B1(n9115), .B2(n9070), .ZN(n9401)
         );
  OAI22_X1 U10338 ( .A1(n9401), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8966), .ZN(n8967) );
  AOI21_X1 U10339 ( .B1(n9406), .B2(n9101), .A(n8967), .ZN(n8968) );
  OAI211_X1 U10340 ( .C1(n9409), .C2(n9105), .A(n8969), .B(n8968), .ZN(
        P1_U3219) );
  INV_X1 U10341 ( .A(n8984), .ZN(n8983) );
  NAND2_X1 U10342 ( .A1(n9258), .A2(n8970), .ZN(n8972) );
  NAND2_X1 U10343 ( .A1(n9108), .A2(n8975), .ZN(n8971) );
  NAND2_X1 U10344 ( .A1(n8972), .A2(n8971), .ZN(n8974) );
  XNOR2_X1 U10345 ( .A(n8974), .B(n8973), .ZN(n8980) );
  NAND2_X1 U10346 ( .A1(n9258), .A2(n8975), .ZN(n8976) );
  OAI21_X1 U10347 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8979) );
  XNOR2_X1 U10348 ( .A(n8980), .B(n8979), .ZN(n8992) );
  INV_X1 U10349 ( .A(n8992), .ZN(n8982) );
  NAND3_X1 U10350 ( .A1(n8984), .A2(n9095), .A3(n8992), .ZN(n8995) );
  OR2_X1 U10351 ( .A1(n9081), .A2(n9082), .ZN(n8987) );
  OR2_X1 U10352 ( .A1(n8985), .A2(n9080), .ZN(n8986) );
  AND2_X1 U10353 ( .A1(n8987), .A2(n8986), .ZN(n9254) );
  INV_X1 U10354 ( .A(n8988), .ZN(n9259) );
  AOI22_X1 U10355 ( .A1(n9259), .A2(n9101), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8989) );
  OAI21_X1 U10356 ( .B1(n9254), .B2(n9098), .A(n8989), .ZN(n8990) );
  AOI21_X1 U10357 ( .B1(n9258), .B2(n9088), .A(n8990), .ZN(n8994) );
  NAND3_X1 U10358 ( .A1(n8992), .A2(n8991), .A3(n9095), .ZN(n8993) );
  NAND4_X1 U10359 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(
        P1_U3220) );
  XOR2_X1 U10360 ( .A(n8998), .B(n8997), .Z(n9003) );
  AOI22_X1 U10361 ( .A1(n9112), .A2(n9069), .B1(n9113), .B2(n9070), .ZN(n9369)
         );
  OAI22_X1 U10362 ( .A1(n9369), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8999), .ZN(n9001) );
  NOR2_X1 U10363 ( .A1(n9575), .A2(n9105), .ZN(n9000) );
  AOI211_X1 U10364 ( .C1(n9373), .C2(n9101), .A(n9001), .B(n9000), .ZN(n9002)
         );
  OAI21_X1 U10365 ( .B1(n9003), .B2(n9075), .A(n9002), .ZN(P1_U3223) );
  OAI21_X1 U10366 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9007) );
  NAND2_X1 U10367 ( .A1(n9007), .A2(n9095), .ZN(n9014) );
  AND2_X1 U10368 ( .A1(n9110), .A2(n9070), .ZN(n9008) );
  AOI21_X1 U10369 ( .B1(n9109), .B2(n9069), .A(n9008), .ZN(n9306) );
  INV_X1 U10370 ( .A(n9306), .ZN(n9012) );
  INV_X1 U10371 ( .A(n9311), .ZN(n9010) );
  OAI22_X1 U10372 ( .A1(n9010), .A2(n9061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9009), .ZN(n9011) );
  AOI21_X1 U10373 ( .B1(n9012), .B2(n9059), .A(n9011), .ZN(n9013) );
  OAI211_X1 U10374 ( .C1(n9566), .C2(n9105), .A(n9014), .B(n9013), .ZN(
        P1_U3225) );
  XOR2_X1 U10375 ( .A(n9016), .B(n9015), .Z(n9024) );
  NAND2_X1 U10376 ( .A1(n9101), .A2(n9017), .ZN(n9019) );
  OAI211_X1 U10377 ( .C1(n9020), .C2(n9098), .A(n9019), .B(n9018), .ZN(n9021)
         );
  AOI21_X1 U10378 ( .B1(n9022), .B2(n9088), .A(n9021), .ZN(n9023) );
  OAI21_X1 U10379 ( .B1(n9024), .B2(n9075), .A(n9023), .ZN(P1_U3226) );
  XOR2_X1 U10380 ( .A(n9026), .B(n9025), .Z(n9034) );
  INV_X1 U10381 ( .A(n9027), .ZN(n9031) );
  NAND2_X1 U10382 ( .A1(n9028), .A2(n9059), .ZN(n9030) );
  OAI211_X1 U10383 ( .C1(n9061), .C2(n9031), .A(n9030), .B(n9029), .ZN(n9032)
         );
  AOI21_X1 U10384 ( .B1(n9521), .B2(n9088), .A(n9032), .ZN(n9033) );
  OAI21_X1 U10385 ( .B1(n9034), .B2(n9075), .A(n9033), .ZN(P1_U3228) );
  OAI21_X1 U10386 ( .B1(n9037), .B2(n9036), .A(n9035), .ZN(n9038) );
  NAND2_X1 U10387 ( .A1(n9038), .A2(n9095), .ZN(n9045) );
  OR2_X1 U10388 ( .A1(n9083), .A2(n9080), .ZN(n9040) );
  NAND2_X1 U10389 ( .A1(n9111), .A2(n9070), .ZN(n9039) );
  AND2_X1 U10390 ( .A1(n9040), .A2(n9039), .ZN(n9321) );
  INV_X1 U10391 ( .A(n9321), .ZN(n9043) );
  OAI22_X1 U10392 ( .A1(n9325), .A2(n9061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9041), .ZN(n9042) );
  AOI21_X1 U10393 ( .B1(n9043), .B2(n9059), .A(n9042), .ZN(n9044) );
  OAI211_X1 U10394 ( .C1(n9329), .C2(n9105), .A(n9045), .B(n9044), .ZN(
        P1_U3229) );
  AOI21_X1 U10395 ( .B1(n9048), .B2(n9047), .A(n9046), .ZN(n9053) );
  OAI22_X1 U10396 ( .A1(n9057), .A2(n9080), .B1(n9049), .B2(n9082), .ZN(n9390)
         );
  AOI22_X1 U10397 ( .A1(n9390), .A2(n9059), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9050) );
  OAI21_X1 U10398 ( .B1(n9061), .B2(n9383), .A(n9050), .ZN(n9051) );
  AOI21_X1 U10399 ( .B1(n9505), .B2(n9088), .A(n9051), .ZN(n9052) );
  OAI21_X1 U10400 ( .B1(n9053), .B2(n9075), .A(n9052), .ZN(P1_U3233) );
  AOI21_X1 U10401 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9064) );
  OAI22_X1 U10402 ( .A1(n9058), .A2(n9080), .B1(n9057), .B2(n9082), .ZN(n9358)
         );
  AOI22_X1 U10403 ( .A1(n9358), .A2(n9059), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9060) );
  OAI21_X1 U10404 ( .B1(n9061), .B2(n9351), .A(n9060), .ZN(n9062) );
  AOI21_X1 U10405 ( .B1(n9349), .B2(n9088), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10406 ( .B1(n9064), .B2(n9075), .A(n9063), .ZN(P1_U3235) );
  XNOR2_X1 U10407 ( .A(n9067), .B(n9066), .ZN(n9068) );
  XNOR2_X1 U10408 ( .A(n9065), .B(n9068), .ZN(n9076) );
  AOI22_X1 U10409 ( .A1(n9070), .A2(n9116), .B1(n9114), .B2(n9069), .ZN(n9415)
         );
  OAI22_X1 U10410 ( .A1(n9415), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9071), .ZN(n9073) );
  NOR2_X1 U10411 ( .A1(n9581), .A2(n9105), .ZN(n9072) );
  AOI211_X1 U10412 ( .C1(n9421), .C2(n9101), .A(n9073), .B(n9072), .ZN(n9074)
         );
  OAI21_X1 U10413 ( .B1(n9076), .B2(n9075), .A(n9074), .ZN(P1_U3238) );
  NAND2_X1 U10414 ( .A1(n9077), .A2(n9095), .ZN(n9091) );
  AOI21_X1 U10415 ( .B1(n9004), .B2(n9079), .A(n9078), .ZN(n9090) );
  OR2_X1 U10416 ( .A1(n9081), .A2(n9080), .ZN(n9085) );
  OR2_X1 U10417 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  AND2_X1 U10418 ( .A1(n9085), .A2(n9084), .ZN(n9289) );
  AOI22_X1 U10419 ( .A1(n9294), .A2(n9101), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9086) );
  OAI21_X1 U10420 ( .B1(n9289), .B2(n9098), .A(n9086), .ZN(n9087) );
  AOI21_X1 U10421 ( .B1(n9293), .B2(n9088), .A(n9087), .ZN(n9089) );
  OAI21_X1 U10422 ( .B1(n9091), .B2(n9090), .A(n9089), .ZN(P1_U3240) );
  OAI21_X1 U10423 ( .B1(n9092), .B2(n9094), .A(n9093), .ZN(n9096) );
  NAND2_X1 U10424 ( .A1(n9096), .A2(n9095), .ZN(n9104) );
  INV_X1 U10425 ( .A(n9097), .ZN(n9099) );
  OAI22_X1 U10426 ( .A1(n9099), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10098), .ZN(n9100) );
  AOI21_X1 U10427 ( .B1(n9102), .B2(n9101), .A(n9100), .ZN(n9103) );
  OAI211_X1 U10428 ( .C1(n9106), .C2(n9105), .A(n9104), .B(n9103), .ZN(
        P1_U3241) );
  MUX2_X1 U10429 ( .A(n9107), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9132), .Z(
        P1_U3584) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9108), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9109), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10432 ( .A(n9110), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9132), .Z(
        P1_U3578) );
  MUX2_X1 U10433 ( .A(n9111), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9132), .Z(
        P1_U3577) );
  MUX2_X1 U10434 ( .A(n9112), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9132), .Z(
        P1_U3576) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9113), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10436 ( .A(n9114), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9132), .Z(
        P1_U3573) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9115), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10438 ( .A(n9116), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9132), .Z(
        P1_U3571) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9117), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10440 ( .A(n9118), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9132), .Z(
        P1_U3569) );
  MUX2_X1 U10441 ( .A(n9119), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9132), .Z(
        P1_U3568) );
  MUX2_X1 U10442 ( .A(n9120), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9132), .Z(
        P1_U3567) );
  MUX2_X1 U10443 ( .A(n9121), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9132), .Z(
        P1_U3566) );
  MUX2_X1 U10444 ( .A(n9122), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9132), .Z(
        P1_U3565) );
  MUX2_X1 U10445 ( .A(n6216), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9132), .Z(
        P1_U3564) );
  MUX2_X1 U10446 ( .A(n9124), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9132), .Z(
        P1_U3563) );
  MUX2_X1 U10447 ( .A(n9125), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9132), .Z(
        P1_U3562) );
  MUX2_X1 U10448 ( .A(n9126), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9132), .Z(
        P1_U3561) );
  MUX2_X1 U10449 ( .A(n9127), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9132), .Z(
        P1_U3560) );
  MUX2_X1 U10450 ( .A(n9128), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9132), .Z(
        P1_U3559) );
  MUX2_X1 U10451 ( .A(n9129), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9132), .Z(
        P1_U3558) );
  MUX2_X1 U10452 ( .A(n9130), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9132), .Z(
        P1_U3557) );
  MUX2_X1 U10453 ( .A(n9131), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9132), .Z(
        P1_U3556) );
  MUX2_X1 U10454 ( .A(n9133), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9132), .Z(
        P1_U3555) );
  OAI211_X1 U10455 ( .C1(n9136), .C2(n9135), .A(n9664), .B(n9134), .ZN(n9144)
         );
  AOI22_X1 U10456 ( .A1(n9597), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9143) );
  NAND2_X1 U10457 ( .A1(n9656), .A2(n9137), .ZN(n9142) );
  OAI211_X1 U10458 ( .C1(n9140), .C2(n9139), .A(n9660), .B(n9138), .ZN(n9141)
         );
  NAND4_X1 U10459 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(
        P1_U3244) );
  NAND2_X1 U10460 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9145) );
  OAI21_X1 U10461 ( .B1(n9676), .B2(n10052), .A(n9145), .ZN(n9146) );
  AOI21_X1 U10462 ( .B1(n9147), .B2(n9656), .A(n9146), .ZN(n9156) );
  OAI211_X1 U10463 ( .C1(n9150), .C2(n9149), .A(n9664), .B(n9148), .ZN(n9155)
         );
  OAI211_X1 U10464 ( .C1(n9153), .C2(n9152), .A(n9660), .B(n9151), .ZN(n9154)
         );
  NAND3_X1 U10465 ( .A1(n9156), .A2(n9155), .A3(n9154), .ZN(P1_U3246) );
  INV_X1 U10466 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U10467 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9157) );
  OAI21_X1 U10468 ( .B1(n9676), .B2(n9158), .A(n9157), .ZN(n9159) );
  AOI21_X1 U10469 ( .B1(n9160), .B2(n9656), .A(n9159), .ZN(n9169) );
  OAI211_X1 U10470 ( .C1(n9163), .C2(n9162), .A(n9664), .B(n9161), .ZN(n9168)
         );
  OAI211_X1 U10471 ( .C1(n9166), .C2(n9165), .A(n9660), .B(n9164), .ZN(n9167)
         );
  NAND3_X1 U10472 ( .A1(n9169), .A2(n9168), .A3(n9167), .ZN(P1_U3248) );
  INV_X1 U10473 ( .A(n9170), .ZN(n9174) );
  INV_X1 U10474 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U10475 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9171) );
  OAI21_X1 U10476 ( .B1(n9676), .B2(n9172), .A(n9171), .ZN(n9173) );
  AOI21_X1 U10477 ( .B1(n9174), .B2(n9656), .A(n9173), .ZN(n9183) );
  OAI211_X1 U10478 ( .C1(n9177), .C2(n9176), .A(n9664), .B(n9175), .ZN(n9182)
         );
  OAI211_X1 U10479 ( .C1(n9180), .C2(n9179), .A(n9660), .B(n9178), .ZN(n9181)
         );
  NAND3_X1 U10480 ( .A1(n9183), .A2(n9182), .A3(n9181), .ZN(P1_U3249) );
  INV_X1 U10481 ( .A(n9184), .ZN(n9188) );
  INV_X1 U10482 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U10483 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9185) );
  OAI21_X1 U10484 ( .B1(n9676), .B2(n9186), .A(n9185), .ZN(n9187) );
  AOI21_X1 U10485 ( .B1(n9188), .B2(n9656), .A(n9187), .ZN(n9197) );
  OAI211_X1 U10486 ( .C1(n9191), .C2(n9190), .A(n9660), .B(n9189), .ZN(n9196)
         );
  OAI211_X1 U10487 ( .C1(n9194), .C2(n9193), .A(n9664), .B(n9192), .ZN(n9195)
         );
  NAND3_X1 U10488 ( .A1(n9197), .A2(n9196), .A3(n9195), .ZN(P1_U3250) );
  INV_X1 U10489 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U10490 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9198) );
  OAI21_X1 U10491 ( .B1(n9676), .B2(n9199), .A(n9198), .ZN(n9200) );
  AOI21_X1 U10492 ( .B1(n9201), .B2(n9656), .A(n9200), .ZN(n9210) );
  OAI211_X1 U10493 ( .C1(n9204), .C2(n9203), .A(n9660), .B(n9202), .ZN(n9209)
         );
  OAI211_X1 U10494 ( .C1(n9207), .C2(n9206), .A(n9664), .B(n9205), .ZN(n9208)
         );
  NAND3_X1 U10495 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(P1_U3251) );
  INV_X1 U10496 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9212) );
  AOI22_X1 U10497 ( .A1(n9214), .A2(n9213), .B1(n9212), .B2(n9211), .ZN(n9667)
         );
  INV_X1 U10498 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9518) );
  AND2_X1 U10499 ( .A1(n9221), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9215) );
  AOI21_X1 U10500 ( .B1(n9518), .B2(n9670), .A(n9215), .ZN(n9666) );
  NAND2_X1 U10501 ( .A1(n9667), .A2(n9666), .ZN(n9665) );
  INV_X1 U10502 ( .A(n9215), .ZN(n9216) );
  NAND2_X1 U10503 ( .A1(n9665), .A2(n9216), .ZN(n9217) );
  XOR2_X1 U10504 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9217), .Z(n9226) );
  OR2_X1 U10505 ( .A1(n9218), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U10506 ( .A1(n9221), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9223) );
  OR2_X1 U10507 ( .A1(n9221), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9222) );
  AND2_X1 U10508 ( .A1(n9223), .A2(n9222), .ZN(n9662) );
  NAND2_X1 U10509 ( .A1(n9663), .A2(n9662), .ZN(n9661) );
  NAND2_X1 U10510 ( .A1(n9661), .A2(n9223), .ZN(n9224) );
  XNOR2_X1 U10511 ( .A(n9224), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9228) );
  INV_X1 U10512 ( .A(n9228), .ZN(n9225) );
  AOI22_X1 U10513 ( .A1(n9226), .A2(n9664), .B1(n9660), .B2(n9225), .ZN(n9231)
         );
  NOR2_X1 U10514 ( .A1(n9226), .A2(n9645), .ZN(n9227) );
  AOI211_X1 U10515 ( .C1(n9660), .C2(n9228), .A(n9656), .B(n9227), .ZN(n9230)
         );
  MUX2_X1 U10516 ( .A(n9231), .B(n9230), .S(n9229), .Z(n9233) );
  NAND2_X1 U10517 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9232) );
  OAI211_X1 U10518 ( .C1(n9234), .C2(n9676), .A(n9233), .B(n9232), .ZN(
        P1_U3262) );
  NAND2_X1 U10519 ( .A1(n9550), .A2(n9243), .ZN(n9241) );
  XNOR2_X1 U10520 ( .A(n9235), .B(n9241), .ZN(n9236) );
  NAND2_X1 U10521 ( .A1(n9457), .A2(n9686), .ZN(n9240) );
  AND2_X1 U10522 ( .A1(n9238), .A2(n9237), .ZN(n9456) );
  INV_X1 U10523 ( .A(n9456), .ZN(n9460) );
  NOR2_X1 U10524 ( .A1(n9460), .A2(n9689), .ZN(n9245) );
  AOI21_X1 U10525 ( .B1(n9689), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9245), .ZN(
        n9239) );
  OAI211_X1 U10526 ( .C1(n9692), .C2(n9546), .A(n9240), .B(n9239), .ZN(
        P1_U3263) );
  OAI211_X1 U10527 ( .C1(n9550), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9461)
         );
  NOR2_X1 U10528 ( .A1(n9550), .A2(n9692), .ZN(n9244) );
  AOI211_X1 U10529 ( .C1(n9709), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9245), .B(
        n9244), .ZN(n9246) );
  OAI21_X1 U10530 ( .B1(n9247), .B2(n9461), .A(n9246), .ZN(P1_U3264) );
  OAI21_X1 U10531 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9466) );
  INV_X1 U10532 ( .A(n9466), .ZN(n9264) );
  XNOR2_X1 U10533 ( .A(n9252), .B(n9251), .ZN(n9253) );
  NAND2_X1 U10534 ( .A1(n9253), .A2(n9391), .ZN(n9255) );
  INV_X1 U10535 ( .A(n9258), .ZN(n9554) );
  INV_X1 U10536 ( .A(n9256), .ZN(n9257) );
  AOI211_X1 U10537 ( .C1(n9258), .C2(n9275), .A(n9418), .B(n9257), .ZN(n9465)
         );
  NAND2_X1 U10538 ( .A1(n9465), .A2(n9686), .ZN(n9261) );
  AOI22_X1 U10539 ( .A1(n9259), .A2(n9703), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9709), .ZN(n9260) );
  OAI211_X1 U10540 ( .C1(n9554), .C2(n9692), .A(n9261), .B(n9260), .ZN(n9262)
         );
  AOI21_X1 U10541 ( .B1(n9464), .B2(n9439), .A(n9262), .ZN(n9263) );
  OAI21_X1 U10542 ( .B1(n9264), .B2(n9426), .A(n9263), .ZN(P1_U3265) );
  XNOR2_X1 U10543 ( .A(n9265), .B(n9268), .ZN(n9471) );
  INV_X1 U10544 ( .A(n9471), .ZN(n9284) );
  OAI21_X1 U10545 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(n9272) );
  INV_X1 U10546 ( .A(n9269), .ZN(n9270) );
  NAND2_X1 U10547 ( .A1(n9266), .A2(n9270), .ZN(n9271) );
  NAND3_X1 U10548 ( .A1(n9272), .A2(n9271), .A3(n9391), .ZN(n9274) );
  NAND2_X1 U10549 ( .A1(n9274), .A2(n9273), .ZN(n9469) );
  INV_X1 U10550 ( .A(n9291), .ZN(n9277) );
  INV_X1 U10551 ( .A(n9275), .ZN(n9276) );
  AOI211_X1 U10552 ( .C1(n9278), .C2(n9277), .A(n9418), .B(n9276), .ZN(n9470)
         );
  NAND2_X1 U10553 ( .A1(n9470), .A2(n9686), .ZN(n9281) );
  AOI22_X1 U10554 ( .A1(n9279), .A2(n9703), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9709), .ZN(n9280) );
  OAI211_X1 U10555 ( .C1(n9558), .C2(n9692), .A(n9281), .B(n9280), .ZN(n9282)
         );
  AOI21_X1 U10556 ( .B1(n9469), .B2(n9439), .A(n9282), .ZN(n9283) );
  OAI21_X1 U10557 ( .B1(n9284), .B2(n9426), .A(n9283), .ZN(P1_U3266) );
  XOR2_X1 U10558 ( .A(n9286), .B(n9285), .Z(n9476) );
  INV_X1 U10559 ( .A(n9476), .ZN(n9299) );
  XNOR2_X1 U10560 ( .A(n9287), .B(n9286), .ZN(n9288) );
  NAND2_X1 U10561 ( .A1(n9288), .A2(n9391), .ZN(n9290) );
  NAND2_X1 U10562 ( .A1(n9290), .A2(n9289), .ZN(n9474) );
  INV_X1 U10563 ( .A(n9308), .ZN(n9292) );
  AOI211_X1 U10564 ( .C1(n9293), .C2(n9292), .A(n9418), .B(n9291), .ZN(n9475)
         );
  NAND2_X1 U10565 ( .A1(n9475), .A2(n9686), .ZN(n9296) );
  AOI22_X1 U10566 ( .A1(n9294), .A2(n9703), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9709), .ZN(n9295) );
  OAI211_X1 U10567 ( .C1(n9562), .C2(n9692), .A(n9296), .B(n9295), .ZN(n9297)
         );
  AOI21_X1 U10568 ( .B1(n9474), .B2(n9439), .A(n9297), .ZN(n9298) );
  OAI21_X1 U10569 ( .B1(n9299), .B2(n9426), .A(n9298), .ZN(P1_U3267) );
  XOR2_X1 U10570 ( .A(n9300), .B(n9301), .Z(n9481) );
  INV_X1 U10571 ( .A(n9481), .ZN(n9316) );
  NAND2_X1 U10572 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  NAND2_X1 U10573 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  NAND2_X1 U10574 ( .A1(n9305), .A2(n9391), .ZN(n9307) );
  NAND2_X1 U10575 ( .A1(n9307), .A2(n9306), .ZN(n9479) );
  INV_X1 U10576 ( .A(n9323), .ZN(n9309) );
  AOI211_X1 U10577 ( .C1(n9310), .C2(n9309), .A(n9418), .B(n9308), .ZN(n9480)
         );
  NAND2_X1 U10578 ( .A1(n9480), .A2(n9686), .ZN(n9313) );
  AOI22_X1 U10579 ( .A1(n9311), .A2(n9703), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9709), .ZN(n9312) );
  OAI211_X1 U10580 ( .C1(n9566), .C2(n9692), .A(n9313), .B(n9312), .ZN(n9314)
         );
  AOI21_X1 U10581 ( .B1(n9479), .B2(n9439), .A(n9314), .ZN(n9315) );
  OAI21_X1 U10582 ( .B1(n9316), .B2(n9426), .A(n9315), .ZN(P1_U3268) );
  XNOR2_X1 U10583 ( .A(n9317), .B(n9319), .ZN(n9488) );
  OAI211_X1 U10584 ( .C1(n9320), .C2(n9319), .A(n9318), .B(n9391), .ZN(n9322)
         );
  NAND2_X1 U10585 ( .A1(n9322), .A2(n9321), .ZN(n9484) );
  INV_X1 U10586 ( .A(n9339), .ZN(n9324) );
  AOI211_X1 U10587 ( .C1(n9486), .C2(n9324), .A(n9418), .B(n9323), .ZN(n9485)
         );
  NAND2_X1 U10588 ( .A1(n9485), .A2(n9686), .ZN(n9328) );
  INV_X1 U10589 ( .A(n9325), .ZN(n9326) );
  AOI22_X1 U10590 ( .A1(n9326), .A2(n9703), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9709), .ZN(n9327) );
  OAI211_X1 U10591 ( .C1(n9329), .C2(n9692), .A(n9328), .B(n9327), .ZN(n9330)
         );
  AOI21_X1 U10592 ( .B1(n9439), .B2(n9484), .A(n9330), .ZN(n9331) );
  OAI21_X1 U10593 ( .B1(n9488), .B2(n9426), .A(n9331), .ZN(P1_U3269) );
  XNOR2_X1 U10594 ( .A(n9332), .B(n9336), .ZN(n9493) );
  INV_X1 U10595 ( .A(n9333), .ZN(n9334) );
  AOI21_X1 U10596 ( .B1(n9336), .B2(n9335), .A(n9334), .ZN(n9338) );
  OAI21_X1 U10597 ( .B1(n9338), .B2(n9715), .A(n9337), .ZN(n9489) );
  INV_X1 U10598 ( .A(n9348), .ZN(n9340) );
  AOI211_X1 U10599 ( .C1(n9491), .C2(n9340), .A(n9418), .B(n9339), .ZN(n9490)
         );
  NAND2_X1 U10600 ( .A1(n9490), .A2(n9686), .ZN(n9343) );
  AOI22_X1 U10601 ( .A1(n9341), .A2(n9703), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9709), .ZN(n9342) );
  OAI211_X1 U10602 ( .C1(n9344), .C2(n9692), .A(n9343), .B(n9342), .ZN(n9345)
         );
  AOI21_X1 U10603 ( .B1(n9489), .B2(n9439), .A(n9345), .ZN(n9346) );
  OAI21_X1 U10604 ( .B1(n9493), .B2(n9426), .A(n9346), .ZN(P1_U3270) );
  XNOR2_X1 U10605 ( .A(n9347), .B(n9357), .ZN(n9496) );
  INV_X1 U10606 ( .A(n9496), .ZN(n9362) );
  AOI211_X1 U10607 ( .C1(n9349), .C2(n4706), .A(n9418), .B(n9348), .ZN(n9495)
         );
  NOR2_X1 U10608 ( .A1(n9571), .A2(n9692), .ZN(n9353) );
  OAI22_X1 U10609 ( .A1(n9351), .A2(n9441), .B1(n9350), .B2(n9439), .ZN(n9352)
         );
  AOI211_X1 U10610 ( .C1(n9495), .C2(n9686), .A(n9353), .B(n9352), .ZN(n9361)
         );
  INV_X1 U10611 ( .A(n9354), .ZN(n9355) );
  AOI211_X1 U10612 ( .C1(n9357), .C2(n9356), .A(n9715), .B(n9355), .ZN(n9359)
         );
  OR2_X1 U10613 ( .A1(n9359), .A2(n9358), .ZN(n9494) );
  NAND2_X1 U10614 ( .A1(n9494), .A2(n9439), .ZN(n9360) );
  OAI211_X1 U10615 ( .C1(n9362), .C2(n9426), .A(n9361), .B(n9360), .ZN(
        P1_U3271) );
  XOR2_X1 U10616 ( .A(n9363), .B(n9365), .Z(n9501) );
  INV_X1 U10617 ( .A(n9501), .ZN(n9378) );
  INV_X1 U10618 ( .A(n9379), .ZN(n9388) );
  NAND2_X1 U10619 ( .A1(n9389), .A2(n9388), .ZN(n9387) );
  NAND2_X1 U10620 ( .A1(n9387), .A2(n9364), .ZN(n9367) );
  INV_X1 U10621 ( .A(n9365), .ZN(n9366) );
  XNOR2_X1 U10622 ( .A(n9367), .B(n9366), .ZN(n9368) );
  NAND2_X1 U10623 ( .A1(n9368), .A2(n9391), .ZN(n9370) );
  NAND2_X1 U10624 ( .A1(n9370), .A2(n9369), .ZN(n9499) );
  AOI211_X1 U10625 ( .C1(n9372), .C2(n9381), .A(n9418), .B(n9371), .ZN(n9500)
         );
  NAND2_X1 U10626 ( .A1(n9500), .A2(n9686), .ZN(n9375) );
  AOI22_X1 U10627 ( .A1(n9373), .A2(n9703), .B1(n9689), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9374) );
  OAI211_X1 U10628 ( .C1(n9575), .C2(n9692), .A(n9375), .B(n9374), .ZN(n9376)
         );
  AOI21_X1 U10629 ( .B1(n9499), .B2(n9439), .A(n9376), .ZN(n9377) );
  OAI21_X1 U10630 ( .B1(n9378), .B2(n9426), .A(n9377), .ZN(P1_U3272) );
  XNOR2_X1 U10631 ( .A(n9380), .B(n9379), .ZN(n9508) );
  INV_X1 U10632 ( .A(n9381), .ZN(n9382) );
  AOI211_X1 U10633 ( .C1(n9505), .C2(n9403), .A(n9418), .B(n9382), .ZN(n9504)
         );
  INV_X1 U10634 ( .A(n9383), .ZN(n9384) );
  AOI22_X1 U10635 ( .A1(n9689), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9384), .B2(
        n9703), .ZN(n9385) );
  OAI21_X1 U10636 ( .B1(n9386), .B2(n9692), .A(n9385), .ZN(n9394) );
  OAI21_X1 U10637 ( .B1(n9389), .B2(n9388), .A(n9387), .ZN(n9392) );
  AOI21_X1 U10638 ( .B1(n9392), .B2(n9391), .A(n9390), .ZN(n9507) );
  NOR2_X1 U10639 ( .A1(n9507), .A2(n9689), .ZN(n9393) );
  AOI211_X1 U10640 ( .C1(n9504), .C2(n9686), .A(n9394), .B(n9393), .ZN(n9395)
         );
  OAI21_X1 U10641 ( .B1(n9508), .B2(n9426), .A(n9395), .ZN(P1_U3273) );
  XOR2_X1 U10642 ( .A(n9396), .B(n9400), .Z(n9514) );
  INV_X1 U10643 ( .A(n9397), .ZN(n9398) );
  AOI21_X1 U10644 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9402) );
  OAI21_X1 U10645 ( .B1(n9402), .B2(n9715), .A(n9401), .ZN(n9510) );
  INV_X1 U10646 ( .A(n9417), .ZN(n9405) );
  INV_X1 U10647 ( .A(n9403), .ZN(n9404) );
  AOI211_X1 U10648 ( .C1(n9512), .C2(n9405), .A(n9418), .B(n9404), .ZN(n9511)
         );
  NAND2_X1 U10649 ( .A1(n9511), .A2(n9450), .ZN(n9408) );
  AOI22_X1 U10650 ( .A1(n9709), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9406), .B2(
        n9703), .ZN(n9407) );
  OAI211_X1 U10651 ( .C1(n9409), .C2(n9692), .A(n9408), .B(n9407), .ZN(n9410)
         );
  AOI21_X1 U10652 ( .B1(n9510), .B2(n9439), .A(n9410), .ZN(n9411) );
  OAI21_X1 U10653 ( .B1(n9514), .B2(n9426), .A(n9411), .ZN(P1_U3274) );
  XNOR2_X1 U10654 ( .A(n9412), .B(n9413), .ZN(n9517) );
  INV_X1 U10655 ( .A(n9517), .ZN(n9427) );
  XNOR2_X1 U10656 ( .A(n9414), .B(n9413), .ZN(n9416) );
  OAI21_X1 U10657 ( .B1(n9416), .B2(n9715), .A(n9415), .ZN(n9515) );
  AOI211_X1 U10658 ( .C1(n9420), .C2(n9419), .A(n9418), .B(n9417), .ZN(n9516)
         );
  NAND2_X1 U10659 ( .A1(n9516), .A2(n9450), .ZN(n9423) );
  AOI22_X1 U10660 ( .A1(n9709), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9421), .B2(
        n9703), .ZN(n9422) );
  OAI211_X1 U10661 ( .C1(n9581), .C2(n9692), .A(n9423), .B(n9422), .ZN(n9424)
         );
  AOI21_X1 U10662 ( .B1(n9439), .B2(n9515), .A(n9424), .ZN(n9425) );
  OAI21_X1 U10663 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(P1_U3275) );
  NAND2_X1 U10664 ( .A1(n9428), .A2(n9439), .ZN(n9438) );
  OAI22_X1 U10665 ( .A1(n9439), .A2(n9430), .B1(n9429), .B2(n9441), .ZN(n9431)
         );
  AOI21_X1 U10666 ( .B1(n9432), .B2(n9678), .A(n9431), .ZN(n9437) );
  NAND2_X1 U10667 ( .A1(n9433), .A2(n9695), .ZN(n9436) );
  NAND2_X1 U10668 ( .A1(n9434), .A2(n9450), .ZN(n9435) );
  NAND4_X1 U10669 ( .A1(n9438), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(
        P1_U3284) );
  NAND2_X1 U10670 ( .A1(n9440), .A2(n9439), .ZN(n9455) );
  OAI22_X1 U10671 ( .A1(n9439), .A2(n9443), .B1(n9442), .B2(n9441), .ZN(n9444)
         );
  AOI21_X1 U10672 ( .B1(n9678), .B2(n9445), .A(n9444), .ZN(n9454) );
  INV_X1 U10673 ( .A(n9446), .ZN(n9447) );
  NOR2_X1 U10674 ( .A1(n9689), .A2(n9447), .ZN(n9449) );
  OAI21_X1 U10675 ( .B1(n9681), .B2(n9449), .A(n9448), .ZN(n9453) );
  NAND2_X1 U10676 ( .A1(n9451), .A2(n9450), .ZN(n9452) );
  NAND4_X1 U10677 ( .A1(n9455), .A2(n9454), .A3(n9453), .A4(n9452), .ZN(
        P1_U3285) );
  INV_X1 U10678 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9458) );
  NOR2_X1 U10679 ( .A1(n9457), .A2(n9456), .ZN(n9543) );
  OAI21_X1 U10680 ( .B1(n9530), .B2(n9546), .A(n9459), .ZN(P1_U3553) );
  AND2_X1 U10681 ( .A1(n9461), .A2(n9460), .ZN(n9547) );
  MUX2_X1 U10682 ( .A(n9462), .B(n9547), .S(n9509), .Z(n9463) );
  OAI21_X1 U10683 ( .B1(n9550), .B2(n9530), .A(n9463), .ZN(P1_U3552) );
  MUX2_X1 U10684 ( .A(n9467), .B(n9551), .S(n9509), .Z(n9468) );
  OAI21_X1 U10685 ( .B1(n9554), .B2(n9530), .A(n9468), .ZN(P1_U3550) );
  AOI211_X1 U10686 ( .C1(n9471), .C2(n9735), .A(n9470), .B(n9469), .ZN(n9555)
         );
  MUX2_X1 U10687 ( .A(n9472), .B(n9555), .S(n9509), .Z(n9473) );
  OAI21_X1 U10688 ( .B1(n9558), .B2(n9530), .A(n9473), .ZN(P1_U3549) );
  AOI211_X1 U10689 ( .C1(n9476), .C2(n9735), .A(n9475), .B(n9474), .ZN(n9559)
         );
  MUX2_X1 U10690 ( .A(n9477), .B(n9559), .S(n9745), .Z(n9478) );
  OAI21_X1 U10691 ( .B1(n9562), .B2(n9530), .A(n9478), .ZN(P1_U3548) );
  AOI211_X1 U10692 ( .C1(n9481), .C2(n9735), .A(n9480), .B(n9479), .ZN(n9563)
         );
  MUX2_X1 U10693 ( .A(n9482), .B(n9563), .S(n9509), .Z(n9483) );
  OAI21_X1 U10694 ( .B1(n9566), .B2(n9530), .A(n9483), .ZN(P1_U3547) );
  AOI211_X1 U10695 ( .C1(n9722), .C2(n9486), .A(n9485), .B(n9484), .ZN(n9487)
         );
  OAI21_X1 U10696 ( .B1(n9488), .B2(n9716), .A(n9487), .ZN(n9567) );
  MUX2_X1 U10697 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9567), .S(n9509), .Z(
        P1_U3546) );
  AOI211_X1 U10698 ( .C1(n9722), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9492)
         );
  OAI21_X1 U10699 ( .B1(n9493), .B2(n9716), .A(n9492), .ZN(n9568) );
  MUX2_X1 U10700 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9568), .S(n9509), .Z(
        P1_U3545) );
  INV_X1 U10701 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9497) );
  AOI211_X1 U10702 ( .C1(n9496), .C2(n9735), .A(n9495), .B(n9494), .ZN(n9569)
         );
  MUX2_X1 U10703 ( .A(n9497), .B(n9569), .S(n9745), .Z(n9498) );
  OAI21_X1 U10704 ( .B1(n9571), .B2(n9530), .A(n9498), .ZN(P1_U3544) );
  INV_X1 U10705 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9502) );
  AOI211_X1 U10706 ( .C1(n9501), .C2(n9735), .A(n9500), .B(n9499), .ZN(n9572)
         );
  MUX2_X1 U10707 ( .A(n9502), .B(n9572), .S(n9509), .Z(n9503) );
  OAI21_X1 U10708 ( .B1(n9575), .B2(n9530), .A(n9503), .ZN(P1_U3543) );
  AOI21_X1 U10709 ( .B1(n9722), .B2(n9505), .A(n9504), .ZN(n9506) );
  OAI211_X1 U10710 ( .C1(n9508), .C2(n9716), .A(n9507), .B(n9506), .ZN(n9576)
         );
  MUX2_X1 U10711 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9576), .S(n9509), .Z(
        P1_U3542) );
  AOI211_X1 U10712 ( .C1(n9722), .C2(n9512), .A(n9511), .B(n9510), .ZN(n9513)
         );
  OAI21_X1 U10713 ( .B1(n9514), .B2(n9716), .A(n9513), .ZN(n9577) );
  MUX2_X1 U10714 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9577), .S(n9745), .Z(
        P1_U3541) );
  AOI211_X1 U10715 ( .C1(n9517), .C2(n9735), .A(n9516), .B(n9515), .ZN(n9578)
         );
  MUX2_X1 U10716 ( .A(n9518), .B(n9578), .S(n9745), .Z(n9519) );
  OAI21_X1 U10717 ( .B1(n9581), .B2(n9530), .A(n9519), .ZN(P1_U3540) );
  AOI21_X1 U10718 ( .B1(n9722), .B2(n9521), .A(n9520), .ZN(n9522) );
  OAI211_X1 U10719 ( .C1(n9524), .C2(n9716), .A(n9523), .B(n9522), .ZN(n9582)
         );
  MUX2_X1 U10720 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9582), .S(n9745), .Z(
        P1_U3539) );
  INV_X1 U10721 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9528) );
  AOI211_X1 U10722 ( .C1(n9527), .C2(n9735), .A(n9526), .B(n9525), .ZN(n9583)
         );
  MUX2_X1 U10723 ( .A(n9528), .B(n9583), .S(n9745), .Z(n9529) );
  OAI21_X1 U10724 ( .B1(n9587), .B2(n9530), .A(n9529), .ZN(P1_U3538) );
  AOI21_X1 U10725 ( .B1(n9722), .B2(n9532), .A(n9531), .ZN(n9533) );
  OAI211_X1 U10726 ( .C1(n9535), .C2(n9716), .A(n9534), .B(n9533), .ZN(n9588)
         );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9588), .S(n9745), .Z(
        P1_U3537) );
  INV_X1 U10728 ( .A(n9726), .ZN(n9542) );
  INV_X1 U10729 ( .A(n9536), .ZN(n9541) );
  AOI21_X1 U10730 ( .B1(n9722), .B2(n9538), .A(n9537), .ZN(n9539) );
  OAI211_X1 U10731 ( .C1(n9542), .C2(n9541), .A(n9540), .B(n9539), .ZN(n9589)
         );
  MUX2_X1 U10732 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9589), .S(n9745), .Z(
        P1_U3536) );
  INV_X1 U10733 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9544) );
  OAI21_X1 U10734 ( .B1(n9586), .B2(n9546), .A(n9545), .ZN(P1_U3521) );
  INV_X1 U10735 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9548) );
  MUX2_X1 U10736 ( .A(n9548), .B(n9547), .S(n9738), .Z(n9549) );
  OAI21_X1 U10737 ( .B1(n9550), .B2(n9586), .A(n9549), .ZN(P1_U3520) );
  INV_X1 U10738 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9552) );
  MUX2_X1 U10739 ( .A(n9552), .B(n9551), .S(n9738), .Z(n9553) );
  INV_X1 U10740 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9556) );
  MUX2_X1 U10741 ( .A(n9556), .B(n9555), .S(n9738), .Z(n9557) );
  OAI21_X1 U10742 ( .B1(n9558), .B2(n9586), .A(n9557), .ZN(P1_U3517) );
  INV_X1 U10743 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9560) );
  MUX2_X1 U10744 ( .A(n9560), .B(n9559), .S(n9738), .Z(n9561) );
  OAI21_X1 U10745 ( .B1(n9562), .B2(n9586), .A(n9561), .ZN(P1_U3516) );
  INV_X1 U10746 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U10747 ( .A(n9564), .B(n9563), .S(n9738), .Z(n9565) );
  OAI21_X1 U10748 ( .B1(n9566), .B2(n9586), .A(n9565), .ZN(P1_U3515) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9567), .S(n9738), .Z(
        P1_U3514) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9568), .S(n9738), .Z(
        P1_U3513) );
  INV_X1 U10751 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10072) );
  MUX2_X1 U10752 ( .A(n10072), .B(n9569), .S(n9738), .Z(n9570) );
  OAI21_X1 U10753 ( .B1(n9571), .B2(n9586), .A(n9570), .ZN(P1_U3512) );
  INV_X1 U10754 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9573) );
  MUX2_X1 U10755 ( .A(n9573), .B(n9572), .S(n9738), .Z(n9574) );
  OAI21_X1 U10756 ( .B1(n9575), .B2(n9586), .A(n9574), .ZN(P1_U3511) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9576), .S(n9738), .Z(
        P1_U3510) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9577), .S(n9738), .Z(
        P1_U3509) );
  INV_X1 U10759 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9579) );
  MUX2_X1 U10760 ( .A(n9579), .B(n9578), .S(n9738), .Z(n9580) );
  OAI21_X1 U10761 ( .B1(n9581), .B2(n9586), .A(n9580), .ZN(P1_U3507) );
  MUX2_X1 U10762 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9582), .S(n9738), .Z(
        P1_U3504) );
  INV_X1 U10763 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9584) );
  MUX2_X1 U10764 ( .A(n9584), .B(n9583), .S(n9738), .Z(n9585) );
  OAI21_X1 U10765 ( .B1(n9587), .B2(n9586), .A(n9585), .ZN(P1_U3501) );
  MUX2_X1 U10766 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9588), .S(n9738), .Z(
        P1_U3498) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9589), .S(n9738), .Z(
        P1_U3495) );
  MUX2_X1 U10768 ( .A(n9590), .B(P1_D_REG_1__SCAN_IN), .S(n9711), .Z(P1_U3440)
         );
  MUX2_X1 U10769 ( .A(n9591), .B(P1_D_REG_0__SCAN_IN), .S(n9711), .Z(P1_U3439)
         );
  MUX2_X1 U10770 ( .A(n9592), .B(n9596), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10771 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10772 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10773 ( .B1(n9594), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9593), .ZN(
        n9595) );
  XOR2_X1 U10774 ( .A(n9596), .B(n9595), .Z(n9600) );
  AOI22_X1 U10775 ( .A1(n9597), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9598) );
  OAI21_X1 U10776 ( .B1(n9600), .B2(n9599), .A(n9598), .ZN(P1_U3243) );
  NOR2_X1 U10777 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  OR3_X1 U10778 ( .A1(n9604), .A2(n9603), .A3(n9645), .ZN(n9610) );
  NOR2_X1 U10779 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  OR3_X1 U10780 ( .A1(n9608), .A2(n9607), .A3(n9649), .ZN(n9609) );
  OAI211_X1 U10781 ( .C1(n9671), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U10782 ( .A(n9612), .ZN(n9614) );
  NAND2_X1 U10783 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9613) );
  OAI211_X1 U10784 ( .C1(n9676), .C2(n9615), .A(n9614), .B(n9613), .ZN(
        P1_U3254) );
  AOI211_X1 U10785 ( .C1(n9618), .C2(n9617), .A(n9616), .B(n9645), .ZN(n9623)
         );
  AOI211_X1 U10786 ( .C1(n9621), .C2(n9620), .A(n9619), .B(n9649), .ZN(n9622)
         );
  AOI211_X1 U10787 ( .C1(n9656), .C2(n9624), .A(n9623), .B(n9622), .ZN(n9626)
         );
  NAND2_X1 U10788 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9625) );
  OAI211_X1 U10789 ( .C1(n9676), .C2(n9627), .A(n9626), .B(n9625), .ZN(
        P1_U3256) );
  INV_X1 U10790 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9644) );
  NAND2_X1 U10791 ( .A1(n9629), .A2(n9628), .ZN(n9632) );
  INV_X1 U10792 ( .A(n9630), .ZN(n9631) );
  NAND2_X1 U10793 ( .A1(n9632), .A2(n9631), .ZN(n9640) );
  NAND2_X1 U10794 ( .A1(n9656), .A2(n9633), .ZN(n9639) );
  AOI21_X1 U10795 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9637) );
  NAND2_X1 U10796 ( .A1(n9660), .A2(n9637), .ZN(n9638) );
  OAI211_X1 U10797 ( .C1(n9645), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9641)
         );
  INV_X1 U10798 ( .A(n9641), .ZN(n9643) );
  NAND2_X1 U10799 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9642) );
  OAI211_X1 U10800 ( .C1(n9676), .C2(n9644), .A(n9643), .B(n9642), .ZN(
        P1_U3257) );
  AOI211_X1 U10801 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n9645), .ZN(n9654)
         );
  AOI211_X1 U10802 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9653)
         );
  AOI211_X1 U10803 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9658)
         );
  NAND2_X1 U10804 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9657) );
  OAI211_X1 U10805 ( .C1(n9676), .C2(n9659), .A(n9658), .B(n9657), .ZN(
        P1_U3258) );
  INV_X1 U10806 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9675) );
  OAI211_X1 U10807 ( .C1(n9663), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9669)
         );
  OAI211_X1 U10808 ( .C1(n9667), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9668)
         );
  OAI211_X1 U10809 ( .C1(n9671), .C2(n9670), .A(n9669), .B(n9668), .ZN(n9672)
         );
  INV_X1 U10810 ( .A(n9672), .ZN(n9674) );
  NAND2_X1 U10811 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9673) );
  OAI211_X1 U10812 ( .C1(n9676), .C2(n9675), .A(n9674), .B(n9673), .ZN(
        P1_U3261) );
  AOI222_X1 U10813 ( .A1(n9679), .A2(n9678), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9689), .C1(n9677), .C2(n9703), .ZN(n9684) );
  AOI22_X1 U10814 ( .A1(n9682), .A2(n9681), .B1(n9686), .B2(n9680), .ZN(n9683)
         );
  OAI211_X1 U10815 ( .C1(n9689), .C2(n9685), .A(n9684), .B(n9683), .ZN(
        P1_U3286) );
  NAND2_X1 U10816 ( .A1(n9687), .A2(n9686), .ZN(n9691) );
  AOI22_X1 U10817 ( .A1(n9689), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9688), .B2(
        n9703), .ZN(n9690) );
  OAI211_X1 U10818 ( .C1(n9693), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9694)
         );
  AOI21_X1 U10819 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(n9697) );
  OAI21_X1 U10820 ( .B1(n9709), .B2(n9698), .A(n9697), .ZN(P1_U3287) );
  NAND2_X1 U10821 ( .A1(n9699), .A2(n9720), .ZN(n9702) );
  INV_X1 U10822 ( .A(n9700), .ZN(n9701) );
  NAND2_X1 U10823 ( .A1(n9702), .A2(n9701), .ZN(n9704) );
  AOI22_X1 U10824 ( .A1(n9719), .A2(n9704), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9703), .ZN(n9705) );
  NAND2_X1 U10825 ( .A1(n9712), .A2(n9705), .ZN(n9706) );
  AOI21_X1 U10826 ( .B1(n9713), .B2(n9707), .A(n9706), .ZN(n9708) );
  AOI22_X1 U10827 ( .A1(n9709), .A2(n9960), .B1(n9708), .B2(n9439), .ZN(
        P1_U3293) );
  AND2_X1 U10828 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9711), .ZN(P1_U3294) );
  AND2_X1 U10829 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9711), .ZN(P1_U3295) );
  AND2_X1 U10830 ( .A1(n9711), .A2(P1_D_REG_29__SCAN_IN), .ZN(P1_U3296) );
  AND2_X1 U10831 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9711), .ZN(P1_U3297) );
  AND2_X1 U10832 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9711), .ZN(P1_U3298) );
  AND2_X1 U10833 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9711), .ZN(P1_U3299) );
  AND2_X1 U10834 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9711), .ZN(P1_U3300) );
  AND2_X1 U10835 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9711), .ZN(P1_U3301) );
  AND2_X1 U10836 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9711), .ZN(P1_U3302) );
  INV_X1 U10837 ( .A(n9711), .ZN(n9710) );
  INV_X1 U10838 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9941) );
  NOR2_X1 U10839 ( .A1(n9710), .A2(n9941), .ZN(P1_U3303) );
  AND2_X1 U10840 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9711), .ZN(P1_U3304) );
  AND2_X1 U10841 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9711), .ZN(P1_U3305) );
  AND2_X1 U10842 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9711), .ZN(P1_U3306) );
  INV_X1 U10843 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U10844 ( .A1(n9710), .A2(n10103), .ZN(P1_U3307) );
  AND2_X1 U10845 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9711), .ZN(P1_U3308) );
  AND2_X1 U10846 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9711), .ZN(P1_U3309) );
  AND2_X1 U10847 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9711), .ZN(P1_U3310) );
  AND2_X1 U10848 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9711), .ZN(P1_U3311) );
  AND2_X1 U10849 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9711), .ZN(P1_U3312) );
  AND2_X1 U10850 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9711), .ZN(P1_U3313) );
  AND2_X1 U10851 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9711), .ZN(P1_U3314) );
  AND2_X1 U10852 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9711), .ZN(P1_U3315) );
  AND2_X1 U10853 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9711), .ZN(P1_U3316) );
  AND2_X1 U10854 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9711), .ZN(P1_U3317) );
  AND2_X1 U10855 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9711), .ZN(P1_U3318) );
  INV_X1 U10856 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U10857 ( .A1(n9710), .A2(n10053), .ZN(P1_U3319) );
  INV_X1 U10858 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U10859 ( .A1(n9710), .A2(n10056), .ZN(P1_U3320) );
  AND2_X1 U10860 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9711), .ZN(P1_U3321) );
  AND2_X1 U10861 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9711), .ZN(P1_U3322) );
  AND2_X1 U10862 ( .A1(n9711), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3323) );
  INV_X1 U10863 ( .A(n9712), .ZN(n9718) );
  INV_X1 U10864 ( .A(n9713), .ZN(n9714) );
  AOI21_X1 U10865 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9717) );
  AOI211_X1 U10866 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9740)
         );
  INV_X1 U10867 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9721) );
  AOI22_X1 U10868 ( .A1(n9738), .A2(n9740), .B1(n9721), .B2(n7727), .ZN(
        P1_U3453) );
  INV_X1 U10869 ( .A(n9722), .ZN(n9732) );
  OAI21_X1 U10870 ( .B1(n9724), .B2(n9732), .A(n9723), .ZN(n9725) );
  AOI21_X1 U10871 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9728) );
  AND2_X1 U10872 ( .A1(n9729), .A2(n9728), .ZN(n9742) );
  INV_X1 U10873 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9730) );
  AOI22_X1 U10874 ( .A1(n9738), .A2(n9742), .B1(n9730), .B2(n7727), .ZN(
        P1_U3456) );
  OAI21_X1 U10875 ( .B1(n6221), .B2(n9732), .A(n9731), .ZN(n9733) );
  AOI211_X1 U10876 ( .C1(n9736), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9744)
         );
  INV_X1 U10877 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9737) );
  AOI22_X1 U10878 ( .A1(n9738), .A2(n9744), .B1(n9737), .B2(n7727), .ZN(
        P1_U3489) );
  INV_X1 U10879 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9739) );
  AOI22_X1 U10880 ( .A1(n9745), .A2(n9740), .B1(n9739), .B2(n9743), .ZN(
        P1_U3522) );
  AOI22_X1 U10881 ( .A1(n9745), .A2(n9742), .B1(n9741), .B2(n9743), .ZN(
        P1_U3523) );
  AOI22_X1 U10882 ( .A1(n9745), .A2(n9744), .B1(n10067), .B2(n9743), .ZN(
        P1_U3534) );
  AOI22_X1 U10883 ( .A1(n9783), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9750) );
  NOR2_X1 U10884 ( .A1(n9746), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9747) );
  OAI22_X1 U10885 ( .A1(n9788), .A2(n9748), .B1(n9762), .B2(n9747), .ZN(n9749)
         );
  OAI211_X1 U10886 ( .C1(n9904), .C2(n9768), .A(n9750), .B(n9749), .ZN(
        P2_U3182) );
  INV_X1 U10887 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U10888 ( .A1(n9768), .A2(n9899), .ZN(n9759) );
  INV_X1 U10889 ( .A(n9751), .ZN(n9752) );
  AOI21_X1 U10890 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9757) );
  XOR2_X1 U10891 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9755), .Z(n9756) );
  OAI22_X1 U10892 ( .A1(n9757), .A2(n9778), .B1(n9779), .B2(n9756), .ZN(n9758)
         );
  AOI211_X1 U10893 ( .C1(n9760), .C2(n9783), .A(n9759), .B(n9758), .ZN(n9765)
         );
  XOR2_X1 U10894 ( .A(n9762), .B(n9761), .Z(n9763) );
  NAND2_X1 U10895 ( .A1(n9788), .A2(n9763), .ZN(n9764) );
  OAI211_X1 U10896 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9766), .A(n9765), .B(
        n9764), .ZN(P2_U3183) );
  INV_X1 U10897 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9767) );
  NOR2_X1 U10898 ( .A1(n9768), .A2(n9767), .ZN(n9782) );
  INV_X1 U10899 ( .A(n9769), .ZN(n9770) );
  AOI21_X1 U10900 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9780) );
  OAI21_X1 U10901 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(n9776) );
  INV_X1 U10902 ( .A(n9776), .ZN(n9777) );
  OAI22_X1 U10903 ( .A1(n9780), .A2(n9779), .B1(n9778), .B2(n9777), .ZN(n9781)
         );
  AOI211_X1 U10904 ( .C1(n9784), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9790)
         );
  XOR2_X1 U10905 ( .A(n9786), .B(n9785), .Z(n9787) );
  NAND2_X1 U10906 ( .A1(n9788), .A2(n9787), .ZN(n9789) );
  OAI211_X1 U10907 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6980), .A(n9790), .B(
        n9789), .ZN(P2_U3184) );
  INV_X1 U10908 ( .A(n9791), .ZN(n9792) );
  AOI21_X1 U10909 ( .B1(n9795), .B2(n9793), .A(n9792), .ZN(n9855) );
  OAI22_X1 U10910 ( .A1(n10129), .A2(n9813), .B1(n10130), .B2(n9794), .ZN(
        n9800) );
  XNOR2_X1 U10911 ( .A(n9796), .B(n9795), .ZN(n9798) );
  NOR2_X1 U10912 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  AOI211_X1 U10913 ( .C1(n9848), .C2(n9855), .A(n9800), .B(n9799), .ZN(n9857)
         );
  INV_X1 U10914 ( .A(n10139), .ZN(n9805) );
  INV_X1 U10915 ( .A(n9801), .ZN(n9803) );
  AOI222_X1 U10916 ( .A1(n9805), .A2(n9804), .B1(n9855), .B2(n9803), .C1(
        n10135), .C2(n9802), .ZN(n9806) );
  OAI221_X1 U10917 ( .B1(n9808), .B2(n9857), .C1(n9807), .C2(n5864), .A(n9806), 
        .ZN(P2_U3224) );
  INV_X1 U10918 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U10919 ( .A1(n9880), .A2(n9810), .B1(n9809), .B2(n9878), .ZN(
        P2_U3390) );
  INV_X1 U10920 ( .A(n9811), .ZN(n9817) );
  OAI22_X1 U10921 ( .A1(n9814), .A2(n9813), .B1(n9812), .B2(n9865), .ZN(n9816)
         );
  AOI211_X1 U10922 ( .C1(n9869), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9882)
         );
  INV_X1 U10923 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10924 ( .A1(n9880), .A2(n9882), .B1(n9818), .B2(n9878), .ZN(
        P2_U3393) );
  INV_X1 U10925 ( .A(n9859), .ZN(n9854) );
  AOI211_X1 U10926 ( .C1(n9854), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9884)
         );
  INV_X1 U10927 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10928 ( .A1(n9880), .A2(n9884), .B1(n9822), .B2(n9878), .ZN(
        P2_U3396) );
  INV_X1 U10929 ( .A(n9823), .ZN(n9827) );
  OAI21_X1 U10930 ( .B1(n9825), .B2(n9865), .A(n9824), .ZN(n9826) );
  AOI21_X1 U10931 ( .B1(n9827), .B2(n9869), .A(n9826), .ZN(n9886) );
  INV_X1 U10932 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10933 ( .A1(n9880), .A2(n9886), .B1(n9828), .B2(n9878), .ZN(
        P2_U3402) );
  AND2_X1 U10934 ( .A1(n9829), .A2(n9869), .ZN(n9832) );
  AND2_X1 U10935 ( .A1(n9830), .A2(n9877), .ZN(n9831) );
  NOR3_X1 U10936 ( .A1(n9833), .A2(n9832), .A3(n9831), .ZN(n9887) );
  INV_X1 U10937 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U10938 ( .A1(n9880), .A2(n9887), .B1(n9834), .B2(n9878), .ZN(
        P2_U3405) );
  NAND2_X1 U10939 ( .A1(n9835), .A2(n9869), .ZN(n9838) );
  NAND2_X1 U10940 ( .A1(n9836), .A2(n9877), .ZN(n9837) );
  INV_X1 U10941 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U10942 ( .A1(n9880), .A2(n9888), .B1(n9840), .B2(n9878), .ZN(
        P2_U3408) );
  AOI22_X1 U10943 ( .A1(n10120), .A2(n9842), .B1(n9877), .B2(n9841), .ZN(n9843) );
  OAI21_X1 U10944 ( .B1(n9844), .B2(n9859), .A(n9843), .ZN(n9846) );
  AOI211_X1 U10945 ( .C1(n9848), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9889)
         );
  INV_X1 U10946 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9849) );
  AOI22_X1 U10947 ( .A1(n9880), .A2(n9889), .B1(n9849), .B2(n9878), .ZN(
        P2_U3411) );
  OAI21_X1 U10948 ( .B1(n9851), .B2(n9865), .A(n9850), .ZN(n9852) );
  AOI21_X1 U10949 ( .B1(n9869), .B2(n9853), .A(n9852), .ZN(n9890) );
  AOI22_X1 U10950 ( .A1(n9880), .A2(n9890), .B1(n5846), .B2(n9878), .ZN(
        P2_U3414) );
  AOI22_X1 U10951 ( .A1(n9855), .A2(n9854), .B1(n9877), .B2(n10135), .ZN(n9856) );
  AND2_X1 U10952 ( .A1(n9857), .A2(n9856), .ZN(n9891) );
  INV_X1 U10953 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10954 ( .A1(n9880), .A2(n9891), .B1(n9858), .B2(n9878), .ZN(
        P2_U3417) );
  NOR2_X1 U10955 ( .A1(n9860), .A2(n9859), .ZN(n9862) );
  AOI211_X1 U10956 ( .C1(n9877), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9892)
         );
  INV_X1 U10957 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9864) );
  AOI22_X1 U10958 ( .A1(n9880), .A2(n9892), .B1(n9864), .B2(n9878), .ZN(
        P2_U3420) );
  NOR2_X1 U10959 ( .A1(n9866), .A2(n9865), .ZN(n9868) );
  AOI211_X1 U10960 ( .C1(n9870), .C2(n9869), .A(n9868), .B(n9867), .ZN(n9893)
         );
  INV_X1 U10961 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9871) );
  AOI22_X1 U10962 ( .A1(n9880), .A2(n9893), .B1(n9871), .B2(n9878), .ZN(
        P2_U3423) );
  NOR2_X1 U10963 ( .A1(n9873), .A2(n9872), .ZN(n9875) );
  AOI211_X1 U10964 ( .C1(n9877), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9896)
         );
  INV_X1 U10965 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U10966 ( .A1(n9880), .A2(n9896), .B1(n9879), .B2(n9878), .ZN(
        P2_U3426) );
  INV_X1 U10967 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U10968 ( .A1(n9897), .A2(n9882), .B1(n9881), .B2(n9894), .ZN(
        P2_U3460) );
  AOI22_X1 U10969 ( .A1(n9897), .A2(n9884), .B1(n9883), .B2(n9894), .ZN(
        P2_U3461) );
  AOI22_X1 U10970 ( .A1(n9897), .A2(n9886), .B1(n9885), .B2(n9894), .ZN(
        P2_U3463) );
  AOI22_X1 U10971 ( .A1(n9897), .A2(n9887), .B1(n6757), .B2(n9894), .ZN(
        P2_U3464) );
  AOI22_X1 U10972 ( .A1(n9897), .A2(n9888), .B1(n6759), .B2(n9894), .ZN(
        P2_U3465) );
  AOI22_X1 U10973 ( .A1(n9897), .A2(n9889), .B1(n5832), .B2(n9894), .ZN(
        P2_U3466) );
  AOI22_X1 U10974 ( .A1(n9897), .A2(n9890), .B1(n7291), .B2(n9894), .ZN(
        P2_U3467) );
  AOI22_X1 U10975 ( .A1(n9897), .A2(n9891), .B1(n5860), .B2(n9894), .ZN(
        P2_U3468) );
  AOI22_X1 U10976 ( .A1(n9897), .A2(n9892), .B1(n7589), .B2(n9894), .ZN(
        P2_U3469) );
  AOI22_X1 U10977 ( .A1(n9897), .A2(n9893), .B1(n7682), .B2(n9894), .ZN(
        P2_U3470) );
  INV_X1 U10978 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U10979 ( .A1(n9897), .A2(n9896), .B1(n9895), .B2(n9894), .ZN(
        P2_U3471) );
  INV_X1 U10980 ( .A(n9898), .ZN(n9901) );
  AOI21_X1 U10981 ( .B1(n9903), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9902), .ZN(
        n9900) );
  OAI22_X1 U10982 ( .A1(n9902), .A2(n9901), .B1(n9900), .B2(n9899), .ZN(
        ADD_1068_U5) );
  AOI21_X1 U10983 ( .B1(n10086), .B2(n9904), .A(n9903), .ZN(ADD_1068_U46) );
  NOR2_X1 U10984 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  XOR2_X1 U10985 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n9907), .Z(ADD_1068_U55) );
  XNOR2_X1 U10986 ( .A(n9909), .B(n9908), .ZN(ADD_1068_U56) );
  XNOR2_X1 U10987 ( .A(n9911), .B(n9910), .ZN(ADD_1068_U57) );
  XNOR2_X1 U10988 ( .A(n9913), .B(n9912), .ZN(ADD_1068_U58) );
  XNOR2_X1 U10989 ( .A(n9915), .B(n9914), .ZN(ADD_1068_U59) );
  XNOR2_X1 U10990 ( .A(n9917), .B(n9916), .ZN(ADD_1068_U60) );
  XNOR2_X1 U10991 ( .A(n9919), .B(n9918), .ZN(ADD_1068_U61) );
  XNOR2_X1 U10992 ( .A(n9921), .B(n9920), .ZN(ADD_1068_U62) );
  XNOR2_X1 U10993 ( .A(n9923), .B(n9922), .ZN(ADD_1068_U63) );
  AOI22_X1 U10994 ( .A1(n10072), .A2(keyinput72), .B1(keyinput95), .B2(n10082), 
        .ZN(n9924) );
  OAI221_X1 U10995 ( .B1(n10072), .B2(keyinput72), .C1(n10082), .C2(keyinput95), .A(n9924), .ZN(n9935) );
  INV_X1 U10996 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U10997 ( .A1(n9927), .A2(keyinput92), .B1(keyinput81), .B2(n9926), 
        .ZN(n9925) );
  OAI221_X1 U10998 ( .B1(n9927), .B2(keyinput92), .C1(n9926), .C2(keyinput81), 
        .A(n9925), .ZN(n9934) );
  AOI22_X1 U10999 ( .A1(n9929), .A2(keyinput67), .B1(keyinput116), .B2(n10088), 
        .ZN(n9928) );
  OAI221_X1 U11000 ( .B1(n9929), .B2(keyinput67), .C1(n10088), .C2(keyinput116), .A(n9928), .ZN(n9933) );
  XNOR2_X1 U11001 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput113), .ZN(n9931) );
  XNOR2_X1 U11002 ( .A(SI_23_), .B(keyinput120), .ZN(n9930) );
  NAND2_X1 U11003 ( .A1(n9931), .A2(n9930), .ZN(n9932) );
  NOR4_X1 U11004 ( .A1(n9935), .A2(n9934), .A3(n9933), .A4(n9932), .ZN(n9973)
         );
  INV_X1 U11005 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11006 ( .A1(n9937), .A2(keyinput124), .B1(keyinput86), .B2(n10052), 
        .ZN(n9936) );
  OAI221_X1 U11007 ( .B1(n9937), .B2(keyinput124), .C1(n10052), .C2(keyinput86), .A(n9936), .ZN(n9947) );
  AOI22_X1 U11008 ( .A1(n10070), .A2(keyinput109), .B1(n9939), .B2(keyinput125), .ZN(n9938) );
  OAI221_X1 U11009 ( .B1(n10070), .B2(keyinput109), .C1(n9939), .C2(
        keyinput125), .A(n9938), .ZN(n9946) );
  AOI22_X1 U11010 ( .A1(n10104), .A2(keyinput126), .B1(n9941), .B2(keyinput68), 
        .ZN(n9940) );
  OAI221_X1 U11011 ( .B1(n10104), .B2(keyinput126), .C1(n9941), .C2(keyinput68), .A(n9940), .ZN(n9945) );
  INV_X1 U11012 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U11013 ( .A1(n9943), .A2(keyinput112), .B1(keyinput84), .B2(n7682), 
        .ZN(n9942) );
  OAI221_X1 U11014 ( .B1(n9943), .B2(keyinput112), .C1(n7682), .C2(keyinput84), 
        .A(n9942), .ZN(n9944) );
  NOR4_X1 U11015 ( .A1(n9947), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n9972)
         );
  INV_X1 U11016 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9949) );
  AOI22_X1 U11017 ( .A1(n9949), .A2(keyinput117), .B1(keyinput78), .B2(n10055), 
        .ZN(n9948) );
  OAI221_X1 U11018 ( .B1(n9949), .B2(keyinput117), .C1(n10055), .C2(keyinput78), .A(n9948), .ZN(n9958) );
  AOI22_X1 U11019 ( .A1(n10089), .A2(keyinput104), .B1(n10053), .B2(keyinput64), .ZN(n9950) );
  OAI221_X1 U11020 ( .B1(n10089), .B2(keyinput104), .C1(n10053), .C2(
        keyinput64), .A(n9950), .ZN(n9957) );
  INV_X1 U11021 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U11022 ( .A1(n10074), .A2(keyinput119), .B1(n9952), .B2(keyinput73), 
        .ZN(n9951) );
  OAI221_X1 U11023 ( .B1(n10074), .B2(keyinput119), .C1(n9952), .C2(keyinput73), .A(n9951), .ZN(n9956) );
  XOR2_X1 U11024 ( .A(n10100), .B(keyinput75), .Z(n9954) );
  XNOR2_X1 U11025 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput99), .ZN(n9953) );
  NAND2_X1 U11026 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NOR4_X1 U11027 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n9971)
         );
  AOI22_X1 U11028 ( .A1(n10056), .A2(keyinput97), .B1(keyinput110), .B2(n9960), 
        .ZN(n9959) );
  OAI221_X1 U11029 ( .B1(n10056), .B2(keyinput97), .C1(n9960), .C2(keyinput110), .A(n9959), .ZN(n9969) );
  AOI22_X1 U11030 ( .A1(n10086), .A2(keyinput94), .B1(n6044), .B2(keyinput69), 
        .ZN(n9961) );
  OAI221_X1 U11031 ( .B1(n10086), .B2(keyinput94), .C1(n6044), .C2(keyinput69), 
        .A(n9961), .ZN(n9968) );
  AOI22_X1 U11032 ( .A1(n9963), .A2(keyinput90), .B1(keyinput105), .B2(n10098), 
        .ZN(n9962) );
  OAI221_X1 U11033 ( .B1(n9963), .B2(keyinput90), .C1(n10098), .C2(keyinput105), .A(n9962), .ZN(n9967) );
  XNOR2_X1 U11034 ( .A(P2_REG1_REG_20__SCAN_IN), .B(keyinput122), .ZN(n9965)
         );
  XNOR2_X1 U11035 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput76), .ZN(n9964) );
  NAND2_X1 U11036 ( .A1(n9965), .A2(n9964), .ZN(n9966) );
  NOR4_X1 U11037 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n9970)
         );
  AND4_X1 U11038 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n10118)
         );
  OAI22_X1 U11039 ( .A1(P1_D_REG_29__SCAN_IN), .A2(keyinput101), .B1(
        keyinput85), .B2(SI_12_), .ZN(n9974) );
  AOI221_X1 U11040 ( .B1(P1_D_REG_29__SCAN_IN), .B2(keyinput101), .C1(SI_12_), 
        .C2(keyinput85), .A(n9974), .ZN(n9981) );
  OAI22_X1 U11041 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(keyinput70), .B1(SI_2_), 
        .B2(keyinput88), .ZN(n9975) );
  AOI221_X1 U11042 ( .B1(P1_DATAO_REG_6__SCAN_IN), .B2(keyinput70), .C1(
        keyinput88), .C2(SI_2_), .A(n9975), .ZN(n9980) );
  OAI22_X1 U11043 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput82), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput89), .ZN(n9976) );
  AOI221_X1 U11044 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput82), .C1(
        keyinput89), .C2(P2_REG0_REG_28__SCAN_IN), .A(n9976), .ZN(n9979) );
  OAI22_X1 U11045 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput100), .B1(
        P1_REG2_REG_6__SCAN_IN), .B2(keyinput91), .ZN(n9977) );
  AOI221_X1 U11046 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput100), .C1(
        keyinput91), .C2(P1_REG2_REG_6__SCAN_IN), .A(n9977), .ZN(n9978) );
  NAND4_X1 U11047 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n10012) );
  OAI22_X1 U11048 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput102), .B1(
        keyinput107), .B2(P1_D_REG_18__SCAN_IN), .ZN(n9982) );
  AOI221_X1 U11049 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput102), .C1(
        P1_D_REG_18__SCAN_IN), .C2(keyinput107), .A(n9982), .ZN(n9989) );
  OAI22_X1 U11050 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput77), .B1(
        P2_D_REG_15__SCAN_IN), .B2(keyinput127), .ZN(n9983) );
  AOI221_X1 U11051 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput77), .C1(
        keyinput127), .C2(P2_D_REG_15__SCAN_IN), .A(n9983), .ZN(n9988) );
  OAI22_X1 U11052 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput80), .B1(
        P2_REG1_REG_31__SCAN_IN), .B2(keyinput121), .ZN(n9984) );
  AOI221_X1 U11053 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput80), .C1(
        keyinput121), .C2(P2_REG1_REG_31__SCAN_IN), .A(n9984), .ZN(n9987) );
  OAI22_X1 U11054 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput93), .B1(
        P2_REG2_REG_29__SCAN_IN), .B2(keyinput123), .ZN(n9985) );
  AOI221_X1 U11055 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput93), .C1(
        keyinput123), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9985), .ZN(n9986) );
  NAND4_X1 U11056 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n10011) );
  OAI22_X1 U11057 ( .A1(n9991), .A2(keyinput115), .B1(keyinput118), .B2(
        P1_WR_REG_SCAN_IN), .ZN(n9990) );
  AOI221_X1 U11058 ( .B1(n9991), .B2(keyinput115), .C1(P1_WR_REG_SCAN_IN), 
        .C2(keyinput118), .A(n9990), .ZN(n10000) );
  OAI22_X1 U11059 ( .A1(SI_14_), .A2(keyinput114), .B1(keyinput108), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9992) );
  AOI221_X1 U11060 ( .B1(SI_14_), .B2(keyinput114), .C1(
        P1_DATAO_REG_14__SCAN_IN), .C2(keyinput108), .A(n9992), .ZN(n9999) );
  OAI22_X1 U11061 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput87), .B1(
        keyinput98), .B2(P2_REG2_REG_3__SCAN_IN), .ZN(n9993) );
  AOI221_X1 U11062 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG2_REG_3__SCAN_IN), .C2(keyinput98), .A(n9993), .ZN(n9998) );
  XOR2_X1 U11063 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput71), .Z(n9996) );
  XNOR2_X1 U11064 ( .A(n9994), .B(keyinput111), .ZN(n9995) );
  NOR2_X1 U11065 ( .A1(n9996), .A2(n9995), .ZN(n9997) );
  NAND4_X1 U11066 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(
        n10010) );
  OAI22_X1 U11067 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput106), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput65), .ZN(n10001) );
  AOI221_X1 U11068 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput106), .C1(
        keyinput65), .C2(P2_D_REG_28__SCAN_IN), .A(n10001), .ZN(n10008) );
  OAI22_X1 U11069 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput74), .B1(
        keyinput103), .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n10002) );
  AOI221_X1 U11070 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput74), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput103), .A(n10002), .ZN(n10007) );
  OAI22_X1 U11071 ( .A1(SI_28_), .A2(keyinput96), .B1(P2_REG2_REG_8__SCAN_IN), 
        .B2(keyinput66), .ZN(n10003) );
  AOI221_X1 U11072 ( .B1(SI_28_), .B2(keyinput96), .C1(keyinput66), .C2(
        P2_REG2_REG_8__SCAN_IN), .A(n10003), .ZN(n10006) );
  OAI22_X1 U11073 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput83), .B1(
        P1_REG1_REG_12__SCAN_IN), .B2(keyinput79), .ZN(n10004) );
  AOI221_X1 U11074 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput83), .C1(keyinput79), .C2(P1_REG1_REG_12__SCAN_IN), .A(n10004), .ZN(n10005) );
  NAND4_X1 U11075 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10009) );
  NOR4_X1 U11076 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10117) );
  AOI22_X1 U11077 ( .A1(P2_D_REG_15__SCAN_IN), .A2(keyinput63), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput37), .ZN(n10013) );
  OAI221_X1 U11078 ( .B1(P2_D_REG_15__SCAN_IN), .B2(keyinput63), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput37), .A(n10013), .ZN(n10020) );
  AOI22_X1 U11079 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput7), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(keyinput61), .ZN(n10014) );
  OAI221_X1 U11080 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput7), .C1(
        P1_DATAO_REG_25__SCAN_IN), .C2(keyinput61), .A(n10014), .ZN(n10019) );
  AOI22_X1 U11081 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput23), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(keyinput28), .ZN(n10015) );
  OAI221_X1 U11082 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput23), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput28), .A(n10015), .ZN(n10018) );
  AOI22_X1 U11083 ( .A1(P1_WR_REG_SCAN_IN), .A2(keyinput54), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput19), .ZN(n10016) );
  OAI221_X1 U11084 ( .B1(P1_WR_REG_SCAN_IN), .B2(keyinput54), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput19), .A(n10016), .ZN(n10017) );
  NOR4_X1 U11085 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10050) );
  AOI22_X1 U11086 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput5), .B1(
        P1_REG0_REG_2__SCAN_IN), .B2(keyinput17), .ZN(n10021) );
  OAI221_X1 U11087 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput5), .C1(
        P1_REG0_REG_2__SCAN_IN), .C2(keyinput17), .A(n10021), .ZN(n10028) );
  AOI22_X1 U11088 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(keyinput20), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput1), .ZN(n10022) );
  OAI221_X1 U11089 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(keyinput20), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput1), .A(n10022), .ZN(n10027) );
  AOI22_X1 U11090 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(keyinput3), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput26), .ZN(n10023) );
  OAI221_X1 U11091 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(keyinput3), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput26), .A(n10023), .ZN(n10026) );
  AOI22_X1 U11092 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(keyinput47), .B1(
        P1_D_REG_22__SCAN_IN), .B2(keyinput4), .ZN(n10024) );
  OAI221_X1 U11093 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(keyinput47), .C1(
        P1_D_REG_22__SCAN_IN), .C2(keyinput4), .A(n10024), .ZN(n10025) );
  NOR4_X1 U11094 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10049) );
  AOI22_X1 U11095 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(keyinput51), .B1(
        P1_REG1_REG_19__SCAN_IN), .B2(keyinput53), .ZN(n10029) );
  OAI221_X1 U11096 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(keyinput51), .C1(
        P1_REG1_REG_19__SCAN_IN), .C2(keyinput53), .A(n10029), .ZN(n10036) );
  AOI22_X1 U11097 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(keyinput2), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput12), .ZN(n10030) );
  OAI221_X1 U11098 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(keyinput2), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput12), .A(n10030), .ZN(n10035) );
  AOI22_X1 U11099 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput46), .B1(
        P1_REG2_REG_21__SCAN_IN), .B2(keyinput60), .ZN(n10031) );
  OAI221_X1 U11100 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput46), .C1(
        P1_REG2_REG_21__SCAN_IN), .C2(keyinput60), .A(n10031), .ZN(n10034) );
  AOI22_X1 U11101 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput57), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput39), .ZN(n10032) );
  OAI221_X1 U11102 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput57), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput39), .A(n10032), .ZN(n10033) );
  NOR4_X1 U11103 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n10048) );
  AOI22_X1 U11104 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(keyinput9), .B1(SI_23_), 
        .B2(keyinput56), .ZN(n10037) );
  OAI221_X1 U11105 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(keyinput9), .C1(SI_23_), 
        .C2(keyinput56), .A(n10037), .ZN(n10046) );
  AOI22_X1 U11106 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput36), .B1(
        P1_REG1_REG_22__SCAN_IN), .B2(keyinput16), .ZN(n10038) );
  OAI221_X1 U11107 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput36), .C1(
        P1_REG1_REG_22__SCAN_IN), .C2(keyinput16), .A(n10038), .ZN(n10045) );
  XNOR2_X1 U11108 ( .A(n10039), .B(keyinput49), .ZN(n10043) );
  XNOR2_X1 U11109 ( .A(SI_2_), .B(keyinput24), .ZN(n10042) );
  XNOR2_X1 U11110 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput6), .ZN(n10041) );
  XNOR2_X1 U11111 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput10), .ZN(n10040)
         );
  NAND4_X1 U11112 ( .A1(n10043), .A2(n10042), .A3(n10041), .A4(n10040), .ZN(
        n10044) );
  NOR3_X1 U11113 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n10047) );
  NAND4_X1 U11114 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10116) );
  AOI22_X1 U11115 ( .A1(n10053), .A2(keyinput0), .B1(keyinput22), .B2(n10052), 
        .ZN(n10051) );
  OAI221_X1 U11116 ( .B1(n10053), .B2(keyinput0), .C1(n10052), .C2(keyinput22), 
        .A(n10051), .ZN(n10065) );
  AOI22_X1 U11117 ( .A1(n10056), .A2(keyinput33), .B1(keyinput14), .B2(n10055), 
        .ZN(n10054) );
  OAI221_X1 U11118 ( .B1(n10056), .B2(keyinput33), .C1(n10055), .C2(keyinput14), .A(n10054), .ZN(n10064) );
  AOI22_X1 U11119 ( .A1(n10059), .A2(keyinput25), .B1(n10058), .B2(keyinput44), 
        .ZN(n10057) );
  OAI221_X1 U11120 ( .B1(n10059), .B2(keyinput25), .C1(n10058), .C2(keyinput44), .A(n10057), .ZN(n10063) );
  XNOR2_X1 U11121 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput38), .ZN(n10061) );
  XNOR2_X1 U11122 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput48), .ZN(n10060)
         );
  NAND2_X1 U11123 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  NOR4_X1 U11124 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        n10114) );
  AOI22_X1 U11125 ( .A1(n4945), .A2(keyinput21), .B1(keyinput15), .B2(n10067), 
        .ZN(n10066) );
  OAI221_X1 U11126 ( .B1(n4945), .B2(keyinput21), .C1(n10067), .C2(keyinput15), 
        .A(n10066), .ZN(n10080) );
  INV_X1 U11127 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U11128 ( .A1(n10070), .A2(keyinput45), .B1(keyinput59), .B2(n10069), 
        .ZN(n10068) );
  OAI221_X1 U11129 ( .B1(n10070), .B2(keyinput45), .C1(n10069), .C2(keyinput59), .A(n10068), .ZN(n10079) );
  AOI22_X1 U11130 ( .A1(n10073), .A2(keyinput32), .B1(keyinput8), .B2(n10072), 
        .ZN(n10071) );
  OAI221_X1 U11131 ( .B1(n10073), .B2(keyinput32), .C1(n10072), .C2(keyinput8), 
        .A(n10071), .ZN(n10078) );
  XOR2_X1 U11132 ( .A(n10074), .B(keyinput55), .Z(n10076) );
  XNOR2_X1 U11133 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput42), .ZN(n10075)
         );
  NAND2_X1 U11134 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  NOR4_X1 U11135 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10113) );
  AOI22_X1 U11136 ( .A1(n10083), .A2(keyinput58), .B1(n10082), .B2(keyinput31), 
        .ZN(n10081) );
  OAI221_X1 U11137 ( .B1(n10083), .B2(keyinput58), .C1(n10082), .C2(keyinput31), .A(n10081), .ZN(n10095) );
  AOI22_X1 U11138 ( .A1(n10086), .A2(keyinput30), .B1(n10085), .B2(keyinput18), 
        .ZN(n10084) );
  OAI221_X1 U11139 ( .B1(n10086), .B2(keyinput30), .C1(n10085), .C2(keyinput18), .A(n10084), .ZN(n10094) );
  AOI22_X1 U11140 ( .A1(n10089), .A2(keyinput40), .B1(keyinput52), .B2(n10088), 
        .ZN(n10087) );
  OAI221_X1 U11141 ( .B1(n10089), .B2(keyinput40), .C1(n10088), .C2(keyinput52), .A(n10087), .ZN(n10093) );
  XNOR2_X1 U11142 ( .A(P1_REG0_REG_15__SCAN_IN), .B(keyinput29), .ZN(n10091)
         );
  XNOR2_X1 U11143 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput13), .ZN(n10090) );
  NAND2_X1 U11144 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  NOR4_X1 U11145 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10112) );
  AOI22_X1 U11146 ( .A1(n10098), .A2(keyinput41), .B1(keyinput27), .B2(n10097), 
        .ZN(n10096) );
  OAI221_X1 U11147 ( .B1(n10098), .B2(keyinput41), .C1(n10097), .C2(keyinput27), .A(n10096), .ZN(n10110) );
  INV_X1 U11148 ( .A(SI_14_), .ZN(n10101) );
  AOI22_X1 U11149 ( .A1(n10101), .A2(keyinput50), .B1(keyinput11), .B2(n10100), 
        .ZN(n10099) );
  OAI221_X1 U11150 ( .B1(n10101), .B2(keyinput50), .C1(n10100), .C2(keyinput11), .A(n10099), .ZN(n10109) );
  AOI22_X1 U11151 ( .A1(n10104), .A2(keyinput62), .B1(n10103), .B2(keyinput43), 
        .ZN(n10102) );
  OAI221_X1 U11152 ( .B1(n10104), .B2(keyinput62), .C1(n10103), .C2(keyinput43), .A(n10102), .ZN(n10108) );
  XOR2_X1 U11153 ( .A(n7301), .B(keyinput34), .Z(n10106) );
  XNOR2_X1 U11154 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput35), .ZN(n10105) );
  NAND2_X1 U11155 ( .A1(n10106), .A2(n10105), .ZN(n10107) );
  NOR4_X1 U11156 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10111) );
  NAND4_X1 U11157 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10115) );
  AOI211_X1 U11158 ( .C1(n10118), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10141) );
  OAI22_X1 U11159 ( .A1(n10121), .A2(n10120), .B1(n7553), .B2(n10119), .ZN(
        n10125) );
  XNOR2_X1 U11160 ( .A(n10123), .B(n10122), .ZN(n10124) );
  XNOR2_X1 U11161 ( .A(n10125), .B(n10124), .ZN(n10127) );
  NAND2_X1 U11162 ( .A1(n10127), .A2(n10126), .ZN(n10137) );
  OAI22_X1 U11163 ( .A1(n10131), .A2(n10130), .B1(n10129), .B2(n10128), .ZN(
        n10132) );
  AOI211_X1 U11164 ( .C1(n10135), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        n10136) );
  OAI211_X1 U11165 ( .C1(n10139), .C2(n10138), .A(n10137), .B(n10136), .ZN(
        n10140) );
  XOR2_X1 U11166 ( .A(n10141), .B(n10140), .Z(P2_U3171) );
  XNOR2_X1 U11167 ( .A(n10143), .B(n10142), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11168 ( .A(n10145), .B(n10144), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11169 ( .A(n10147), .B(n10146), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11170 ( .A(n10149), .B(n10148), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11171 ( .A(n10151), .B(n10150), .ZN(ADD_1068_U48) );
  XOR2_X1 U11172 ( .A(n10153), .B(n10152), .Z(ADD_1068_U54) );
  XOR2_X1 U11173 ( .A(n10155), .B(n10154), .Z(ADD_1068_U53) );
  XNOR2_X1 U11174 ( .A(n10157), .B(n10156), .ZN(ADD_1068_U52) );
  AND2_X1 U6553 ( .A1(n5079), .A2(n7883), .ZN(n5430) );
  CLKBUF_X2 U4857 ( .A(n5431), .Z(n5463) );
  AND2_X1 U6556 ( .A1(n8270), .A2(n7883), .ZN(n5431) );
  CLKBUF_X2 U4920 ( .A(n4891), .Z(n6376) );
  CLKBUF_X1 U4935 ( .A(n5779), .Z(n6094) );
  CLKBUF_X2 U4971 ( .A(n5785), .Z(n8055) );
  CLKBUF_X1 U5029 ( .A(n5428), .Z(n5464) );
  CLKBUF_X1 U5757 ( .A(n5429), .Z(n5362) );
  CLKBUF_X1 U5849 ( .A(n9509), .Z(n9745) );
endmodule

