

module b22_C_gen_AntiSAT_k_256_6 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710;

  INV_X4 U7419 ( .A(n13155), .ZN(P3_U3897) );
  INV_X4 U7420 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  AND2_X1 U7421 ( .A1(n14584), .A2(n8492), .ZN(n14601) );
  NAND2_X1 U7422 ( .A1(n13748), .A2(n6813), .ZN(n13704) );
  NAND2_X1 U7423 ( .A1(n8306), .A2(n8305), .ZN(n14877) );
  NAND2_X1 U7424 ( .A1(n7225), .A2(n7229), .ZN(n9581) );
  OAI21_X1 U7425 ( .B1(n13527), .B2(n9823), .A(n10137), .ZN(n12486) );
  NAND2_X1 U7426 ( .A1(n10304), .A2(n10303), .ZN(n11471) );
  AND2_X1 U7427 ( .A1(n6871), .A2(n11846), .ZN(n11848) );
  CLKBUF_X2 U7428 ( .A(n8031), .Z(n6677) );
  NAND2_X1 U7429 ( .A1(n11485), .A2(n11487), .ZN(n12624) );
  INV_X4 U7430 ( .A(n8580), .ZN(n6678) );
  CLKBUF_X1 U7431 ( .A(n10024), .Z(n6994) );
  CLKBUF_X2 U7432 ( .A(n8655), .Z(n12882) );
  INV_X2 U7433 ( .A(n10701), .ZN(n10448) );
  OR2_X1 U7434 ( .A1(n8646), .A2(n10496), .ZN(n8632) );
  INV_X1 U7435 ( .A(n12926), .ZN(n13871) );
  NOR2_X2 U7436 ( .A1(n8611), .A2(n10971), .ZN(n8613) );
  INV_X2 U7437 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9493) );
  OR2_X2 U7438 ( .A1(n11061), .A2(n11059), .ZN(n10283) );
  OR2_X1 U7439 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U7440 ( .A1(n13739), .A2(n13738), .ZN(n6672) );
  CLKBUF_X1 U7441 ( .A(n11020), .Z(n6673) );
  NAND2_X1 U7442 ( .A1(n13739), .A2(n13738), .ZN(n13737) );
  OAI21_X1 U7443 ( .B1(n7678), .B2(n12822), .A(n7677), .ZN(n12833) );
  AND2_X1 U7444 ( .A1(n10444), .A2(n14710), .ZN(n10417) );
  CLKBUF_X3 U7445 ( .A(n9646), .Z(n10000) );
  INV_X1 U7446 ( .A(n10024), .ZN(n9951) );
  XNOR2_X1 U7447 ( .A(n7042), .B(n13288), .ZN(n13267) );
  INV_X1 U7448 ( .A(n8458), .ZN(n8483) );
  NOR2_X2 U7449 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7921) );
  AND4_X1 U7450 ( .A1(n9675), .A2(n9674), .A3(n9673), .A4(n9672), .ZN(n12094)
         );
  NOR2_X1 U7451 ( .A1(n9997), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10012) );
  INV_X2 U7452 ( .A(n12624), .ZN(n11532) );
  INV_X1 U7453 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U7454 ( .A1(n10938), .A2(n6675), .ZN(n8867) );
  INV_X1 U7455 ( .A(n12868), .ZN(n12883) );
  AND2_X1 U7456 ( .A1(n13992), .A2(n7341), .ZN(n13952) );
  CLKBUF_X2 U7457 ( .A(n12846), .Z(n6675) );
  NAND2_X1 U7458 ( .A1(n7011), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8589) );
  INV_X1 U7459 ( .A(n6967), .ZN(n10458) );
  AOI21_X1 U7460 ( .B1(n12376), .B2(P1_REG1_REG_16__SCAN_IN), .A(n12375), .ZN(
        n12379) );
  AND2_X1 U7461 ( .A1(n14634), .A2(n14625), .ZN(n14618) );
  INV_X2 U7463 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7784) );
  OR2_X1 U7464 ( .A1(n15005), .A2(n15006), .ZN(n6923) );
  INV_X1 U7465 ( .A(n15591), .ZN(n15622) );
  NAND2_X1 U7466 ( .A1(n8740), .A2(n8739), .ZN(n15434) );
  NAND2_X1 U7467 ( .A1(n12852), .A2(n12851), .ZN(n14145) );
  INV_X1 U7468 ( .A(n12882), .ZN(n12866) );
  NAND2_X2 U7469 ( .A1(n8555), .A2(n14947), .ZN(n10562) );
  XNOR2_X1 U7470 ( .A(n14692), .B(n14548), .ZN(n14685) );
  XNOR2_X1 U7471 ( .A(n7872), .B(n7871), .ZN(n12179) );
  INV_X2 U7472 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9392) );
  AOI21_X1 U7473 ( .B1(n13299), .B2(n15503), .A(n13280), .ZN(n13281) );
  INV_X1 U7474 ( .A(n15389), .ZN(n13800) );
  AND3_X1 U7475 ( .A1(n8352), .A2(n6817), .A3(n8351), .ZN(n6674) );
  NAND2_X2 U7476 ( .A1(n11408), .A2(n15384), .ZN(n15392) );
  OR2_X2 U7477 ( .A1(n13174), .A2(n13175), .ZN(n7332) );
  OR2_X2 U7478 ( .A1(n9983), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9997) );
  NAND2_X2 U7479 ( .A1(n14631), .A2(n14630), .ZN(n14629) );
  NAND2_X2 U7480 ( .A1(n14642), .A2(n7750), .ZN(n14631) );
  NAND2_X2 U7483 ( .A1(n11106), .A2(n11105), .ZN(n11104) );
  AOI21_X2 U7484 ( .B1(n7431), .B2(n7435), .A(n7432), .ZN(n13986) );
  OAI21_X2 U7485 ( .B1(n11775), .B2(n11459), .A(n11460), .ZN(n11830) );
  NAND2_X2 U7486 ( .A1(n7440), .A2(n11458), .ZN(n11775) );
  XNOR2_X2 U7487 ( .A(n8589), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8590) );
  AOI21_X2 U7488 ( .B1(n9160), .B2(n9155), .A(n9159), .ZN(n9156) );
  OAI21_X2 U7489 ( .B1(n8204), .B2(n7546), .A(n7544), .ZN(n7858) );
  OAI222_X1 U7490 ( .A1(n12975), .A2(P3_U3151), .B1(n13672), .B2(n12974), .C1(
        n12973), .C2(n12971), .ZN(P3_U3265) );
  XNOR2_X2 U7491 ( .A(n9606), .B(n9605), .ZN(n12975) );
  AOI21_X2 U7492 ( .B1(n14341), .B2(n14342), .A(n6969), .ZN(n14294) );
  OR2_X2 U7493 ( .A1(n15030), .A2(n10013), .ZN(n13337) );
  NAND2_X2 U7494 ( .A1(n8719), .A2(n8718), .ZN(n15429) );
  OAI21_X2 U7495 ( .B1(n10381), .B2(n10380), .A(n14287), .ZN(n14341) );
  OAI21_X2 U7496 ( .B1(n14629), .B2(n7385), .A(n7381), .ZN(n14586) );
  NAND2_X1 U7497 ( .A1(n10537), .A2(n8484), .ZN(n7965) );
  AOI21_X2 U7498 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n9174), .A(n14963), .ZN(
        n15706) );
  NAND2_X2 U7499 ( .A1(n8496), .A2(n8495), .ZN(n11143) );
  NAND2_X2 U7500 ( .A1(n8983), .A2(n8982), .ZN(n13748) );
  NAND2_X2 U7501 ( .A1(n11002), .A2(n8715), .ZN(n11009) );
  NAND2_X2 U7502 ( .A1(n11003), .A2(n11004), .ZN(n11002) );
  INV_X2 U7503 ( .A(n8597), .ZN(n12606) );
  INV_X4 U7504 ( .A(n12674), .ZN(n12844) );
  NAND2_X4 U7505 ( .A1(n12645), .A2(n12926), .ZN(n12674) );
  XNOR2_X2 U7506 ( .A(n7907), .B(n7906), .ZN(n10598) );
  XNOR2_X2 U7507 ( .A(n13203), .B(n13204), .ZN(n13176) );
  AND2_X2 U7508 ( .A1(n7330), .A2(n7329), .ZN(n13203) );
  XNOR2_X2 U7509 ( .A(n9568), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9810) );
  INV_X1 U7510 ( .A(n12857), .ZN(n12846) );
  XNOR2_X2 U7511 ( .A(n8158), .B(n8110), .ZN(n10938) );
  XNOR2_X2 U7512 ( .A(n8109), .B(n10577), .ZN(n8158) );
  XNOR2_X2 U7513 ( .A(n9581), .B(n12212), .ZN(n9956) );
  AOI21_X2 U7514 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(n9137), .A(n9136), .ZN(
        n9139) );
  NAND2_X1 U7515 ( .A1(n14259), .A2(n14260), .ZN(n14258) );
  AND2_X1 U7516 ( .A1(n10196), .A2(n10195), .ZN(n13376) );
  CLKBUF_X1 U7517 ( .A(n14378), .Z(n6996) );
  OR2_X1 U7518 ( .A1(n7625), .A2(n9967), .ZN(n7624) );
  OR2_X1 U7519 ( .A1(n14993), .A2(n15130), .ZN(n12404) );
  NAND2_X1 U7520 ( .A1(n7830), .A2(n7829), .ZN(n8066) );
  INV_X4 U7521 ( .A(n13030), .ZN(n12598) );
  INV_X2 U7522 ( .A(n15120), .ZN(n6676) );
  NAND4_X1 U7523 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n15612)
         );
  INV_X2 U7524 ( .A(n8031), .ZN(n8442) );
  INV_X2 U7525 ( .A(n12844), .ZN(n12787) );
  NAND4_X2 U7526 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n14411)
         );
  AND2_X2 U7527 ( .A1(n10702), .A2(n12018), .ZN(n15209) );
  INV_X1 U7528 ( .A(n13794), .ZN(n12706) );
  AND2_X1 U7529 ( .A1(n10969), .A2(n10967), .ZN(n12899) );
  INV_X1 U7530 ( .A(n13796), .ZN(n12692) );
  INV_X1 U7531 ( .A(n14953), .ZN(n10479) );
  INV_X2 U7532 ( .A(n8457), .ZN(n8484) );
  INV_X1 U7533 ( .A(n14806), .ZN(n11046) );
  BUF_X1 U7534 ( .A(n7789), .Z(n12638) );
  BUF_X2 U7535 ( .A(n8656), .Z(n12868) );
  INV_X1 U7536 ( .A(n10698), .ZN(n6679) );
  NOR2_X1 U7538 ( .A1(n7873), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7785) );
  OAI21_X1 U7539 ( .B1(n8545), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7876) );
  OR2_X1 U7540 ( .A1(n9764), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9777) );
  INV_X4 U7541 ( .A(n10501), .ZN(n10497) );
  AOI22_X1 U7542 ( .A1(n7335), .A2(P3_IR_REG_0__SCAN_IN), .B1(n6873), .B2(
        n7334), .ZN(n7333) );
  CLKBUF_X2 U7543 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14955) );
  OAI21_X1 U7544 ( .B1(n10060), .B2(n11498), .A(n6943), .ZN(n7637) );
  NAND2_X1 U7545 ( .A1(n6945), .A2(n10067), .ZN(n13347) );
  AOI21_X1 U7546 ( .B1(n13029), .B2(n13028), .A(n6786), .ZN(n13032) );
  XNOR2_X1 U7547 ( .A(n12979), .B(n12982), .ZN(n13103) );
  OAI21_X1 U7548 ( .B1(n9955), .B2(n10190), .A(n7648), .ZN(n13375) );
  INV_X1 U7549 ( .A(n13020), .ZN(n6890) );
  NAND2_X1 U7550 ( .A1(n13123), .A2(n6822), .ZN(n13020) );
  AOI21_X1 U7551 ( .B1(n7302), .B2(n7306), .A(n6778), .ZN(n7300) );
  OR2_X1 U7552 ( .A1(n6851), .A2(n6850), .ZN(n6849) );
  NAND2_X1 U7553 ( .A1(n10011), .A2(n10010), .ZN(n12515) );
  AND2_X1 U7554 ( .A1(n7562), .A2(n7561), .ZN(n7560) );
  NAND2_X1 U7555 ( .A1(n8460), .A2(n8459), .ZN(n14533) );
  NAND2_X1 U7556 ( .A1(n12861), .A2(n12860), .ZN(n13876) );
  NAND2_X1 U7557 ( .A1(n13077), .A2(n12585), .ZN(n13125) );
  NAND2_X1 U7558 ( .A1(n13958), .A2(n13957), .ZN(n13956) );
  NAND2_X1 U7559 ( .A1(n13068), .A2(n12582), .ZN(n13079) );
  NAND2_X1 U7561 ( .A1(n13070), .A2(n13069), .ZN(n13068) );
  AOI21_X1 U7562 ( .B1(n13306), .B2(n15550), .A(n13305), .ZN(n7561) );
  XNOR2_X1 U7563 ( .A(n8448), .B(n8447), .ZN(n14239) );
  NAND2_X1 U7564 ( .A1(n13000), .A2(n12576), .ZN(n13147) );
  NAND2_X1 U7565 ( .A1(n9053), .A2(n9052), .ZN(n14149) );
  XNOR2_X1 U7566 ( .A(n8437), .B(n8436), .ZN(n14242) );
  AND2_X1 U7567 ( .A1(n7158), .A2(n7160), .ZN(n8260) );
  NAND2_X1 U7568 ( .A1(n9836), .A2(n10142), .ZN(n13519) );
  OAI21_X1 U7569 ( .B1(n8415), .B2(n8414), .A(n8417), .ZN(n8437) );
  NAND2_X1 U7570 ( .A1(n7244), .A2(n8364), .ZN(n8381) );
  NAND2_X1 U7571 ( .A1(n7048), .A2(n8987), .ZN(n14180) );
  NAND2_X1 U7572 ( .A1(n11620), .A2(n8830), .ZN(n11938) );
  OR2_X1 U7573 ( .A1(n8074), .A2(n8075), .ZN(n8076) );
  NAND2_X1 U7574 ( .A1(n9006), .A2(n9005), .ZN(n14175) );
  XNOR2_X1 U7575 ( .A(n8363), .B(SI_24_), .ZN(n8360) );
  NAND2_X1 U7576 ( .A1(n7636), .A2(n9577), .ZN(n9578) );
  NAND2_X1 U7577 ( .A1(n12246), .A2(n6908), .ZN(n12566) );
  NAND2_X1 U7578 ( .A1(n9762), .A2(n7745), .ZN(n7660) );
  XNOR2_X1 U7579 ( .A(n8165), .B(n8164), .ZN(n11015) );
  NAND2_X1 U7580 ( .A1(n7017), .A2(n7015), .ZN(n9889) );
  NAND2_X1 U7581 ( .A1(n8113), .A2(n8112), .ZN(n14921) );
  NAND2_X1 U7582 ( .A1(n9716), .A2(n10107), .ZN(n11958) );
  AND2_X1 U7583 ( .A1(n7859), .A2(n7055), .ZN(n7054) );
  AND2_X1 U7584 ( .A1(n15558), .A2(n11723), .ZN(n11725) );
  OAI21_X1 U7585 ( .B1(n14978), .B2(n14979), .A(n7279), .ZN(n6920) );
  NAND2_X1 U7586 ( .A1(n7058), .A2(n7056), .ZN(n8204) );
  AND2_X2 U7587 ( .A1(n15392), .A2(n13871), .ZN(n14108) );
  NAND2_X1 U7588 ( .A1(n8093), .A2(n8092), .ZN(n15284) );
  NAND2_X1 U7589 ( .A1(n8777), .A2(n8776), .ZN(n15449) );
  NAND2_X1 U7590 ( .A1(n8066), .A2(n7831), .ZN(n7834) );
  AOI21_X1 U7591 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n9143), .A(n9142), .ZN(
        n9196) );
  AND2_X1 U7592 ( .A1(n10087), .A2(n10091), .ZN(n11502) );
  NAND2_X1 U7593 ( .A1(n10095), .A2(n10098), .ZN(n15576) );
  NAND2_X2 U7594 ( .A1(n14590), .A2(n15117), .ZN(n15120) );
  NAND2_X2 U7595 ( .A1(n10488), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15090) );
  XNOR2_X1 U7596 ( .A(n12169), .B(n12083), .ZN(n12057) );
  INV_X1 U7597 ( .A(n15491), .ZN(n15595) );
  INV_X1 U7598 ( .A(n15596), .ZN(n15573) );
  NAND2_X1 U7599 ( .A1(n6877), .A2(n6875), .ZN(n11394) );
  XNOR2_X1 U7600 ( .A(n8653), .B(n14213), .ZN(n8638) );
  CLKBUF_X3 U7601 ( .A(n8653), .Z(n13693) );
  NAND2_X1 U7602 ( .A1(n8684), .A2(n8683), .ZN(n15417) );
  NAND4_X2 U7603 ( .A1(n7958), .A2(n7957), .A3(n7956), .A4(n7955), .ZN(n14406)
         );
  NAND2_X1 U7604 ( .A1(n6966), .A2(n15209), .ZN(n14710) );
  INV_X1 U7605 ( .A(n11393), .ZN(n15588) );
  INV_X1 U7606 ( .A(n6976), .ZN(n15239) );
  NOR2_X1 U7607 ( .A1(n11594), .A2(n11606), .ZN(n11760) );
  NAND4_X1 U7608 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n14408)
         );
  BUF_X1 U7609 ( .A(n10241), .Z(n14410) );
  NAND2_X1 U7610 ( .A1(n8669), .A2(n6846), .ZN(n15410) );
  AND2_X4 U7611 ( .A1(n9612), .A2(n9611), .ZN(n9816) );
  NAND2_X2 U7612 ( .A1(n10699), .A2(n10698), .ZN(n10701) );
  CLKBUF_X1 U7613 ( .A(n8198), .Z(n8465) );
  INV_X2 U7614 ( .A(n8468), .ZN(n8461) );
  NAND2_X1 U7615 ( .A1(n15380), .A2(n12897), .ZN(n14018) );
  INV_X1 U7617 ( .A(n8466), .ZN(n8198) );
  NAND2_X1 U7618 ( .A1(n11566), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11677) );
  NAND2_X2 U7619 ( .A1(n12638), .A2(n7790), .ZN(n8468) );
  NAND2_X1 U7620 ( .A1(n14953), .A2(n6966), .ZN(n10699) );
  NAND2_X1 U7621 ( .A1(n11362), .A2(n12621), .ZN(n11361) );
  MUX2_X1 U7622 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9609), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9610) );
  NAND2_X1 U7623 ( .A1(n11578), .A2(n11577), .ZN(n11681) );
  CLKBUF_X1 U7624 ( .A(n8611), .Z(n12862) );
  AND2_X1 U7625 ( .A1(n11565), .A2(n11675), .ZN(n11566) );
  MUX2_X1 U7626 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10033), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n10036) );
  OAI21_X1 U7627 ( .B1(n10219), .B2(n9595), .A(n7014), .ZN(n10222) );
  NAND2_X1 U7628 ( .A1(n9065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U7629 ( .A1(n13664), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9606) );
  NOR2_X1 U7630 ( .A1(n10218), .A2(n10217), .ZN(n11329) );
  NAND2_X1 U7631 ( .A1(n8537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7890) );
  AND2_X1 U7632 ( .A1(n8551), .A2(n6716), .ZN(n10463) );
  XNOR2_X1 U7633 ( .A(n7883), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10703) );
  XNOR2_X1 U7634 ( .A(n7810), .B(n7242), .ZN(n7809) );
  XNOR2_X1 U7635 ( .A(n7787), .B(n7786), .ZN(n7788) );
  NAND2_X1 U7636 ( .A1(n7243), .A2(n7807), .ZN(n7810) );
  XNOR2_X1 U7637 ( .A(n7888), .B(P1_IR_REG_19__SCAN_IN), .ZN(n8263) );
  AOI21_X1 U7638 ( .B1(n10224), .B2(P3_IR_REG_24__SCAN_IN), .A(n7035), .ZN(
        n7034) );
  XNOR2_X1 U7639 ( .A(n7876), .B(n7782), .ZN(n14947) );
  OAI21_X1 U7640 ( .B1(n8166), .B2(n7195), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7888) );
  XNOR2_X1 U7641 ( .A(n8620), .B(P2_IR_REG_19__SCAN_IN), .ZN(n12926) );
  XNOR2_X1 U7642 ( .A(n9598), .B(n9597), .ZN(n12561) );
  OAI21_X1 U7643 ( .B1(n6911), .B2(n6779), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9598) );
  OR2_X1 U7645 ( .A1(n8606), .A2(n8588), .ZN(n8608) );
  OR2_X1 U7646 ( .A1(n7885), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U7647 ( .A1(n9857), .A2(n9856), .ZN(n9859) );
  NAND2_X1 U7648 ( .A1(n7925), .A2(n7924), .ZN(n14429) );
  AND2_X1 U7649 ( .A1(n9800), .A2(n6807), .ZN(n9857) );
  CLKBUF_X1 U7650 ( .A(n7884), .Z(n7885) );
  INV_X1 U7651 ( .A(n7884), .ZN(n7777) );
  AND2_X1 U7652 ( .A1(n8585), .A2(n7692), .ZN(n8615) );
  AND2_X1 U7653 ( .A1(n7776), .A2(n7588), .ZN(n7587) );
  AND2_X1 U7654 ( .A1(n8585), .A2(n8586), .ZN(n8606) );
  NAND2_X1 U7655 ( .A1(n7802), .A2(n7803), .ZN(n7808) );
  AND3_X1 U7656 ( .A1(n8584), .A2(n6844), .A3(n6801), .ZN(n8586) );
  AND2_X1 U7657 ( .A1(n6889), .A2(n6888), .ZN(n6884) );
  AND2_X1 U7658 ( .A1(n6880), .A2(n6879), .ZN(n6882) );
  AND3_X1 U7659 ( .A1(n8618), .A2(n6859), .A3(n6858), .ZN(n8584) );
  AND4_X1 U7660 ( .A1(n10061), .A2(n10034), .A3(n10032), .A4(n10031), .ZN(
        n9592) );
  AND2_X1 U7661 ( .A1(n8647), .A2(n8562), .ZN(n8667) );
  AND4_X1 U7662 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8569), .ZN(n6844)
         );
  AND4_X1 U7663 ( .A1(n7772), .A2(n7771), .A3(n8089), .A4(n7770), .ZN(n7773)
         );
  AND2_X1 U7664 ( .A1(n9546), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9652) );
  AND4_X1 U7665 ( .A1(n7775), .A2(n7774), .A3(n9493), .A4(n9298), .ZN(n7776)
         );
  AND4_X1 U7666 ( .A1(n8565), .A2(n8564), .A3(n8736), .A4(n8563), .ZN(n8566)
         );
  NAND4_X1 U7667 ( .A1(n7798), .A2(n7797), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7803) );
  AND4_X1 U7668 ( .A1(n8561), .A2(n8560), .A3(n8680), .A4(n8559), .ZN(n8567)
         );
  XNOR2_X1 U7669 ( .A(n6919), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n9167) );
  NOR2_X1 U7670 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n7765) );
  NOR2_X1 U7671 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7766) );
  INV_X1 U7672 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6873) );
  XNOR2_X1 U7673 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9653) );
  INV_X1 U7674 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7801) );
  INV_X1 U7675 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7798) );
  INV_X1 U7676 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7797) );
  NOR2_X1 U7677 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9689) );
  INV_X1 U7678 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6919) );
  INV_X1 U7679 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n6918) );
  INV_X1 U7680 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6917) );
  NOR2_X1 U7681 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7774) );
  NOR2_X1 U7682 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n7775) );
  INV_X1 U7683 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7881) );
  NOR2_X1 U7684 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n6916) );
  NOR2_X1 U7685 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n6889) );
  NOR2_X1 U7686 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n6888) );
  CLKBUF_X1 U7687 ( .A(P2_IR_REG_22__SCAN_IN), .Z(n9066) );
  INV_X1 U7688 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U7689 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6880) );
  INV_X1 U7690 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n10034) );
  INV_X1 U7691 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8736) );
  INV_X4 U7692 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7693 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6879) );
  NOR2_X1 U7694 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8561) );
  INV_X1 U7695 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n10061) );
  NOR2_X2 U7696 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8618) );
  OAI21_X2 U7697 ( .B1(n7630), .B2(n7228), .A(n7226), .ZN(n9582) );
  AND2_X1 U7698 ( .A1(n8579), .A2(n8578), .ZN(n10971) );
  NAND2_X1 U7699 ( .A1(n15187), .A2(n15186), .ZN(n15185) );
  NAND2_X1 U7700 ( .A1(n8613), .A2(n8612), .ZN(n12644) );
  OAI21_X2 U7701 ( .B1(n7680), .B2(n7682), .A(n7681), .ZN(n12820) );
  OR2_X1 U7702 ( .A1(n12758), .A2(n7143), .ZN(n7138) );
  NAND2_X2 U7703 ( .A1(n11938), .A2(n11939), .ZN(n11937) );
  NOR2_X2 U7704 ( .A1(n11795), .A2(n15423), .ZN(n11837) );
  INV_X1 U7705 ( .A(n8031), .ZN(n6680) );
  NAND2_X2 U7706 ( .A1(n7788), .A2(n7694), .ZN(n8469) );
  NAND2_X2 U7707 ( .A1(n13704), .A2(n9002), .ZN(n9015) );
  AND2_X1 U7708 ( .A1(n8612), .A2(n12862), .ZN(n15380) );
  NOR2_X2 U7709 ( .A1(n12500), .A2(n14207), .ZN(n14112) );
  NOR2_X4 U7710 ( .A1(n14707), .A2(n14872), .ZN(n14687) );
  NOR2_X2 U7711 ( .A1(n14016), .A2(n14165), .ZN(n14007) );
  XNOR2_X2 U7712 ( .A(n8605), .B(n8604), .ZN(n10782) );
  NAND2_X1 U7713 ( .A1(n14866), .A2(n14576), .ZN(n7713) );
  AND2_X1 U7714 ( .A1(n8568), .A2(n7693), .ZN(n7692) );
  INV_X1 U7715 ( .A(n12641), .ZN(n9611) );
  NAND2_X1 U7716 ( .A1(n10371), .A2(n10370), .ZN(n7609) );
  NAND2_X1 U7717 ( .A1(n14674), .A2(n6756), .ZN(n7378) );
  AOI21_X1 U7718 ( .B1(n6686), .B2(n7709), .A(n6785), .ZN(n7708) );
  NOR2_X1 U7719 ( .A1(n14655), .A2(n6717), .ZN(n7709) );
  NAND2_X1 U7720 ( .A1(n6686), .A2(n14661), .ZN(n7710) );
  NAND2_X1 U7721 ( .A1(n7845), .A2(n7844), .ZN(n8129) );
  NAND2_X1 U7722 ( .A1(n12566), .A2(n12565), .ZN(n12569) );
  INV_X1 U7723 ( .A(n13126), .ZN(n6991) );
  INV_X1 U7724 ( .A(n13125), .ZN(n6912) );
  NAND2_X1 U7725 ( .A1(n9611), .A2(n12975), .ZN(n10024) );
  NOR2_X1 U7726 ( .A1(n13267), .A2(n13266), .ZN(n13284) );
  AND2_X1 U7727 ( .A1(n13775), .A2(n9047), .ZN(n7481) );
  CLKBUF_X1 U7728 ( .A(n8430), .Z(n6972) );
  CLKBUF_X1 U7729 ( .A(n8469), .Z(n6973) );
  NAND2_X1 U7730 ( .A1(n14978), .A2(n14979), .ZN(n14977) );
  AOI21_X1 U7731 ( .B1(n12727), .B2(n6698), .A(n12733), .ZN(n7125) );
  NAND2_X1 U7732 ( .A1(n7118), .A2(n7117), .ZN(n7116) );
  INV_X1 U7733 ( .A(n12776), .ZN(n7117) );
  NAND2_X1 U7734 ( .A1(n7119), .A2(n12777), .ZN(n7118) );
  NAND2_X1 U7735 ( .A1(n7675), .A2(n7115), .ZN(n7114) );
  INV_X1 U7736 ( .A(n12777), .ZN(n7115) );
  INV_X1 U7737 ( .A(n7113), .ZN(n7112) );
  INV_X1 U7738 ( .A(n12792), .ZN(n7149) );
  INV_X1 U7739 ( .A(n12808), .ZN(n7688) );
  INV_X1 U7740 ( .A(n12809), .ZN(n7689) );
  AOI21_X1 U7741 ( .B1(n6763), .B2(n10207), .A(n6982), .ZN(n10209) );
  NAND2_X1 U7742 ( .A1(n7633), .A2(n12624), .ZN(n7632) );
  NAND2_X1 U7743 ( .A1(n15040), .A2(n12545), .ZN(n7633) );
  INV_X1 U7744 ( .A(n9570), .ZN(n7622) );
  OAI21_X1 U7745 ( .B1(n7703), .B2(n7701), .A(n12343), .ZN(n7700) );
  OAI21_X1 U7746 ( .B1(n9175), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6726), .ZN(
        n6926) );
  NAND2_X1 U7747 ( .A1(n6684), .A2(n12590), .ZN(n6894) );
  AOI21_X1 U7748 ( .B1(n6684), .B2(n7394), .A(n6820), .ZN(n7393) );
  INV_X1 U7749 ( .A(n13085), .ZN(n7394) );
  OR2_X1 U7750 ( .A1(n13378), .A2(n12992), .ZN(n10196) );
  AND2_X1 U7751 ( .A1(n7651), .A2(n10185), .ZN(n7650) );
  AND2_X1 U7752 ( .A1(n10162), .A2(n13508), .ZN(n7659) );
  NOR2_X1 U7753 ( .A1(n13477), .A2(n7656), .ZN(n7655) );
  INV_X1 U7754 ( .A(n7658), .ZN(n7656) );
  AND3_X1 U7755 ( .A1(n9637), .A2(n6915), .A3(n6797), .ZN(n11393) );
  NAND2_X1 U7756 ( .A1(n9805), .A2(n10521), .ZN(n6915) );
  NAND2_X1 U7757 ( .A1(n15608), .A2(n15491), .ZN(n10080) );
  OR2_X1 U7758 ( .A1(n9859), .A2(n6906), .ZN(n10038) );
  NAND2_X1 U7759 ( .A1(n7397), .A2(n6907), .ZN(n6906) );
  INV_X1 U7760 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6907) );
  AND2_X1 U7761 ( .A1(n6789), .A2(n10031), .ZN(n7397) );
  NOR2_X1 U7762 ( .A1(n9859), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U7763 ( .A1(n6775), .A2(n12828), .ZN(n7677) );
  OAI211_X1 U7764 ( .C1(n12893), .C2(n12936), .A(n6724), .B(n12937), .ZN(
        n12943) );
  NOR2_X1 U7765 ( .A1(n14180), .A2(n14031), .ZN(n7427) );
  NOR2_X1 U7766 ( .A1(n7427), .A2(n7424), .ZN(n7423) );
  INV_X1 U7767 ( .A(n7425), .ZN(n7424) );
  AND2_X1 U7768 ( .A1(n11444), .A2(n6861), .ZN(n7492) );
  NAND2_X1 U7769 ( .A1(n11829), .A2(n11443), .ZN(n6861) );
  AND2_X1 U7770 ( .A1(n12909), .A2(n11464), .ZN(n7444) );
  OR2_X1 U7771 ( .A1(n9079), .A2(n14255), .ZN(n9095) );
  OR2_X1 U7772 ( .A1(n9065), .A2(n9066), .ZN(n9082) );
  XNOR2_X1 U7773 ( .A(n14837), .B(n14550), .ZN(n14583) );
  NOR2_X1 U7774 ( .A1(n14537), .A2(n7742), .ZN(n7741) );
  INV_X1 U7775 ( .A(n12408), .ZN(n7742) );
  OR2_X1 U7776 ( .A1(n14921), .A2(n14560), .ZN(n14535) );
  INV_X1 U7777 ( .A(n14983), .ZN(n7355) );
  INV_X1 U7778 ( .A(n12351), .ZN(n7361) );
  NOR2_X1 U7779 ( .A1(n12033), .A2(n6687), .ZN(n7703) );
  AND2_X1 U7780 ( .A1(n14583), .A2(n14581), .ZN(n7387) );
  OAI21_X1 U7781 ( .B1(n11207), .B2(n7729), .A(n7727), .ZN(n11304) );
  INV_X1 U7782 ( .A(n7728), .ZN(n7727) );
  OAI21_X1 U7783 ( .B1(n7730), .B2(n7729), .A(n11305), .ZN(n7728) );
  INV_X1 U7784 ( .A(n11277), .ZN(n7729) );
  AND2_X1 U7785 ( .A1(n7780), .A2(n7781), .ZN(n7743) );
  OAI21_X2 U7786 ( .B1(n8381), .B2(n8380), .A(n8382), .ZN(n8397) );
  INV_X1 U7787 ( .A(n7779), .ZN(n7588) );
  AOI21_X1 U7788 ( .B1(n7060), .B2(n7062), .A(n7057), .ZN(n7056) );
  NAND2_X1 U7789 ( .A1(n8129), .A2(n7060), .ZN(n7058) );
  INV_X1 U7790 ( .A(n7061), .ZN(n7060) );
  AND2_X1 U7791 ( .A1(n7538), .A2(n7840), .ZN(n7537) );
  XNOR2_X1 U7792 ( .A(n6926), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U7793 ( .A(n9132), .B(n9133), .ZN(n9179) );
  NOR2_X1 U7794 ( .A1(n12101), .A2(n7389), .ZN(n7392) );
  XNOR2_X1 U7795 ( .A(n12045), .B(n11394), .ZN(n12046) );
  XNOR2_X1 U7796 ( .A(n12598), .B(n15581), .ZN(n12049) );
  NAND2_X1 U7797 ( .A1(n10057), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U7798 ( .A1(n12549), .A2(n10204), .ZN(n7663) );
  AND4_X1 U7799 ( .A1(n6733), .A2(n10057), .A3(n10210), .A4(n7747), .ZN(n10058) );
  AND2_X1 U7800 ( .A1(n9587), .A2(n6886), .ZN(n6885) );
  INV_X1 U7801 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U7802 ( .A1(n15517), .A2(n11857), .ZN(n7339) );
  OR2_X1 U7803 ( .A1(n13191), .A2(n13192), .ZN(n7551) );
  NAND2_X1 U7804 ( .A1(n7551), .A2(n7550), .ZN(n15543) );
  INV_X1 U7805 ( .A(n15545), .ZN(n7550) );
  XNOR2_X1 U7806 ( .A(n13200), .B(n13204), .ZN(n13194) );
  INV_X1 U7807 ( .A(n12541), .ZN(n7312) );
  OAI21_X1 U7808 ( .B1(n13436), .B2(n7290), .A(n7286), .ZN(n13411) );
  AOI21_X1 U7809 ( .B1(n7289), .B2(n13443), .A(n6762), .ZN(n7286) );
  NAND2_X1 U7810 ( .A1(n12517), .A2(n12516), .ZN(n12519) );
  AND4_X1 U7811 ( .A1(n9659), .A2(n9660), .A3(n9658), .A4(n9657), .ZN(n15596)
         );
  NAND2_X1 U7812 ( .A1(n11532), .A2(n10230), .ZN(n15594) );
  NAND2_X1 U7813 ( .A1(n10724), .A2(n11329), .ZN(n11344) );
  AOI21_X1 U7814 ( .B1(n10009), .B2(n7236), .A(n7234), .ZN(n7233) );
  NAND2_X1 U7815 ( .A1(n7235), .A2(n9618), .ZN(n7234) );
  NAND2_X1 U7816 ( .A1(n7236), .A2(n7237), .ZN(n7235) );
  NAND2_X1 U7817 ( .A1(n9800), .A2(n6910), .ZN(n6911) );
  NOR2_X1 U7818 ( .A1(n9593), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n6910) );
  OAI22_X1 U7819 ( .A1(n9980), .A2(n9583), .B1(P1_DATAO_REG_26__SCAN_IN), .B2(
        n14950), .ZN(n9994) );
  OR2_X1 U7820 ( .A1(n9936), .A2(n9935), .ZN(n7630) );
  OR2_X1 U7821 ( .A1(n9032), .A2(n9033), .ZN(n7485) );
  INV_X1 U7822 ( .A(n12839), .ZN(n7674) );
  AND2_X1 U7823 ( .A1(n8590), .A2(n12606), .ZN(n8655) );
  INV_X1 U7824 ( .A(n7414), .ZN(n7413) );
  OAI22_X1 U7825 ( .A1(n13940), .A2(n7419), .B1(n13903), .B2(n13937), .ZN(
        n7414) );
  NAND2_X1 U7826 ( .A1(n13939), .A2(n13927), .ZN(n7506) );
  INV_X1 U7827 ( .A(n7433), .ZN(n7432) );
  AOI21_X1 U7828 ( .B1(n7435), .B2(n7434), .A(n6791), .ZN(n7433) );
  AOI21_X1 U7829 ( .B1(n7496), .B2(n6842), .A(n6703), .ZN(n7072) );
  NOR2_X1 U7830 ( .A1(n14075), .A2(n7493), .ZN(n6842) );
  BUF_X1 U7831 ( .A(n8646), .Z(n12879) );
  AOI21_X1 U7832 ( .B1(n7496), .B2(n7495), .A(n6771), .ZN(n7494) );
  INV_X1 U7833 ( .A(n7501), .ZN(n7495) );
  NAND2_X1 U7834 ( .A1(n14075), .A2(n7501), .ZN(n7498) );
  OR2_X1 U7835 ( .A1(n14191), .A2(n13892), .ZN(n7428) );
  NAND2_X1 U7836 ( .A1(n14073), .A2(n6749), .ZN(n13891) );
  NAND2_X1 U7837 ( .A1(n7507), .A2(n7518), .ZN(n7517) );
  NAND2_X1 U7838 ( .A1(n7521), .A2(n7520), .ZN(n7507) );
  INV_X2 U7839 ( .A(n8916), .ZN(n10747) );
  OR2_X1 U7840 ( .A1(n11817), .A2(n11463), .ZN(n11465) );
  INV_X1 U7841 ( .A(n14090), .ZN(n14124) );
  INV_X1 U7842 ( .A(n7411), .ZN(n7408) );
  NOR2_X1 U7843 ( .A1(n10964), .A2(n10963), .ZN(n12122) );
  OR2_X1 U7844 ( .A1(n12176), .A2(n9084), .ZN(n15396) );
  INV_X1 U7845 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8607) );
  AND2_X1 U7846 ( .A1(n10386), .A2(n10387), .ZN(n6969) );
  NAND2_X1 U7847 ( .A1(n6794), .A2(n7609), .ZN(n7605) );
  NAND2_X1 U7848 ( .A1(n7609), .A2(n7607), .ZN(n7606) );
  INV_X1 U7849 ( .A(n14318), .ZN(n7607) );
  CLKBUF_X1 U7850 ( .A(n8468), .Z(n6970) );
  AND4_X1 U7851 ( .A1(n8084), .A2(n8083), .A3(n8082), .A4(n8081), .ZN(n15096)
         );
  AND4_X1 U7852 ( .A1(n8023), .A2(n8022), .A3(n8021), .A4(n8020), .ZN(n11518)
         );
  NAND2_X1 U7853 ( .A1(n8441), .A2(n8440), .ZN(n14822) );
  OR2_X1 U7854 ( .A1(n7266), .A2(n14579), .ZN(n7750) );
  XNOR2_X1 U7855 ( .A(n14843), .B(n14309), .ZN(n14630) );
  INV_X1 U7856 ( .A(n7713), .ZN(n7711) );
  NAND2_X1 U7857 ( .A1(n14673), .A2(n14672), .ZN(n14674) );
  OR2_X1 U7858 ( .A1(n14877), .A2(n14546), .ZN(n14547) );
  AOI21_X1 U7859 ( .B1(n7753), .B2(n7375), .A(n6769), .ZN(n7374) );
  OAI21_X1 U7860 ( .B1(n14561), .B2(n14560), .A(n14559), .ZN(n14786) );
  INV_X1 U7861 ( .A(n10562), .ZN(n8264) );
  NAND2_X1 U7862 ( .A1(n12514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7783) );
  INV_X2 U7863 ( .A(n7808), .ZN(n10501) );
  XNOR2_X1 U7864 ( .A(n8025), .B(n8024), .ZN(n10564) );
  NAND2_X1 U7865 ( .A1(n7529), .A2(n7825), .ZN(n8025) );
  NAND2_X1 U7866 ( .A1(n7993), .A2(n7823), .ZN(n7529) );
  XOR2_X1 U7867 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9172) );
  OAI21_X1 U7868 ( .B1(n9197), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n9147), .ZN(
        n9165) );
  AOI21_X1 U7869 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n13218), .A(n9154), .ZN(
        n9160) );
  NOR2_X1 U7870 ( .A1(n9163), .A2(n9162), .ZN(n9154) );
  NAND2_X1 U7871 ( .A1(n6898), .A2(n6897), .ZN(n13029) );
  AOI21_X1 U7872 ( .B1(n6900), .B2(n6903), .A(n6770), .ZN(n6897) );
  NAND2_X1 U7873 ( .A1(n13060), .A2(n6900), .ZN(n6898) );
  NAND2_X1 U7874 ( .A1(n9948), .A2(n9947), .ZN(n13015) );
  NOR2_X1 U7875 ( .A1(n12248), .A2(n6909), .ZN(n6908) );
  INV_X1 U7876 ( .A(n12245), .ZN(n6909) );
  INV_X1 U7877 ( .A(n13018), .ZN(n12588) );
  NAND2_X1 U7878 ( .A1(n15539), .A2(n6834), .ZN(n7324) );
  AOI21_X1 U7879 ( .B1(n7083), .B2(n15550), .A(n7080), .ZN(n7079) );
  OR2_X1 U7880 ( .A1(n9050), .A2(n9051), .ZN(n7003) );
  NAND2_X1 U7881 ( .A1(n14159), .A2(n13783), .ZN(n7031) );
  NAND2_X1 U7882 ( .A1(n6920), .A2(n14977), .ZN(n15145) );
  INV_X1 U7883 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U7884 ( .A1(n15157), .A2(n6939), .ZN(n15162) );
  OAI21_X1 U7885 ( .B1(n15158), .B2(n15159), .A(n6940), .ZN(n6939) );
  INV_X1 U7886 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6940) );
  OAI21_X1 U7887 ( .B1(n6734), .B2(n7133), .A(n7132), .ZN(n12699) );
  NAND2_X1 U7888 ( .A1(n6776), .A2(n12693), .ZN(n7132) );
  NAND2_X1 U7889 ( .A1(n8057), .A2(n8054), .ZN(n7167) );
  AND2_X1 U7890 ( .A1(n8056), .A2(n7169), .ZN(n7168) );
  INV_X1 U7891 ( .A(n8054), .ZN(n7169) );
  OR2_X1 U7892 ( .A1(n12722), .A2(n12721), .ZN(n12728) );
  OAI21_X1 U7893 ( .B1(n12732), .B2(n7124), .A(n7123), .ZN(n7122) );
  INV_X1 U7894 ( .A(n7128), .ZN(n7124) );
  INV_X1 U7895 ( .A(n7125), .ZN(n7123) );
  AND2_X1 U7896 ( .A1(n7131), .A2(n7129), .ZN(n7126) );
  NAND2_X1 U7897 ( .A1(n7126), .A2(n7128), .ZN(n7127) );
  INV_X1 U7898 ( .A(n12757), .ZN(n7144) );
  NAND2_X1 U7899 ( .A1(n12773), .A2(n6700), .ZN(n7675) );
  NOR2_X1 U7900 ( .A1(n6722), .A2(n7144), .ZN(n7143) );
  OAI22_X1 U7901 ( .A1(n12752), .A2(n7691), .B1(n12750), .B2(n12751), .ZN(
        n12758) );
  AND2_X1 U7902 ( .A1(n12750), .A2(n12751), .ZN(n7691) );
  NAND2_X1 U7903 ( .A1(n6722), .A2(n7144), .ZN(n7142) );
  NAND2_X1 U7904 ( .A1(n7558), .A2(n7557), .ZN(n8288) );
  NAND2_X1 U7905 ( .A1(n14571), .A2(n7944), .ZN(n7557) );
  NAND2_X1 U7906 ( .A1(n10382), .A2(n6677), .ZN(n7558) );
  OAI21_X1 U7907 ( .B1(n7110), .B2(n6725), .A(n7111), .ZN(n12782) );
  OR2_X1 U7908 ( .A1(n6812), .A2(n7113), .ZN(n7111) );
  AND2_X1 U7909 ( .A1(n7570), .A2(n7180), .ZN(n7179) );
  OR2_X1 U7910 ( .A1(n8307), .A2(n7181), .ZN(n7180) );
  NOR2_X1 U7911 ( .A1(n6723), .A2(n7149), .ZN(n7148) );
  INV_X1 U7912 ( .A(n7552), .ZN(n7170) );
  NAND2_X1 U7913 ( .A1(n8370), .A2(n7553), .ZN(n7552) );
  NAND2_X1 U7914 ( .A1(n7891), .A2(n10699), .ZN(n8473) );
  NAND2_X1 U7915 ( .A1(n12803), .A2(n7154), .ZN(n7153) );
  OR2_X1 U7916 ( .A1(n12799), .A2(n12798), .ZN(n12804) );
  NAND2_X1 U7917 ( .A1(n12805), .A2(n7152), .ZN(n7151) );
  INV_X1 U7918 ( .A(n12803), .ZN(n7152) );
  NAND2_X1 U7919 ( .A1(n7687), .A2(n12814), .ZN(n7686) );
  INV_X1 U7920 ( .A(n7690), .ZN(n7687) );
  AND2_X1 U7921 ( .A1(n12808), .A2(n12809), .ZN(n7690) );
  AND2_X1 U7922 ( .A1(n6810), .A2(n7685), .ZN(n7684) );
  NAND2_X1 U7923 ( .A1(n6788), .A2(n12814), .ZN(n7685) );
  NOR2_X1 U7924 ( .A1(n12814), .A2(n6788), .ZN(n7683) );
  NAND2_X1 U7925 ( .A1(n13623), .A2(n13371), .ZN(n10187) );
  INV_X1 U7926 ( .A(n7516), .ZN(n7510) );
  AND2_X1 U7927 ( .A1(n8444), .A2(n8446), .ZN(n7536) );
  AOI21_X1 U7928 ( .B1(n7191), .B2(n7194), .A(n7189), .ZN(n7188) );
  INV_X1 U7929 ( .A(n8478), .ZN(n7189) );
  NOR2_X1 U7930 ( .A1(n8477), .A2(n7194), .ZN(n7193) );
  INV_X1 U7931 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U7932 ( .A1(n8342), .A2(n8341), .ZN(n8363) );
  NAND2_X1 U7933 ( .A1(n7860), .A2(n10831), .ZN(n7863) );
  INV_X1 U7934 ( .A(n7545), .ZN(n7544) );
  OAI21_X1 U7935 ( .B1(n8203), .B2(n7546), .A(n7856), .ZN(n7545) );
  INV_X1 U7936 ( .A(n7063), .ZN(n7062) );
  NAND2_X1 U7937 ( .A1(n7846), .A2(n10569), .ZN(n7063) );
  OR2_X1 U7938 ( .A1(n7846), .A2(n10569), .ZN(n7064) );
  AOI21_X1 U7939 ( .B1(n7992), .B2(n7825), .A(n8024), .ZN(n7530) );
  OAI21_X1 U7940 ( .B1(n10502), .B2(n10558), .A(n6963), .ZN(n7824) );
  NAND2_X1 U7941 ( .A1(n10502), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6963) );
  OR2_X1 U7942 ( .A1(n10209), .A2(n7632), .ZN(n7631) );
  OAI21_X1 U7943 ( .B1(n10209), .B2(n10208), .A(n11532), .ZN(n7634) );
  INV_X1 U7944 ( .A(n7564), .ZN(n11575) );
  NAND2_X1 U7945 ( .A1(n7043), .A2(n11606), .ZN(n6874) );
  NAND2_X1 U7946 ( .A1(n6874), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7526) );
  NOR2_X1 U7947 ( .A1(n7094), .A2(n11989), .ZN(n7093) );
  INV_X1 U7948 ( .A(n7093), .ZN(n7088) );
  NOR2_X1 U7949 ( .A1(n13245), .A2(n13246), .ZN(n13247) );
  INV_X1 U7950 ( .A(n13327), .ZN(n7082) );
  OR2_X1 U7951 ( .A1(n12515), .A2(n12996), .ZN(n10065) );
  OR2_X1 U7952 ( .A1(n13552), .A2(n9991), .ZN(n10068) );
  INV_X1 U7953 ( .A(n12532), .ZN(n7307) );
  OR2_X1 U7954 ( .A1(n13430), .A2(n13439), .ZN(n10176) );
  INV_X1 U7955 ( .A(n12520), .ZN(n7296) );
  NOR2_X1 U7956 ( .A1(n7295), .A2(n7294), .ZN(n7293) );
  INV_X1 U7957 ( .A(n7298), .ZN(n7294) );
  INV_X1 U7958 ( .A(n12526), .ZN(n7295) );
  AND2_X1 U7959 ( .A1(n13459), .A2(n10161), .ZN(n10159) );
  NAND2_X1 U7960 ( .A1(n15563), .A2(n12102), .ZN(n10098) );
  NAND2_X1 U7961 ( .A1(n10223), .A2(n7670), .ZN(n9602) );
  NAND2_X1 U7962 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), 
        .ZN(n7000) );
  AOI21_X1 U7963 ( .B1(n7620), .B2(n7622), .A(n6825), .ZN(n7618) );
  NOR2_X1 U7964 ( .A1(n7621), .A2(n7215), .ZN(n7213) );
  NAND2_X1 U7965 ( .A1(n7614), .A2(n7612), .ZN(n9568) );
  NAND2_X1 U7966 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7613), .ZN(n7612) );
  NOR2_X1 U7967 ( .A1(n7218), .A2(n6685), .ZN(n7217) );
  INV_X1 U7968 ( .A(n7221), .ZN(n7220) );
  OAI21_X1 U7969 ( .B1(n7222), .B2(n6685), .A(n9726), .ZN(n7221) );
  XNOR2_X1 U7970 ( .A(n12761), .B(n9007), .ZN(n8876) );
  INV_X1 U7971 ( .A(n8793), .ZN(n7461) );
  INV_X1 U7972 ( .A(n7480), .ZN(n7476) );
  OR4_X1 U7973 ( .A1(n14074), .A2(n14093), .A3(n12920), .A4(n12919), .ZN(
        n12921) );
  AND2_X1 U7974 ( .A1(n13928), .A2(n7023), .ZN(n7022) );
  NOR2_X1 U7975 ( .A1(n13902), .A2(n7024), .ZN(n7023) );
  NOR2_X1 U7976 ( .A1(n13998), .A2(n7070), .ZN(n7069) );
  INV_X1 U7977 ( .A(n13919), .ZN(n7070) );
  OR2_X1 U7978 ( .A1(n13998), .A2(n6739), .ZN(n7068) );
  NOR2_X1 U7979 ( .A1(n14068), .A2(n14074), .ZN(n7501) );
  INV_X1 U7980 ( .A(n7513), .ZN(n7511) );
  NAND2_X1 U7981 ( .A1(n15074), .A2(n13789), .ZN(n7516) );
  NOR2_X1 U7982 ( .A1(n15074), .A2(n13789), .ZN(n7514) );
  INV_X1 U7983 ( .A(n11443), .ZN(n6860) );
  NAND2_X1 U7984 ( .A1(n11405), .A2(n11437), .ZN(n7489) );
  AOI21_X1 U7985 ( .B1(n7599), .B2(n14350), .A(n7598), .ZN(n7597) );
  INV_X1 U7986 ( .A(n14275), .ZN(n7598) );
  NAND2_X1 U7987 ( .A1(n7188), .A2(n7190), .ZN(n7184) );
  INV_X1 U7988 ( .A(n7191), .ZN(n7190) );
  NAND2_X1 U7989 ( .A1(n7193), .A2(n7536), .ZN(n7183) );
  INV_X1 U7990 ( .A(n7188), .ZN(n7187) );
  INV_X1 U7991 ( .A(n7193), .ZN(n7186) );
  INV_X1 U7992 ( .A(n7789), .ZN(n7694) );
  INV_X1 U7993 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7772) );
  OR2_X1 U7994 ( .A1(n7708), .A2(n14643), .ZN(n7704) );
  NOR2_X1 U7995 ( .A1(n14754), .A2(n7723), .ZN(n7722) );
  INV_X1 U7996 ( .A(n14770), .ZN(n7723) );
  NOR2_X1 U7997 ( .A1(n7366), .A2(n14569), .ZN(n7365) );
  INV_X1 U7998 ( .A(n7369), .ZN(n7366) );
  NOR2_X1 U7999 ( .A1(n14754), .A2(n7721), .ZN(n7720) );
  NOR2_X1 U8000 ( .A1(n14893), .A2(n7271), .ZN(n7270) );
  NAND2_X1 U8001 ( .A1(n8244), .A2(n7272), .ZN(n7271) );
  OR2_X1 U8002 ( .A1(n11205), .A2(n11204), .ZN(n11207) );
  OR2_X1 U8003 ( .A1(n14408), .A2(n15232), .ZN(n11151) );
  AND2_X1 U8004 ( .A1(n6693), .A2(n7265), .ZN(n7264) );
  NAND2_X1 U8005 ( .A1(n14687), .A2(n6693), .ZN(n14648) );
  OAI21_X1 U8006 ( .B1(n12021), .B2(n7701), .A(n7699), .ZN(n12346) );
  INV_X1 U8007 ( .A(n7700), .ZN(n7699) );
  NAND2_X1 U8008 ( .A1(n8439), .A2(n8438), .ZN(n8448) );
  INV_X1 U8009 ( .A(n8436), .ZN(n7254) );
  INV_X1 U8010 ( .A(n8302), .ZN(n7865) );
  NAND2_X1 U8011 ( .A1(n7053), .A2(n7050), .ZN(n8298) );
  AOI21_X1 U8012 ( .B1(n7859), .B2(n7052), .A(n7051), .ZN(n7050) );
  NAND2_X1 U8013 ( .A1(n7054), .A2(n8250), .ZN(n7053) );
  INV_X1 U8014 ( .A(n7863), .ZN(n7051) );
  NAND2_X1 U8015 ( .A1(n7858), .A2(SI_18_), .ZN(n7859) );
  XNOR2_X1 U8016 ( .A(n7858), .B(SI_18_), .ZN(n8250) );
  NAND2_X1 U8017 ( .A1(n7822), .A2(n7821), .ZN(n7993) );
  XNOR2_X1 U8018 ( .A(n7814), .B(SI_3_), .ZN(n7935) );
  INV_X1 U8019 ( .A(n7005), .ZN(n9132) );
  OAI21_X1 U8020 ( .B1(n9166), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6702), .ZN(
        n7005) );
  INV_X1 U8021 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9133) );
  AOI21_X1 U8022 ( .B1(n9805), .B2(n10503), .A(n6957), .ZN(n6956) );
  NOR2_X1 U8023 ( .A1(n10229), .A2(n11569), .ZN(n6957) );
  INV_X1 U8024 ( .A(n12593), .ZN(n7395) );
  NOR2_X2 U8025 ( .A1(n15614), .A2(n12637), .ZN(n11369) );
  AOI21_X1 U8026 ( .B1(n12089), .B2(n7391), .A(n12053), .ZN(n7390) );
  INV_X1 U8027 ( .A(n12050), .ZN(n7391) );
  INV_X1 U8028 ( .A(n13540), .ZN(n11485) );
  INV_X1 U8029 ( .A(n10212), .ZN(n10211) );
  AND2_X1 U8030 ( .A1(n10027), .A2(n10026), .ZN(n13033) );
  AND4_X1 U8031 ( .A1(n9756), .A2(n9755), .A3(n9754), .A4(n9753), .ZN(n12243)
         );
  AND4_X1 U8032 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n12054)
         );
  NAND2_X1 U8033 ( .A1(n9816), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9648) );
  OAI21_X1 U8034 ( .B1(n11569), .B2(n15501), .A(n11561), .ZN(n13162) );
  XNOR2_X1 U8035 ( .A(n7564), .B(n11562), .ZN(n11740) );
  XNOR2_X1 U8036 ( .A(n7564), .B(n11574), .ZN(n11743) );
  INV_X1 U8037 ( .A(n11590), .ZN(n7103) );
  AND2_X1 U8038 ( .A1(n6692), .A2(n7102), .ZN(n7095) );
  OR2_X1 U8039 ( .A1(n11768), .A2(n11767), .ZN(n6871) );
  INV_X1 U8040 ( .A(n11762), .ZN(n7336) );
  AND2_X1 U8041 ( .A1(n7526), .A2(n7525), .ZN(n11768) );
  NAND2_X1 U8042 ( .A1(n11872), .A2(n7093), .ZN(n7090) );
  NAND2_X1 U8043 ( .A1(n6870), .A2(n6720), .ZN(n7039) );
  NAND2_X1 U8044 ( .A1(n7039), .A2(n7038), .ZN(n12257) );
  INV_X1 U8045 ( .A(n12002), .ZN(n7038) );
  NAND2_X1 U8046 ( .A1(n7332), .A2(n7331), .ZN(n7330) );
  INV_X1 U8047 ( .A(n15540), .ZN(n7331) );
  NAND2_X1 U8048 ( .A1(n15534), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U8049 ( .A1(n15549), .A2(n13183), .ZN(n13184) );
  AND2_X1 U8050 ( .A1(n15543), .A2(n13193), .ZN(n13200) );
  OR2_X1 U8051 ( .A1(n13194), .A2(n9815), .ZN(n6869) );
  OR2_X1 U8052 ( .A1(n15019), .A2(n13237), .ZN(n7078) );
  NOR2_X1 U8053 ( .A1(n13300), .A2(n13301), .ZN(n13304) );
  INV_X1 U8054 ( .A(n6872), .ZN(n13298) );
  NAND2_X1 U8055 ( .A1(n12540), .A2(n12539), .ZN(n13343) );
  INV_X1 U8056 ( .A(n7649), .ZN(n7648) );
  OAI21_X1 U8057 ( .B1(n7650), .B2(n10190), .A(n13376), .ZN(n7649) );
  NAND2_X1 U8058 ( .A1(n9955), .A2(n7650), .ZN(n13384) );
  NAND2_X1 U8059 ( .A1(n9930), .A2(n9929), .ZN(n9939) );
  AOI21_X1 U8060 ( .B1(n7655), .B2(n7653), .A(n6781), .ZN(n7652) );
  INV_X1 U8061 ( .A(n7655), .ZN(n7654) );
  NAND2_X1 U8062 ( .A1(n13457), .A2(n12528), .ZN(n13436) );
  NAND2_X1 U8063 ( .A1(n10162), .A2(n6751), .ZN(n7658) );
  NAND2_X1 U8064 ( .A1(n13509), .A2(n7659), .ZN(n7657) );
  NAND2_X1 U8065 ( .A1(n7657), .A2(n7655), .ZN(n13474) );
  AND4_X1 U8066 ( .A1(n9869), .A2(n9868), .A3(n9867), .A4(n9866), .ZN(n13517)
         );
  AND2_X1 U8067 ( .A1(n10146), .A2(n10150), .ZN(n13518) );
  NAND2_X1 U8068 ( .A1(n12481), .A2(n12480), .ZN(n12517) );
  AND4_X1 U8069 ( .A1(n9797), .A2(n9796), .A3(n9795), .A4(n9794), .ZN(n13531)
         );
  AOI21_X1 U8070 ( .B1(n7647), .B2(n12165), .A(n7643), .ZN(n7642) );
  INV_X1 U8071 ( .A(n10117), .ZN(n7643) );
  AND2_X1 U8072 ( .A1(n12217), .A2(n12216), .ZN(n12219) );
  AND2_X1 U8073 ( .A1(n9732), .A2(n9731), .ZN(n9750) );
  NAND2_X1 U8074 ( .A1(n11721), .A2(n11720), .ZN(n15577) );
  INV_X1 U8075 ( .A(n11362), .ZN(n11487) );
  OR2_X1 U8076 ( .A1(n13660), .A2(n10495), .ZN(n11529) );
  AND2_X1 U8077 ( .A1(n11532), .A2(n11354), .ZN(n15613) );
  INV_X1 U8078 ( .A(n15599), .ZN(n15619) );
  AND2_X1 U8079 ( .A1(n7207), .A2(n6839), .ZN(n15036) );
  NAND2_X1 U8080 ( .A1(n13663), .A2(n9805), .ZN(n7207) );
  AND2_X1 U8081 ( .A1(n15029), .A2(n15028), .ZN(n15039) );
  INV_X1 U8082 ( .A(n15607), .ZN(n15650) );
  NOR2_X1 U8083 ( .A1(n11481), .A2(n11346), .ZN(n12610) );
  INV_X1 U8084 ( .A(n15613), .ZN(n15597) );
  NAND2_X1 U8085 ( .A1(n13540), .A2(n11362), .ZN(n15607) );
  NAND2_X1 U8086 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7617), .ZN(n7616) );
  NAND2_X1 U8087 ( .A1(n7623), .A2(n7206), .ZN(n9980) );
  NAND2_X1 U8088 ( .A1(n7624), .A2(n7627), .ZN(n7206) );
  INV_X1 U8089 ( .A(n10227), .ZN(n10226) );
  INV_X1 U8090 ( .A(n7671), .ZN(n7669) );
  INV_X1 U8091 ( .A(n7229), .ZN(n7228) );
  AOI21_X1 U8092 ( .B1(n7229), .B2(n7227), .A(n12212), .ZN(n7226) );
  INV_X1 U8093 ( .A(n7230), .ZN(n7227) );
  NAND2_X1 U8094 ( .A1(n10223), .A2(n9594), .ZN(n10227) );
  NAND2_X1 U8095 ( .A1(n12040), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U8096 ( .A1(n7204), .A2(n7202), .ZN(n9936) );
  NAND2_X1 U8097 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n7203), .ZN(n7202) );
  NAND2_X1 U8098 ( .A1(n10035), .A2(n10034), .ZN(n10213) );
  XNOR2_X1 U8099 ( .A(n9578), .B(n7635), .ZN(n9913) );
  AND2_X1 U8100 ( .A1(n10041), .A2(n10040), .ZN(n12621) );
  MUX2_X1 U8101 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10039), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n10041) );
  NAND2_X1 U8102 ( .A1(n6691), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U8103 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n11133), .ZN(n9574) );
  NAND2_X1 U8104 ( .A1(n7214), .A2(n9569), .ZN(n9825) );
  NAND2_X1 U8105 ( .A1(n9810), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7214) );
  INV_X1 U8106 ( .A(n9679), .ZN(n7666) );
  AND3_X1 U8107 ( .A1(n6884), .A2(n6916), .A3(n6881), .ZN(n7667) );
  INV_X1 U8108 ( .A(n7668), .ZN(n6881) );
  NOR2_X1 U8109 ( .A1(n9556), .A2(n7223), .ZN(n7222) );
  AND2_X1 U8110 ( .A1(n10558), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9556) );
  INV_X1 U8111 ( .A(n9555), .ZN(n7223) );
  XNOR2_X1 U8112 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9726) );
  CLKBUF_X1 U8113 ( .A(n9697), .Z(n6979) );
  AND2_X1 U8114 ( .A1(n9683), .A2(n9682), .ZN(n11596) );
  NAND2_X1 U8115 ( .A1(n9633), .A2(n9587), .ZN(n9664) );
  INV_X1 U8116 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7334) );
  OR3_X1 U8117 ( .A1(n14255), .A2(n12210), .A3(n12330), .ZN(n10494) );
  AND2_X1 U8118 ( .A1(n8879), .A2(n8878), .ZN(n12199) );
  OR2_X1 U8119 ( .A1(n8876), .A2(n8877), .ZN(n8878) );
  AND2_X1 U8120 ( .A1(n12010), .A2(n8848), .ZN(n7480) );
  AND2_X1 U8121 ( .A1(n12199), .A2(n6737), .ZN(n7478) );
  INV_X1 U8122 ( .A(n13799), .ZN(n11021) );
  INV_X1 U8123 ( .A(n8934), .ZN(n7453) );
  NAND2_X1 U8124 ( .A1(n7473), .A2(n7472), .ZN(n13719) );
  AND2_X1 U8125 ( .A1(n8891), .A2(n8911), .ZN(n7472) );
  NAND2_X1 U8126 ( .A1(n13719), .A2(n8912), .ZN(n13730) );
  NAND2_X1 U8127 ( .A1(n13730), .A2(n13731), .ZN(n13729) );
  INV_X1 U8128 ( .A(n7451), .ZN(n7450) );
  OAI21_X1 U8129 ( .B1(n6718), .B2(n7452), .A(n13682), .ZN(n7451) );
  INV_X1 U8130 ( .A(n8955), .ZN(n7452) );
  AND2_X1 U8131 ( .A1(n7458), .A2(n7455), .ZN(n7454) );
  INV_X1 U8132 ( .A(n11622), .ZN(n7455) );
  AOI21_X1 U8134 ( .B1(n12836), .B2(n12835), .A(n6787), .ZN(n7134) );
  XNOR2_X1 U8135 ( .A(n12856), .B(n13879), .ZN(n12937) );
  NAND2_X1 U8136 ( .A1(n12882), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6853) );
  INV_X1 U8137 ( .A(n7343), .ZN(n7341) );
  NAND2_X1 U8138 ( .A1(n13992), .A2(n13974), .ZN(n13968) );
  NOR2_X1 U8139 ( .A1(n13897), .A2(n7439), .ZN(n7438) );
  INV_X1 U8140 ( .A(n13896), .ZN(n7436) );
  NOR2_X1 U8141 ( .A1(n6746), .A2(n7426), .ZN(n7425) );
  INV_X1 U8142 ( .A(n7428), .ZN(n7426) );
  INV_X1 U8143 ( .A(n7500), .ZN(n7499) );
  OAI21_X1 U8144 ( .B1(n14068), .B2(n7503), .A(n6699), .ZN(n7500) );
  NAND2_X1 U8145 ( .A1(n6843), .A2(n6740), .ZN(n14075) );
  NAND2_X1 U8146 ( .A1(n14094), .A2(n6743), .ZN(n6843) );
  OR2_X1 U8147 ( .A1(n14195), .A2(n14127), .ZN(n6984) );
  OR2_X1 U8148 ( .A1(n13909), .A2(n13887), .ZN(n7754) );
  NAND2_X1 U8149 ( .A1(n7517), .A2(n7516), .ZN(n7515) );
  INV_X1 U8150 ( .A(n7514), .ZN(n7512) );
  OR2_X1 U8151 ( .A1(n12736), .A2(n13790), .ZN(n7430) );
  AOI21_X1 U8152 ( .B1(n11654), .B2(n11653), .A(n6735), .ZN(n11887) );
  AND2_X1 U8153 ( .A1(n7442), .A2(n12910), .ZN(n7441) );
  OR2_X1 U8154 ( .A1(n7444), .A2(n7443), .ZN(n7442) );
  INV_X1 U8155 ( .A(n11466), .ZN(n7443) );
  NAND2_X1 U8156 ( .A1(n11465), .A2(n7444), .ZN(n11802) );
  NAND2_X1 U8157 ( .A1(n11777), .A2(n11442), .ZN(n11832) );
  NAND2_X1 U8158 ( .A1(n11832), .A2(n12904), .ZN(n11831) );
  NAND2_X1 U8159 ( .A1(n11790), .A2(n11440), .ZN(n11778) );
  INV_X1 U8160 ( .A(n13795), .ZN(n11779) );
  INV_X1 U8161 ( .A(n15388), .ZN(n14126) );
  NAND2_X1 U8162 ( .A1(n12016), .A2(n6675), .ZN(n7048) );
  NAND2_X1 U8163 ( .A1(n8919), .A2(n8918), .ZN(n14200) );
  INV_X1 U8164 ( .A(n15467), .ZN(n15450) );
  AND2_X1 U8165 ( .A1(n9081), .A2(n9080), .ZN(n10964) );
  AND2_X1 U8166 ( .A1(n9086), .A2(n9085), .ZN(n12119) );
  NAND2_X1 U8167 ( .A1(n14235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6845) );
  NOR2_X1 U8168 ( .A1(n9082), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U8169 ( .A1(n9070), .A2(n9067), .ZN(n9076) );
  INV_X1 U8170 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9067) );
  XNOR2_X1 U8171 ( .A(n9083), .B(P2_IR_REG_23__SCAN_IN), .ZN(n12176) );
  INV_X1 U8172 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8565) );
  AND2_X1 U8173 ( .A1(n10463), .A2(n10477), .ZN(n8552) );
  INV_X1 U8174 ( .A(n14396), .ZN(n14571) );
  NAND2_X1 U8175 ( .A1(n10462), .A2(n10456), .ZN(n7580) );
  NAND2_X1 U8176 ( .A1(n7592), .A2(n6947), .ZN(n14304) );
  AND2_X1 U8177 ( .A1(n7591), .A2(n14305), .ZN(n6947) );
  AND2_X1 U8178 ( .A1(n8195), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U8179 ( .A1(n8209), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8269) );
  AND2_X1 U8180 ( .A1(n15083), .A2(n10336), .ZN(n7585) );
  NAND2_X1 U8181 ( .A1(n10333), .A2(n10332), .ZN(n15103) );
  AOI21_X1 U8182 ( .B1(n7605), .B2(n7606), .A(n7603), .ZN(n7602) );
  INV_X1 U8183 ( .A(n14361), .ZN(n7603) );
  AND4_X1 U8184 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n14579)
         );
  AND2_X1 U8185 ( .A1(n7796), .A2(n7795), .ZN(n14576) );
  AND4_X1 U8186 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n14570)
         );
  AND4_X1 U8187 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n12412)
         );
  NAND2_X2 U8188 ( .A1(n7694), .A2(n7790), .ZN(n8430) );
  NAND2_X1 U8189 ( .A1(n7199), .A2(n7887), .ZN(n7198) );
  INV_X1 U8190 ( .A(n7200), .ZN(n7199) );
  NAND2_X1 U8191 ( .A1(n14603), .A2(n14594), .ZN(n14587) );
  OAI22_X1 U8192 ( .A1(n14628), .A2(n14630), .B1(n7265), .B2(n14580), .ZN(
        n14617) );
  NOR2_X1 U8193 ( .A1(n7380), .A2(n7751), .ZN(n7377) );
  AOI21_X1 U8194 ( .B1(n14686), .B2(n14685), .A(n7760), .ZN(n14673) );
  OR2_X1 U8195 ( .A1(n14571), .A2(n10382), .ZN(n7748) );
  NAND2_X1 U8196 ( .A1(n14769), .A2(n7722), .ZN(n7718) );
  NAND2_X1 U8197 ( .A1(n8244), .A2(n14565), .ZN(n7721) );
  NAND2_X1 U8198 ( .A1(n7718), .A2(n7716), .ZN(n14752) );
  INV_X1 U8199 ( .A(n7720), .ZN(n7716) );
  AOI21_X1 U8200 ( .B1(n7374), .B2(n7371), .A(n7370), .ZN(n7369) );
  NOR2_X1 U8201 ( .A1(n8244), .A2(n14566), .ZN(n7370) );
  NOR2_X1 U8202 ( .A1(n7375), .A2(n14567), .ZN(n7371) );
  NAND2_X1 U8203 ( .A1(n7374), .A2(n7373), .ZN(n7372) );
  INV_X1 U8204 ( .A(n14567), .ZN(n7373) );
  INV_X1 U8205 ( .A(n14781), .ZN(n7375) );
  NAND2_X1 U8206 ( .A1(n7735), .A2(n7734), .ZN(n7733) );
  NOR2_X1 U8207 ( .A1(n14540), .A2(n7737), .ZN(n7736) );
  NAND2_X1 U8208 ( .A1(n12409), .A2(n7741), .ZN(n7740) );
  AND2_X1 U8209 ( .A1(n14539), .A2(n8493), .ZN(n14787) );
  NAND2_X1 U8210 ( .A1(n6793), .A2(n7361), .ZN(n7357) );
  OR2_X1 U8211 ( .A1(n12033), .A2(n7360), .ZN(n7359) );
  NAND2_X1 U8212 ( .A1(n12349), .A2(n7361), .ZN(n7358) );
  NAND2_X1 U8213 ( .A1(n12021), .A2(n7703), .ZN(n12342) );
  NAND2_X1 U8214 ( .A1(n12034), .A2(n12033), .ZN(n12350) );
  INV_X1 U8215 ( .A(n7198), .ZN(n7197) );
  NAND2_X1 U8216 ( .A1(n6792), .A2(n6696), .ZN(n7696) );
  OR2_X1 U8217 ( .A1(n14403), .A2(n15263), .ZN(n11512) );
  NAND2_X1 U8218 ( .A1(n15209), .A2(n6681), .ZN(n11140) );
  AND2_X1 U8219 ( .A1(n7986), .A2(n7985), .ZN(n11276) );
  OAI21_X1 U8220 ( .B1(n11199), .B2(n6752), .A(n11200), .ZN(n7388) );
  OR2_X1 U8221 ( .A1(n11322), .A2(n11138), .ZN(n14590) );
  NAND2_X1 U8222 ( .A1(n8402), .A2(n8401), .ZN(n14837) );
  OAI21_X1 U8223 ( .B1(n14684), .B2(n7710), .A(n7708), .ZN(n14650) );
  INV_X1 U8224 ( .A(n10382), .ZN(n14883) );
  NAND2_X1 U8225 ( .A1(n8266), .A2(n8265), .ZN(n14888) );
  OAI21_X1 U8226 ( .B1(n8452), .B2(n7250), .A(n7246), .ZN(n7245) );
  INV_X1 U8227 ( .A(n7249), .ZN(n7246) );
  OAI22_X1 U8228 ( .A1(n7252), .A2(n7250), .B1(n8479), .B2(n7251), .ZN(n7249)
         );
  NAND2_X1 U8229 ( .A1(n7251), .A2(n8479), .ZN(n7250) );
  AND2_X1 U8230 ( .A1(n7253), .A2(n8451), .ZN(n7252) );
  INV_X1 U8231 ( .A(n8454), .ZN(n7253) );
  NAND2_X1 U8232 ( .A1(n8448), .A2(n8447), .ZN(n8452) );
  INV_X1 U8233 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U8234 ( .A1(n8399), .A2(n8398), .ZN(n8415) );
  OAI21_X1 U8235 ( .B1(n8397), .B2(n13670), .A(n8396), .ZN(n8399) );
  NAND2_X1 U8236 ( .A1(n8397), .A2(n13670), .ZN(n8398) );
  XNOR2_X1 U8237 ( .A(n8397), .B(n8383), .ZN(n14251) );
  XNOR2_X1 U8238 ( .A(n8129), .B(n8128), .ZN(n10745) );
  OAI21_X1 U8239 ( .B1(n7834), .B2(n8085), .A(n7541), .ZN(n8103) );
  XNOR2_X1 U8240 ( .A(n9166), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U8241 ( .A1(n15697), .A2(n9182), .ZN(n9186) );
  OR2_X1 U8242 ( .A1(n15701), .A2(n9191), .ZN(n6925) );
  NAND2_X1 U8243 ( .A1(n15148), .A2(n6924), .ZN(n9201) );
  OAI21_X1 U8244 ( .B1(n15150), .B2(n15149), .A(n6927), .ZN(n6924) );
  NAND2_X1 U8245 ( .A1(n13094), .A2(n13092), .ZN(n6914) );
  INV_X1 U8246 ( .A(n13423), .ZN(n13403) );
  NAND2_X1 U8247 ( .A1(n12044), .A2(n12043), .ZN(n12110) );
  NAND2_X1 U8248 ( .A1(n13110), .A2(n12570), .ZN(n13049) );
  OAI21_X1 U8249 ( .B1(n13020), .B2(n6893), .A(n6891), .ZN(n12989) );
  NAND2_X1 U8250 ( .A1(n7392), .A2(n12111), .ZN(n12098) );
  XNOR2_X1 U8251 ( .A(n12052), .B(n15574), .ZN(n12089) );
  NOR2_X1 U8252 ( .A1(n6697), .A2(n13142), .ZN(n7400) );
  NOR2_X1 U8253 ( .A1(n12980), .A2(n13390), .ZN(n7402) );
  AOI21_X1 U8254 ( .B1(n12980), .B2(n13412), .A(n12596), .ZN(n7403) );
  NAND2_X1 U8255 ( .A1(n12047), .A2(n15573), .ZN(n12048) );
  CLKBUF_X1 U8256 ( .A(n13151), .Z(n13135) );
  INV_X1 U8257 ( .A(n12243), .ZN(n12305) );
  INV_X1 U8258 ( .A(n12051), .ZN(n15574) );
  NAND2_X1 U8259 ( .A1(n7104), .A2(n7101), .ZN(n7100) );
  INV_X1 U8260 ( .A(n11690), .ZN(n7101) );
  NAND2_X1 U8261 ( .A1(n11550), .A2(n6692), .ZN(n7099) );
  NAND2_X1 U8262 ( .A1(n6954), .A2(n6953), .ZN(n15517) );
  INV_X1 U8263 ( .A(n15513), .ZN(n6953) );
  OR2_X1 U8264 ( .A1(n11851), .A2(n9752), .ZN(n6870) );
  XNOR2_X1 U8265 ( .A(n11996), .B(n11997), .ZN(n11851) );
  INV_X1 U8266 ( .A(n11985), .ZN(n7045) );
  NOR2_X1 U8267 ( .A1(n12258), .A2(n12259), .ZN(n13191) );
  NOR2_X1 U8268 ( .A1(n13202), .A2(n13211), .ZN(n13245) );
  NOR2_X1 U8269 ( .A1(n13304), .A2(n13303), .ZN(n13313) );
  NAND2_X1 U8270 ( .A1(n13313), .A2(n6863), .ZN(n6862) );
  AND2_X1 U8271 ( .A1(n6865), .A2(n13321), .ZN(n6863) );
  INV_X1 U8272 ( .A(n7042), .ZN(n13283) );
  AOI21_X1 U8273 ( .B1(n12547), .B2(n15599), .A(n12546), .ZN(n13541) );
  NAND2_X1 U8274 ( .A1(n10020), .A2(n10019), .ZN(n13606) );
  NAND2_X1 U8275 ( .A1(n12640), .A2(n9805), .ZN(n10020) );
  AND2_X1 U8276 ( .A1(n13606), .A2(n13639), .ZN(n6958) );
  AND2_X1 U8277 ( .A1(n11331), .A2(n11330), .ZN(n13659) );
  OR2_X1 U8278 ( .A1(n11344), .A2(P3_D_REG_1__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U8279 ( .A1(n8957), .A2(n8956), .ZN(n14191) );
  AND2_X1 U8280 ( .A1(n7466), .A2(n7464), .ZN(n7463) );
  INV_X1 U8281 ( .A(n7469), .ZN(n7464) );
  AND2_X1 U8282 ( .A1(n7467), .A2(n9100), .ZN(n7466) );
  AOI21_X1 U8283 ( .B1(n9102), .B2(n7469), .A(n7468), .ZN(n7467) );
  AND2_X1 U8284 ( .A1(n7470), .A2(n13691), .ZN(n7468) );
  OR2_X1 U8285 ( .A1(n9102), .A2(n13696), .ZN(n7471) );
  NAND2_X1 U8286 ( .A1(n6672), .A2(n7485), .ZN(n13715) );
  INV_X1 U8287 ( .A(n13717), .ZN(n7030) );
  NOR2_X1 U8288 ( .A1(n13716), .A2(n7484), .ZN(n7483) );
  INV_X1 U8289 ( .A(n7485), .ZN(n7484) );
  INV_X1 U8290 ( .A(n13892), .ZN(n14092) );
  NAND2_X1 U8291 ( .A1(n9104), .A2(n15384), .ZN(n13783) );
  OAI21_X1 U8292 ( .B1(n7413), .B2(n7418), .A(n7412), .ZN(n7411) );
  NAND2_X1 U8293 ( .A1(n6784), .A2(n7413), .ZN(n7412) );
  NAND2_X1 U8294 ( .A1(n7410), .A2(n6750), .ZN(n7409) );
  INV_X1 U8295 ( .A(n13951), .ZN(n7410) );
  NAND2_X1 U8296 ( .A1(n13951), .A2(n7405), .ZN(n7404) );
  NOR2_X1 U8297 ( .A1(n13928), .A2(n7406), .ZN(n7405) );
  INV_X1 U8298 ( .A(n7415), .ZN(n7406) );
  AOI21_X1 U8299 ( .B1(n14139), .B2(n14108), .A(n13931), .ZN(n7076) );
  AOI21_X1 U8300 ( .B1(n6847), .B2(n14129), .A(n6826), .ZN(n14142) );
  XNOR2_X1 U8301 ( .A(n7506), .B(n7418), .ZN(n6847) );
  NAND2_X1 U8302 ( .A1(n13929), .A2(n13930), .ZN(n7504) );
  XNOR2_X1 U8303 ( .A(n13932), .B(n13940), .ZN(n14147) );
  AOI21_X1 U8304 ( .B1(n13951), .B2(n7024), .A(n7416), .ZN(n13932) );
  AOI21_X1 U8305 ( .B1(n13961), .B2(n14129), .A(n6985), .ZN(n14151) );
  NAND2_X1 U8306 ( .A1(n6987), .A2(n6986), .ZN(n6985) );
  NAND2_X1 U8307 ( .A1(n13960), .A2(n14124), .ZN(n6986) );
  NAND2_X1 U8308 ( .A1(n9035), .A2(n9034), .ZN(n14159) );
  NAND2_X1 U8309 ( .A1(n8628), .A2(n8627), .ZN(n14165) );
  NAND2_X1 U8310 ( .A1(n15401), .A2(n10963), .ZN(n15384) );
  NOR2_X1 U8311 ( .A1(n7577), .A2(n15101), .ZN(n7576) );
  NOR2_X1 U8312 ( .A1(n7578), .A2(n7581), .ZN(n7577) );
  NOR2_X1 U8313 ( .A1(n10462), .A2(n10456), .ZN(n7581) );
  INV_X1 U8314 ( .A(n7580), .ZN(n7578) );
  NAND2_X1 U8315 ( .A1(n7580), .A2(n7582), .ZN(n7579) );
  INV_X1 U8316 ( .A(n10462), .ZN(n7582) );
  OAI21_X1 U8317 ( .B1(n14610), .B2(n14388), .A(n10491), .ZN(n10492) );
  NAND2_X1 U8318 ( .A1(n8053), .A2(n8052), .ZN(n11705) );
  NAND2_X1 U8319 ( .A1(n8208), .A2(n8207), .ZN(n14905) );
  AND4_X1 U8320 ( .A1(n8119), .A2(n8118), .A3(n8117), .A4(n8116), .ZN(n14560)
         );
  NOR2_X1 U8321 ( .A1(n8166), .A2(n7200), .ZN(n8220) );
  AOI21_X1 U8322 ( .B1(n7384), .B2(n7383), .A(n7382), .ZN(n7381) );
  INV_X1 U8323 ( .A(n14584), .ZN(n7382) );
  AOI21_X1 U8324 ( .B1(n14558), .B2(n15253), .A(n7761), .ZN(n14826) );
  NAND2_X1 U8325 ( .A1(n8147), .A2(n8146), .ZN(n15087) );
  NAND2_X1 U8326 ( .A1(n8071), .A2(n8070), .ZN(n12030) );
  OR2_X1 U8327 ( .A1(n11140), .A2(n11139), .ZN(n15117) );
  NOR2_X1 U8328 ( .A1(n9171), .A2(n15708), .ZN(n14965) );
  INV_X1 U8329 ( .A(n7007), .ZN(n9173) );
  XNOR2_X1 U8330 ( .A(n6925), .B(n6728), .ZN(n14972) );
  AND2_X1 U8331 ( .A1(n6925), .A2(n6728), .ZN(n9194) );
  INV_X1 U8332 ( .A(n15146), .ZN(n6974) );
  INV_X1 U8333 ( .A(n15163), .ZN(n7008) );
  INV_X1 U8334 ( .A(n15162), .ZN(n7009) );
  NAND2_X1 U8335 ( .A1(n9205), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8336 ( .A1(n6929), .A2(n6928), .ZN(n7044) );
  NAND2_X1 U8337 ( .A1(n15004), .A2(n6930), .ZN(n6928) );
  AND2_X1 U8338 ( .A1(n12656), .A2(n12655), .ZN(n12659) );
  AND2_X1 U8339 ( .A1(n12662), .A2(n12661), .ZN(n12668) );
  OR2_X1 U8340 ( .A1(n12701), .A2(n12700), .ZN(n12709) );
  INV_X1 U8341 ( .A(n6698), .ZN(n7131) );
  NAND2_X1 U8342 ( .A1(n6698), .A2(n12727), .ZN(n7128) );
  OR2_X1 U8343 ( .A1(n8055), .A2(n7168), .ZN(n7163) );
  NAND2_X1 U8344 ( .A1(n8095), .A2(n7178), .ZN(n7177) );
  NAND2_X1 U8345 ( .A1(n7166), .A2(n7164), .ZN(n8073) );
  AOI21_X1 U8346 ( .B1(n7168), .B2(n7167), .A(n7165), .ZN(n7164) );
  INV_X1 U8347 ( .A(n8075), .ZN(n7165) );
  NAND2_X1 U8348 ( .A1(n7121), .A2(n7120), .ZN(n12741) );
  AOI21_X1 U8349 ( .B1(n6690), .B2(n7130), .A(n6727), .ZN(n7120) );
  INV_X1 U8350 ( .A(n7675), .ZN(n7119) );
  NAND2_X1 U8351 ( .A1(n7161), .A2(n8248), .ZN(n7160) );
  NAND2_X1 U8352 ( .A1(n7141), .A2(n7139), .ZN(n12765) );
  AND2_X1 U8353 ( .A1(n12766), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U8354 ( .A1(n7143), .A2(n7142), .ZN(n7140) );
  OAI22_X1 U8355 ( .A1(n7116), .A2(n6754), .B1(n6683), .B2(n7114), .ZN(n7113)
         );
  INV_X1 U8356 ( .A(n6700), .ZN(n7676) );
  INV_X1 U8357 ( .A(n8308), .ZN(n7181) );
  NAND2_X1 U8358 ( .A1(n7568), .A2(n7571), .ZN(n7567) );
  INV_X1 U8359 ( .A(n8319), .ZN(n7571) );
  AND2_X1 U8360 ( .A1(n7146), .A2(n7145), .ZN(n12797) );
  NAND2_X1 U8361 ( .A1(n6790), .A2(n7147), .ZN(n7145) );
  NAND2_X1 U8362 ( .A1(n6723), .A2(n7149), .ZN(n7147) );
  NAND2_X1 U8363 ( .A1(n10194), .A2(n10193), .ZN(n6981) );
  NAND2_X1 U8364 ( .A1(n10207), .A2(n10206), .ZN(n6983) );
  NOR2_X1 U8365 ( .A1(n7175), .A2(n8387), .ZN(n7172) );
  NAND2_X1 U8366 ( .A1(n7174), .A2(n7552), .ZN(n7173) );
  INV_X1 U8367 ( .A(n8387), .ZN(n7174) );
  INV_X1 U8368 ( .A(n8446), .ZN(n7535) );
  NAND2_X1 U8369 ( .A1(n6827), .A2(n7854), .ZN(n7546) );
  NOR2_X1 U8370 ( .A1(n12521), .A2(n7299), .ZN(n7298) );
  INV_X1 U8371 ( .A(n12518), .ZN(n7299) );
  NOR2_X1 U8372 ( .A1(n12828), .A2(n6775), .ZN(n7679) );
  NOR2_X1 U8373 ( .A1(n7683), .A2(n7684), .ZN(n7682) );
  AOI22_X1 U8374 ( .A1(n7684), .A2(n7686), .B1(n7683), .B2(n7690), .ZN(n7681)
         );
  OR4_X1 U8375 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n12912) );
  AND2_X1 U8376 ( .A1(n7192), .A2(n8477), .ZN(n7191) );
  NAND2_X1 U8377 ( .A1(n7534), .A2(n7536), .ZN(n7192) );
  INV_X1 U8378 ( .A(n12341), .ZN(n7701) );
  INV_X1 U8379 ( .A(n8261), .ZN(n7055) );
  NOR2_X1 U8380 ( .A1(n8261), .A2(n8249), .ZN(n7052) );
  OAI21_X1 U8381 ( .B1(n7064), .B2(n7062), .A(n7849), .ZN(n7061) );
  INV_X1 U8382 ( .A(n7852), .ZN(n7057) );
  INV_X1 U8383 ( .A(n8102), .ZN(n7540) );
  NAND2_X1 U8384 ( .A1(n7935), .A2(n7815), .ZN(n7002) );
  OAI21_X1 U8385 ( .B1(n10502), .B2(n10540), .A(n6962), .ZN(n7817) );
  NAND2_X1 U8386 ( .A1(n10502), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6962) );
  OAI21_X1 U8387 ( .B1(n10502), .B2(n7026), .A(n7025), .ZN(n7814) );
  NAND2_X1 U8388 ( .A1(n10497), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7025) );
  INV_X1 U8389 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7799) );
  NAND2_X1 U8390 ( .A1(n6878), .A2(n13661), .ZN(n6877) );
  NAND2_X1 U8391 ( .A1(n6876), .A2(n11483), .ZN(n6875) );
  INV_X1 U8392 ( .A(n11361), .ZN(n6878) );
  NAND2_X1 U8393 ( .A1(n15031), .A2(n10208), .ZN(n7662) );
  NOR2_X1 U8394 ( .A1(n13376), .A2(n7303), .ZN(n7302) );
  INV_X1 U8395 ( .A(n12534), .ZN(n7303) );
  NAND2_X1 U8396 ( .A1(n12533), .A2(n7305), .ZN(n7304) );
  OR2_X1 U8397 ( .A1(n9949), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9959) );
  AND2_X1 U8398 ( .A1(n10176), .A2(n10175), .ZN(n12530) );
  INV_X1 U8399 ( .A(n7659), .ZN(n7653) );
  NAND2_X1 U8400 ( .A1(n7297), .A2(n12520), .ZN(n13499) );
  NAND2_X1 U8401 ( .A1(n12519), .A2(n7298), .ZN(n7297) );
  OAI21_X1 U8402 ( .B1(n11957), .B2(n7647), .A(n12165), .ZN(n7641) );
  INV_X1 U8403 ( .A(n9730), .ZN(n7647) );
  OR2_X1 U8404 ( .A1(n15560), .A2(n15561), .ZN(n15558) );
  NAND2_X1 U8405 ( .A1(n15573), .A2(n12115), .ZN(n10091) );
  OR2_X1 U8406 ( .A1(n11344), .A2(n11343), .ZN(n11480) );
  XNOR2_X1 U8407 ( .A(n7106), .B(P3_IR_REG_27__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U8408 ( .A1(n9602), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7106) );
  INV_X1 U8409 ( .A(n9582), .ZN(n7625) );
  NAND2_X1 U8410 ( .A1(n9595), .A2(n9594), .ZN(n7671) );
  NOR2_X1 U8411 ( .A1(n7232), .A2(n7231), .ZN(n7230) );
  INV_X1 U8412 ( .A(n7629), .ZN(n7231) );
  NAND2_X1 U8413 ( .A1(n9945), .A2(n7628), .ZN(n7229) );
  INV_X1 U8414 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7398) );
  INV_X1 U8415 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9571) );
  INV_X1 U8416 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9875) );
  INV_X1 U8417 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U8418 ( .A1(n6917), .A2(n6918), .ZN(n7668) );
  NOR2_X1 U8419 ( .A1(n8922), .A2(n8921), .ZN(n8920) );
  NOR2_X1 U8420 ( .A1(n8781), .A2(n8780), .ZN(n8779) );
  AND2_X1 U8421 ( .A1(n8779), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8800) );
  INV_X1 U8422 ( .A(n12943), .ZN(n12949) );
  OR2_X1 U8423 ( .A1(n14145), .A2(n13903), .ZN(n13927) );
  NOR2_X1 U8424 ( .A1(n14145), .A2(n7343), .ZN(n7342) );
  NAND2_X1 U8425 ( .A1(n7344), .A2(n13974), .ZN(n7343) );
  INV_X1 U8426 ( .A(n7438), .ZN(n7434) );
  NOR2_X1 U8427 ( .A1(n14049), .A2(n14175), .ZN(n7349) );
  AND2_X1 U8428 ( .A1(n14200), .A2(n13889), .ZN(n13890) );
  OAI21_X1 U8429 ( .B1(n7511), .B2(n6782), .A(n7508), .ZN(n6855) );
  AOI21_X1 U8430 ( .B1(n7513), .B2(n7510), .A(n7509), .ZN(n7508) );
  INV_X1 U8431 ( .A(n12287), .ZN(n7509) );
  INV_X1 U8432 ( .A(n12913), .ZN(n7520) );
  NOR2_X1 U8433 ( .A1(n11838), .A2(n15434), .ZN(n7348) );
  NOR2_X1 U8434 ( .A1(n8724), .A2(n8723), .ZN(n8722) );
  AND2_X1 U8435 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8685) );
  NAND2_X1 U8436 ( .A1(n13799), .A2(n6951), .ZN(n10966) );
  NAND2_X1 U8437 ( .A1(n7351), .A2(n12497), .ZN(n12500) );
  INV_X1 U8438 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8604) );
  NOR2_X1 U8439 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6859) );
  NOR2_X1 U8440 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6858) );
  NAND2_X1 U8441 ( .A1(n8584), .A2(n8615), .ZN(n8576) );
  INV_X1 U8442 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8568) );
  INV_X1 U8443 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8559) );
  INV_X1 U8444 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8560) );
  OR2_X1 U8445 ( .A1(n8716), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8735) );
  INV_X1 U8446 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8562) );
  NOR2_X2 U8447 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8647) );
  AND2_X1 U8448 ( .A1(n10481), .A2(n6679), .ZN(n10368) );
  INV_X1 U8449 ( .A(n7741), .ZN(n7737) );
  INV_X1 U8450 ( .A(n7738), .ZN(n7735) );
  INV_X1 U8451 ( .A(n14540), .ZN(n7734) );
  OR2_X1 U8452 ( .A1(n14911), .A2(n14562), .ZN(n14539) );
  OR2_X1 U8453 ( .A1(n12030), .A2(n11705), .ZN(n7259) );
  INV_X1 U8454 ( .A(n11519), .ZN(n7697) );
  NOR2_X1 U8455 ( .A1(n11208), .A2(n7731), .ZN(n7730) );
  INV_X1 U8456 ( .A(n11206), .ZN(n7731) );
  NAND2_X1 U8457 ( .A1(n14687), .A2(n6688), .ZN(n14665) );
  NAND2_X1 U8458 ( .A1(n14687), .A2(n14679), .ZN(n14678) );
  OR2_X1 U8459 ( .A1(n14877), .A2(n14720), .ZN(n14707) );
  OR2_X1 U8460 ( .A1(n14883), .A2(n14571), .ZN(n14545) );
  AND2_X1 U8461 ( .A1(n10479), .A2(n11885), .ZN(n10702) );
  INV_X1 U8462 ( .A(n8482), .ZN(n7251) );
  INV_X1 U8463 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7782) );
  INV_X1 U8464 ( .A(n8360), .ZN(n8362) );
  AND2_X1 U8465 ( .A1(n7776), .A2(n7590), .ZN(n7589) );
  NOR2_X1 U8466 ( .A1(n7779), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n7590) );
  INV_X1 U8467 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U8468 ( .A1(n7059), .A2(n7063), .ZN(n8109) );
  AOI21_X1 U8469 ( .B1(n7835), .B2(n7542), .A(n6768), .ZN(n7541) );
  INV_X1 U8470 ( .A(n7833), .ZN(n7542) );
  AND2_X1 U8471 ( .A1(n7769), .A2(n7959), .ZN(n8087) );
  AOI21_X1 U8472 ( .B1(n7530), .B2(n7531), .A(n6777), .ZN(n7527) );
  INV_X1 U8473 ( .A(n7825), .ZN(n7531) );
  OR2_X1 U8474 ( .A1(n7983), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7994) );
  INV_X1 U8475 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7768) );
  OAI21_X1 U8476 ( .B1(n7808), .B2(n10496), .A(n7804), .ZN(n7806) );
  AOI21_X1 U8477 ( .B1(n7007), .B2(n7006), .A(n7281), .ZN(n9131) );
  AND2_X1 U8478 ( .A1(n14426), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7281) );
  INV_X1 U8479 ( .A(n9172), .ZN(n7006) );
  NOR2_X1 U8480 ( .A1(n9141), .A2(n9140), .ZN(n9193) );
  OAI21_X1 U8481 ( .B1(n9317), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9144), .ZN(
        n9146) );
  OR2_X1 U8482 ( .A1(n9196), .A2(n9195), .ZN(n9144) );
  AND2_X1 U8483 ( .A1(n6901), .A2(n6904), .ZN(n6900) );
  INV_X1 U8484 ( .A(n13133), .ZN(n6904) );
  NAND2_X1 U8485 ( .A1(n6902), .A2(n6710), .ZN(n6901) );
  INV_X1 U8486 ( .A(n13061), .ZN(n6902) );
  INV_X1 U8487 ( .A(n6710), .ZN(n6903) );
  AND2_X1 U8488 ( .A1(n12978), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U8489 ( .A1(n6894), .A2(n7393), .ZN(n6892) );
  INV_X1 U8490 ( .A(n7393), .ZN(n6893) );
  AND2_X1 U8491 ( .A1(n9864), .A2(n9863), .ZN(n9881) );
  INV_X1 U8492 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U8493 ( .A1(n9750), .A2(n9749), .ZN(n9764) );
  NOR2_X1 U8494 ( .A1(n9792), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9817) );
  OR2_X1 U8495 ( .A1(n9829), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U8496 ( .A1(n9844), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9864) );
  AND2_X1 U8497 ( .A1(n9978), .A2(n9977), .ZN(n12992) );
  AND4_X1 U8498 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n13128)
         );
  AND4_X1 U8499 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9692), .ZN(n12051)
         );
  NAND2_X1 U8500 ( .A1(n9816), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9639) );
  OR2_X1 U8501 ( .A1(n11564), .A2(n11577), .ZN(n11565) );
  NAND2_X1 U8502 ( .A1(n11579), .A2(n11681), .ZN(n11580) );
  NAND2_X1 U8503 ( .A1(n7549), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11682) );
  INV_X1 U8504 ( .A(n11580), .ZN(n7549) );
  NOR2_X1 U8505 ( .A1(n11765), .A2(n7526), .ZN(n11764) );
  INV_X1 U8506 ( .A(n7087), .ZN(n7086) );
  AOI21_X1 U8507 ( .B1(n7089), .B2(n7088), .A(n12260), .ZN(n7087) );
  NOR2_X1 U8508 ( .A1(n13184), .A2(n13185), .ZN(n13213) );
  OR2_X1 U8509 ( .A1(n13213), .A2(n7105), .ZN(n13235) );
  OR2_X1 U8510 ( .A1(n13214), .A2(n13212), .ZN(n7105) );
  NAND2_X1 U8511 ( .A1(n7077), .A2(n13271), .ZN(n13272) );
  NAND2_X1 U8512 ( .A1(n7078), .A2(n13270), .ZN(n7077) );
  OR2_X1 U8513 ( .A1(n13273), .A2(n13272), .ZN(n13291) );
  NAND2_X1 U8514 ( .A1(n6866), .A2(n13312), .ZN(n6865) );
  XNOR2_X1 U8515 ( .A(n13324), .B(n7084), .ZN(n7083) );
  INV_X1 U8516 ( .A(n13323), .ZN(n7084) );
  NAND2_X1 U8517 ( .A1(n7322), .A2(n7081), .ZN(n7080) );
  NAND2_X1 U8518 ( .A1(n15539), .A2(n7323), .ZN(n7322) );
  NOR2_X1 U8519 ( .A1(n6831), .A2(n7082), .ZN(n7081) );
  INV_X1 U8520 ( .A(n10065), .ZN(n7664) );
  INV_X1 U8521 ( .A(n7310), .ZN(n7308) );
  AOI21_X1 U8522 ( .B1(n7311), .B2(n13346), .A(n7313), .ZN(n7310) );
  AND2_X1 U8523 ( .A1(n12515), .A2(n13345), .ZN(n7313) );
  NAND2_X1 U8524 ( .A1(n10065), .A2(n10064), .ZN(n13328) );
  AND2_X1 U8525 ( .A1(n10068), .A2(n10067), .ZN(n13362) );
  NAND2_X1 U8526 ( .A1(n7304), .A2(n7302), .ZN(n13369) );
  NAND2_X1 U8527 ( .A1(n12533), .A2(n12532), .ZN(n13388) );
  NAND2_X1 U8528 ( .A1(n9955), .A2(n10185), .ZN(n13386) );
  INV_X1 U8529 ( .A(n12530), .ZN(n13429) );
  NOR2_X1 U8530 ( .A1(n7288), .A2(n7287), .ZN(n13422) );
  INV_X1 U8531 ( .A(n12529), .ZN(n7287) );
  INV_X1 U8532 ( .A(n13435), .ZN(n7288) );
  NAND2_X1 U8533 ( .A1(n13435), .A2(n7289), .ZN(n13421) );
  NAND2_X1 U8534 ( .A1(n13436), .A2(n13437), .ZN(n13435) );
  AND2_X1 U8535 ( .A1(n9917), .A2(n9916), .ZN(n9930) );
  NAND2_X1 U8536 ( .A1(n12526), .A2(n6765), .ZN(n7291) );
  AND2_X1 U8537 ( .A1(n10166), .A2(n10167), .ZN(n13460) );
  NOR2_X1 U8538 ( .A1(n9906), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U8539 ( .A1(n9881), .A2(n9880), .ZN(n9893) );
  OR2_X1 U8540 ( .A1(n9893), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9906) );
  OR2_X1 U8541 ( .A1(n13499), .A2(n13467), .ZN(n13484) );
  AND2_X1 U8542 ( .A1(n10145), .A2(n13492), .ZN(n13508) );
  NAND2_X1 U8543 ( .A1(n13509), .A2(n13508), .ZN(n13507) );
  INV_X1 U8544 ( .A(n12473), .ZN(n12450) );
  AND3_X1 U8545 ( .A1(n9776), .A2(n9775), .A3(n9774), .ZN(n12442) );
  AND2_X1 U8546 ( .A1(n10044), .A2(n12301), .ZN(n12218) );
  NOR2_X1 U8547 ( .A1(n12165), .A2(n7315), .ZN(n7314) );
  INV_X1 U8548 ( .A(n12162), .ZN(n7315) );
  NAND2_X1 U8549 ( .A1(n12163), .A2(n12162), .ZN(n12166) );
  INV_X1 U8550 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9731) );
  NOR2_X1 U8551 ( .A1(n9717), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9732) );
  OR2_X1 U8552 ( .A1(n9704), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9717) );
  INV_X1 U8553 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9688) );
  AND2_X1 U8554 ( .A1(n10100), .A2(n10096), .ZN(n15561) );
  AND3_X1 U8555 ( .A1(n9703), .A2(n9702), .A3(n9701), .ZN(n15567) );
  AND3_X1 U8556 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(n15581) );
  AND3_X1 U8557 ( .A1(n9669), .A2(n9668), .A3(n9667), .ZN(n12045) );
  CLKBUF_X1 U8558 ( .A(n11495), .Z(n15593) );
  AND2_X1 U8559 ( .A1(n11491), .A2(n11490), .ZN(n15602) );
  INV_X1 U8560 ( .A(n11364), .ZN(n15608) );
  INV_X1 U8561 ( .A(n15675), .ZN(n15051) );
  AND2_X1 U8562 ( .A1(n15602), .A2(n15654), .ZN(n15675) );
  OR2_X1 U8563 ( .A1(n6709), .A2(n9586), .ZN(n7236) );
  NAND2_X1 U8564 ( .A1(n7240), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U8565 ( .A1(n7239), .A2(n7241), .ZN(n7237) );
  NOR2_X1 U8566 ( .A1(n7671), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7670) );
  CLKBUF_X1 U8567 ( .A(n11533), .Z(n6997) );
  NAND2_X1 U8568 ( .A1(n10225), .A2(n9596), .ZN(n6998) );
  NAND2_X1 U8569 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n7016), .ZN(n7015) );
  NAND2_X1 U8570 ( .A1(n9876), .A2(n9875), .ZN(n9901) );
  AOI21_X1 U8571 ( .B1(n7210), .B2(n7620), .A(n7209), .ZN(n7211) );
  INV_X1 U8572 ( .A(n7618), .ZN(n7209) );
  XNOR2_X1 U8573 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9787) );
  INV_X1 U8574 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9562) );
  XNOR2_X1 U8575 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9770) );
  XNOR2_X1 U8576 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9758) );
  NAND2_X1 U8577 ( .A1(n9559), .A2(n9558), .ZN(n9745) );
  INV_X1 U8578 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9557) );
  XNOR2_X1 U8579 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9743) );
  INV_X1 U8580 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9723) );
  INV_X1 U8581 ( .A(n13696), .ZN(n7470) );
  NOR2_X1 U8582 ( .A1(n7470), .A2(n13691), .ZN(n7469) );
  OR2_X1 U8583 ( .A1(n8762), .A2(n8761), .ZN(n8781) );
  NAND2_X1 U8584 ( .A1(n8940), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8974) );
  AND2_X1 U8585 ( .A1(n13871), .A2(n12897), .ZN(n12863) );
  NOR2_X1 U8586 ( .A1(n8988), .A2(n13708), .ZN(n9008) );
  NAND2_X1 U8587 ( .A1(n8800), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8854) );
  AOI21_X1 U8588 ( .B1(n7460), .B2(n7459), .A(n6780), .ZN(n7458) );
  NOR2_X1 U8589 ( .A1(n11166), .A2(n7461), .ZN(n7459) );
  INV_X1 U8590 ( .A(n11268), .ZN(n7460) );
  NAND2_X1 U8591 ( .A1(n8638), .A2(n8637), .ZN(n8645) );
  INV_X1 U8592 ( .A(n8879), .ZN(n7475) );
  AND2_X1 U8593 ( .A1(n12961), .A2(n12925), .ZN(n10748) );
  NOR2_X1 U8594 ( .A1(n7021), .A2(n6960), .ZN(n12927) );
  NAND2_X1 U8595 ( .A1(n12937), .A2(n6730), .ZN(n6960) );
  AND2_X1 U8596 ( .A1(n12945), .A2(n12949), .ZN(n7673) );
  INV_X1 U8597 ( .A(n12952), .ZN(n6959) );
  INV_X1 U8598 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12201) );
  NOR2_X1 U8599 ( .A1(n13940), .A2(n13957), .ZN(n7415) );
  NAND2_X1 U8600 ( .A1(n13959), .A2(n14124), .ZN(n7505) );
  NAND2_X1 U8601 ( .A1(n13956), .A2(n6736), .ZN(n13939) );
  OAI21_X1 U8602 ( .B1(n13965), .B2(n13925), .A(n13924), .ZN(n13958) );
  NAND2_X1 U8603 ( .A1(n13959), .A2(n14126), .ZN(n6987) );
  AND2_X1 U8604 ( .A1(n7068), .A2(n6800), .ZN(n7065) );
  NAND2_X1 U8605 ( .A1(n9008), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U8606 ( .A1(n7349), .A2(n14020), .ZN(n14016) );
  INV_X1 U8607 ( .A(n7349), .ZN(n14039) );
  OAI21_X1 U8608 ( .B1(n14054), .B2(n6689), .A(n7421), .ZN(n7420) );
  INV_X1 U8609 ( .A(n7427), .ZN(n7421) );
  NAND2_X1 U8610 ( .A1(n7350), .A2(n14053), .ZN(n14049) );
  AOI22_X1 U8611 ( .A1(n12498), .A2(n12920), .B1(n12497), .B2(n12496), .ZN(
        n12499) );
  NAND2_X1 U8612 ( .A1(n8870), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8902) );
  OAI22_X1 U8613 ( .A1(n12312), .A2(n12917), .B1(n12334), .B2(n13788), .ZN(
        n12493) );
  NAND2_X1 U8614 ( .A1(n6856), .A2(n6854), .ZN(n12312) );
  NAND2_X1 U8615 ( .A1(n6857), .A2(n11887), .ZN(n6856) );
  INV_X1 U8616 ( .A(n6855), .ZN(n6854) );
  NOR2_X1 U8617 ( .A1(n7511), .A2(n7519), .ZN(n6857) );
  NAND2_X1 U8618 ( .A1(n7352), .A2(n12284), .ZN(n12316) );
  AOI21_X1 U8619 ( .B1(n12126), .B2(n12125), .A(n12124), .ZN(n12281) );
  INV_X1 U8620 ( .A(n7352), .ZN(n12133) );
  NAND2_X1 U8621 ( .A1(n15457), .A2(n11647), .ZN(n11659) );
  NAND2_X1 U8622 ( .A1(n11640), .A2(n11639), .ZN(n11654) );
  NOR2_X1 U8623 ( .A1(n11810), .A2(n15449), .ZN(n11647) );
  NAND2_X1 U8624 ( .A1(n7492), .A2(n6860), .ZN(n7490) );
  NAND2_X1 U8625 ( .A1(n7348), .A2(n7347), .ZN(n11810) );
  INV_X1 U8626 ( .A(n7348), .ZN(n11822) );
  INV_X1 U8627 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U8628 ( .A1(n11778), .A2(n12906), .ZN(n11777) );
  NAND2_X1 U8629 ( .A1(n7346), .A2(n7345), .ZN(n11795) );
  NAND2_X1 U8630 ( .A1(n11437), .A2(n7489), .ZN(n7486) );
  AND2_X1 U8631 ( .A1(n11437), .A2(n11415), .ZN(n7488) );
  INV_X1 U8632 ( .A(n7489), .ZN(n12901) );
  NAND2_X1 U8633 ( .A1(n11416), .A2(n11415), .ZN(n11417) );
  INV_X1 U8634 ( .A(n7445), .ZN(n12900) );
  NAND2_X1 U8635 ( .A1(n10970), .A2(n12900), .ZN(n11416) );
  CLKBUF_X1 U8636 ( .A(n10979), .Z(n15471) );
  NAND2_X1 U8637 ( .A1(n8665), .A2(n12846), .ZN(n6846) );
  OR2_X1 U8638 ( .A1(n8575), .A2(n8571), .ZN(n6989) );
  OR2_X1 U8639 ( .A1(n8754), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8756) );
  OR2_X1 U8640 ( .A1(n8756), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8794) );
  OR2_X1 U8641 ( .A1(n8677), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U8642 ( .A1(n6993), .A2(n6992), .ZN(n14266) );
  INV_X1 U8643 ( .A(n14269), .ZN(n6992) );
  NAND2_X1 U8644 ( .A1(n8312), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8327) );
  NOR2_X1 U8645 ( .A1(n8058), .A2(n11950), .ZN(n8078) );
  OR2_X1 U8647 ( .A1(n6996), .A2(n14318), .ZN(n7608) );
  INV_X1 U8648 ( .A(n8327), .ZN(n8328) );
  NAND2_X1 U8649 ( .A1(n7593), .A2(n7597), .ZN(n14334) );
  NAND2_X1 U8650 ( .A1(n14352), .A2(n7599), .ZN(n7593) );
  OR2_X1 U8651 ( .A1(n7596), .A2(n14332), .ZN(n6694) );
  INV_X1 U8652 ( .A(n7597), .ZN(n7596) );
  AOI21_X1 U8653 ( .B1(n7597), .B2(n7600), .A(n7595), .ZN(n7594) );
  INV_X1 U8654 ( .A(n14333), .ZN(n7595) );
  INV_X4 U8655 ( .A(n10457), .ZN(n10444) );
  OR2_X1 U8656 ( .A1(n8269), .A2(n7763), .ZN(n8280) );
  OR2_X1 U8657 ( .A1(n8280), .A2(n14346), .ZN(n8292) );
  NOR2_X1 U8658 ( .A1(n8292), .A2(n14299), .ZN(n8310) );
  OR2_X1 U8659 ( .A1(n8096), .A2(n15092), .ZN(n8136) );
  OR2_X1 U8660 ( .A1(n8121), .A2(n8114), .ZN(n8172) );
  NOR2_X1 U8661 ( .A1(n8172), .A2(n8171), .ZN(n8195) );
  AND2_X1 U8662 ( .A1(n8491), .A2(n8490), .ZN(n7759) );
  NAND2_X1 U8663 ( .A1(n7187), .A2(n7186), .ZN(n7185) );
  NAND2_X1 U8664 ( .A1(n7184), .A2(n7183), .ZN(n7182) );
  AND4_X1 U8665 ( .A1(n8007), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(n11279)
         );
  AOI21_X1 U8666 ( .B1(n10592), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14458), .ZN(
        n10595) );
  AOI21_X1 U8667 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10636), .A(n10635), .ZN(
        n10639) );
  INV_X1 U8668 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11950) );
  OR2_X1 U8669 ( .A1(n8130), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8144) );
  AOI21_X1 U8670 ( .B1(n12141), .B2(P1_REG1_REG_13__SCAN_IN), .A(n12140), .ZN(
        n14481) );
  XNOR2_X1 U8671 ( .A(n12142), .B(n12153), .ZN(n15187) );
  NAND2_X1 U8672 ( .A1(n7886), .A2(n9493), .ZN(n7200) );
  NOR2_X1 U8673 ( .A1(n6701), .A2(n14830), .ZN(n7261) );
  INV_X1 U8674 ( .A(n7387), .ZN(n7383) );
  AND4_X1 U8675 ( .A1(n8379), .A2(n8378), .A3(n8377), .A4(n8376), .ZN(n14309)
         );
  INV_X1 U8676 ( .A(n14583), .ZN(n14616) );
  INV_X1 U8677 ( .A(n7705), .ZN(n14628) );
  OAI211_X1 U8678 ( .C1(n14684), .C2(n7706), .A(n7704), .B(n6783), .ZN(n7705)
         );
  OR2_X1 U8679 ( .A1(n7710), .A2(n14643), .ZN(n7706) );
  INV_X1 U8680 ( .A(n8353), .ZN(n8354) );
  OR2_X1 U8681 ( .A1(n14877), .A2(n14573), .ZN(n14574) );
  NAND2_X1 U8682 ( .A1(n7270), .A2(n14742), .ZN(n7269) );
  OR2_X1 U8683 ( .A1(n14883), .A2(n6715), .ZN(n14720) );
  INV_X1 U8684 ( .A(n7717), .ZN(n7715) );
  NOR2_X1 U8685 ( .A1(n7724), .A2(n7720), .ZN(n7717) );
  NAND2_X1 U8686 ( .A1(n7726), .A2(n7725), .ZN(n7724) );
  INV_X1 U8687 ( .A(n14733), .ZN(n7725) );
  AOI21_X1 U8688 ( .B1(n7365), .B2(n7372), .A(n7363), .ZN(n7362) );
  INV_X1 U8689 ( .A(n14568), .ZN(n7363) );
  NOR2_X1 U8690 ( .A1(n14789), .A2(n7268), .ZN(n14747) );
  INV_X1 U8691 ( .A(n7270), .ZN(n7268) );
  NOR2_X1 U8692 ( .A1(n14789), .A2(n7271), .ZN(n14761) );
  OR2_X1 U8693 ( .A1(n14788), .A2(n14911), .ZN(n14789) );
  NOR2_X1 U8694 ( .A1(n14789), .A2(n14905), .ZN(n14776) );
  NOR2_X1 U8695 ( .A1(n14797), .A2(n7739), .ZN(n7738) );
  INV_X1 U8696 ( .A(n14536), .ZN(n7739) );
  NOR2_X1 U8697 ( .A1(n8136), .A2(n10953), .ZN(n8137) );
  AOI21_X1 U8698 ( .B1(n6695), .B2(n7358), .A(n6774), .ZN(n7353) );
  NOR3_X1 U8699 ( .A1(n11522), .A2(n15284), .A3(n7257), .ZN(n15113) );
  NAND2_X1 U8700 ( .A1(n15116), .A2(n7258), .ZN(n7257) );
  INV_X1 U8701 ( .A(n7259), .ZN(n7258) );
  NOR3_X1 U8702 ( .A1(n11522), .A2(n7259), .A3(n15284), .ZN(n15115) );
  OR2_X1 U8703 ( .A1(n8017), .A2(n8016), .ZN(n8039) );
  OR2_X1 U8704 ( .A1(n8039), .A2(n8038), .ZN(n8058) );
  NAND2_X1 U8705 ( .A1(n11514), .A2(n11704), .ZN(n11698) );
  NOR2_X1 U8706 ( .A1(n7975), .A2(n7974), .ZN(n8001) );
  INV_X1 U8707 ( .A(n11276), .ZN(n11281) );
  OR2_X1 U8708 ( .A1(n11217), .A2(n11281), .ZN(n11313) );
  NAND2_X1 U8709 ( .A1(n11201), .A2(n11208), .ZN(n11283) );
  NAND2_X1 U8710 ( .A1(n11207), .A2(n11206), .ZN(n11209) );
  OAI21_X1 U8711 ( .B1(n15201), .B2(n15200), .A(n11151), .ZN(n11176) );
  NAND2_X1 U8712 ( .A1(n11047), .A2(n11046), .ZN(n15207) );
  NOR2_X1 U8713 ( .A1(n15207), .A2(n15206), .ZN(n15208) );
  INV_X1 U8714 ( .A(n14533), .ZN(n14818) );
  NAND2_X1 U8715 ( .A1(n7386), .A2(n7384), .ZN(n14600) );
  AND2_X1 U8716 ( .A1(n7386), .A2(n6729), .ZN(n14602) );
  NAND2_X1 U8717 ( .A1(n7999), .A2(n7998), .ZN(n11314) );
  INV_X1 U8718 ( .A(n15283), .ZN(n15246) );
  INV_X1 U8719 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7786) );
  XNOR2_X1 U8720 ( .A(n8546), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U8721 ( .A1(n6824), .A2(n6707), .ZN(n7256) );
  XNOR2_X1 U8722 ( .A(n8336), .B(SI_22_), .ZN(n9004) );
  NAND2_X1 U8723 ( .A1(n6965), .A2(n6964), .ZN(n8537) );
  INV_X1 U8724 ( .A(n7889), .ZN(n6965) );
  AOI21_X1 U8725 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8304) );
  XNOR2_X1 U8726 ( .A(n7880), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U8727 ( .A1(n7859), .A2(n7049), .ZN(n8262) );
  OR2_X1 U8728 ( .A1(n8250), .A2(n7857), .ZN(n7049) );
  NAND2_X1 U8729 ( .A1(n7543), .A2(n7854), .ZN(n8219) );
  NAND2_X1 U8730 ( .A1(n8204), .A2(n8203), .ZN(n7543) );
  XNOR2_X1 U8731 ( .A(n7993), .B(n7992), .ZN(n10555) );
  INV_X1 U8732 ( .A(n7809), .ZN(n7919) );
  INV_X1 U8733 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U8734 ( .A1(n9169), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9168) );
  XNOR2_X1 U8735 ( .A(n9167), .B(n7004), .ZN(n9170) );
  INV_X1 U8736 ( .A(n9168), .ZN(n7004) );
  OAI21_X1 U8737 ( .B1(n9167), .B2(n9168), .A(n7280), .ZN(n7007) );
  NAND2_X1 U8738 ( .A1(n9130), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7280) );
  INV_X1 U8739 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U8740 ( .A(n9131), .B(n9335), .ZN(n9175) );
  XNOR2_X1 U8741 ( .A(n9179), .B(n7037), .ZN(n9181) );
  INV_X1 U8742 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7037) );
  NOR2_X1 U8743 ( .A1(n15694), .A2(n9178), .ZN(n9180) );
  NOR2_X1 U8744 ( .A1(n9135), .A2(n9134), .ZN(n9184) );
  NOR2_X1 U8745 ( .A1(n14967), .A2(n9187), .ZN(n9189) );
  XOR2_X1 U8746 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9139), .Z(n9188) );
  OAI21_X1 U8747 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n9194), .A(n6936), .ZN(
        n6935) );
  AOI21_X1 U8748 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n9149), .A(n9148), .ZN(
        n9200) );
  NOR2_X1 U8749 ( .A1(n9165), .A2(n9164), .ZN(n9148) );
  OAI22_X1 U8750 ( .A1(n9202), .A2(n9153), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n9152), .ZN(n9162) );
  NAND2_X1 U8751 ( .A1(n9996), .A2(n9995), .ZN(n13352) );
  NAND2_X1 U8752 ( .A1(n12246), .A2(n12245), .ZN(n12247) );
  NAND2_X1 U8753 ( .A1(n13123), .A2(n12587), .ZN(n13019) );
  NAND2_X1 U8754 ( .A1(n13084), .A2(n12593), .ZN(n13040) );
  NAND2_X1 U8755 ( .A1(n9928), .A2(n9927), .ZN(n13430) );
  AND4_X1 U8756 ( .A1(n9782), .A2(n9781), .A3(n9780), .A4(n9779), .ZN(n13055)
         );
  NAND2_X1 U8757 ( .A1(n13145), .A2(n12579), .ZN(n13070) );
  NAND2_X1 U8758 ( .A1(n13079), .A2(n13078), .ZN(n13077) );
  AND4_X1 U8759 ( .A1(n9738), .A2(n9737), .A3(n9736), .A4(n9735), .ZN(n12215)
         );
  NAND2_X1 U8760 ( .A1(n12186), .A2(n12185), .ZN(n12189) );
  INV_X1 U8761 ( .A(n13138), .ZN(n15492) );
  NAND2_X1 U8762 ( .A1(n13086), .A2(n13085), .ZN(n13084) );
  NAND2_X1 U8763 ( .A1(n13020), .A2(n12590), .ZN(n13086) );
  OAI21_X1 U8764 ( .B1(n13049), .B2(n13114), .A(n13047), .ZN(n6913) );
  AND2_X1 U8765 ( .A1(n9933), .A2(n9932), .ZN(n13439) );
  NAND2_X1 U8766 ( .A1(n9938), .A2(n9937), .ZN(n13107) );
  AND4_X1 U8767 ( .A1(n9769), .A2(n9768), .A3(n9767), .A4(n9766), .ZN(n13116)
         );
  NAND2_X1 U8768 ( .A1(n6895), .A2(n6896), .ZN(n12068) );
  INV_X1 U8769 ( .A(n13359), .ZN(n13139) );
  NAND2_X1 U8770 ( .A1(n6899), .A2(n6710), .ZN(n6905) );
  NAND2_X1 U8771 ( .A1(n13060), .A2(n13061), .ZN(n6899) );
  NAND2_X1 U8772 ( .A1(n9982), .A2(n9981), .ZN(n13552) );
  INV_X1 U8773 ( .A(n15490), .ZN(n13154) );
  NAND2_X1 U8774 ( .A1(n11353), .A2(n12608), .ZN(n13149) );
  OAI211_X1 U8775 ( .C1(n11352), .C2(P3_U3151), .A(n11351), .B(n11528), .ZN(
        n13151) );
  NAND2_X1 U8776 ( .A1(n13147), .A2(n13146), .ZN(n13145) );
  AND2_X1 U8777 ( .A1(n7638), .A2(n7640), .ZN(n6943) );
  OR2_X1 U8778 ( .A1(n13660), .A2(n11348), .ZN(n13155) );
  AND2_X1 U8779 ( .A1(n10027), .A2(n9617), .ZN(n12545) );
  INV_X1 U8780 ( .A(n12992), .ZN(n13391) );
  NAND2_X1 U8781 ( .A1(n9966), .A2(n9965), .ZN(n13371) );
  AND4_X1 U8782 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n13491)
         );
  INV_X1 U8783 ( .A(n13128), .ZN(n13504) );
  INV_X1 U8784 ( .A(n13531), .ZN(n13114) );
  INV_X1 U8785 ( .A(n13055), .ZN(n13111) );
  INV_X1 U8786 ( .A(n13116), .ZN(n12563) );
  INV_X1 U8787 ( .A(n12215), .ZN(n12220) );
  INV_X1 U8788 ( .A(n12054), .ZN(n15562) );
  NAND2_X1 U8789 ( .A1(n9646), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U8790 ( .A1(n9646), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U8791 ( .A1(n9847), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U8792 ( .A1(n11550), .A2(n11551), .ZN(n11691) );
  NAND2_X1 U8793 ( .A1(n7098), .A2(n7096), .ZN(n11754) );
  INV_X1 U8794 ( .A(n7097), .ZN(n7096) );
  OAI21_X1 U8795 ( .B1(n6719), .B2(n11753), .A(n11752), .ZN(n7097) );
  INV_X1 U8796 ( .A(n6871), .ZN(n11847) );
  NAND2_X1 U8797 ( .A1(n7090), .A2(n7091), .ZN(n11992) );
  INV_X1 U8798 ( .A(n7039), .ZN(n12003) );
  INV_X1 U8799 ( .A(n7339), .ZN(n11979) );
  INV_X1 U8800 ( .A(n7551), .ZN(n15546) );
  NAND2_X1 U8801 ( .A1(n15552), .A2(n15551), .ZN(n15549) );
  INV_X1 U8802 ( .A(n7332), .ZN(n15541) );
  INV_X1 U8803 ( .A(n7330), .ZN(n15542) );
  INV_X1 U8804 ( .A(n6869), .ZN(n13201) );
  INV_X1 U8805 ( .A(n7078), .ZN(n13269) );
  AND2_X1 U8806 ( .A1(n13267), .A2(n13266), .ZN(n6955) );
  OAI21_X1 U8807 ( .B1(n13313), .B2(n7563), .A(n15500), .ZN(n7562) );
  AND2_X1 U8808 ( .A1(n13304), .A2(n13303), .ZN(n7563) );
  NAND2_X1 U8809 ( .A1(n6865), .A2(n6867), .ZN(n6864) );
  NAND2_X1 U8810 ( .A1(n13321), .A2(n13311), .ZN(n6867) );
  NOR2_X1 U8811 ( .A1(n7328), .A2(n13310), .ZN(n7321) );
  NAND2_X1 U8812 ( .A1(n9601), .A2(n9600), .ZN(n15040) );
  AND2_X1 U8813 ( .A1(n10012), .A2(n13034), .ZN(n15030) );
  OAI21_X1 U8814 ( .B1(n13334), .B2(n13333), .A(n13336), .ZN(n13545) );
  AND2_X1 U8815 ( .A1(n13343), .A2(n7311), .ZN(n13333) );
  NAND2_X1 U8816 ( .A1(n13384), .A2(n10189), .ZN(n13377) );
  NAND2_X1 U8817 ( .A1(n7657), .A2(n7658), .ZN(n13476) );
  NAND2_X1 U8818 ( .A1(n12519), .A2(n12518), .ZN(n13515) );
  INV_X1 U8819 ( .A(n13539), .ZN(n13524) );
  NAND2_X1 U8820 ( .A1(n7660), .A2(n9763), .ZN(n12300) );
  NAND2_X1 U8821 ( .A1(n7645), .A2(n9730), .ZN(n12160) );
  NAND2_X1 U8822 ( .A1(n11958), .A2(n11957), .ZN(n7645) );
  OR2_X1 U8823 ( .A1(n11529), .A2(n11357), .ZN(n15591) );
  AND2_X1 U8824 ( .A1(n11483), .A2(n13325), .ZN(n15609) );
  AOI21_X1 U8825 ( .B1(n9805), .B2(n10531), .A(n6949), .ZN(n6948) );
  NOR2_X1 U8826 ( .A1(n10229), .A2(n6887), .ZN(n6949) );
  NAND2_X1 U8827 ( .A1(n11505), .A2(n15591), .ZN(n15625) );
  AND3_X2 U8828 ( .A1(n12633), .A2(n12632), .A3(n12631), .ZN(n15693) );
  AND2_X1 U8829 ( .A1(n15038), .A2(n15037), .ZN(n15060) );
  INV_X1 U8830 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n7012) );
  INV_X1 U8831 ( .A(n12602), .ZN(n13623) );
  INV_X1 U8832 ( .A(n13015), .ZN(n13627) );
  NAND2_X1 U8833 ( .A1(n9915), .A2(n9914), .ZN(n13638) );
  NAND2_X1 U8834 ( .A1(n9904), .A2(n9903), .ZN(n13644) );
  AND2_X1 U8835 ( .A1(n12617), .A2(n12616), .ZN(n15681) );
  INV_X2 U8836 ( .A(n15681), .ZN(n15679) );
  OR2_X1 U8837 ( .A1(n15681), .A2(n15607), .ZN(n13657) );
  NAND2_X1 U8838 ( .A1(n11531), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13660) );
  NAND2_X1 U8839 ( .A1(n10217), .A2(n9604), .ZN(n13664) );
  XNOR2_X1 U8840 ( .A(n9623), .B(n7208), .ZN(n13663) );
  INV_X1 U8841 ( .A(n9622), .ZN(n7208) );
  XNOR2_X1 U8842 ( .A(n10018), .B(n10017), .ZN(n12640) );
  NAND2_X1 U8843 ( .A1(n10222), .A2(n10221), .ZN(n12280) );
  NAND2_X1 U8844 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n9595), .ZN(n7014) );
  NAND2_X1 U8845 ( .A1(n9956), .A2(n12209), .ZN(n7626) );
  AND2_X1 U8846 ( .A1(n10225), .A2(n9594), .ZN(n7035) );
  INV_X1 U8847 ( .A(SI_23_), .ZN(n11511) );
  AND2_X1 U8848 ( .A1(n7630), .A2(n7629), .ZN(n9946) );
  XNOR2_X1 U8849 ( .A(n10062), .B(n10061), .ZN(n13540) );
  INV_X1 U8850 ( .A(SI_19_), .ZN(n10831) );
  INV_X1 U8851 ( .A(n13325), .ZN(n13314) );
  INV_X1 U8852 ( .A(SI_16_), .ZN(n10693) );
  NAND2_X1 U8853 ( .A1(n7619), .A2(n9570), .ZN(n9839) );
  NAND2_X1 U8854 ( .A1(n9825), .A2(n9824), .ZN(n7619) );
  NAND2_X1 U8855 ( .A1(n9800), .A2(n9588), .ZN(n9840) );
  INV_X1 U8856 ( .A(SI_13_), .ZN(n10569) );
  NAND2_X1 U8857 ( .A1(n7667), .A2(n7666), .ZN(n9798) );
  INV_X1 U8858 ( .A(SI_12_), .ZN(n10546) );
  INV_X1 U8859 ( .A(SI_11_), .ZN(n10519) );
  INV_X1 U8860 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9783) );
  INV_X1 U8861 ( .A(n12007), .ZN(n11999) );
  INV_X1 U8862 ( .A(n7219), .ZN(n9727) );
  AOI21_X1 U8863 ( .B1(n7224), .B2(n7222), .A(n6685), .ZN(n7219) );
  NAND2_X1 U8864 ( .A1(n7224), .A2(n9555), .ZN(n9713) );
  INV_X1 U8865 ( .A(n11588), .ZN(n11577) );
  NAND2_X1 U8866 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7566) );
  NAND2_X1 U8867 ( .A1(n10225), .A2(n9587), .ZN(n7565) );
  AND2_X1 U8868 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7335) );
  NAND2_X1 U8869 ( .A1(n7479), .A2(n7478), .ZN(n12197) );
  AND2_X1 U8870 ( .A1(n7479), .A2(n6737), .ZN(n12198) );
  NAND2_X1 U8871 ( .A1(n11937), .A2(n7480), .ZN(n7479) );
  NAND2_X1 U8872 ( .A1(n11164), .A2(n8793), .ZN(n11269) );
  AND4_X1 U8873 ( .A1(n8690), .A2(n8689), .A3(n8688), .A4(n8687), .ZN(n12678)
         );
  NAND2_X1 U8874 ( .A1(n6990), .A2(n6718), .ZN(n7449) );
  NAND2_X1 U8875 ( .A1(n13748), .A2(n8986), .ZN(n13703) );
  NAND2_X1 U8876 ( .A1(n7473), .A2(n8891), .ZN(n13721) );
  NAND2_X1 U8877 ( .A1(n8900), .A2(n8899), .ZN(n14207) );
  NAND2_X1 U8878 ( .A1(n11165), .A2(n11166), .ZN(n11164) );
  AOI21_X1 U8879 ( .B1(n7450), .B2(n7452), .A(n7448), .ZN(n7447) );
  INV_X1 U8880 ( .A(n13681), .ZN(n7448) );
  AND2_X1 U8881 ( .A1(n11937), .A2(n8848), .ZN(n12011) );
  NAND2_X1 U8882 ( .A1(n7456), .A2(n7458), .ZN(n11623) );
  NAND2_X1 U8883 ( .A1(n8816), .A2(n8815), .ZN(n12736) );
  AND4_X1 U8884 ( .A1(n8670), .A2(n8672), .A3(n8671), .A4(n8673), .ZN(n11404)
         );
  NAND2_X1 U8885 ( .A1(n6990), .A2(n8934), .ZN(n13765) );
  NAND2_X1 U8886 ( .A1(n8939), .A2(n8938), .ZN(n14195) );
  NAND2_X1 U8887 ( .A1(n8610), .A2(n8609), .ZN(n14154) );
  NAND2_X1 U8888 ( .A1(n10890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13781) );
  NAND2_X1 U8889 ( .A1(n7136), .A2(n7137), .ZN(n12941) );
  NAND2_X1 U8890 ( .A1(n12838), .A2(n7674), .ZN(n7137) );
  NAND2_X1 U8891 ( .A1(n7135), .A2(n7134), .ZN(n7136) );
  INV_X1 U8892 ( .A(n8612), .ZN(n12961) );
  AND2_X1 U8893 ( .A1(n8727), .A2(n6853), .ZN(n6852) );
  INV_X1 U8894 ( .A(n11404), .ZN(n13798) );
  AND2_X1 U8895 ( .A1(n15366), .A2(n15365), .ZN(n15367) );
  INV_X1 U8896 ( .A(n13876), .ZN(n14138) );
  NAND2_X1 U8897 ( .A1(n7437), .A2(n13896), .ZN(n14003) );
  NAND2_X1 U8898 ( .A1(n6995), .A2(n7438), .ZN(n7437) );
  AND2_X1 U8899 ( .A1(n7067), .A2(n6739), .ZN(n13999) );
  OAI21_X1 U8900 ( .B1(n14075), .B2(n7497), .A(n7494), .ZN(n14029) );
  AOI21_X1 U8901 ( .B1(n13891), .B2(n7425), .A(n6689), .ZN(n14055) );
  NAND2_X1 U8902 ( .A1(n7498), .A2(n7499), .ZN(n14045) );
  NAND2_X1 U8903 ( .A1(n13891), .A2(n7428), .ZN(n14067) );
  AOI21_X1 U8904 ( .B1(n14075), .B2(n14072), .A(n7502), .ZN(n14059) );
  NAND2_X1 U8905 ( .A1(n7515), .A2(n7512), .ZN(n12289) );
  INV_X1 U8906 ( .A(n7517), .ZN(n12128) );
  NAND2_X1 U8907 ( .A1(n11802), .A2(n11466), .ZN(n11467) );
  AND2_X1 U8908 ( .A1(n11465), .A2(n11464), .ZN(n11803) );
  NAND2_X1 U8909 ( .A1(n11831), .A2(n11443), .ZN(n11818) );
  AND2_X1 U8910 ( .A1(n12926), .A2(n12897), .ZN(n15385) );
  AND3_X2 U8911 ( .A1(n10965), .A2(n12121), .A3(n12122), .ZN(n15489) );
  NOR2_X1 U8912 ( .A1(n7408), .A2(n15454), .ZN(n7407) );
  NOR2_X1 U8913 ( .A1(n14144), .A2(n6849), .ZN(n14146) );
  AND2_X1 U8914 ( .A1(n14145), .A2(n15450), .ZN(n6850) );
  AND3_X2 U8915 ( .A1(n12122), .A2(n12121), .A3(n12120), .ZN(n15475) );
  INV_X1 U8916 ( .A(n15396), .ZN(n15401) );
  AND2_X1 U8917 ( .A1(n8607), .A2(n8587), .ZN(n7522) );
  XNOR2_X1 U8918 ( .A(n9078), .B(n9077), .ZN(n14255) );
  OAI21_X1 U8919 ( .B1(n9076), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9078) );
  INV_X1 U8920 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12332) );
  XNOR2_X1 U8921 ( .A(n9069), .B(n9068), .ZN(n12330) );
  NAND2_X1 U8922 ( .A1(n9073), .A2(n9076), .ZN(n12210) );
  INV_X1 U8923 ( .A(n9072), .ZN(n9073) );
  INV_X1 U8924 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12040) );
  INV_X1 U8925 ( .A(n10971), .ZN(n12897) );
  INV_X1 U8926 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10927) );
  INV_X1 U8927 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10691) );
  INV_X1 U8928 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10544) );
  INV_X1 U8929 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10509) );
  NAND2_X1 U8930 ( .A1(n7573), .A2(n10260), .ZN(n10930) );
  AND2_X1 U8931 ( .A1(n10588), .A2(n10560), .ZN(n14986) );
  NAND2_X1 U8932 ( .A1(n15103), .A2(n7585), .ZN(n15082) );
  INV_X1 U8933 ( .A(n7608), .ZN(n14317) );
  OAI21_X1 U8934 ( .B1(n14352), .B2(n6694), .A(n6682), .ZN(n14336) );
  OAI21_X1 U8935 ( .B1(n10333), .B2(n7584), .A(n7583), .ZN(n12394) );
  AOI21_X1 U8936 ( .B1(n7585), .B2(n15099), .A(n6741), .ZN(n7583) );
  INV_X1 U8937 ( .A(n7585), .ZN(n7584) );
  AOI21_X1 U8938 ( .B1(n14352), .B2(n14351), .A(n14350), .ZN(n14354) );
  INV_X1 U8939 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n15092) );
  NAND2_X1 U8940 ( .A1(n7601), .A2(n7605), .ZN(n14360) );
  OR2_X1 U8941 ( .A1(n6996), .A2(n7606), .ZN(n7601) );
  OR2_X1 U8942 ( .A1(n15093), .A2(n15246), .ZN(n14388) );
  AOI21_X1 U8943 ( .B1(n10620), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10664), .ZN(
        n10618) );
  AOI21_X1 U8944 ( .B1(n10833), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10832), .ZN(
        n10836) );
  NOR2_X1 U8945 ( .A1(n14505), .A2(n14504), .ZN(n14506) );
  XNOR2_X1 U8946 ( .A(n7263), .B(n7262), .ZN(n14814) );
  INV_X1 U8947 ( .A(n7376), .ZN(n14659) );
  NAND2_X1 U8948 ( .A1(n14674), .A2(n6721), .ZN(n14660) );
  NAND2_X1 U8949 ( .A1(n7707), .A2(n6686), .ZN(n14656) );
  NAND2_X1 U8950 ( .A1(n14684), .A2(n6717), .ZN(n7707) );
  OAI21_X1 U8951 ( .B1(n14684), .B2(n14685), .A(n6712), .ZN(n14671) );
  NAND2_X1 U8952 ( .A1(n14954), .A2(n10562), .ZN(n14692) );
  NAND2_X1 U8953 ( .A1(n14725), .A2(n7748), .ZN(n14700) );
  AND2_X1 U8954 ( .A1(n7559), .A2(n8286), .ZN(n10382) );
  NAND2_X1 U8955 ( .A1(n11884), .A2(n8484), .ZN(n7559) );
  INV_X1 U8956 ( .A(n14888), .ZN(n14742) );
  AOI21_X1 U8957 ( .B1(n14769), .B2(n14770), .A(n7719), .ZN(n14753) );
  INV_X1 U8958 ( .A(n7721), .ZN(n7719) );
  NAND2_X1 U8959 ( .A1(n7367), .A2(n7369), .ZN(n14746) );
  OR2_X1 U8960 ( .A1(n14785), .A2(n7372), .ZN(n7367) );
  NAND2_X1 U8961 ( .A1(n7368), .A2(n7374), .ZN(n14760) );
  NAND2_X1 U8962 ( .A1(n14785), .A2(n7375), .ZN(n7368) );
  AND2_X1 U8963 ( .A1(n7740), .A2(n7738), .ZN(n14915) );
  NAND2_X1 U8964 ( .A1(n7740), .A2(n14536), .ZN(n14798) );
  NAND2_X1 U8965 ( .A1(n12409), .A2(n12408), .ZN(n14538) );
  NAND2_X1 U8966 ( .A1(n8133), .A2(n8132), .ZN(n15130) );
  NAND2_X1 U8967 ( .A1(n7356), .A2(n7357), .ZN(n14982) );
  OR2_X1 U8968 ( .A1(n12034), .A2(n7358), .ZN(n7356) );
  NAND2_X1 U8969 ( .A1(n8106), .A2(n8105), .ZN(n15122) );
  NAND2_X1 U8970 ( .A1(n12342), .A2(n12341), .ZN(n15108) );
  NAND2_X1 U8971 ( .A1(n12350), .A2(n12349), .ZN(n15111) );
  NOR2_X1 U8972 ( .A1(n7702), .A2(n6687), .ZN(n12023) );
  INV_X1 U8973 ( .A(n12021), .ZN(n7702) );
  NAND2_X1 U8974 ( .A1(n7197), .A2(n7196), .ZN(n7195) );
  INV_X1 U8975 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8976 ( .A1(n7698), .A2(n11519), .ZN(n11703) );
  NAND2_X1 U8977 ( .A1(n11517), .A2(n11516), .ZN(n7698) );
  NAND2_X1 U8978 ( .A1(n8030), .A2(n8029), .ZN(n15263) );
  NOR2_X1 U8979 ( .A1(n6676), .A2(n11141), .ZN(n15126) );
  NAND2_X1 U8980 ( .A1(n15120), .A2(n11157), .ZN(n14780) );
  OAI211_X2 U8981 ( .C1(n10562), .C2(n14456), .A(n7965), .B(n7964), .ZN(n11203) );
  INV_X1 U8982 ( .A(n11047), .ZN(n15216) );
  INV_X1 U8983 ( .A(n14780), .ZN(n15215) );
  AND2_X1 U8984 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  AND3_X1 U8985 ( .A1(n14852), .A2(n14851), .A3(n14850), .ZN(n14854) );
  NAND2_X1 U8986 ( .A1(n7248), .A2(n7247), .ZN(n14237) );
  NAND2_X1 U8987 ( .A1(n8452), .A2(n6836), .ZN(n7247) );
  INV_X1 U8988 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n12508) );
  INV_X1 U8989 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7874) );
  XNOR2_X1 U8990 ( .A(n8415), .B(n8400), .ZN(n14945) );
  CLKBUF_X1 U8991 ( .A(n14947), .Z(n6988) );
  INV_X1 U8992 ( .A(n10465), .ZN(n14952) );
  INV_X1 U8993 ( .A(n10463), .ZN(n12207) );
  XNOR2_X1 U8994 ( .A(n8318), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14954) );
  OR2_X1 U8995 ( .A1(n9004), .A2(n10501), .ZN(n8318) );
  INV_X1 U8996 ( .A(n8486), .ZN(n11885) );
  NOR2_X1 U8997 ( .A1(n8166), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8205) );
  INV_X1 U8998 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11016) );
  INV_X1 U8999 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10689) );
  INV_X1 U9000 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10653) );
  OR3_X1 U9001 ( .A1(n8067), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n8068) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10572) );
  INV_X1 U9003 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10556) );
  XNOR2_X1 U9004 ( .A(n9170), .B(n10877), .ZN(n15709) );
  XNOR2_X1 U9005 ( .A(n9186), .B(n9185), .ZN(n14968) );
  NOR2_X1 U9006 ( .A1(n14968), .A2(n14969), .ZN(n14967) );
  NOR2_X1 U9007 ( .A1(n15702), .A2(n15703), .ZN(n15701) );
  NOR2_X1 U9008 ( .A1(n6922), .A2(n6921), .ZN(n14978) );
  NOR2_X1 U9009 ( .A1(n6937), .A2(n6938), .ZN(n6921) );
  NAND2_X1 U9010 ( .A1(n6935), .A2(n6933), .ZN(n6922) );
  INV_X1 U9011 ( .A(n9194), .ZN(n6937) );
  AND2_X1 U9012 ( .A1(n7018), .A2(n7019), .ZN(n15150) );
  NAND2_X1 U9013 ( .A1(n15150), .A2(n15149), .ZN(n15148) );
  OR2_X1 U9014 ( .A1(n7273), .A2(n9201), .ZN(n15155) );
  NAND2_X1 U9015 ( .A1(n15152), .A2(n15154), .ZN(n15158) );
  AND2_X1 U9016 ( .A1(n7278), .A2(n7276), .ZN(n15166) );
  NAND2_X1 U9017 ( .A1(n7274), .A2(n15165), .ZN(n15005) );
  OAI21_X1 U9018 ( .B1(n15166), .B2(n15167), .A(n7275), .ZN(n7274) );
  INV_X1 U9019 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7275) );
  INV_X1 U9020 ( .A(n6923), .ZN(n15004) );
  NAND2_X1 U9021 ( .A1(n12098), .A2(n12050), .ZN(n12088) );
  NAND2_X1 U9022 ( .A1(n6823), .A2(n15494), .ZN(n7401) );
  NAND2_X1 U9023 ( .A1(n12048), .A2(n12111), .ZN(n12100) );
  NAND2_X1 U9024 ( .A1(n7099), .A2(n7100), .ZN(n11693) );
  INV_X1 U9025 ( .A(n6870), .ZN(n11998) );
  OAI211_X1 U9026 ( .C1(n13313), .C2(n6864), .A(n15500), .B(n6862), .ZN(n6868)
         );
  AOI21_X1 U9027 ( .B1(n13606), .B2(n13582), .A(n7317), .ZN(n7316) );
  NAND2_X1 U9028 ( .A1(n7013), .A2(n6942), .ZN(P3_U3456) );
  NOR2_X1 U9029 ( .A1(n6958), .A2(n6833), .ZN(n6942) );
  NOR2_X1 U9030 ( .A1(n9103), .A2(n9102), .ZN(n13692) );
  NAND2_X1 U9031 ( .A1(n7466), .A2(n7471), .ZN(n7465) );
  AOI21_X1 U9032 ( .B1(n7482), .B2(n7032), .A(n7029), .ZN(n13718) );
  NAND2_X1 U9033 ( .A1(n7031), .A2(n7030), .ZN(n7029) );
  AOI21_X1 U9034 ( .B1(n13715), .B2(n13716), .A(n13785), .ZN(n7032) );
  OAI21_X1 U9035 ( .B1(n14142), .B2(n15394), .A(n7074), .ZN(P2_U3236) );
  INV_X1 U9036 ( .A(n7075), .ZN(n7074) );
  OAI21_X1 U9037 ( .B1(n14143), .B2(n14133), .A(n7076), .ZN(n7075) );
  NAND2_X1 U9038 ( .A1(n6848), .A2(n15392), .ZN(n13949) );
  NOR2_X1 U9039 ( .A1(n14151), .A2(n15394), .ZN(n13962) );
  NAND2_X1 U9040 ( .A1(n7579), .A2(n15081), .ZN(n7575) );
  NOR2_X1 U9041 ( .A1(n14970), .A2(n9194), .ZN(n14975) );
  INV_X1 U9042 ( .A(n7019), .ZN(n15144) );
  INV_X1 U9043 ( .A(n7278), .ZN(n15161) );
  INV_X1 U9044 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7010) );
  NOR2_X1 U9045 ( .A1(n7044), .A2(n6932), .ZN(n14958) );
  AND2_X1 U9046 ( .A1(n6744), .A2(n14957), .ZN(n6932) );
  XNOR2_X1 U9047 ( .A(n9545), .B(n6841), .ZN(n7282) );
  NAND2_X1 U9048 ( .A1(n7283), .A2(n7284), .ZN(n6941) );
  CLKBUF_X3 U9049 ( .A(n12844), .Z(n12825) );
  OR2_X1 U9050 ( .A1(n7594), .A2(n14332), .ZN(n6682) );
  NAND2_X1 U9051 ( .A1(n12772), .A2(n7676), .ZN(n6683) );
  NOR2_X1 U9052 ( .A1(n13041), .A2(n7395), .ZN(n6684) );
  INV_X2 U9053 ( .A(n14018), .ZN(n8580) );
  INV_X1 U9054 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6887) );
  INV_X1 U9055 ( .A(n13957), .ZN(n7024) );
  AND2_X1 U9056 ( .A1(n10556), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6685) );
  OR2_X2 U9057 ( .A1(n7712), .A2(n7711), .ZN(n6686) );
  INV_X1 U9058 ( .A(n14643), .ZN(n7380) );
  NAND2_X1 U9059 ( .A1(n11404), .A2(n15410), .ZN(n11437) );
  AND2_X1 U9060 ( .A1(n12030), .A2(n12020), .ZN(n6687) );
  AND2_X1 U9061 ( .A1(n14679), .A2(n7267), .ZN(n6688) );
  AND2_X1 U9062 ( .A1(n14185), .A2(n13914), .ZN(n6689) );
  NAND2_X1 U9063 ( .A1(n7127), .A2(n12733), .ZN(n6690) );
  NAND2_X1 U9064 ( .A1(n9876), .A2(n6789), .ZN(n6691) );
  AND2_X1 U9065 ( .A1(n7104), .A2(n11551), .ZN(n6692) );
  AND2_X1 U9066 ( .A1(n6688), .A2(n7266), .ZN(n6693) );
  AND2_X1 U9067 ( .A1(n7357), .A2(n7355), .ZN(n6695) );
  INV_X1 U9068 ( .A(n13443), .ZN(n13437) );
  NAND2_X1 U9069 ( .A1(n8882), .A2(n8881), .ZN(n12771) );
  OR2_X1 U9070 ( .A1(n11705), .A2(n11709), .ZN(n6696) );
  XOR2_X1 U9071 ( .A(n6711), .B(n7402), .Z(n6697) );
  NAND2_X1 U9072 ( .A1(n10204), .A2(n10203), .ZN(n12548) );
  NAND2_X1 U9073 ( .A1(n8223), .A2(n8222), .ZN(n14899) );
  AND2_X1 U9074 ( .A1(n12724), .A2(n12723), .ZN(n6698) );
  OR2_X1 U9075 ( .A1(n14066), .A2(n13914), .ZN(n6699) );
  NAND2_X1 U9076 ( .A1(n8443), .A2(n7535), .ZN(n7534) );
  INV_X1 U9077 ( .A(n7534), .ZN(n7194) );
  AND2_X1 U9078 ( .A1(n12770), .A2(n12769), .ZN(n6700) );
  INV_X1 U9079 ( .A(n7306), .ZN(n7305) );
  OR2_X1 U9080 ( .A1(n12535), .A2(n7307), .ZN(n7306) );
  OR2_X1 U9081 ( .A1(n14533), .A2(n14822), .ZN(n6701) );
  NAND2_X1 U9082 ( .A1(n6926), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6702) );
  NOR2_X1 U9083 ( .A1(n14175), .A2(n13894), .ZN(n6703) );
  AND2_X1 U9084 ( .A1(n14325), .A2(n14324), .ZN(n6704) );
  INV_X1 U9085 ( .A(n14957), .ZN(n6930) );
  AND2_X1 U9086 ( .A1(n12789), .A2(n12788), .ZN(n6705) );
  OR2_X1 U9087 ( .A1(n7103), .A2(n11696), .ZN(n6706) );
  XNOR2_X1 U9088 ( .A(n9902), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U9089 ( .A1(n8585), .A2(n8568), .ZN(n8833) );
  INV_X1 U9090 ( .A(n14031), .ZN(n7047) );
  NOR2_X1 U9091 ( .A1(n7092), .A2(n11993), .ZN(n7089) );
  OR2_X1 U9092 ( .A1(n7865), .A2(SI_21_), .ZN(n6707) );
  OR2_X1 U9093 ( .A1(n11522), .A2(n7259), .ZN(n6708) );
  INV_X1 U9094 ( .A(n15539), .ZN(n15515) );
  INV_X1 U9095 ( .A(n13142), .ZN(n15494) );
  INV_X1 U9096 ( .A(n15417), .ZN(n7345) );
  AND2_X1 U9097 ( .A1(n12605), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7615) );
  INV_X1 U9098 ( .A(n13322), .ZN(n7328) );
  AND2_X1 U9099 ( .A1(n7238), .A2(n10017), .ZN(n6709) );
  INV_X2 U9100 ( .A(n8646), .ZN(n8666) );
  NAND2_X1 U9101 ( .A1(n12991), .A2(n12992), .ZN(n6710) );
  INV_X1 U9102 ( .A(n9847), .ZN(n9943) );
  XOR2_X1 U9103 ( .A(n12987), .B(n13402), .Z(n6711) );
  NAND2_X1 U9104 ( .A1(n9633), .A2(n6885), .ZN(n9679) );
  NAND2_X1 U9105 ( .A1(n6979), .A2(n9696), .ZN(n7224) );
  XNOR2_X1 U9106 ( .A(n7890), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14953) );
  OR2_X1 U9107 ( .A1(n14692), .A2(n14548), .ZN(n6712) );
  NAND2_X1 U9108 ( .A1(n9958), .A2(n9957), .ZN(n12602) );
  OR2_X1 U9109 ( .A1(n10024), .A2(n11534), .ZN(n6713) );
  NAND2_X1 U9110 ( .A1(n10213), .A2(n10036), .ZN(n11362) );
  XOR2_X1 U9111 ( .A(n11596), .B(P3_REG1_REG_4__SCAN_IN), .Z(n6714) );
  OR2_X1 U9112 ( .A1(n14789), .A2(n7269), .ZN(n6715) );
  OAI21_X1 U9113 ( .B1(n9064), .B2(n9063), .A(n13690), .ZN(n9102) );
  NAND2_X1 U9114 ( .A1(n9970), .A2(n9969), .ZN(n13378) );
  NAND4_X1 U9115 ( .A1(n9641), .A2(n9640), .A3(n9639), .A4(n9638), .ZN(n15614)
         );
  INV_X1 U9116 ( .A(n12094), .ZN(n15563) );
  AOI22_X1 U9117 ( .A1(n14237), .A2(n8484), .B1(n8483), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n14522) );
  INV_X1 U9118 ( .A(n14522), .ZN(n7262) );
  NAND2_X1 U9119 ( .A1(n7777), .A2(n7589), .ZN(n6716) );
  NAND2_X1 U9120 ( .A1(n8836), .A2(n8835), .ZN(n12749) );
  INV_X1 U9121 ( .A(n9602), .ZN(n10217) );
  AND2_X1 U9122 ( .A1(n7713), .A2(n6712), .ZN(n6717) );
  INV_X1 U9123 ( .A(n7519), .ZN(n7518) );
  NOR2_X1 U9124 ( .A1(n15468), .A2(n13790), .ZN(n7519) );
  NOR2_X1 U9125 ( .A1(n13764), .A2(n7453), .ZN(n6718) );
  AND2_X1 U9126 ( .A1(n7100), .A2(n6706), .ZN(n6719) );
  OR2_X1 U9127 ( .A1(n11997), .A2(n11996), .ZN(n6720) );
  NAND2_X1 U9128 ( .A1(n7499), .A2(n6758), .ZN(n7497) );
  NAND2_X1 U9129 ( .A1(n13405), .A2(n10181), .ZN(n9955) );
  INV_X1 U9130 ( .A(n14830), .ZN(n14610) );
  OR2_X1 U9131 ( .A1(n14679), .A2(n14576), .ZN(n6721) );
  AND2_X1 U9132 ( .A1(n12754), .A2(n12753), .ZN(n6722) );
  AND2_X1 U9133 ( .A1(n12791), .A2(n12790), .ZN(n6723) );
  NAND2_X1 U9134 ( .A1(n12939), .A2(n12938), .ZN(n6724) );
  AND2_X1 U9135 ( .A1(n12765), .A2(n12764), .ZN(n6725) );
  OR2_X1 U9136 ( .A1(n9131), .A2(n9335), .ZN(n6726) );
  AND2_X1 U9137 ( .A1(n7125), .A2(n7126), .ZN(n6727) );
  AND2_X2 U9138 ( .A1(n6887), .A2(n6873), .ZN(n9633) );
  XNOR2_X1 U9139 ( .A(n9193), .B(n9192), .ZN(n6728) );
  NAND2_X1 U9140 ( .A1(n6948), .A2(n9645), .ZN(n11366) );
  NAND2_X1 U9141 ( .A1(n11021), .A2(n12663), .ZN(n11415) );
  OR2_X1 U9142 ( .A1(n14837), .A2(n14582), .ZN(n6729) );
  NAND2_X1 U9143 ( .A1(n6912), .A2(n6991), .ZN(n13123) );
  NOR4_X1 U9144 ( .A1(n13976), .A2(n13985), .A3(n13998), .A4(n12923), .ZN(
        n6730) );
  INV_X1 U9145 ( .A(n8085), .ZN(n7835) );
  XNOR2_X1 U9146 ( .A(n7836), .B(SI_10_), .ZN(n8085) );
  NAND2_X1 U9147 ( .A1(n8369), .A2(n8368), .ZN(n14647) );
  INV_X1 U9148 ( .A(n14647), .ZN(n7266) );
  AND2_X1 U9149 ( .A1(n7608), .A2(n7611), .ZN(n6731) );
  NAND2_X1 U9150 ( .A1(n8851), .A2(n8850), .ZN(n12756) );
  OR2_X1 U9151 ( .A1(n13204), .A2(n13200), .ZN(n6732) );
  NAND2_X1 U9152 ( .A1(n9018), .A2(n9017), .ZN(n14170) );
  INV_X1 U9153 ( .A(n14180), .ZN(n14053) );
  INV_X1 U9154 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9335) );
  INV_X1 U9155 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14233) );
  NAND2_X1 U9156 ( .A1(n8344), .A2(n8343), .ZN(n14857) );
  INV_X1 U9157 ( .A(n14857), .ZN(n7267) );
  XOR2_X1 U9158 ( .A(n15040), .B(n12545), .Z(n6733) );
  NAND2_X1 U9159 ( .A1(n10465), .A2(n8552), .ZN(n10481) );
  INV_X1 U9160 ( .A(n14732), .ZN(n7726) );
  XNOR2_X1 U9161 ( .A(n13352), .B(n13359), .ZN(n13346) );
  NOR3_X1 U9162 ( .A1(n12684), .A2(n12683), .A3(n12682), .ZN(n6734) );
  AND2_X1 U9163 ( .A1(n12731), .A2(n11658), .ZN(n6735) );
  XNOR2_X1 U9164 ( .A(n14647), .B(n14579), .ZN(n14643) );
  INV_X1 U9165 ( .A(n13928), .ZN(n7418) );
  AND2_X1 U9166 ( .A1(n13940), .A2(n13941), .ZN(n6736) );
  NAND2_X1 U9167 ( .A1(n8863), .A2(n8862), .ZN(n6737) );
  INV_X1 U9168 ( .A(n8404), .ZN(n7556) );
  INV_X1 U9169 ( .A(n8371), .ZN(n7553) );
  OR2_X1 U9170 ( .A1(n13916), .A2(n13894), .ZN(n6738) );
  NAND2_X1 U9171 ( .A1(n14170), .A2(n13918), .ZN(n6739) );
  NAND2_X1 U9172 ( .A1(n12881), .A2(n12880), .ZN(n14140) );
  INV_X1 U9173 ( .A(n14140), .ZN(n7340) );
  OR2_X1 U9174 ( .A1(n14103), .A2(n14127), .ZN(n6740) );
  INV_X1 U9175 ( .A(n7600), .ZN(n7599) );
  OAI21_X1 U9176 ( .B1(n14350), .B2(n14351), .A(n10404), .ZN(n7600) );
  AND2_X1 U9177 ( .A1(n10343), .A2(n10342), .ZN(n6741) );
  AND3_X1 U9178 ( .A1(n10197), .A2(n6980), .A3(n13362), .ZN(n6742) );
  OR2_X1 U9179 ( .A1(n14195), .A2(n13913), .ZN(n6743) );
  AND4_X1 U9180 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .ZN(n11709)
         );
  AND2_X1 U9181 ( .A1(n6931), .A2(n6923), .ZN(n6744) );
  AND2_X1 U9182 ( .A1(n14543), .A2(n7722), .ZN(n6745) );
  AND2_X1 U9183 ( .A1(n14066), .A2(n13893), .ZN(n6746) );
  AND2_X1 U9184 ( .A1(n7376), .A2(n7379), .ZN(n6747) );
  INV_X1 U9185 ( .A(n14893), .ZN(n14751) );
  NAND2_X1 U9186 ( .A1(n8253), .A2(n8252), .ZN(n14893) );
  INV_X1 U9187 ( .A(n7350), .ZN(n14062) );
  NOR2_X1 U9188 ( .A1(n14078), .A2(n14185), .ZN(n7350) );
  AND2_X1 U9189 ( .A1(n10117), .A2(n10116), .ZN(n12165) );
  AND2_X1 U9190 ( .A1(n7437), .A2(n7435), .ZN(n6748) );
  OR2_X1 U9191 ( .A1(n14084), .A2(n14092), .ZN(n6749) );
  AND2_X1 U9192 ( .A1(n7413), .A2(n13928), .ZN(n6750) );
  NAND2_X1 U9193 ( .A1(n13492), .A2(n10157), .ZN(n6751) );
  NOR2_X1 U9194 ( .A1(n9679), .A2(n7668), .ZN(n9699) );
  NOR2_X1 U9195 ( .A1(n14406), .A2(n11203), .ZN(n6752) );
  OR2_X1 U9196 ( .A1(n7990), .A2(n7989), .ZN(n6753) );
  AND2_X1 U9197 ( .A1(n6683), .A2(n12777), .ZN(n6754) );
  OR2_X1 U9198 ( .A1(n7175), .A2(n7170), .ZN(n6755) );
  AND2_X1 U9199 ( .A1(n6721), .A2(n14655), .ZN(n6756) );
  AND2_X1 U9200 ( .A1(n13084), .A2(n6684), .ZN(n6757) );
  NAND2_X1 U9201 ( .A1(n14180), .A2(n7047), .ZN(n6758) );
  AND2_X1 U9202 ( .A1(n7744), .A2(n7782), .ZN(n6759) );
  INV_X1 U9203 ( .A(n14822), .ZN(n14594) );
  INV_X1 U9204 ( .A(n7419), .ZN(n7416) );
  NAND2_X1 U9205 ( .A1(n14149), .A2(n13942), .ZN(n7419) );
  NOR2_X1 U9206 ( .A1(n8403), .A2(n7556), .ZN(n6760) );
  NAND2_X1 U9207 ( .A1(n7718), .A2(n7717), .ZN(n6761) );
  NOR2_X1 U9208 ( .A1(n13430), .A2(n13087), .ZN(n6762) );
  AND2_X1 U9209 ( .A1(n13330), .A2(n10202), .ZN(n6763) );
  AND2_X1 U9210 ( .A1(n7523), .A2(n7524), .ZN(n6764) );
  OR2_X1 U9211 ( .A1(n12527), .A2(n7296), .ZN(n6765) );
  AND2_X1 U9212 ( .A1(n7304), .A2(n12534), .ZN(n6766) );
  AND2_X1 U9213 ( .A1(n8073), .A2(n8072), .ZN(n6767) );
  AND2_X1 U9214 ( .A1(n7836), .A2(SI_10_), .ZN(n6768) );
  NOR2_X1 U9215 ( .A1(n14905), .A2(n14564), .ZN(n6769) );
  NOR2_X1 U9216 ( .A1(n12993), .A2(n13372), .ZN(n6770) );
  NOR2_X1 U9217 ( .A1(n14180), .A2(n7047), .ZN(n6771) );
  INV_X1 U9218 ( .A(n7751), .ZN(n7379) );
  AND2_X1 U9219 ( .A1(n14685), .A2(n6712), .ZN(n6772) );
  AND2_X1 U9220 ( .A1(n7138), .A2(n7142), .ZN(n6773) );
  NOR2_X1 U9221 ( .A1(n15087), .A2(n14399), .ZN(n6774) );
  AND2_X1 U9222 ( .A1(n12824), .A2(n12823), .ZN(n6775) );
  AND2_X1 U9223 ( .A1(n12690), .A2(n12689), .ZN(n6776) );
  AND2_X1 U9224 ( .A1(n7826), .A2(SI_7_), .ZN(n6777) );
  INV_X1 U9225 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9588) );
  INV_X1 U9226 ( .A(n7611), .ZN(n7610) );
  AND2_X1 U9227 ( .A1(n13378), .A2(n13391), .ZN(n6778) );
  NAND2_X1 U9228 ( .A1(n7670), .A2(n9599), .ZN(n6779) );
  NOR2_X1 U9229 ( .A1(n9679), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9681) );
  INV_X1 U9230 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10540) );
  INV_X1 U9231 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10496) );
  INV_X1 U9232 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10558) );
  INV_X1 U9233 ( .A(n7290), .ZN(n7289) );
  NAND2_X1 U9234 ( .A1(n13429), .A2(n12529), .ZN(n7290) );
  AND2_X1 U9235 ( .A1(n8812), .A2(n8811), .ZN(n6780) );
  NAND2_X1 U9236 ( .A1(n10167), .A2(n13459), .ZN(n6781) );
  OR2_X1 U9237 ( .A1(n7520), .A2(n7519), .ZN(n6782) );
  INV_X1 U9238 ( .A(n7503), .ZN(n7502) );
  NAND2_X1 U9239 ( .A1(n14191), .A2(n14092), .ZN(n7503) );
  NAND2_X1 U9240 ( .A1(n14647), .A2(n14579), .ZN(n6783) );
  OR2_X1 U9241 ( .A1(n7418), .A2(n7415), .ZN(n6784) );
  NOR2_X1 U9242 ( .A1(n7267), .A2(n14577), .ZN(n6785) );
  AND2_X1 U9243 ( .A1(n13027), .A2(n13139), .ZN(n6786) );
  INV_X1 U9244 ( .A(n7482), .ZN(n13714) );
  INV_X1 U9245 ( .A(n7497), .ZN(n7496) );
  NOR2_X1 U9246 ( .A1(n12838), .A2(n7674), .ZN(n6787) );
  AND2_X1 U9247 ( .A1(n7689), .A2(n7688), .ZN(n6788) );
  INV_X1 U9248 ( .A(n12349), .ZN(n7360) );
  INV_X1 U9249 ( .A(n12805), .ZN(n7154) );
  AND2_X1 U9250 ( .A1(n9875), .A2(n7398), .ZN(n6789) );
  OAI21_X1 U9251 ( .B1(n8191), .B2(n7162), .A(n8230), .ZN(n7161) );
  OR2_X1 U9252 ( .A1(n7148), .A2(n6705), .ZN(n6790) );
  AND2_X1 U9253 ( .A1(n14165), .A2(n13920), .ZN(n6791) );
  OR2_X1 U9254 ( .A1(n11704), .A2(n7697), .ZN(n6792) );
  NAND2_X1 U9255 ( .A1(n7359), .A2(n12352), .ZN(n6793) );
  OR2_X1 U9256 ( .A1(n6704), .A2(n7610), .ZN(n6794) );
  INV_X1 U9257 ( .A(n13917), .ZN(n7493) );
  AND2_X1 U9258 ( .A1(n7073), .A2(n7072), .ZN(n6795) );
  AND3_X1 U9259 ( .A1(n10210), .A2(n10203), .A3(n10029), .ZN(n6796) );
  NAND2_X1 U9260 ( .A1(n8385), .A2(n8384), .ZN(n14843) );
  INV_X1 U9261 ( .A(n14843), .ZN(n7265) );
  OR2_X1 U9262 ( .A1(n10229), .A2(n11575), .ZN(n6797) );
  AND2_X1 U9263 ( .A1(n7541), .A2(n7540), .ZN(n6798) );
  OR2_X1 U9264 ( .A1(n12788), .A2(n12789), .ZN(n6799) );
  OR2_X1 U9265 ( .A1(n13921), .A2(n13920), .ZN(n6800) );
  AND3_X1 U9266 ( .A1(n7693), .A2(n8568), .A3(n8604), .ZN(n6801) );
  NOR2_X1 U9267 ( .A1(n14004), .A2(n7436), .ZN(n7435) );
  AND2_X1 U9268 ( .A1(n7342), .A2(n7340), .ZN(n6802) );
  OR2_X1 U9269 ( .A1(n15468), .A2(n12738), .ZN(n6803) );
  OR2_X1 U9270 ( .A1(n15457), .A2(n11658), .ZN(n6804) );
  NOR2_X1 U9271 ( .A1(n11268), .A2(n7461), .ZN(n6805) );
  NOR2_X1 U9272 ( .A1(n13330), .A2(n7312), .ZN(n7311) );
  XNOR2_X1 U9273 ( .A(n9202), .B(n9203), .ZN(n7273) );
  AND2_X1 U9274 ( .A1(n10124), .A2(n9763), .ZN(n6806) );
  AND2_X1 U9275 ( .A1(n9588), .A2(n7396), .ZN(n6807) );
  AND2_X1 U9276 ( .A1(n14572), .A2(n7748), .ZN(n6808) );
  AND2_X1 U9277 ( .A1(n14827), .A2(n14825), .ZN(n6809) );
  NAND2_X1 U9278 ( .A1(n12813), .A2(n12812), .ZN(n6810) );
  AND2_X1 U9279 ( .A1(n7156), .A2(n7155), .ZN(n6811) );
  NAND2_X1 U9280 ( .A1(n7116), .A2(n7114), .ZN(n6812) );
  AND2_X1 U9281 ( .A1(n8997), .A2(n8986), .ZN(n6813) );
  AND2_X1 U9282 ( .A1(n12187), .A2(n12185), .ZN(n6814) );
  OR2_X1 U9283 ( .A1(n8309), .A2(n8308), .ZN(n6815) );
  AND2_X1 U9284 ( .A1(n6696), .A2(n11516), .ZN(n6816) );
  OR2_X1 U9285 ( .A1(n7553), .A2(n8370), .ZN(n6817) );
  AND2_X1 U9286 ( .A1(n7743), .A2(n6759), .ZN(n6818) );
  INV_X1 U9287 ( .A(n11753), .ZN(n7102) );
  INV_X1 U9288 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9594) );
  INV_X1 U9289 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9599) );
  INV_X1 U9290 ( .A(n8193), .ZN(n7162) );
  AND2_X1 U9291 ( .A1(n7173), .A2(n6755), .ZN(n6819) );
  OR2_X1 U9292 ( .A1(n15036), .A2(n15029), .ZN(n10057) );
  INV_X1 U9293 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9587) );
  INV_X1 U9294 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8571) );
  INV_X1 U9295 ( .A(n7385), .ZN(n7384) );
  NAND2_X1 U9296 ( .A1(n14601), .A2(n6729), .ZN(n7385) );
  INV_X1 U9297 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6964) );
  INV_X1 U9298 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7026) );
  INV_X1 U9299 ( .A(n14149), .ZN(n7344) );
  INV_X1 U9300 ( .A(SI_2_), .ZN(n7242) );
  OAI21_X1 U9301 ( .B1(n9824), .B2(n7622), .A(n9837), .ZN(n7621) );
  AND2_X1 U9302 ( .A1(n12594), .A2(n13439), .ZN(n6820) );
  INV_X1 U9303 ( .A(n8585), .ZN(n8831) );
  NAND2_X1 U9304 ( .A1(n7449), .A2(n8955), .ZN(n13683) );
  NOR2_X1 U9305 ( .A1(n14785), .A2(n7753), .ZN(n6821) );
  XNOR2_X1 U9306 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9696) );
  INV_X1 U9307 ( .A(n9696), .ZN(n7218) );
  AND4_X1 U9308 ( .A1(n8064), .A2(n8063), .A3(n8062), .A4(n8061), .ZN(n12020)
         );
  INV_X1 U9309 ( .A(n7714), .ZN(n14716) );
  AOI22_X1 U9310 ( .A1(n14769), .A2(n6745), .B1(n14543), .B2(n7715), .ZN(n7714) );
  INV_X1 U9311 ( .A(n7092), .ZN(n7091) );
  INV_X1 U9312 ( .A(n7621), .ZN(n7620) );
  INV_X1 U9313 ( .A(n11596), .ZN(n11696) );
  AND2_X1 U9314 ( .A1(n12588), .A2(n12587), .ZN(n6822) );
  XOR2_X1 U9315 ( .A(n6711), .B(n7403), .Z(n6823) );
  OR2_X1 U9316 ( .A1(n8300), .A2(SI_20_), .ZN(n6824) );
  AND2_X1 U9317 ( .A1(n11016), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U9318 ( .A1(n7505), .A2(n7504), .ZN(n6826) );
  OR2_X1 U9319 ( .A1(n7855), .A2(SI_17_), .ZN(n6827) );
  INV_X1 U9320 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10721) );
  INV_X1 U9321 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7613) );
  INV_X1 U9322 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7016) );
  AND2_X1 U9323 ( .A1(n13037), .A2(n13038), .ZN(n6828) );
  OR2_X1 U9324 ( .A1(n8166), .A2(n7198), .ZN(n6829) );
  AND2_X1 U9325 ( .A1(n15103), .A2(n10336), .ZN(n6830) );
  INV_X1 U9326 ( .A(n15296), .ZN(n15300) );
  AND2_X1 U9327 ( .A1(n11568), .A2(n13268), .ZN(n15500) );
  NOR2_X1 U9328 ( .A1(n11522), .A2(n11705), .ZN(n7260) );
  INV_X1 U9329 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7203) );
  INV_X1 U9330 ( .A(n14905), .ZN(n7272) );
  AND2_X1 U9331 ( .A1(n15503), .A2(n13325), .ZN(n6831) );
  INV_X1 U9332 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7396) );
  INV_X1 U9333 ( .A(n13412), .ZN(n13390) );
  AND2_X1 U9334 ( .A1(n7090), .A2(n7089), .ZN(n6832) );
  NOR2_X1 U9335 ( .A1(n15679), .A2(n7012), .ZN(n6833) );
  INV_X1 U9336 ( .A(n7628), .ZN(n7232) );
  NAND2_X1 U9337 ( .A1(n12178), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7628) );
  INV_X1 U9338 ( .A(n7351), .ZN(n12317) );
  NOR2_X1 U9339 ( .A1(n12316), .A2(n12761), .ZN(n7351) );
  INV_X1 U9340 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12017) );
  INV_X1 U9341 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10960) );
  INV_X1 U9342 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9343 ( .A1(n8759), .A2(n8758), .ZN(n12717) );
  INV_X1 U9344 ( .A(n12717), .ZN(n7347) );
  INV_X1 U9345 ( .A(n12663), .ZN(n6951) );
  AND2_X1 U9346 ( .A1(n7328), .A2(n7327), .ZN(n6834) );
  INV_X1 U9347 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7635) );
  AND2_X1 U9348 ( .A1(n7099), .A2(n6719), .ZN(n6835) );
  NAND2_X1 U9349 ( .A1(n11374), .A2(n12614), .ZN(n13142) );
  NAND2_X1 U9350 ( .A1(n11413), .A2(n11410), .ZN(n11797) );
  INV_X1 U9351 ( .A(n11797), .ZN(n7346) );
  AND2_X1 U9352 ( .A1(n7252), .A2(n8482), .ZN(n6836) );
  AND2_X1 U9353 ( .A1(n13286), .A2(n13309), .ZN(n6837) );
  NAND2_X1 U9354 ( .A1(n12332), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7627) );
  INV_X1 U9355 ( .A(n7615), .ZN(n7239) );
  INV_X1 U9356 ( .A(n13321), .ZN(n6866) );
  AND2_X1 U9357 ( .A1(n6896), .A2(n7390), .ZN(n6838) );
  NAND2_X1 U9358 ( .A1(n9651), .A2(SI_31_), .ZN(n6839) );
  AND2_X1 U9359 ( .A1(n7627), .A2(n12209), .ZN(n6840) );
  AND2_X1 U9360 ( .A1(n11599), .A2(n11598), .ZN(n11765) );
  INV_X1 U9361 ( .A(n9585), .ZN(n7240) );
  INV_X1 U9362 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6938) );
  INV_X1 U9363 ( .A(n9586), .ZN(n7241) );
  AND2_X1 U9364 ( .A1(n14944), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9586) );
  INV_X1 U9365 ( .A(n11997), .ZN(n7338) );
  INV_X1 U9366 ( .A(n13286), .ZN(n7327) );
  INV_X1 U9367 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7771) );
  XNOR2_X1 U9368 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(n9211), .ZN(n6841) );
  INV_X1 U9369 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14426) );
  INV_X1 U9370 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7215) );
  INV_X1 U9371 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6927) );
  INV_X1 U9372 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7157) );
  XNOR2_X1 U9373 ( .A(n13189), .B(n13190), .ZN(n12258) );
  NAND2_X1 U9374 ( .A1(n8584), .A2(n6844), .ZN(n8603) );
  XNOR2_X2 U9376 ( .A(n6845), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8597) );
  NAND3_X1 U9377 ( .A1(n7487), .A2(n7486), .A3(n11792), .ZN(n11790) );
  NAND3_X1 U9378 ( .A1(n7417), .A2(n14142), .A3(n14141), .ZN(n14219) );
  OR2_X1 U9379 ( .A1(n6851), .A2(n13948), .ZN(n6848) );
  OAI21_X1 U9380 ( .B1(n13946), .B2(n13945), .A(n13944), .ZN(n6851) );
  NAND3_X1 U9381 ( .A1(n8728), .A2(n6852), .A3(n8729), .ZN(n13795) );
  NAND3_X1 U9382 ( .A1(n7040), .A2(n7320), .A3(n6868), .ZN(P3_U3201) );
  AND2_X2 U9383 ( .A1(n6869), .A2(n6732), .ZN(n13202) );
  NOR2_X2 U9384 ( .A1(n11931), .A2(n11860), .ZN(n11930) );
  XNOR2_X2 U9385 ( .A(n11848), .B(n11861), .ZN(n11931) );
  XNOR2_X2 U9386 ( .A(n6872), .B(n13288), .ZN(n13263) );
  NAND2_X2 U9387 ( .A1(n13262), .A2(n13261), .ZN(n6872) );
  OR2_X2 U9388 ( .A1(n13254), .A2(n13253), .ZN(n13262) );
  NOR2_X1 U9389 ( .A1(n15013), .A2(n13249), .ZN(n13254) );
  AND3_X1 U9390 ( .A1(n6917), .A2(n6918), .A3(n6873), .ZN(n6883) );
  NAND2_X1 U9391 ( .A1(n7525), .A2(n6874), .ZN(n11600) );
  OAI211_X2 U9392 ( .C1(n9633), .C2(n7566), .A(n7565), .B(n9664), .ZN(n7564)
         );
  NAND2_X1 U9393 ( .A1(n13002), .A2(n13001), .ZN(n13000) );
  INV_X2 U9394 ( .A(n11394), .ZN(n13030) );
  INV_X1 U9395 ( .A(n12621), .ZN(n11483) );
  NAND2_X1 U9396 ( .A1(n11362), .A2(n13325), .ZN(n6876) );
  AND4_X2 U9397 ( .A1(n6884), .A2(n6916), .A3(n6883), .A4(n6882), .ZN(n9800)
         );
  OAI21_X2 U9398 ( .B1(n6890), .B2(n6894), .A(n7393), .ZN(n12979) );
  AND2_X1 U9399 ( .A1(n7390), .A2(n12069), .ZN(n6895) );
  NAND3_X1 U9400 ( .A1(n7392), .A2(n12111), .A3(n12089), .ZN(n6896) );
  XNOR2_X1 U9401 ( .A(n6905), .B(n13133), .ZN(n13143) );
  INV_X1 U9402 ( .A(n10038), .ZN(n10037) );
  INV_X2 U9403 ( .A(n6911), .ZN(n10223) );
  NAND2_X1 U9404 ( .A1(n6913), .A2(n12572), .ZN(n13094) );
  NAND2_X1 U9405 ( .A1(n6914), .A2(n13093), .ZN(n13002) );
  NAND2_X1 U9406 ( .A1(n12186), .A2(n6814), .ZN(n12246) );
  NAND2_X1 U9407 ( .A1(n11397), .A2(n11398), .ZN(n12044) );
  XNOR2_X1 U9408 ( .A(n11394), .B(n11393), .ZN(n12042) );
  OAI211_X1 U9409 ( .C1(n6838), .C2(n12069), .A(n12068), .B(n15494), .ZN(
        n12075) );
  XNOR2_X1 U9410 ( .A(n9189), .B(n9190), .ZN(n15702) );
  NAND3_X1 U9411 ( .A1(n6930), .A2(n9205), .A3(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n6929) );
  NAND2_X1 U9412 ( .A1(n14970), .A2(n6934), .ZN(n6933) );
  NAND2_X1 U9413 ( .A1(n14974), .A2(n6938), .ZN(n6934) );
  INV_X1 U9414 ( .A(n14974), .ZN(n6936) );
  NOR2_X1 U9415 ( .A1(n14975), .A2(n14974), .ZN(n14973) );
  NAND2_X1 U9416 ( .A1(n6975), .A2(n6974), .ZN(n7019) );
  NOR2_X2 U9417 ( .A1(n14972), .A2(n14971), .ZN(n14970) );
  XNOR2_X1 U9418 ( .A(n9177), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15695) );
  XNOR2_X1 U9419 ( .A(n6941), .B(n7282), .ZN(SUB_1596_U4) );
  NAND2_X1 U9420 ( .A1(n11371), .A2(n6950), .ZN(n11396) );
  NAND2_X1 U9421 ( .A1(n10037), .A2(n10032), .ZN(n10040) );
  NAND2_X4 U9422 ( .A1(n13320), .A2(n12561), .ZN(n10229) );
  NAND2_X1 U9423 ( .A1(n12078), .A2(n12059), .ZN(n12061) );
  NAND2_X1 U9424 ( .A1(n12068), .A2(n12056), .ZN(n12080) );
  NAND2_X1 U9425 ( .A1(n12989), .A2(n12988), .ZN(n13060) );
  NAND2_X1 U9426 ( .A1(n12080), .A2(n12079), .ZN(n12078) );
  NAND2_X1 U9427 ( .A1(n9687), .A2(n10095), .ZN(n15557) );
  OAI21_X1 U9428 ( .B1(n13444), .B2(n13437), .A(n9923), .ZN(n13428) );
  NAND2_X1 U9429 ( .A1(n14088), .A2(n6984), .ZN(n14073) );
  NAND2_X1 U9430 ( .A1(n13984), .A2(n13899), .ZN(n13975) );
  NAND2_X1 U9431 ( .A1(n14034), .A2(n7493), .ZN(n14033) );
  NAND2_X1 U9432 ( .A1(n6944), .A2(n11403), .ZN(n11455) );
  NAND2_X1 U9433 ( .A1(n11457), .A2(n11456), .ZN(n11789) );
  AOI21_X1 U9434 ( .B1(n14111), .B2(n14110), .A(n13890), .ZN(n14089) );
  AOI21_X1 U9435 ( .B1(n7665), .B2(n10064), .A(n7664), .ZN(n12549) );
  NAND2_X1 U9436 ( .A1(n10006), .A2(n10063), .ZN(n13329) );
  NAND2_X1 U9437 ( .A1(n9670), .A2(n10087), .ZN(n15572) );
  AOI21_X1 U9438 ( .B1(n7663), .B2(n6796), .A(n7661), .ZN(n10030) );
  NAND2_X1 U9439 ( .A1(n6946), .A2(n10100), .ZN(n11719) );
  NAND2_X1 U9440 ( .A1(n7422), .A2(n7420), .ZN(n14034) );
  NAND2_X1 U9441 ( .A1(n11402), .A2(n7445), .ZN(n6944) );
  NAND2_X1 U9442 ( .A1(n13361), .A2(n10068), .ZN(n6945) );
  NAND2_X1 U9443 ( .A1(n15557), .A2(n15561), .ZN(n6946) );
  OR2_X1 U9444 ( .A1(n13542), .A2(n15675), .ZN(n7319) );
  AND3_X2 U9445 ( .A1(n8567), .A2(n8566), .A3(n8667), .ZN(n8585) );
  NAND2_X1 U9446 ( .A1(n9944), .A2(n10070), .ZN(n13405) );
  OAI21_X1 U9447 ( .B1(n13509), .B2(n7654), .A(n7652), .ZN(n9912) );
  NAND2_X1 U9448 ( .A1(n14304), .A2(n10432), .ZN(n14369) );
  NAND2_X1 U9449 ( .A1(n10277), .A2(n10276), .ZN(n11061) );
  OAI21_X1 U9450 ( .B1(n11471), .B2(n11472), .A(n10311), .ZN(n10317) );
  NAND2_X1 U9451 ( .A1(n7873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U9452 ( .A1(n8548), .A2(n6818), .ZN(n7873) );
  NAND2_X1 U9453 ( .A1(n10791), .A2(n10792), .ZN(n10253) );
  XNOR2_X1 U9454 ( .A(n10249), .B(n10250), .ZN(n10792) );
  NAND2_X1 U9455 ( .A1(n10883), .A2(n10882), .ZN(n7573) );
  OR2_X1 U9456 ( .A1(n12857), .A2(n10499), .ZN(n8631) );
  INV_X1 U9457 ( .A(n12654), .ZN(n14213) );
  NAND2_X1 U9458 ( .A1(n11367), .A2(n11368), .ZN(n6950) );
  NAND2_X1 U9459 ( .A1(n13112), .A2(n13111), .ZN(n13110) );
  OAI21_X1 U9460 ( .B1(n12284), .B2(n12283), .A(n12282), .ZN(n12315) );
  AND2_X2 U9461 ( .A1(n12538), .A2(n12537), .ZN(n12540) );
  NAND3_X2 U9462 ( .A1(n8660), .A2(n8659), .A3(n6952), .ZN(n13799) );
  AND2_X1 U9463 ( .A1(n8657), .A2(n8658), .ZN(n6952) );
  AND2_X2 U9464 ( .A1(n15526), .A2(n11850), .ZN(n11996) );
  NOR2_X2 U9465 ( .A1(n15008), .A2(n13227), .ZN(n13231) );
  NAND2_X1 U9466 ( .A1(n7046), .A2(n7045), .ZN(n12269) );
  NOR2_X1 U9467 ( .A1(n11928), .A2(n11929), .ZN(n11927) );
  NOR2_X1 U9468 ( .A1(n11595), .A2(n15570), .ZN(n11759) );
  OAI21_X1 U9469 ( .B1(n13287), .B2(n7324), .A(n7079), .ZN(n7041) );
  INV_X1 U9470 ( .A(n15514), .ZN(n6954) );
  NAND2_X1 U9471 ( .A1(n13164), .A2(n11561), .ZN(n11739) );
  NOR2_X1 U9472 ( .A1(n6955), .A2(n13284), .ZN(n13279) );
  AOI21_X2 U9473 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n11696), .A(n11679), .ZN(
        n11594) );
  INV_X1 U9474 ( .A(n12975), .ZN(n9612) );
  NAND2_X1 U9475 ( .A1(n6956), .A2(n9654), .ZN(n11364) );
  OR2_X1 U9476 ( .A1(n10220), .A2(n7000), .ZN(n6999) );
  OAI21_X1 U9477 ( .B1(n11344), .B2(P3_D_REG_0__SCAN_IN), .A(n11332), .ZN(
        n7033) );
  AOI21_X1 U9478 ( .B1(n12945), .B2(n12951), .A(n6959), .ZN(n12953) );
  INV_X4 U9479 ( .A(n10501), .ZN(n10502) );
  NAND2_X1 U9480 ( .A1(n7539), .A2(n7537), .ZN(n8143) );
  NAND2_X1 U9481 ( .A1(n6961), .A2(n7818), .ZN(n7982) );
  NAND3_X1 U9482 ( .A1(n7816), .A2(n7020), .A3(n7002), .ZN(n6961) );
  NAND2_X1 U9483 ( .A1(n10227), .A2(n7034), .ZN(n12233) );
  NAND2_X1 U9484 ( .A1(n8129), .A2(n7064), .ZN(n7059) );
  OAI21_X2 U9485 ( .B1(n11937), .B2(n7477), .A(n7474), .ZN(n8890) );
  NAND2_X1 U9486 ( .A1(n6999), .A2(n6998), .ZN(n10218) );
  NAND2_X1 U9487 ( .A1(n11396), .A2(n11395), .ZN(n11397) );
  NAND2_X1 U9488 ( .A1(n9610), .A2(n13664), .ZN(n12641) );
  NAND2_X1 U9489 ( .A1(n7812), .A2(n7532), .ZN(n7020) );
  NAND2_X1 U9490 ( .A1(n8362), .A2(n8361), .ZN(n7244) );
  INV_X1 U9491 ( .A(n8437), .ZN(n7255) );
  NAND2_X1 U9492 ( .A1(n8480), .A2(n8456), .ZN(n12858) );
  NAND2_X1 U9493 ( .A1(n7672), .A2(n12953), .ZN(n12964) );
  INV_X1 U9494 ( .A(n12950), .ZN(n12951) );
  NAND2_X1 U9495 ( .A1(n7009), .A2(n7008), .ZN(n7278) );
  NAND2_X1 U9496 ( .A1(n15155), .A2(n15156), .ZN(n15152) );
  OR2_X1 U9497 ( .A1(n8662), .A2(n8661), .ZN(n8664) );
  OAI21_X2 U9498 ( .B1(n11020), .B2(n11019), .A(n8676), .ZN(n10987) );
  AOI22_X2 U9499 ( .A1(n8666), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n10747), .B2(
        n10775), .ZN(n8652) );
  OAI21_X2 U9500 ( .B1(n11009), .B2(n11008), .A(n8734), .ZN(n11039) );
  INV_X1 U9501 ( .A(n8615), .ZN(n8864) );
  NAND2_X1 U9502 ( .A1(n8697), .A2(n8696), .ZN(n10984) );
  NOR2_X1 U9503 ( .A1(n13714), .A2(n9048), .ZN(n13776) );
  NAND2_X1 U9504 ( .A1(n7457), .A2(n6805), .ZN(n7456) );
  NAND2_X1 U9505 ( .A1(n10992), .A2(n8664), .ZN(n11020) );
  INV_X1 U9506 ( .A(n7033), .ZN(n13661) );
  OAI21_X1 U9508 ( .B1(n8637), .B2(n8638), .A(n8645), .ZN(n10898) );
  NOR2_X1 U9509 ( .A1(n12288), .A2(n7514), .ZN(n7513) );
  INV_X1 U9510 ( .A(n7302), .ZN(n7301) );
  NAND2_X1 U9511 ( .A1(n13343), .A2(n12541), .ZN(n13331) );
  NAND2_X1 U9512 ( .A1(n9872), .A2(n9870), .ZN(n7017) );
  NAND2_X1 U9513 ( .A1(n9554), .A2(n9553), .ZN(n9697) );
  OAI22_X1 U9514 ( .A1(n12493), .A2(n12492), .B1(n12496), .B2(n12771), .ZN(
        n13911) );
  OR2_X1 U9515 ( .A1(n8035), .A2(n8034), .ZN(n8036) );
  NAND2_X1 U9516 ( .A1(n7163), .A2(n7167), .ZN(n8074) );
  OAI21_X1 U9517 ( .B1(n8260), .B2(n14568), .A(n8259), .ZN(n8276) );
  OAI22_X1 U9518 ( .A1(n7176), .A2(n6767), .B1(n8095), .B2(n7178), .ZN(n8152)
         );
  OAI21_X1 U9519 ( .B1(n6674), .B2(n6819), .A(n7171), .ZN(n7554) );
  OR3_X1 U9520 ( .A1(n8192), .A2(n7757), .A3(n7159), .ZN(n7158) );
  AOI21_X1 U9521 ( .B1(n8445), .B2(n7185), .A(n7182), .ZN(n8536) );
  INV_X1 U9522 ( .A(n8263), .ZN(n6966) );
  NAND2_X1 U9523 ( .A1(n14384), .A2(n14382), .ZN(n14379) );
  INV_X2 U9524 ( .A(n10296), .ZN(n10288) );
  NAND2_X1 U9525 ( .A1(n6968), .A2(n7179), .ZN(n7569) );
  NAND3_X1 U9526 ( .A1(n8291), .A2(n8290), .A3(n6815), .ZN(n6968) );
  NAND2_X2 U9527 ( .A1(n14294), .A2(n14293), .ZN(n14352) );
  NAND2_X1 U9528 ( .A1(n14379), .A2(n14380), .ZN(n14378) );
  NAND2_X1 U9529 ( .A1(n10362), .A2(n10363), .ZN(n14384) );
  NAND2_X1 U9530 ( .A1(n7604), .A2(n7602), .ZN(n14359) );
  INV_X1 U9531 ( .A(n7991), .ZN(n6971) );
  NAND2_X1 U9532 ( .A1(n6971), .A2(n6753), .ZN(n8010) );
  NAND2_X1 U9533 ( .A1(n12392), .A2(n10351), .ZN(n14268) );
  NAND2_X1 U9534 ( .A1(n11363), .A2(n15595), .ZN(n11395) );
  NAND2_X1 U9535 ( .A1(n11151), .A2(n8500), .ZN(n15200) );
  NAND2_X1 U9536 ( .A1(n7378), .A2(n7377), .ZN(n14642) );
  NAND2_X1 U9537 ( .A1(n11150), .A2(n11149), .ZN(n11199) );
  NAND2_X1 U9538 ( .A1(n14727), .A2(n14726), .ZN(n14725) );
  NAND2_X1 U9539 ( .A1(n14826), .A2(n6809), .ZN(n14927) );
  NAND2_X1 U9540 ( .A1(n7364), .A2(n7362), .ZN(n14731) );
  NAND2_X1 U9541 ( .A1(n7354), .A2(n7353), .ZN(n12402) );
  INV_X1 U9542 ( .A(n7388), .ZN(n11201) );
  NAND2_X1 U9543 ( .A1(n8466), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7916) );
  AND2_X4 U9544 ( .A1(n7789), .A2(n7788), .ZN(n8466) );
  NAND2_X1 U9545 ( .A1(n14266), .A2(n10358), .ZN(n10362) );
  NAND2_X1 U9546 ( .A1(n7936), .A2(n7813), .ZN(n7533) );
  NAND2_X1 U9547 ( .A1(n7533), .A2(n7815), .ZN(n7963) );
  XNOR2_X1 U9548 ( .A(n7036), .B(n9180), .ZN(n15699) );
  INV_X1 U9549 ( .A(n15145), .ZN(n6975) );
  OAI21_X2 U9550 ( .B1(n10510), .B2(n8457), .A(n6977), .ZN(n6976) );
  AND2_X1 U9551 ( .A1(n7939), .A2(n7938), .ZN(n6977) );
  NAND2_X1 U9552 ( .A1(n7812), .A2(n7811), .ZN(n7936) );
  NAND2_X1 U9553 ( .A1(n6978), .A2(n10210), .ZN(n10212) );
  NAND3_X1 U9554 ( .A1(n7631), .A2(n7634), .A3(n10057), .ZN(n6978) );
  NAND2_X1 U9555 ( .A1(n9573), .A2(n9572), .ZN(n9872) );
  NAND2_X1 U9556 ( .A1(n7205), .A2(n9579), .ZN(n9926) );
  NAND2_X1 U9557 ( .A1(n9575), .A2(n9574), .ZN(n9900) );
  NAND2_X1 U9558 ( .A1(n7637), .A2(n10216), .ZN(n10234) );
  NAND2_X1 U9559 ( .A1(n7626), .A2(n9582), .ZN(n9968) );
  NAND2_X1 U9560 ( .A1(n7212), .A2(n7211), .ZN(n9855) );
  NAND2_X1 U9561 ( .A1(n6981), .A2(n6742), .ZN(n10198) );
  NAND2_X1 U9562 ( .A1(n10192), .A2(n13376), .ZN(n6980) );
  NAND3_X1 U9563 ( .A1(n6983), .A2(n10205), .A3(n6733), .ZN(n6982) );
  NOR2_X1 U9564 ( .A1(n12270), .A2(n12463), .ZN(n13174) );
  NOR2_X2 U9565 ( .A1(n13205), .A2(n13206), .ZN(n13225) );
  NOR2_X2 U9566 ( .A1(n13176), .A2(n13177), .ZN(n13205) );
  AOI21_X2 U9567 ( .B1(n11677), .B2(n11675), .A(n11676), .ZN(n11679) );
  XNOR2_X1 U9568 ( .A(n13287), .B(n7327), .ZN(n13307) );
  NAND2_X1 U9569 ( .A1(n8606), .A2(n8607), .ZN(n7011) );
  OR2_X1 U9570 ( .A1(n12885), .A2(n8654), .ZN(n8659) );
  NAND2_X1 U9571 ( .A1(n7066), .A2(n7065), .ZN(n13981) );
  AND2_X1 U9572 ( .A1(n10264), .A2(n10260), .ZN(n7572) );
  NAND2_X1 U9573 ( .A1(n13375), .A2(n10195), .ZN(n13361) );
  NAND2_X1 U9574 ( .A1(n9852), .A2(n10150), .ZN(n13509) );
  INV_X1 U9575 ( .A(n7641), .ZN(n7646) );
  AND2_X4 U9576 ( .A1(n10229), .A2(n10501), .ZN(n9651) );
  INV_X1 U9577 ( .A(n11533), .ZN(n13320) );
  INV_X1 U9578 ( .A(n14268), .ZN(n6993) );
  NAND2_X1 U9579 ( .A1(n9103), .A2(n9102), .ZN(n9101) );
  INV_X1 U9580 ( .A(n10987), .ZN(n8697) );
  OAI211_X1 U9581 ( .C1(P2_IR_REG_21__SCAN_IN), .C2(P2_IR_REG_31__SCAN_IN), 
        .A(n6989), .B(n9065), .ZN(n8611) );
  AOI21_X2 U9582 ( .B1(n11039), .B2(n11038), .A(n8753), .ZN(n11106) );
  INV_X1 U9583 ( .A(n10481), .ZN(n7586) );
  NAND2_X1 U9584 ( .A1(n13605), .A2(n15679), .ZN(n7013) );
  NAND2_X1 U9585 ( .A1(n9656), .A2(n10086), .ZN(n11478) );
  OR2_X2 U9586 ( .A1(n15524), .A2(n15523), .ZN(n15526) );
  NOR2_X1 U9587 ( .A1(n11930), .A2(n11849), .ZN(n15524) );
  NAND2_X1 U9588 ( .A1(n7319), .A2(n13541), .ZN(n13605) );
  NAND2_X1 U9589 ( .A1(n7644), .A2(n7642), .ZN(n12213) );
  NAND2_X1 U9590 ( .A1(n9809), .A2(n10132), .ZN(n13527) );
  INV_X1 U9591 ( .A(n12486), .ZN(n9835) );
  NAND4_X2 U9592 ( .A1(n6713), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n15491)
         );
  NAND2_X1 U9593 ( .A1(n12061), .A2(n12060), .ZN(n12186) );
  OAI21_X1 U9594 ( .B1(n11465), .B2(n7443), .A(n7441), .ZN(n11644) );
  NAND2_X1 U9595 ( .A1(n7429), .A2(n6803), .ZN(n12123) );
  OAI22_X2 U9596 ( .A1(n13975), .A2(n13901), .B1(n13900), .B2(n13974), .ZN(
        n13951) );
  NAND2_X1 U9597 ( .A1(n7255), .A2(n7254), .ZN(n8439) );
  INV_X1 U9598 ( .A(n12123), .ZN(n12126) );
  NAND2_X1 U9599 ( .A1(n8336), .A2(n8335), .ZN(n8342) );
  NAND2_X1 U9600 ( .A1(n11889), .A2(n7430), .ZN(n7429) );
  NAND2_X1 U9601 ( .A1(n12924), .A2(n7022), .ZN(n7021) );
  AOI22_X2 U9602 ( .A1(n12315), .A2(n12917), .B1(n12761), .B2(n13788), .ZN(
        n12498) );
  OAI21_X2 U9603 ( .B1(n12899), .B2(n11610), .A(n10978), .ZN(n11402) );
  NOR2_X2 U9604 ( .A1(n11980), .A2(n11981), .ZN(n11986) );
  NAND2_X1 U9605 ( .A1(n7028), .A2(n7027), .ZN(n11595) );
  NAND2_X4 U9606 ( .A1(n8867), .A2(n8866), .ZN(n12761) );
  NAND2_X2 U9607 ( .A1(n13774), .A2(n7003), .ZN(n9103) );
  NAND2_X2 U9608 ( .A1(n13737), .A2(n7483), .ZN(n7482) );
  INV_X1 U9609 ( .A(n7478), .ZN(n7477) );
  NAND2_X1 U9610 ( .A1(n7528), .A2(n7527), .ZN(n8047) );
  NAND2_X1 U9611 ( .A1(n15145), .A2(n15146), .ZN(n9198) );
  INV_X1 U9612 ( .A(n9181), .ZN(n7036) );
  INV_X1 U9613 ( .A(n7044), .ZN(n7283) );
  XNOR2_X1 U9614 ( .A(n14958), .B(n7010), .ZN(SUB_1596_U62) );
  AOI21_X2 U9615 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14494), .A(n14493), .ZN(
        n14503) );
  XNOR2_X2 U9616 ( .A(n9392), .B(n7937), .ZN(n14446) );
  NAND2_X1 U9617 ( .A1(n11369), .A2(n10080), .ZN(n11368) );
  AND2_X1 U9618 ( .A1(n11395), .A2(n11365), .ZN(n11371) );
  NAND2_X1 U9619 ( .A1(n15389), .A2(n12654), .ZN(n10969) );
  AND3_X2 U9620 ( .A1(n6764), .A2(n8635), .A3(n8636), .ZN(n15389) );
  AND2_X4 U9621 ( .A1(n10229), .A2(n10502), .ZN(n9805) );
  NAND3_X1 U9622 ( .A1(n14241), .A2(n12606), .A3(P2_REG0_REG_1__SCAN_IN), .ZN(
        n7523) );
  NAND2_X1 U9623 ( .A1(n15577), .A2(n15576), .ZN(n15575) );
  NAND2_X1 U9624 ( .A1(n15595), .A2(n11364), .ZN(n10078) );
  AND2_X4 U9625 ( .A1(n12975), .A2(n12641), .ZN(n9847) );
  NAND2_X1 U9626 ( .A1(n11497), .A2(n11496), .ZN(n11501) );
  OAI21_X2 U9627 ( .B1(n12533), .B2(n7301), .A(n7300), .ZN(n13358) );
  NAND2_X1 U9628 ( .A1(n7292), .A2(n7291), .ZN(n13457) );
  AOI21_X1 U9629 ( .B1(n7309), .B2(n7311), .A(n7308), .ZN(n12542) );
  OAI21_X1 U9630 ( .B1(n13039), .B2(n13142), .A(n6828), .ZN(P3_U3160) );
  NAND2_X1 U9631 ( .A1(n10284), .A2(n10283), .ZN(n11112) );
  NAND2_X1 U9632 ( .A1(n7777), .A2(n7776), .ZN(n7879) );
  INV_X1 U9633 ( .A(n7879), .ZN(n7882) );
  AOI22_X1 U9634 ( .A1(n14410), .A2(n10417), .B1(n15216), .B2(n10288), .ZN(
        n10250) );
  NOR2_X1 U9635 ( .A1(n14672), .A2(n6772), .ZN(n7712) );
  OAI21_X2 U9636 ( .B1(n8298), .B2(n7256), .A(n7867), .ZN(n8336) );
  INV_X1 U9637 ( .A(n13387), .ZN(n7651) );
  NAND2_X1 U9638 ( .A1(n9913), .A2(n11886), .ZN(n7205) );
  NAND2_X1 U9639 ( .A1(n9926), .A2(n9924), .ZN(n7204) );
  NAND2_X1 U9640 ( .A1(n9900), .A2(n9899), .ZN(n7636) );
  NAND2_X1 U9641 ( .A1(n9566), .A2(n9565), .ZN(n9788) );
  NAND2_X1 U9642 ( .A1(n7201), .A2(n9567), .ZN(n9804) );
  NOR2_X1 U9643 ( .A1(n11927), .A2(n11856), .ZN(n15514) );
  NOR2_X2 U9644 ( .A1(n15009), .A2(n15010), .ZN(n15008) );
  XNOR2_X1 U9645 ( .A(n11855), .B(n11861), .ZN(n11928) );
  NAND3_X2 U9646 ( .A1(n8631), .A2(n8632), .A3(n8633), .ZN(n12654) );
  NAND2_X1 U9647 ( .A1(n7456), .A2(n7454), .ZN(n11620) );
  NAND2_X1 U9648 ( .A1(n9101), .A2(n9100), .ZN(n9129) );
  NAND2_X1 U9649 ( .A1(n9198), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7018) );
  NAND2_X1 U9650 ( .A1(n15162), .A2(n15163), .ZN(n7277) );
  NOR2_X1 U9651 ( .A1(n9179), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U9652 ( .A1(n12941), .A2(n7673), .ZN(n7672) );
  NOR2_X1 U9653 ( .A1(n9200), .A2(n9199), .ZN(n9150) );
  NOR2_X1 U9654 ( .A1(n9193), .A2(n9192), .ZN(n9142) );
  NOR2_X1 U9655 ( .A1(n9184), .A2(n9183), .ZN(n9136) );
  NAND2_X1 U9656 ( .A1(n11594), .A2(n11606), .ZN(n7027) );
  INV_X1 U9657 ( .A(n11760), .ZN(n7028) );
  INV_X1 U9658 ( .A(n7041), .ZN(n7040) );
  INV_X1 U9659 ( .A(n13329), .ZN(n7665) );
  INV_X4 U9660 ( .A(n13693), .ZN(n9007) );
  INV_X1 U9661 ( .A(n10986), .ZN(n8696) );
  NOR2_X1 U9662 ( .A1(n15695), .A2(n15696), .ZN(n15694) );
  NAND2_X1 U9663 ( .A1(n7277), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U9664 ( .A1(n11657), .A2(n6804), .ZN(n11889) );
  NAND2_X1 U9665 ( .A1(n13888), .A2(n7754), .ZN(n14111) );
  NAND2_X1 U9666 ( .A1(n11789), .A2(n12903), .ZN(n7440) );
  NOR2_X2 U9667 ( .A1(n13263), .A2(n13595), .ZN(n13300) );
  INV_X1 U9668 ( .A(n11599), .ZN(n7043) );
  NAND2_X2 U9669 ( .A1(n13265), .A2(n13264), .ZN(n7042) );
  NOR2_X2 U9670 ( .A1(n13285), .A2(n13284), .ZN(n13287) );
  NOR2_X1 U9671 ( .A1(n15014), .A2(n15015), .ZN(n15013) );
  XNOR2_X1 U9672 ( .A(n13247), .B(n13248), .ZN(n15014) );
  NAND2_X2 U9673 ( .A1(n9650), .A2(n7333), .ZN(n11569) );
  OAI21_X1 U9674 ( .B1(n11579), .B2(n7548), .A(n7547), .ZN(n11684) );
  NAND2_X1 U9675 ( .A1(n15699), .A2(n15698), .ZN(n15697) );
  AND2_X2 U9676 ( .A1(n12269), .A2(n12268), .ZN(n13173) );
  INV_X1 U9677 ( .A(n11986), .ZN(n7046) );
  OAI21_X1 U9678 ( .B1(n13307), .B2(n15515), .A(n7560), .ZN(P3_U3200) );
  NAND3_X1 U9679 ( .A1(n7072), .A2(n7069), .A3(n7073), .ZN(n7066) );
  NAND3_X1 U9680 ( .A1(n7072), .A2(n7073), .A3(n13919), .ZN(n7067) );
  NAND2_X1 U9681 ( .A1(n7071), .A2(n13917), .ZN(n7073) );
  INV_X1 U9682 ( .A(n7494), .ZN(n7071) );
  INV_X1 U9683 ( .A(n11872), .ZN(n7085) );
  AOI21_X1 U9684 ( .B1(n7085), .B2(n7089), .A(n7086), .ZN(n12261) );
  NAND2_X1 U9685 ( .A1(n11872), .A2(n11871), .ZN(n11990) );
  NOR2_X1 U9686 ( .A1(n11991), .A2(n11989), .ZN(n7092) );
  INV_X1 U9687 ( .A(n11871), .ZN(n7094) );
  NAND2_X1 U9688 ( .A1(n11550), .A2(n7095), .ZN(n7098) );
  INV_X1 U9689 ( .A(n11689), .ZN(n7104) );
  NAND3_X1 U9690 ( .A1(n7108), .A2(n12666), .A3(n7107), .ZN(n7109) );
  NAND2_X1 U9691 ( .A1(n12658), .A2(n12659), .ZN(n7107) );
  OAI21_X1 U9692 ( .B1(n12658), .B2(n12659), .A(n12660), .ZN(n7108) );
  AOI21_X1 U9693 ( .B1(n12677), .B2(n12676), .A(n12675), .ZN(n12684) );
  NAND2_X1 U9694 ( .A1(n7109), .A2(n12671), .ZN(n12677) );
  NAND2_X1 U9695 ( .A1(n12768), .A2(n7112), .ZN(n7110) );
  NAND2_X1 U9696 ( .A1(n12728), .A2(n7122), .ZN(n7121) );
  INV_X1 U9697 ( .A(n12727), .ZN(n7129) );
  INV_X1 U9698 ( .A(n12732), .ZN(n7130) );
  OAI21_X1 U9699 ( .B1(n6776), .B2(n12693), .A(n12694), .ZN(n7133) );
  INV_X1 U9700 ( .A(n12834), .ZN(n7135) );
  NAND2_X1 U9701 ( .A1(n12758), .A2(n7142), .ZN(n7141) );
  NAND4_X1 U9702 ( .A1(n12784), .A2(n12783), .A3(n6799), .A4(n7147), .ZN(n7146) );
  NAND2_X1 U9703 ( .A1(n12804), .A2(n7153), .ZN(n7150) );
  NAND2_X1 U9704 ( .A1(n7150), .A2(n7151), .ZN(n7680) );
  NAND3_X1 U9705 ( .A1(n8642), .A2(n8641), .A3(n6811), .ZN(n10891) );
  NAND3_X1 U9706 ( .A1(n8597), .A2(n8590), .A3(P2_REG3_REG_0__SCAN_IN), .ZN(
        n7155) );
  NAND2_X2 U9707 ( .A1(n14241), .A2(n12606), .ZN(n12885) );
  NAND3_X1 U9708 ( .A1(n14241), .A2(n12606), .A3(P2_REG0_REG_0__SCAN_IN), .ZN(
        n7156) );
  MUX2_X1 U9709 ( .A(n11885), .B(n10703), .S(n8473), .Z(n8031) );
  NAND2_X1 U9710 ( .A1(n8193), .A2(n8248), .ZN(n7159) );
  NAND2_X1 U9711 ( .A1(n8055), .A2(n7167), .ZN(n7166) );
  NOR2_X1 U9712 ( .A1(n6760), .A2(n7172), .ZN(n7171) );
  INV_X1 U9713 ( .A(n8386), .ZN(n7175) );
  NAND2_X1 U9714 ( .A1(n8076), .A2(n7177), .ZN(n7176) );
  INV_X1 U9715 ( .A(n8094), .ZN(n7178) );
  NAND2_X1 U9716 ( .A1(n9804), .A2(n9802), .ZN(n7614) );
  NAND2_X1 U9717 ( .A1(n9788), .A2(n9787), .ZN(n7201) );
  INV_X1 U9718 ( .A(n9569), .ZN(n7210) );
  NAND2_X1 U9719 ( .A1(n9810), .A2(n7213), .ZN(n7212) );
  NAND2_X1 U9720 ( .A1(n7216), .A2(n7220), .ZN(n9559) );
  NAND2_X1 U9721 ( .A1(n9697), .A2(n7217), .ZN(n7216) );
  NAND2_X1 U9722 ( .A1(n7630), .A2(n7230), .ZN(n7225) );
  AOI21_X1 U9723 ( .B1(n10009), .B2(n9585), .A(n7615), .ZN(n10018) );
  OAI21_X1 U9724 ( .B1(n10009), .B2(n7237), .A(n7236), .ZN(n9619) );
  INV_X1 U9725 ( .A(n7233), .ZN(n9620) );
  OR2_X1 U9726 ( .A1(n7905), .A2(n7904), .ZN(n7243) );
  NAND2_X1 U9727 ( .A1(n8452), .A2(n7252), .ZN(n8480) );
  INV_X1 U9728 ( .A(n7245), .ZN(n7248) );
  NAND2_X1 U9729 ( .A1(n8452), .A2(n8451), .ZN(n8455) );
  NAND2_X1 U9730 ( .A1(n12937), .A2(n12893), .ZN(n12940) );
  AND2_X2 U9731 ( .A1(n14618), .A2(n14610), .ZN(n14603) );
  NAND2_X1 U9732 ( .A1(n14618), .A2(n7261), .ZN(n7263) );
  AND2_X2 U9733 ( .A1(n14687), .A2(n7264), .ZN(n14634) );
  AND3_X2 U9734 ( .A1(n7910), .A2(n7908), .A3(n7909), .ZN(n11047) );
  INV_X1 U9735 ( .A(n15154), .ZN(n15153) );
  NAND2_X1 U9736 ( .A1(n9201), .A2(n7273), .ZN(n15154) );
  NAND2_X1 U9737 ( .A1(n7285), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7284) );
  NAND2_X1 U9738 ( .A1(n6744), .A2(n14957), .ZN(n7285) );
  NAND2_X1 U9739 ( .A1(n12519), .A2(n7293), .ZN(n7292) );
  OR2_X2 U9740 ( .A1(n11501), .A2(n11502), .ZN(n11721) );
  INV_X1 U9741 ( .A(n12540), .ZN(n7309) );
  NAND2_X1 U9742 ( .A1(n12163), .A2(n7314), .ZN(n12217) );
  NAND2_X1 U9743 ( .A1(n7318), .A2(n7316), .ZN(P3_U3488) );
  NOR2_X1 U9744 ( .A1(n15693), .A2(n10023), .ZN(n7317) );
  NAND2_X1 U9745 ( .A1(n13605), .A2(n15693), .ZN(n7318) );
  NAND3_X1 U9746 ( .A1(n13287), .A2(n7321), .A3(n15539), .ZN(n7320) );
  INV_X1 U9747 ( .A(n7325), .ZN(n7323) );
  OAI21_X1 U9748 ( .B1(n7328), .B2(n6837), .A(n7326), .ZN(n7325) );
  NAND2_X1 U9749 ( .A1(n7328), .A2(n13309), .ZN(n7326) );
  INV_X1 U9750 ( .A(n7337), .ZN(n11763) );
  NOR2_X2 U9751 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  AND2_X2 U9752 ( .A1(n7337), .A2(n7336), .ZN(n11854) );
  OR2_X1 U9753 ( .A1(n11759), .A2(n11760), .ZN(n7337) );
  NOR2_X2 U9754 ( .A1(n11858), .A2(n11873), .ZN(n11980) );
  XNOR2_X2 U9755 ( .A(n7339), .B(n7338), .ZN(n11858) );
  XNOR2_X2 U9756 ( .A(n13226), .B(n15012), .ZN(n15009) );
  OAI21_X2 U9757 ( .B1(n13225), .B2(n13224), .A(n13233), .ZN(n13226) );
  NAND2_X1 U9758 ( .A1(n13992), .A2(n7342), .ZN(n13933) );
  AND2_X2 U9759 ( .A1(n13992), .A2(n6802), .ZN(n13904) );
  NOR2_X2 U9760 ( .A1(n11609), .A2(n12663), .ZN(n11410) );
  NOR2_X2 U9761 ( .A1(n11890), .A2(n12749), .ZN(n7352) );
  NAND2_X1 U9762 ( .A1(n12034), .A2(n6695), .ZN(n7354) );
  NAND2_X1 U9763 ( .A1(n14785), .A2(n7365), .ZN(n7364) );
  CLKBUF_X1 U9764 ( .A(n7378), .Z(n7376) );
  NAND2_X1 U9765 ( .A1(n14629), .A2(n7387), .ZN(n7386) );
  AND2_X1 U9766 ( .A1(n14629), .A2(n14581), .ZN(n14615) );
  NAND2_X1 U9767 ( .A1(n14725), .A2(n6808), .ZN(n14698) );
  INV_X1 U9768 ( .A(n12048), .ZN(n7389) );
  NAND2_X1 U9769 ( .A1(n12597), .A2(n7400), .ZN(n7399) );
  OAI211_X1 U9770 ( .C1(n12597), .C2(n7401), .A(n7399), .B(n12603), .ZN(
        P3_U3169) );
  XNOR2_X1 U9771 ( .A(n12597), .B(n12980), .ZN(n13011) );
  NAND2_X1 U9772 ( .A1(n11513), .A2(n11512), .ZN(n11514) );
  AND2_X2 U9773 ( .A1(n7777), .A2(n7587), .ZN(n8548) );
  NAND3_X1 U9774 ( .A1(n8597), .A2(n8590), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n7524) );
  NAND3_X1 U9775 ( .A1(n7409), .A2(n7411), .A3(n7404), .ZN(n14143) );
  NAND3_X1 U9776 ( .A1(n7409), .A2(n7407), .A3(n7404), .ZN(n7417) );
  NAND2_X1 U9777 ( .A1(n13891), .A2(n7423), .ZN(n7422) );
  INV_X1 U9778 ( .A(n14033), .ZN(n7431) );
  NAND2_X1 U9779 ( .A1(n6995), .A2(n6738), .ZN(n14015) );
  INV_X1 U9780 ( .A(n6738), .ZN(n7439) );
  NAND2_X1 U9781 ( .A1(n10966), .A2(n11415), .ZN(n7445) );
  NAND2_X1 U9782 ( .A1(n13729), .A2(n7450), .ZN(n7446) );
  NAND2_X1 U9783 ( .A1(n7446), .A2(n7447), .ZN(n13750) );
  INV_X1 U9784 ( .A(n11165), .ZN(n7457) );
  NAND2_X1 U9785 ( .A1(n9103), .A2(n7463), .ZN(n7462) );
  OAI211_X1 U9786 ( .C1(n9103), .C2(n7465), .A(n13701), .B(n7462), .ZN(
        P2_U3192) );
  NAND2_X1 U9787 ( .A1(n12363), .A2(n12362), .ZN(n7473) );
  AOI21_X2 U9788 ( .B1(n7478), .B2(n7476), .A(n7475), .ZN(n7474) );
  NAND2_X1 U9789 ( .A1(n11416), .A2(n7488), .ZN(n7487) );
  NAND2_X1 U9790 ( .A1(n11438), .A2(n11437), .ZN(n11791) );
  NAND2_X1 U9791 ( .A1(n11417), .A2(n12901), .ZN(n11438) );
  NAND2_X1 U9792 ( .A1(n11832), .A2(n7492), .ZN(n7491) );
  NAND3_X1 U9793 ( .A1(n7491), .A2(n11445), .A3(n7490), .ZN(n11805) );
  INV_X1 U9794 ( .A(n11887), .ZN(n7521) );
  NAND2_X1 U9795 ( .A1(n8606), .A2(n7522), .ZN(n14235) );
  INV_X1 U9796 ( .A(n11765), .ZN(n7525) );
  NAND2_X1 U9797 ( .A1(n7993), .A2(n7530), .ZN(n7528) );
  AND2_X1 U9798 ( .A1(n7815), .A2(n7811), .ZN(n7532) );
  NAND2_X1 U9799 ( .A1(n7834), .A2(n6798), .ZN(n7539) );
  NAND2_X1 U9800 ( .A1(n7834), .A2(n7833), .ZN(n8086) );
  NAND3_X1 U9801 ( .A1(n7541), .A2(n8085), .A3(n7540), .ZN(n7538) );
  INV_X1 U9802 ( .A(n11681), .ZN(n7548) );
  AOI21_X2 U9803 ( .B1(n11681), .B2(n11545), .A(n6714), .ZN(n7547) );
  NAND2_X1 U9804 ( .A1(n7554), .A2(n7555), .ZN(n8424) );
  NAND2_X1 U9805 ( .A1(n8403), .A2(n7556), .ZN(n7555) );
  NAND2_X1 U9806 ( .A1(n7569), .A2(n7567), .ZN(n8324) );
  INV_X1 U9807 ( .A(n8320), .ZN(n7568) );
  NAND2_X1 U9808 ( .A1(n8320), .A2(n8319), .ZN(n7570) );
  NAND2_X1 U9809 ( .A1(n8324), .A2(n8325), .ZN(n8322) );
  NAND2_X1 U9810 ( .A1(n7573), .A2(n7572), .ZN(n11027) );
  NAND2_X1 U9811 ( .A1(n14258), .A2(n7576), .ZN(n7574) );
  OAI211_X1 U9812 ( .C1(n14258), .C2(n7575), .A(n7574), .B(n10493), .ZN(
        P1_U3220) );
  NAND3_X1 U9813 ( .A1(n10444), .A2(n14710), .A3(n14411), .ZN(n10243) );
  OR2_X2 U9814 ( .A1(n7586), .A2(n6679), .ZN(n10457) );
  NAND3_X1 U9815 ( .A1(n6682), .A2(n6694), .A3(n10424), .ZN(n7591) );
  NAND3_X1 U9816 ( .A1(n14352), .A2(n6682), .A3(n10424), .ZN(n7592) );
  NAND2_X1 U9817 ( .A1(n14378), .A2(n7605), .ZN(n7604) );
  NAND2_X1 U9818 ( .A1(n10366), .A2(n10367), .ZN(n7611) );
  OAI21_X2 U9819 ( .B1(n9994), .B2(n9584), .A(n7616), .ZN(n10009) );
  NAND2_X1 U9820 ( .A1(n9956), .A2(n6840), .ZN(n7623) );
  AOI21_X1 U9821 ( .B1(n10212), .B2(n11488), .A(n7639), .ZN(n7638) );
  NOR2_X1 U9822 ( .A1(n10059), .A2(n11361), .ZN(n7639) );
  NAND2_X1 U9823 ( .A1(n10211), .A2(n15609), .ZN(n7640) );
  NAND2_X1 U9824 ( .A1(n11958), .A2(n7646), .ZN(n7644) );
  NAND2_X1 U9825 ( .A1(n7660), .A2(n6806), .ZN(n12457) );
  AND2_X1 U9826 ( .A1(n10223), .A2(n7669), .ZN(n10220) );
  OR2_X1 U9827 ( .A1(n12821), .A2(n7679), .ZN(n7678) );
  INV_X1 U9828 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9829 ( .A1(n11517), .A2(n6816), .ZN(n7695) );
  NAND2_X1 U9830 ( .A1(n7695), .A2(n7696), .ZN(n11707) );
  NAND3_X1 U9831 ( .A1(n7769), .A2(n7773), .A3(n7959), .ZN(n7884) );
  NAND2_X1 U9832 ( .A1(n11278), .A2(n11277), .ZN(n11306) );
  NAND2_X1 U9833 ( .A1(n11207), .A2(n7730), .ZN(n11278) );
  NAND2_X1 U9834 ( .A1(n12409), .A2(n7736), .ZN(n7732) );
  NAND2_X1 U9835 ( .A1(n7732), .A2(n7733), .ZN(n14773) );
  NAND2_X1 U9836 ( .A1(n8548), .A2(n7743), .ZN(n8545) );
  AOI22_X1 U9837 ( .A1(n13911), .A2(n13910), .B1(n13909), .B2(n14125), .ZN(
        n14122) );
  OAI21_X1 U9838 ( .B1(n8613), .B2(n8612), .A(n12644), .ZN(n8621) );
  NAND2_X1 U9839 ( .A1(n8150), .A2(n8149), .ZN(n8192) );
  NAND2_X1 U9840 ( .A1(n8424), .A2(n8425), .ZN(n8429) );
  NAND2_X1 U9841 ( .A1(n11700), .A2(n11699), .ZN(n12032) );
  NAND2_X1 U9842 ( .A1(n11698), .A2(n11697), .ZN(n11700) );
  NAND2_X1 U9843 ( .A1(n8536), .A2(n7759), .ZN(n8533) );
  OAI21_X1 U9844 ( .B1(n9129), .B2(n13692), .A(n7749), .ZN(P2_U3186) );
  XNOR2_X1 U9845 ( .A(n15612), .B(n15588), .ZN(n11495) );
  INV_X1 U9846 ( .A(n10040), .ZN(n10035) );
  INV_X1 U9847 ( .A(n9876), .ZN(n9873) );
  NAND2_X1 U9848 ( .A1(n8572), .A2(n8571), .ZN(n9065) );
  OR2_X2 U9849 ( .A1(n10317), .A2(n10316), .ZN(n11947) );
  NAND2_X1 U9850 ( .A1(n10241), .A2(n11047), .ZN(n8495) );
  INV_X1 U9851 ( .A(n12644), .ZN(n12645) );
  INV_X1 U9852 ( .A(n8578), .ZN(n8572) );
  OR2_X1 U9853 ( .A1(n12858), .A2(n8457), .ZN(n8460) );
  AND2_X1 U9854 ( .A1(n10891), .A2(n15381), .ZN(n12647) );
  NAND2_X1 U9855 ( .A1(n7948), .A2(n8495), .ZN(n15201) );
  INV_X1 U9856 ( .A(n12885), .ZN(n12840) );
  OAI222_X1 U9857 ( .A1(P3_U3151), .A2(n13268), .B1(n12971), .B2(n12970), .C1(
        n13672), .C2(n12969), .ZN(P3_U3268) );
  OR2_X1 U9858 ( .A1(n7785), .A2(n7784), .ZN(n7787) );
  OR2_X1 U9859 ( .A1(n8430), .A2(n7898), .ZN(n7901) );
  OR2_X1 U9860 ( .A1(n8430), .A2(n7892), .ZN(n7895) );
  XNOR2_X1 U9861 ( .A(n12569), .B(n12567), .ZN(n13112) );
  NAND2_X1 U9862 ( .A1(n14705), .A2(n14547), .ZN(n14684) );
  AND2_X1 U9863 ( .A1(n10972), .A2(n12930), .ZN(n14095) );
  OR2_X1 U9864 ( .A1(n12305), .A2(n12223), .ZN(n7745) );
  AND2_X1 U9865 ( .A1(n7844), .A2(n7843), .ZN(n7746) );
  AND4_X1 U9866 ( .A1(n13346), .A2(n13362), .A3(n10056), .A4(n10055), .ZN(
        n7747) );
  NOR2_X1 U9867 ( .A1(n9128), .A2(n9127), .ZN(n7749) );
  AND2_X1 U9868 ( .A1(n7267), .A2(n14578), .ZN(n7751) );
  OR2_X1 U9869 ( .A1(n12977), .A2(n13403), .ZN(n7752) );
  AND2_X1 U9870 ( .A1(n14563), .A2(n14562), .ZN(n7753) );
  INV_X1 U9871 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12967) );
  INV_X1 U9872 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11135) );
  AND2_X1 U9873 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7755) );
  AND2_X1 U9874 ( .A1(n8292), .A2(n14299), .ZN(n7756) );
  NOR2_X1 U9875 ( .A1(n8152), .A2(n8151), .ZN(n7757) );
  AND2_X1 U9876 ( .A1(n9030), .A2(n9029), .ZN(n7758) );
  INV_X1 U9877 ( .A(n14702), .ZN(n14572) );
  AND2_X1 U9878 ( .A1(n14692), .A2(n14575), .ZN(n7760) );
  AND2_X1 U9879 ( .A1(n14557), .A2(n14986), .ZN(n7761) );
  OR2_X1 U9880 ( .A1(n8557), .A2(n8556), .ZN(n7762) );
  INV_X1 U9881 ( .A(n12165), .ZN(n12164) );
  OR2_X1 U9882 ( .A1(n11152), .A2(n6680), .ZN(n7947) );
  INV_X1 U9883 ( .A(n7969), .ZN(n7970) );
  NAND2_X1 U9884 ( .A1(n7971), .A2(n7970), .ZN(n7972) );
  INV_X1 U9885 ( .A(n8011), .ZN(n8012) );
  NAND2_X1 U9886 ( .A1(n8037), .A2(n8036), .ZN(n8055) );
  NAND2_X1 U9887 ( .A1(n8188), .A2(n8493), .ZN(n8189) );
  NOR2_X1 U9888 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  INV_X1 U9889 ( .A(n14899), .ZN(n8244) );
  AND2_X1 U9890 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  AOI21_X1 U9891 ( .B1(n12820), .B2(n12819), .A(n12818), .ZN(n12822) );
  INV_X1 U9892 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7770) );
  INV_X1 U9893 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9298) );
  AOI22_X1 U9894 ( .A1(n8429), .A2(n8428), .B1(n8427), .B2(n8426), .ZN(n8445)
         );
  INV_X1 U9895 ( .A(n13346), .ZN(n12539) );
  NOR2_X1 U9896 ( .A1(n9959), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9972) );
  INV_X1 U9897 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9576) );
  INV_X1 U9898 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U9899 ( .A1(n14610), .A2(n14557), .ZN(n14553) );
  INV_X1 U9900 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7780) );
  INV_X1 U9901 ( .A(n8217), .ZN(n7855) );
  OR2_X1 U9902 ( .A1(n9939), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U9903 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  NAND2_X1 U9904 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n9576), .ZN(n9577) );
  AND2_X1 U9905 ( .A1(n8920), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8940) );
  INV_X1 U9906 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8780) );
  NOR2_X1 U9907 ( .A1(n8871), .A2(n12201), .ZN(n8870) );
  NOR2_X1 U9908 ( .A1(n12749), .A2(n13789), .ZN(n12124) );
  INV_X1 U9909 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7781) );
  AND2_X1 U9910 ( .A1(n12981), .A2(n7752), .ZN(n12978) );
  INV_X1 U9911 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U9912 ( .A1(n11479), .A2(n11346), .ZN(n12608) );
  OAI22_X1 U9913 ( .A1(n13411), .A2(n12531), .B1(n13403), .B2(n13631), .ZN(
        n13400) );
  NAND2_X1 U9914 ( .A1(n9835), .A2(n10143), .ZN(n9836) );
  NAND2_X1 U9915 ( .A1(n15575), .A2(n11722), .ZN(n15560) );
  INV_X1 U9916 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9596) );
  INV_X1 U9917 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U9918 ( .A1(n8916), .A2(n10502), .ZN(n8646) );
  NAND2_X2 U9919 ( .A1(n10979), .A2(n12651), .ZN(n8653) );
  INV_X1 U9920 ( .A(n13751), .ZN(n8982) );
  INV_X1 U9921 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8852) );
  BUF_X4 U9922 ( .A(n12825), .Z(n12837) );
  NOR2_X1 U9923 ( .A1(n9020), .A2(n8592), .ZN(n9021) );
  OR2_X1 U9924 ( .A1(n8974), .A2(n8973), .ZN(n8988) );
  INV_X1 U9925 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8853) );
  OR2_X1 U9926 ( .A1(n14159), .A2(n13898), .ZN(n13899) );
  INV_X1 U9927 ( .A(n10296), .ZN(n10451) );
  INV_X1 U9928 ( .A(n10296), .ZN(n10437) );
  NAND2_X1 U9929 ( .A1(n8328), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8353) );
  OR2_X1 U9930 ( .A1(n15284), .A2(n14400), .ZN(n12349) );
  NAND2_X1 U9931 ( .A1(n7837), .A2(n10519), .ZN(n7840) );
  NAND2_X1 U9932 ( .A1(n7808), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7804) );
  NOR2_X1 U9933 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9188), .ZN(n9140) );
  NAND2_X1 U9934 ( .A1(n9817), .A2(n13096), .ZN(n9829) );
  OR2_X1 U9935 ( .A1(n11356), .A2(n11355), .ZN(n13138) );
  AND2_X1 U9936 ( .A1(n11329), .A2(n10228), .ZN(n10495) );
  AND2_X1 U9937 ( .A1(n11556), .A2(n11555), .ZN(n11568) );
  INV_X1 U9938 ( .A(n13371), .ZN(n13402) );
  INV_X1 U9939 ( .A(n10159), .ZN(n13477) );
  INV_X1 U9940 ( .A(n15033), .ZN(n13522) );
  INV_X1 U9941 ( .A(n13659), .ZN(n12626) );
  INV_X1 U9942 ( .A(n10229), .ZN(n11530) );
  INV_X1 U9943 ( .A(n13097), .ZN(n13532) );
  OAI21_X1 U9944 ( .B1(n10213), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10215) );
  OR2_X1 U9945 ( .A1(n9739), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U9946 ( .A1(n9126), .A2(n9125), .ZN(n9127) );
  OR3_X1 U9947 ( .A1(n8854), .A2(n8852), .A3(n8853), .ZN(n8871) );
  OR2_X1 U9948 ( .A1(n13742), .A2(n14090), .ZN(n13759) );
  OR2_X1 U9949 ( .A1(n8902), .A2(n8901), .ZN(n8922) );
  OR2_X1 U9950 ( .A1(n11904), .A2(n11903), .ZN(n12431) );
  INV_X1 U9951 ( .A(n13960), .ZN(n13900) );
  NAND2_X1 U9952 ( .A1(n15392), .A2(n11412), .ZN(n14102) );
  NAND2_X1 U9953 ( .A1(n10748), .A2(n10752), .ZN(n15388) );
  INV_X1 U9954 ( .A(n9118), .ZN(n10963) );
  INV_X1 U9955 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8680) );
  INV_X1 U9956 ( .A(n10929), .ZN(n10264) );
  AND2_X1 U9957 ( .A1(n14953), .A2(n10703), .ZN(n10560) );
  OR3_X1 U9958 ( .A1(n15283), .A2(n10560), .A3(n11139), .ZN(n10482) );
  AOI21_X1 U9959 ( .B1(n8531), .B2(n10480), .A(n8530), .ZN(n8532) );
  AND2_X1 U9960 ( .A1(n8310), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8312) );
  INV_X1 U9961 ( .A(n7788), .ZN(n7790) );
  OR2_X1 U9962 ( .A1(n8468), .A2(n7899), .ZN(n7900) );
  INV_X1 U9963 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10953) );
  AND2_X1 U9964 ( .A1(n11096), .A2(n11095), .ZN(n11098) );
  NAND2_X1 U9965 ( .A1(n14698), .A2(n14574), .ZN(n14686) );
  INV_X1 U9966 ( .A(n14987), .ZN(n15097) );
  NAND2_X1 U9967 ( .A1(n12032), .A2(n12031), .ZN(n12034) );
  XNOR2_X1 U9968 ( .A(n7853), .B(SI_16_), .ZN(n8203) );
  AND3_X1 U9969 ( .A1(n9954), .A2(n9953), .A3(n9952), .ZN(n13412) );
  INV_X1 U9970 ( .A(n13149), .ZN(n13134) );
  NAND2_X1 U9971 ( .A1(n15591), .A2(n11359), .ZN(n15490) );
  NAND2_X1 U9972 ( .A1(n9990), .A2(n9989), .ZN(n13372) );
  INV_X1 U9973 ( .A(n13517), .ZN(n13488) );
  INV_X1 U9974 ( .A(n15520), .ZN(n15550) );
  AND2_X1 U9975 ( .A1(n11568), .A2(n11560), .ZN(n15539) );
  NAND2_X1 U9976 ( .A1(n10005), .A2(n10004), .ZN(n13359) );
  INV_X1 U9977 ( .A(n15594), .ZN(n15615) );
  NAND2_X1 U9978 ( .A1(n11499), .A2(n11498), .ZN(n15599) );
  NOR2_X1 U9979 ( .A1(n12488), .A2(n15607), .ZN(n15033) );
  NOR2_X1 U9980 ( .A1(n11529), .A2(n11482), .ZN(n12633) );
  INV_X1 U9981 ( .A(n15602), .ZN(n15656) );
  INV_X1 U9982 ( .A(n15654), .ZN(n15672) );
  INV_X1 U9983 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9605) );
  INV_X1 U9984 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9597) );
  XNOR2_X1 U9985 ( .A(n10215), .B(n10214), .ZN(n11531) );
  OR2_X1 U9986 ( .A1(n9741), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9772) );
  INV_X1 U9987 ( .A(n13785), .ZN(n9100) );
  INV_X1 U9988 ( .A(n15381), .ZN(n12648) );
  NOR2_X1 U9989 ( .A1(n15400), .A2(n9120), .ZN(n9105) );
  OR2_X1 U9990 ( .A1(n8721), .A2(n13953), .ZN(n9060) );
  INV_X1 U9991 ( .A(n15364), .ZN(n11902) );
  AND2_X1 U9992 ( .A1(n10782), .A2(n10783), .ZN(n15364) );
  INV_X1 U9993 ( .A(n13902), .ZN(n13940) );
  AND2_X1 U9994 ( .A1(n15471), .A2(n15470), .ZN(n15454) );
  AND2_X1 U9995 ( .A1(n10962), .A2(n10961), .ZN(n12121) );
  INV_X1 U9996 ( .A(n14388), .ZN(n15088) );
  AND4_X1 U9997 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n14550)
         );
  OR2_X1 U9998 ( .A1(n15180), .A2(n15169), .ZN(n12377) );
  INV_X1 U9999 ( .A(n12377), .ZN(n15188) );
  INV_X1 U10000 ( .A(n15193), .ZN(n14489) );
  INV_X1 U10001 ( .A(n15209), .ZN(n14862) );
  INV_X1 U10002 ( .A(n15289), .ZN(n15248) );
  NAND2_X1 U10003 ( .A1(n15274), .A2(n15266), .ZN(n15289) );
  NAND2_X1 U10004 ( .A1(n8544), .A2(n8543), .ZN(n15253) );
  OR2_X1 U10005 ( .A1(n10486), .A2(P1_U3086), .ZN(n11322) );
  OR2_X1 U10006 ( .A1(n10466), .A2(n14952), .ZN(n10708) );
  XNOR2_X1 U10007 ( .A(n7963), .B(n7962), .ZN(n10537) );
  AND2_X1 U10008 ( .A1(n11557), .A2(n11556), .ZN(n15538) );
  INV_X1 U10009 ( .A(n13151), .ZN(n13121) );
  OR2_X1 U10010 ( .A1(n13155), .A2(n12543), .ZN(n15520) );
  INV_X1 U10011 ( .A(n15500), .ZN(n15547) );
  AND2_X1 U10012 ( .A1(n13442), .A2(n13441), .ZN(n13580) );
  AND2_X1 U10013 ( .A1(n13351), .A2(n11718), .ZN(n13539) );
  INV_X2 U10014 ( .A(n15625), .ZN(n15627) );
  INV_X1 U10015 ( .A(n15693), .ZN(n15691) );
  INV_X1 U10016 ( .A(n13582), .ZN(n13604) );
  NAND2_X1 U10017 ( .A1(n10725), .A2(n11344), .ZN(n10726) );
  INV_X1 U10018 ( .A(SI_25_), .ZN(n12277) );
  INV_X1 U10019 ( .A(SI_14_), .ZN(n10577) );
  INV_X1 U10020 ( .A(n13783), .ZN(n13747) );
  NAND2_X1 U10021 ( .A1(n9105), .A2(n9099), .ZN(n13785) );
  NAND2_X1 U10022 ( .A1(n15302), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15379) );
  INV_X1 U10023 ( .A(n15371), .ZN(n15363) );
  NAND2_X1 U10024 ( .A1(n15392), .A2(n11409), .ZN(n14133) );
  INV_X1 U10025 ( .A(n15489), .ZN(n15487) );
  AND3_X1 U10026 ( .A1(n15464), .A2(n15463), .A3(n15462), .ZN(n15486) );
  INV_X1 U10027 ( .A(n15475), .ZN(n15474) );
  OR2_X1 U10028 ( .A1(n15396), .A2(n15395), .ZN(n15397) );
  INV_X1 U10029 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14250) );
  INV_X1 U10030 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11017) );
  INV_X1 U10031 ( .A(n14866), .ZN(n14679) );
  AND4_X1 U10032 ( .A1(n8177), .A2(n8176), .A3(n8175), .A4(n8174), .ZN(n14562)
         );
  OR2_X1 U10033 ( .A1(n15180), .A2(n10588), .ZN(n15193) );
  OR2_X1 U10034 ( .A1(n15180), .A2(n10596), .ZN(n15183) );
  INV_X1 U10035 ( .A(n15177), .ZN(n15197) );
  INV_X1 U10036 ( .A(n15126), .ZN(n14802) );
  INV_X1 U10037 ( .A(n15300), .ZN(n15140) );
  OR2_X1 U10038 ( .A1(n11322), .A2(n11321), .ZN(n15290) );
  AND2_X1 U10039 ( .A1(n10559), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10552) );
  INV_X1 U10040 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12329) );
  INV_X1 U10041 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10790) );
  XNOR2_X1 U10042 ( .A(n9544), .B(n9543), .ZN(n9545) );
  AND2_X1 U10043 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10750), .ZN(P2_U3947) );
  NAND2_X1 U10044 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7975) );
  INV_X1 U10045 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10046 ( .A1(n8001), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8017) );
  INV_X1 U10047 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8016) );
  INV_X1 U10048 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10049 ( .A1(n8078), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10050 ( .A1(n8137), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8121) );
  INV_X1 U10051 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8114) );
  INV_X1 U10052 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U10053 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7763) );
  INV_X1 U10054 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14346) );
  INV_X1 U10055 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14299) );
  OR2_X1 U10056 ( .A1(n8312), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U10057 ( .A1(n7764), .A2(n8327), .ZN(n14282) );
  INV_X1 U10058 ( .A(n14282), .ZN(n14675) );
  NOR2_X1 U10059 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7767) );
  AND4_X2 U10060 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n9392), .ZN(n7769)
         );
  AND2_X2 U10061 ( .A1(n7921), .A2(n7768), .ZN(n7959) );
  INV_X2 U10062 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8089) );
  NAND4_X1 U10063 ( .A1(n7778), .A2(n7881), .A3(n6964), .A4(n8538), .ZN(n7779)
         );
  NAND2_X1 U10064 ( .A1(n7785), .A2(n7786), .ZN(n12514) );
  XNOR2_X2 U10065 ( .A(n7783), .B(n12508), .ZN(n7789) );
  INV_X1 U10066 ( .A(n6972), .ZN(n8293) );
  NAND2_X1 U10067 ( .A1(n14675), .A2(n8293), .ZN(n7796) );
  INV_X1 U10068 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n7793) );
  INV_X2 U10069 ( .A(n8469), .ZN(n7929) );
  NAND2_X1 U10070 ( .A1(n7929), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10071 ( .A1(n8461), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7791) );
  OAI211_X1 U10072 ( .C1(n7793), .C2(n8465), .A(n7792), .B(n7791), .ZN(n7794)
         );
  INV_X1 U10073 ( .A(n7794), .ZN(n7795) );
  INV_X1 U10074 ( .A(n14576), .ZN(n14395) );
  INV_X1 U10075 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7800) );
  NAND4_X1 U10076 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7802) );
  XNOR2_X1 U10077 ( .A(n7806), .B(SI_1_), .ZN(n7905) );
  MUX2_X1 U10078 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n7808), .Z(n7805) );
  NAND2_X1 U10079 ( .A1(n7805), .A2(SI_0_), .ZN(n7904) );
  NAND2_X1 U10080 ( .A1(n7806), .A2(SI_1_), .ZN(n7807) );
  MUX2_X1 U10081 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n10502), .Z(n7920) );
  NAND2_X1 U10082 ( .A1(n7809), .A2(n7920), .ZN(n7812) );
  NAND2_X1 U10083 ( .A1(n7810), .A2(SI_2_), .ZN(n7811) );
  INV_X1 U10084 ( .A(n7935), .ZN(n7813) );
  NAND2_X1 U10085 ( .A1(n7814), .A2(SI_3_), .ZN(n7815) );
  XNOR2_X1 U10086 ( .A(n7817), .B(SI_4_), .ZN(n7962) );
  INV_X1 U10087 ( .A(n7962), .ZN(n7816) );
  NAND2_X1 U10088 ( .A1(n7817), .A2(SI_4_), .ZN(n7818) );
  MUX2_X1 U10089 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n10502), .Z(n7820) );
  XNOR2_X1 U10090 ( .A(n7820), .B(SI_5_), .ZN(n7981) );
  INV_X1 U10091 ( .A(n7981), .ZN(n7819) );
  NAND2_X1 U10092 ( .A1(n7982), .A2(n7819), .ZN(n7822) );
  NAND2_X1 U10093 ( .A1(n7820), .A2(SI_5_), .ZN(n7821) );
  XNOR2_X1 U10094 ( .A(n7824), .B(SI_6_), .ZN(n7992) );
  INV_X1 U10095 ( .A(n7992), .ZN(n7823) );
  NAND2_X1 U10096 ( .A1(n7824), .A2(SI_6_), .ZN(n7825) );
  MUX2_X1 U10097 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n10497), .Z(n7826) );
  XNOR2_X1 U10098 ( .A(n7826), .B(SI_7_), .ZN(n8024) );
  MUX2_X1 U10099 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n10502), .Z(n7828) );
  XNOR2_X1 U10100 ( .A(n7828), .B(SI_8_), .ZN(n8046) );
  INV_X1 U10101 ( .A(n8046), .ZN(n7827) );
  NAND2_X1 U10102 ( .A1(n8047), .A2(n7827), .ZN(n7830) );
  NAND2_X1 U10103 ( .A1(n7828), .A2(SI_8_), .ZN(n7829) );
  MUX2_X1 U10104 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n10497), .Z(n7832) );
  XNOR2_X1 U10105 ( .A(n7832), .B(SI_9_), .ZN(n8065) );
  INV_X1 U10106 ( .A(n8065), .ZN(n7831) );
  NAND2_X1 U10107 ( .A1(n7832), .A2(SI_9_), .ZN(n7833) );
  MUX2_X1 U10108 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n10502), .Z(n7836) );
  MUX2_X1 U10109 ( .A(n10691), .B(n10689), .S(n10497), .Z(n7837) );
  INV_X1 U10110 ( .A(n7837), .ZN(n7838) );
  NAND2_X1 U10111 ( .A1(n7838), .A2(SI_11_), .ZN(n7839) );
  NAND2_X1 U10112 ( .A1(n7840), .A2(n7839), .ZN(n8102) );
  MUX2_X1 U10113 ( .A(n10721), .B(n7613), .S(n10502), .Z(n7841) );
  NAND2_X1 U10114 ( .A1(n7841), .A2(n10546), .ZN(n7844) );
  INV_X1 U10115 ( .A(n7841), .ZN(n7842) );
  NAND2_X1 U10116 ( .A1(n7842), .A2(SI_12_), .ZN(n7843) );
  NAND2_X1 U10117 ( .A1(n8143), .A2(n7746), .ZN(n7845) );
  MUX2_X1 U10118 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n10497), .Z(n8127) );
  INV_X1 U10119 ( .A(n8127), .ZN(n7846) );
  MUX2_X1 U10120 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n10502), .Z(n8110) );
  INV_X1 U10121 ( .A(n8110), .ZN(n8159) );
  MUX2_X1 U10122 ( .A(n11017), .B(n11016), .S(n10497), .Z(n8163) );
  INV_X1 U10123 ( .A(n8163), .ZN(n7847) );
  NAND2_X1 U10124 ( .A1(n7847), .A2(SI_15_), .ZN(n7850) );
  OAI21_X1 U10125 ( .B1(n10577), .B2(n8159), .A(n7850), .ZN(n7848) );
  INV_X1 U10126 ( .A(n7848), .ZN(n7849) );
  NOR2_X1 U10127 ( .A1(n8110), .A2(SI_14_), .ZN(n7851) );
  INV_X1 U10128 ( .A(SI_15_), .ZN(n10647) );
  AOI22_X1 U10129 ( .A1(n7851), .A2(n7850), .B1(n8163), .B2(n10647), .ZN(n7852) );
  MUX2_X1 U10130 ( .A(n10927), .B(n9571), .S(n10502), .Z(n7853) );
  NAND2_X1 U10131 ( .A1(n7853), .A2(n10693), .ZN(n7854) );
  MUX2_X1 U10132 ( .A(n10960), .B(n7016), .S(n10497), .Z(n8217) );
  NAND2_X1 U10133 ( .A1(n7855), .A2(SI_17_), .ZN(n7856) );
  MUX2_X1 U10134 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n10502), .Z(n8249) );
  INV_X1 U10135 ( .A(n8249), .ZN(n7857) );
  MUX2_X1 U10136 ( .A(n12967), .B(n9576), .S(n10497), .Z(n7860) );
  INV_X1 U10137 ( .A(n7860), .ZN(n7861) );
  NAND2_X1 U10138 ( .A1(n7861), .A2(SI_19_), .ZN(n7862) );
  NAND2_X1 U10139 ( .A1(n7863), .A2(n7862), .ZN(n8261) );
  MUX2_X1 U10140 ( .A(n12017), .B(n7203), .S(n10497), .Z(n8302) );
  MUX2_X1 U10141 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n10497), .Z(n8300) );
  INV_X1 U10142 ( .A(n8300), .ZN(n7864) );
  INV_X1 U10143 ( .A(SI_20_), .ZN(n11085) );
  NOR2_X1 U10144 ( .A1(n7864), .A2(n11085), .ZN(n7866) );
  AOI22_X1 U10145 ( .A1(n7866), .A2(n6707), .B1(n7865), .B2(SI_21_), .ZN(n7867) );
  INV_X1 U10146 ( .A(n9004), .ZN(n7868) );
  MUX2_X1 U10147 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n10502), .Z(n9003) );
  NAND2_X1 U10148 ( .A1(n7868), .A2(n9003), .ZN(n7870) );
  NAND2_X1 U10149 ( .A1(n8336), .A2(SI_22_), .ZN(n7869) );
  NAND2_X1 U10150 ( .A1(n7870), .A2(n7869), .ZN(n7872) );
  MUX2_X1 U10151 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n10497), .Z(n8339) );
  XNOR2_X1 U10152 ( .A(n8339), .B(SI_23_), .ZN(n7871) );
  XNOR2_X2 U10153 ( .A(n7875), .B(n7874), .ZN(n8555) );
  NAND2_X2 U10154 ( .A1(n10562), .A2(n10502), .ZN(n8457) );
  NAND2_X1 U10155 ( .A1(n12179), .A2(n8484), .ZN(n7878) );
  NAND2_X4 U10156 ( .A1(n10562), .A2(n10501), .ZN(n8458) );
  INV_X1 U10157 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12182) );
  OR2_X1 U10158 ( .A1(n8458), .A2(n12182), .ZN(n7877) );
  NAND2_X2 U10159 ( .A1(n7878), .A2(n7877), .ZN(n14866) );
  NAND2_X1 U10160 ( .A1(n7879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U10161 ( .A1(n7882), .A2(n7881), .ZN(n7889) );
  NAND2_X1 U10162 ( .A1(n7889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7883) );
  INV_X1 U10163 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7886) );
  INV_X1 U10164 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10165 ( .A1(n6681), .A2(n10479), .ZN(n7891) );
  MUX2_X1 U10166 ( .A(n14395), .B(n14866), .S(n7944), .Z(n8325) );
  NAND2_X1 U10167 ( .A1(n7929), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7896) );
  INV_X1 U10168 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10169 ( .A1(n8466), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7894) );
  INV_X1 U10170 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10244) );
  OR2_X1 U10171 ( .A1(n8468), .A2(n10244), .ZN(n7893) );
  NAND2_X1 U10172 ( .A1(n10497), .A2(SI_0_), .ZN(n7897) );
  XNOR2_X1 U10173 ( .A(n7897), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14956) );
  MUX2_X1 U10174 ( .A(n14955), .B(n14956), .S(n10562), .Z(n14806) );
  OR2_X2 U10175 ( .A1(n14411), .A2(n11046), .ZN(n8498) );
  NAND2_X1 U10176 ( .A1(n10703), .A2(n11885), .ZN(n10698) );
  NAND2_X1 U10177 ( .A1(n8498), .A2(n10698), .ZN(n7911) );
  NAND2_X1 U10178 ( .A1(n14411), .A2(n11046), .ZN(n8497) );
  NAND2_X1 U10179 ( .A1(n8466), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7903) );
  INV_X1 U10180 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10599) );
  OR2_X1 U10181 ( .A1(n8469), .A2(n10599), .ZN(n7902) );
  INV_X1 U10182 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7898) );
  INV_X1 U10183 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7899) );
  NAND4_X1 U10184 ( .A1(n7903), .A2(n7900), .A3(n7901), .A4(n7902), .ZN(n10241) );
  INV_X1 U10185 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10498) );
  OR2_X1 U10186 ( .A1(n8458), .A2(n10498), .ZN(n7910) );
  XNOR2_X1 U10187 ( .A(n7905), .B(n7904), .ZN(n10499) );
  OR2_X1 U10188 ( .A1(n8457), .A2(n10499), .ZN(n7909) );
  INV_X1 U10189 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U10190 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14955), .ZN(n7906) );
  OR2_X1 U10191 ( .A1(n10562), .A2(n10598), .ZN(n7908) );
  NAND3_X1 U10192 ( .A1(n7911), .A2(n8497), .A3(n8495), .ZN(n7912) );
  OR2_X1 U10193 ( .A1(n10241), .A2(n11047), .ZN(n8496) );
  NAND2_X1 U10194 ( .A1(n7912), .A2(n8496), .ZN(n7940) );
  NAND2_X1 U10195 ( .A1(n7929), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7918) );
  INV_X1 U10196 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7913) );
  OR2_X1 U10197 ( .A1(n8430), .A2(n7913), .ZN(n7917) );
  INV_X1 U10198 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7914) );
  INV_X1 U10199 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10590) );
  OR2_X1 U10200 ( .A1(n8468), .A2(n10590), .ZN(n7915) );
  XNOR2_X1 U10201 ( .A(n7919), .B(n7920), .ZN(n8650) );
  INV_X1 U10202 ( .A(n8650), .ZN(n10508) );
  OR2_X1 U10203 ( .A1(n8457), .A2(n10508), .ZN(n7928) );
  INV_X1 U10204 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10500) );
  OR2_X1 U10205 ( .A1(n8458), .A2(n10500), .ZN(n7927) );
  NOR2_X1 U10206 ( .A1(n7921), .A2(n7784), .ZN(n7922) );
  MUX2_X1 U10207 ( .A(n7784), .B(n7922), .S(P1_IR_REG_2__SCAN_IN), .Z(n7923)
         );
  INV_X1 U10208 ( .A(n7923), .ZN(n7925) );
  INV_X1 U10209 ( .A(n7959), .ZN(n7924) );
  OR2_X1 U10210 ( .A1(n10562), .A2(n14429), .ZN(n7926) );
  AND3_X2 U10211 ( .A1(n7928), .A2(n7927), .A3(n7926), .ZN(n15232) );
  NAND2_X1 U10212 ( .A1(n14408), .A2(n15232), .ZN(n8500) );
  NAND2_X1 U10213 ( .A1(n7929), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7934) );
  OR2_X1 U10214 ( .A1(n8430), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7933) );
  INV_X1 U10215 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7930) );
  OR2_X1 U10216 ( .A1(n8198), .A2(n7930), .ZN(n7932) );
  INV_X1 U10217 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10591) );
  OR2_X1 U10218 ( .A1(n8468), .A2(n10591), .ZN(n7931) );
  NAND4_X2 U10219 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n14407) );
  XNOR2_X1 U10220 ( .A(n7936), .B(n7935), .ZN(n8665) );
  INV_X1 U10221 ( .A(n8665), .ZN(n10510) );
  INV_X1 U10222 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10511) );
  OR2_X1 U10223 ( .A1(n8458), .A2(n10511), .ZN(n7939) );
  OR2_X1 U10224 ( .A1(n7959), .A2(n7784), .ZN(n7937) );
  OR2_X1 U10225 ( .A1(n10562), .A2(n14446), .ZN(n7938) );
  NAND2_X1 U10226 ( .A1(n14407), .A2(n15239), .ZN(n8499) );
  NAND4_X1 U10227 ( .A1(n7940), .A2(n8031), .A3(n8500), .A4(n8499), .ZN(n7952)
         );
  INV_X1 U10228 ( .A(n11151), .ZN(n7941) );
  NAND3_X1 U10229 ( .A1(n7941), .A2(n8031), .A3(n8499), .ZN(n7943) );
  OR2_X1 U10230 ( .A1(n8499), .A2(n8031), .ZN(n7942) );
  AND2_X1 U10231 ( .A1(n7943), .A2(n7942), .ZN(n7951) );
  OR2_X2 U10232 ( .A1(n14407), .A2(n15239), .ZN(n11152) );
  INV_X1 U10233 ( .A(n6677), .ZN(n7944) );
  INV_X1 U10234 ( .A(n8500), .ZN(n7945) );
  NAND3_X1 U10235 ( .A1(n7945), .A2(n6680), .A3(n11152), .ZN(n7946) );
  AND2_X1 U10236 ( .A1(n7947), .A2(n7946), .ZN(n7950) );
  NAND2_X1 U10237 ( .A1(n8496), .A2(n8498), .ZN(n7948) );
  NAND4_X1 U10238 ( .A1(n15201), .A2(n8442), .A3(n11152), .A4(n11151), .ZN(
        n7949) );
  NAND4_X1 U10239 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n7968)
         );
  NAND2_X1 U10240 ( .A1(n8461), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7958) );
  INV_X1 U10241 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7953) );
  OR2_X1 U10242 ( .A1(n8469), .A2(n7953), .ZN(n7957) );
  OAI21_X1 U10243 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7975), .ZN(n11158) );
  OR2_X1 U10244 ( .A1(n8430), .A2(n11158), .ZN(n7956) );
  INV_X1 U10245 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7954) );
  OR2_X1 U10246 ( .A1(n8198), .A2(n7954), .ZN(n7955) );
  NAND2_X1 U10247 ( .A1(n7959), .A2(n9392), .ZN(n7983) );
  NAND2_X1 U10248 ( .A1(n7983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7961) );
  INV_X1 U10249 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7960) );
  XNOR2_X1 U10250 ( .A(n7961), .B(n7960), .ZN(n14456) );
  INV_X1 U10251 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10538) );
  OR2_X1 U10252 ( .A1(n8458), .A2(n10538), .ZN(n7964) );
  MUX2_X1 U10253 ( .A(n14406), .B(n11203), .S(n8031), .Z(n7969) );
  NAND2_X1 U10254 ( .A1(n7968), .A2(n7969), .ZN(n7967) );
  MUX2_X1 U10255 ( .A(n14406), .B(n11203), .S(n8442), .Z(n7966) );
  NAND2_X1 U10256 ( .A1(n7967), .A2(n7966), .ZN(n7973) );
  INV_X1 U10257 ( .A(n7968), .ZN(n7971) );
  NAND2_X1 U10258 ( .A1(n7973), .A2(n7972), .ZN(n7990) );
  NAND2_X1 U10259 ( .A1(n8466), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7980) );
  INV_X1 U10260 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11215) );
  OR2_X1 U10261 ( .A1(n8469), .A2(n11215), .ZN(n7979) );
  INV_X1 U10262 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10593) );
  OR2_X1 U10263 ( .A1(n8468), .A2(n10593), .ZN(n7978) );
  AND2_X1 U10264 ( .A1(n7975), .A2(n7974), .ZN(n7976) );
  OR2_X1 U10265 ( .A1(n7976), .A2(n8001), .ZN(n11218) );
  OR2_X1 U10266 ( .A1(n8430), .A2(n11218), .ZN(n7977) );
  NAND4_X1 U10267 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n14405) );
  XNOR2_X1 U10268 ( .A(n7982), .B(n7981), .ZN(n10541) );
  NAND2_X1 U10269 ( .A1(n10541), .A2(n8484), .ZN(n7986) );
  NAND2_X1 U10270 ( .A1(n7994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7984) );
  XNOR2_X1 U10271 ( .A(n7984), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U10272 ( .A1(n8483), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8264), .B2(
        n10619), .ZN(n7985) );
  MUX2_X1 U10273 ( .A(n14405), .B(n11281), .S(n8442), .Z(n7989) );
  INV_X1 U10274 ( .A(n14405), .ZN(n7987) );
  MUX2_X1 U10275 ( .A(n11276), .B(n7987), .S(n8442), .Z(n7988) );
  AOI21_X1 U10276 ( .B1(n7990), .B2(n7989), .A(n7988), .ZN(n7991) );
  NAND2_X1 U10277 ( .A1(n10555), .A2(n8484), .ZN(n7999) );
  INV_X1 U10278 ( .A(n7994), .ZN(n7996) );
  INV_X1 U10279 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10280 ( .A1(n7996), .A2(n7995), .ZN(n8026) );
  NAND2_X1 U10281 ( .A1(n8026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7997) );
  XNOR2_X1 U10282 ( .A(n7997), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U10283 ( .A1(n8483), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8264), .B2(
        n10620), .ZN(n7998) );
  NAND2_X1 U10284 ( .A1(n8461), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8007) );
  INV_X1 U10285 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8000) );
  OR2_X1 U10286 ( .A1(n6973), .A2(n8000), .ZN(n8006) );
  OR2_X1 U10287 ( .A1(n8001), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U10288 ( .A1(n8017), .A2(n8002), .ZN(n11381) );
  OR2_X1 U10289 ( .A1(n8430), .A2(n11381), .ZN(n8005) );
  INV_X1 U10290 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8003) );
  OR2_X1 U10291 ( .A1(n8198), .A2(n8003), .ZN(n8004) );
  INV_X1 U10292 ( .A(n11279), .ZN(n14404) );
  MUX2_X1 U10293 ( .A(n11314), .B(n14404), .S(n8442), .Z(n8011) );
  NAND2_X1 U10294 ( .A1(n8010), .A2(n8011), .ZN(n8009) );
  MUX2_X1 U10295 ( .A(n11314), .B(n14404), .S(n6677), .Z(n8008) );
  NAND2_X1 U10296 ( .A1(n8009), .A2(n8008), .ZN(n8015) );
  INV_X1 U10297 ( .A(n8010), .ZN(n8013) );
  NAND2_X1 U10298 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  NAND2_X1 U10299 ( .A1(n8015), .A2(n8014), .ZN(n8035) );
  NAND2_X1 U10300 ( .A1(n8461), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8023) );
  INV_X1 U10301 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10621) );
  OR2_X1 U10302 ( .A1(n6973), .A2(n10621), .ZN(n8022) );
  NAND2_X1 U10303 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  NAND2_X1 U10304 ( .A1(n8039), .A2(n8018), .ZN(n11288) );
  OR2_X1 U10305 ( .A1(n6972), .A2(n11288), .ZN(n8021) );
  INV_X1 U10306 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8019) );
  OR2_X1 U10307 ( .A1(n8465), .A2(n8019), .ZN(n8020) );
  INV_X1 U10308 ( .A(n11518), .ZN(n14403) );
  NAND2_X1 U10309 ( .A1(n10564), .A2(n8484), .ZN(n8030) );
  INV_X1 U10310 ( .A(n8026), .ZN(n8028) );
  INV_X1 U10311 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U10312 ( .A1(n8028), .A2(n8027), .ZN(n8067) );
  NAND2_X1 U10313 ( .A1(n8067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8049) );
  XNOR2_X1 U10314 ( .A(n8049), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U10315 ( .A1(n8483), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8264), .B2(
        n10636), .ZN(n8029) );
  MUX2_X1 U10316 ( .A(n14403), .B(n15263), .S(n8442), .Z(n8034) );
  NAND2_X1 U10317 ( .A1(n8035), .A2(n8034), .ZN(n8033) );
  MUX2_X1 U10318 ( .A(n14403), .B(n15263), .S(n6677), .Z(n8032) );
  NAND2_X1 U10319 ( .A1(n8033), .A2(n8032), .ZN(n8037) );
  NAND2_X1 U10320 ( .A1(n7929), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8045) );
  INV_X1 U10321 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10637) );
  OR2_X1 U10322 ( .A1(n6970), .A2(n10637), .ZN(n8044) );
  NAND2_X1 U10323 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  NAND2_X1 U10324 ( .A1(n8058), .A2(n8040), .ZN(n11523) );
  OR2_X1 U10325 ( .A1(n6972), .A2(n11523), .ZN(n8043) );
  INV_X1 U10326 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8041) );
  OR2_X1 U10327 ( .A1(n8198), .A2(n8041), .ZN(n8042) );
  INV_X1 U10328 ( .A(n11709), .ZN(n14402) );
  XNOR2_X1 U10329 ( .A(n8047), .B(n8046), .ZN(n10571) );
  NAND2_X1 U10330 ( .A1(n10571), .A2(n8484), .ZN(n8053) );
  INV_X1 U10331 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10332 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U10333 ( .A1(n8050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8051) );
  XNOR2_X1 U10334 ( .A(n8051), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U10335 ( .A1(n8483), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8264), .B2(
        n10671), .ZN(n8052) );
  MUX2_X1 U10336 ( .A(n14402), .B(n11705), .S(n6677), .Z(n8056) );
  MUX2_X1 U10337 ( .A(n14402), .B(n11705), .S(n8442), .Z(n8054) );
  INV_X1 U10338 ( .A(n8056), .ZN(n8057) );
  NAND2_X1 U10339 ( .A1(n8466), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8064) );
  INV_X1 U10340 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11701) );
  OR2_X1 U10341 ( .A1(n6973), .A2(n11701), .ZN(n8063) );
  INV_X1 U10342 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10669) );
  OR2_X1 U10343 ( .A1(n6970), .A2(n10669), .ZN(n8062) );
  INV_X1 U10344 ( .A(n8078), .ZN(n8060) );
  NAND2_X1 U10345 ( .A1(n8058), .A2(n11950), .ZN(n8059) );
  NAND2_X1 U10346 ( .A1(n8060), .A2(n8059), .ZN(n11951) );
  OR2_X1 U10347 ( .A1(n6972), .A2(n11951), .ZN(n8061) );
  INV_X1 U10348 ( .A(n12020), .ZN(n14401) );
  XNOR2_X1 U10349 ( .A(n8066), .B(n8065), .ZN(n10575) );
  NAND2_X1 U10350 ( .A1(n10575), .A2(n8484), .ZN(n8071) );
  NAND2_X1 U10351 ( .A1(n8068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8069) );
  XNOR2_X1 U10352 ( .A(n8069), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U10353 ( .A1(n8483), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8264), .B2(
        n10731), .ZN(n8070) );
  MUX2_X1 U10354 ( .A(n14401), .B(n12030), .S(n8442), .Z(n8075) );
  MUX2_X1 U10355 ( .A(n14401), .B(n12030), .S(n6677), .Z(n8072) );
  NAND2_X1 U10356 ( .A1(n8461), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8084) );
  INV_X1 U10357 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8077) );
  OR2_X1 U10358 ( .A1(n6973), .A2(n8077), .ZN(n8083) );
  OR2_X1 U10359 ( .A1(n8078), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U10360 ( .A1(n8096), .A2(n8079), .ZN(n12025) );
  OR2_X1 U10361 ( .A1(n6972), .A2(n12025), .ZN(n8082) );
  INV_X1 U10362 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8080) );
  OR2_X1 U10363 ( .A1(n8198), .A2(n8080), .ZN(n8081) );
  INV_X1 U10364 ( .A(n15096), .ZN(n14400) );
  XNOR2_X1 U10365 ( .A(n8086), .B(n8085), .ZN(n10650) );
  NAND2_X1 U10366 ( .A1(n10650), .A2(n8484), .ZN(n8093) );
  NOR2_X1 U10367 ( .A1(n8087), .A2(n7784), .ZN(n8088) );
  MUX2_X1 U10368 ( .A(n7784), .B(n8088), .S(P1_IR_REG_10__SCAN_IN), .Z(n8091)
         );
  NAND2_X1 U10369 ( .A1(n8087), .A2(n8089), .ZN(n8130) );
  INV_X1 U10370 ( .A(n8130), .ZN(n8090) );
  NOR2_X1 U10371 ( .A1(n8091), .A2(n8090), .ZN(n10833) );
  AOI22_X1 U10372 ( .A1(n8483), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8264), 
        .B2(n10833), .ZN(n8092) );
  MUX2_X1 U10373 ( .A(n14400), .B(n15284), .S(n6677), .Z(n8095) );
  MUX2_X1 U10374 ( .A(n14400), .B(n15284), .S(n8442), .Z(n8094) );
  NAND2_X1 U10375 ( .A1(n8466), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10376 ( .A1(n8096), .A2(n15092), .ZN(n8097) );
  NAND2_X1 U10377 ( .A1(n8136), .A2(n8097), .ZN(n15118) );
  OR2_X1 U10378 ( .A1(n6972), .A2(n15118), .ZN(n8100) );
  INV_X1 U10379 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n15119) );
  OR2_X1 U10380 ( .A1(n6973), .A2(n15119), .ZN(n8099) );
  INV_X1 U10381 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10834) );
  OR2_X1 U10382 ( .A1(n6970), .A2(n10834), .ZN(n8098) );
  NAND4_X1 U10383 ( .A1(n8101), .A2(n8100), .A3(n8099), .A4(n8098), .ZN(n14985) );
  XNOR2_X1 U10384 ( .A(n8103), .B(n8102), .ZN(n10688) );
  NAND2_X1 U10385 ( .A1(n10688), .A2(n8484), .ZN(n8106) );
  NAND2_X1 U10386 ( .A1(n8130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8104) );
  XNOR2_X1 U10387 ( .A(n8104), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U10388 ( .A1(n8483), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8264), 
        .B2(n10949), .ZN(n8105) );
  MUX2_X1 U10389 ( .A(n14985), .B(n15122), .S(n7944), .Z(n8151) );
  NAND2_X1 U10390 ( .A1(n8152), .A2(n8151), .ZN(n8108) );
  MUX2_X1 U10391 ( .A(n14985), .B(n15122), .S(n6677), .Z(n8107) );
  NAND2_X1 U10392 ( .A1(n8108), .A2(n8107), .ZN(n8150) );
  NAND2_X1 U10393 ( .A1(n10938), .A2(n8484), .ZN(n8113) );
  NAND2_X1 U10394 ( .A1(n7885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8111) );
  XNOR2_X1 U10395 ( .A(n8111), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U10396 ( .A1(n8483), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8264), 
        .B2(n14475), .ZN(n8112) );
  NAND2_X1 U10397 ( .A1(n8466), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8119) );
  INV_X1 U10398 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12139) );
  OR2_X1 U10399 ( .A1(n6970), .A2(n12139), .ZN(n8118) );
  INV_X1 U10400 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12151) );
  OR2_X1 U10401 ( .A1(n6973), .A2(n12151), .ZN(n8117) );
  NAND2_X1 U10402 ( .A1(n8121), .A2(n8114), .ZN(n8115) );
  NAND2_X1 U10403 ( .A1(n8172), .A2(n8115), .ZN(n14271) );
  OR2_X1 U10404 ( .A1(n6972), .A2(n14271), .ZN(n8116) );
  NAND2_X1 U10405 ( .A1(n14921), .A2(n14560), .ZN(n14536) );
  NAND2_X1 U10406 ( .A1(n8461), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8126) );
  INV_X1 U10407 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12353) );
  OR2_X1 U10408 ( .A1(n6973), .A2(n12353), .ZN(n8125) );
  OR2_X1 U10409 ( .A1(n8137), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10410 ( .A1(n8121), .A2(n8120), .ZN(n12396) );
  OR2_X1 U10411 ( .A1(n6972), .A2(n12396), .ZN(n8124) );
  INV_X1 U10412 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8122) );
  OR2_X1 U10413 ( .A1(n8198), .A2(n8122), .ZN(n8123) );
  INV_X1 U10414 ( .A(n12412), .ZN(n14988) );
  XNOR2_X1 U10415 ( .A(n8127), .B(n10569), .ZN(n8128) );
  NAND2_X1 U10416 ( .A1(n10745), .A2(n8484), .ZN(n8133) );
  OAI21_X1 U10417 ( .B1(n8144), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8131) );
  XNOR2_X1 U10418 ( .A(n8131), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U10419 ( .A1(n8483), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8264), 
        .B2(n12141), .ZN(n8132) );
  MUX2_X1 U10420 ( .A(n14988), .B(n15130), .S(n8442), .Z(n8178) );
  NAND2_X1 U10421 ( .A1(n12412), .A2(n8442), .ZN(n8134) );
  OAI21_X1 U10422 ( .B1(n15130), .B2(n8442), .A(n8134), .ZN(n8179) );
  OR2_X1 U10423 ( .A1(n8178), .A2(n8179), .ZN(n8135) );
  AND3_X1 U10424 ( .A1(n14535), .A2(n14536), .A3(n8135), .ZN(n8153) );
  NAND2_X1 U10425 ( .A1(n8466), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8142) );
  AND2_X1 U10426 ( .A1(n8136), .A2(n10953), .ZN(n8138) );
  OR2_X1 U10427 ( .A1(n8138), .A2(n8137), .ZN(n15091) );
  OR2_X1 U10428 ( .A1(n6972), .A2(n15091), .ZN(n8141) );
  INV_X1 U10429 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n14981) );
  OR2_X1 U10430 ( .A1(n6973), .A2(n14981), .ZN(n8140) );
  INV_X1 U10431 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10947) );
  OR2_X1 U10432 ( .A1(n6970), .A2(n10947), .ZN(n8139) );
  NAND4_X1 U10433 ( .A1(n8142), .A2(n8141), .A3(n8140), .A4(n8139), .ZN(n14399) );
  INV_X1 U10434 ( .A(n14399), .ZN(n15098) );
  XNOR2_X1 U10435 ( .A(n8143), .B(n7746), .ZN(n10720) );
  NAND2_X1 U10436 ( .A1(n10720), .A2(n8484), .ZN(n8147) );
  NAND2_X1 U10437 ( .A1(n8144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8145) );
  XNOR2_X1 U10438 ( .A(n8145), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U10439 ( .A1(n8483), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8264), 
        .B2(n11093), .ZN(n8146) );
  INV_X1 U10440 ( .A(n15087), .ZN(n14998) );
  MUX2_X1 U10441 ( .A(n15098), .B(n14998), .S(n8442), .Z(n8155) );
  MUX2_X1 U10442 ( .A(n14399), .B(n15087), .S(n6677), .Z(n8154) );
  NAND2_X1 U10443 ( .A1(n8155), .A2(n8154), .ZN(n8148) );
  AND2_X1 U10444 ( .A1(n8153), .A2(n8148), .ZN(n8149) );
  INV_X1 U10445 ( .A(n8153), .ZN(n8184) );
  INV_X1 U10446 ( .A(n8154), .ZN(n8157) );
  INV_X1 U10447 ( .A(n8155), .ZN(n8156) );
  NAND2_X1 U10448 ( .A1(n8157), .A2(n8156), .ZN(n8183) );
  INV_X1 U10449 ( .A(n8158), .ZN(n8160) );
  NAND2_X1 U10450 ( .A1(n8160), .A2(n8159), .ZN(n8162) );
  NAND2_X1 U10451 ( .A1(n8109), .A2(n10577), .ZN(n8161) );
  NAND2_X1 U10452 ( .A1(n8162), .A2(n8161), .ZN(n8165) );
  XNOR2_X1 U10453 ( .A(n8163), .B(SI_15_), .ZN(n8164) );
  NAND2_X1 U10454 ( .A1(n11015), .A2(n8484), .ZN(n8169) );
  NAND2_X1 U10455 ( .A1(n8166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8167) );
  XNOR2_X1 U10456 ( .A(n8167), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U10457 ( .A1(n8483), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8264), 
        .B2(n12153), .ZN(n8168) );
  NAND2_X2 U10458 ( .A1(n8169), .A2(n8168), .ZN(n14911) );
  NAND2_X1 U10459 ( .A1(n8466), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8177) );
  INV_X1 U10460 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8170) );
  OR2_X1 U10461 ( .A1(n6973), .A2(n8170), .ZN(n8176) );
  INV_X1 U10462 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15186) );
  OR2_X1 U10463 ( .A1(n6970), .A2(n15186), .ZN(n8175) );
  AND2_X1 U10464 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  OR2_X1 U10465 ( .A1(n8173), .A2(n8195), .ZN(n14792) );
  OR2_X1 U10466 ( .A1(n6972), .A2(n14792), .ZN(n8174) );
  NAND2_X1 U10467 ( .A1(n14535), .A2(n14536), .ZN(n12410) );
  INV_X1 U10468 ( .A(n8178), .ZN(n8181) );
  INV_X1 U10469 ( .A(n8179), .ZN(n8180) );
  OR3_X1 U10470 ( .A1(n12410), .A2(n8181), .A3(n8180), .ZN(n8182) );
  OAI211_X1 U10471 ( .C1(n8184), .C2(n8183), .A(n14539), .B(n8182), .ZN(n8190)
         );
  NOR2_X1 U10472 ( .A1(n14560), .A2(n7944), .ZN(n8187) );
  NAND2_X1 U10473 ( .A1(n14560), .A2(n7944), .ZN(n8185) );
  NAND2_X1 U10474 ( .A1(n14921), .A2(n8185), .ZN(n8186) );
  OAI21_X1 U10475 ( .B1(n14921), .B2(n8187), .A(n8186), .ZN(n8188) );
  NAND2_X1 U10476 ( .A1(n14911), .A2(n14562), .ZN(n8493) );
  MUX2_X1 U10477 ( .A(n8493), .B(n14539), .S(n7944), .Z(n8193) );
  NAND2_X1 U10478 ( .A1(n8461), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8202) );
  INV_X1 U10479 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8194) );
  OR2_X1 U10480 ( .A1(n6973), .A2(n8194), .ZN(n8201) );
  NOR2_X1 U10481 ( .A1(n8195), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8196) );
  OR2_X1 U10482 ( .A1(n8209), .A2(n8196), .ZN(n14777) );
  OR2_X1 U10483 ( .A1(n6972), .A2(n14777), .ZN(n8200) );
  INV_X1 U10484 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8197) );
  OR2_X1 U10485 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  NAND4_X1 U10486 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8199), .ZN(n14564) );
  XNOR2_X1 U10487 ( .A(n8204), .B(n8203), .ZN(n10880) );
  NAND2_X1 U10488 ( .A1(n10880), .A2(n8484), .ZN(n8208) );
  OR2_X1 U10489 ( .A1(n8205), .A2(n7784), .ZN(n8206) );
  XNOR2_X1 U10490 ( .A(n8206), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U10491 ( .A1(n8483), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8264), 
        .B2(n12376), .ZN(n8207) );
  MUX2_X1 U10492 ( .A(n14564), .B(n14905), .S(n6677), .Z(n8242) );
  OR2_X1 U10493 ( .A1(n8209), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U10494 ( .A1(n8269), .A2(n8210), .ZN(n14763) );
  OR2_X1 U10495 ( .A1(n6972), .A2(n14763), .ZN(n8216) );
  INV_X1 U10496 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8211) );
  OR2_X1 U10497 ( .A1(n6970), .A2(n8211), .ZN(n8215) );
  INV_X1 U10498 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14767) );
  OR2_X1 U10499 ( .A1(n6973), .A2(n14767), .ZN(n8214) );
  INV_X1 U10500 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8212) );
  OR2_X1 U10501 ( .A1(n8465), .A2(n8212), .ZN(n8213) );
  NAND4_X1 U10502 ( .A1(n8216), .A2(n8215), .A3(n8214), .A4(n8213), .ZN(n14565) );
  NOR2_X1 U10503 ( .A1(n14564), .A2(n7944), .ZN(n8231) );
  AOI21_X1 U10504 ( .B1(n8242), .B2(n14565), .A(n8231), .ZN(n8229) );
  XNOR2_X1 U10505 ( .A(n8217), .B(SI_17_), .ZN(n8218) );
  XNOR2_X1 U10506 ( .A(n8219), .B(n8218), .ZN(n10958) );
  NAND2_X1 U10507 ( .A1(n10958), .A2(n8484), .ZN(n8223) );
  OR2_X1 U10508 ( .A1(n8220), .A2(n7784), .ZN(n8221) );
  XNOR2_X1 U10509 ( .A(n8221), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U10510 ( .A1(n8483), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8264), 
        .B2(n14494), .ZN(n8222) );
  NAND2_X1 U10511 ( .A1(n14565), .A2(n8442), .ZN(n8239) );
  OR2_X1 U10512 ( .A1(n14905), .A2(n8239), .ZN(n8225) );
  NOR2_X1 U10513 ( .A1(n14565), .A2(n8442), .ZN(n8232) );
  INV_X1 U10514 ( .A(n14564), .ZN(n14541) );
  NAND2_X1 U10515 ( .A1(n8232), .A2(n14541), .ZN(n8224) );
  AND2_X1 U10516 ( .A1(n8225), .A2(n8224), .ZN(n8235) );
  INV_X1 U10517 ( .A(n14565), .ZN(n14566) );
  NAND2_X1 U10518 ( .A1(n8242), .A2(n14566), .ZN(n8226) );
  OR2_X1 U10519 ( .A1(n14905), .A2(n6677), .ZN(n8238) );
  NAND2_X1 U10520 ( .A1(n8226), .A2(n8238), .ZN(n8227) );
  NAND2_X1 U10521 ( .A1(n8227), .A2(n8244), .ZN(n8228) );
  OAI211_X1 U10522 ( .C1(n8229), .C2(n8244), .A(n8235), .B(n8228), .ZN(n8230)
         );
  NAND2_X1 U10523 ( .A1(n8242), .A2(n8231), .ZN(n8234) );
  INV_X1 U10524 ( .A(n8232), .ZN(n8233) );
  NAND2_X1 U10525 ( .A1(n8234), .A2(n8233), .ZN(n8237) );
  INV_X1 U10526 ( .A(n8235), .ZN(n8236) );
  AOI22_X1 U10527 ( .A1(n8237), .A2(n14899), .B1(n8242), .B2(n8236), .ZN(n8247) );
  INV_X1 U10528 ( .A(n8238), .ZN(n8241) );
  INV_X1 U10529 ( .A(n8239), .ZN(n8240) );
  AOI21_X1 U10530 ( .B1(n8242), .B2(n8241), .A(n8240), .ZN(n8243) );
  INV_X1 U10531 ( .A(n8243), .ZN(n8245) );
  NAND2_X1 U10532 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  XNOR2_X1 U10533 ( .A(n8250), .B(n8249), .ZN(n11132) );
  NAND2_X1 U10534 ( .A1(n11132), .A2(n8484), .ZN(n8253) );
  NAND2_X1 U10535 ( .A1(n6829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8251) );
  XNOR2_X1 U10536 ( .A(n8251), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14508) );
  AOI22_X1 U10537 ( .A1(n8483), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8264), 
        .B2(n14508), .ZN(n8252) );
  XNOR2_X1 U10538 ( .A(n8269), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U10539 ( .A1(n14749), .A2(n8293), .ZN(n8258) );
  NAND2_X1 U10540 ( .A1(n8466), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8257) );
  INV_X1 U10541 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14496) );
  OR2_X1 U10542 ( .A1(n6970), .A2(n14496), .ZN(n8256) );
  INV_X1 U10543 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8254) );
  OR2_X1 U10544 ( .A1(n6973), .A2(n8254), .ZN(n8255) );
  NAND4_X1 U10545 ( .A1(n8258), .A2(n8257), .A3(n8256), .A4(n8255), .ZN(n14398) );
  OR2_X1 U10546 ( .A1(n14893), .A2(n14398), .ZN(n14568) );
  INV_X1 U10547 ( .A(n14398), .ZN(n14542) );
  MUX2_X1 U10548 ( .A(n14542), .B(n14751), .S(n7944), .Z(n8259) );
  AND2_X1 U10549 ( .A1(n14893), .A2(n14398), .ZN(n14569) );
  NAND2_X1 U10550 ( .A1(n8260), .A2(n14569), .ZN(n8275) );
  XNOR2_X1 U10551 ( .A(n8262), .B(n8261), .ZN(n11299) );
  NAND2_X1 U10552 ( .A1(n11299), .A2(n8484), .ZN(n8266) );
  AOI22_X1 U10553 ( .A1(n8483), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8264), 
        .B2(n6681), .ZN(n8265) );
  INV_X1 U10554 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8268) );
  INV_X1 U10555 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8267) );
  OAI21_X1 U10556 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8270) );
  NAND2_X1 U10557 ( .A1(n8270), .A2(n8280), .ZN(n14738) );
  OR2_X1 U10558 ( .A1(n14738), .A2(n6972), .ZN(n8274) );
  NAND2_X1 U10559 ( .A1(n7929), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10560 ( .A1(n8466), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10561 ( .A1(n8461), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8271) );
  OR2_X1 U10562 ( .A1(n14888), .A2(n14570), .ZN(n8277) );
  NAND2_X1 U10563 ( .A1(n14888), .A2(n14570), .ZN(n14543) );
  NAND2_X1 U10564 ( .A1(n8277), .A2(n14543), .ZN(n14732) );
  NAND3_X1 U10565 ( .A1(n8276), .A2(n8275), .A3(n7726), .ZN(n8279) );
  MUX2_X1 U10566 ( .A(n14543), .B(n8277), .S(n6677), .Z(n8278) );
  NAND2_X1 U10567 ( .A1(n8279), .A2(n8278), .ZN(n8289) );
  NAND2_X1 U10568 ( .A1(n8280), .A2(n14346), .ZN(n8281) );
  NAND2_X1 U10569 ( .A1(n8292), .A2(n8281), .ZN(n14722) );
  NAND2_X1 U10570 ( .A1(n8461), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10571 ( .A1(n7929), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8282) );
  AND2_X1 U10572 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  NAND2_X1 U10573 ( .A1(n8466), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8284) );
  OAI211_X1 U10574 ( .C1(n14722), .C2(n6972), .A(n8285), .B(n8284), .ZN(n14396) );
  XNOR2_X1 U10575 ( .A(n8298), .B(n11085), .ZN(n8297) );
  XNOR2_X1 U10576 ( .A(n8297), .B(n8300), .ZN(n11884) );
  INV_X1 U10577 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11886) );
  OR2_X1 U10578 ( .A1(n8458), .A2(n11886), .ZN(n8286) );
  MUX2_X1 U10579 ( .A(n14396), .B(n14883), .S(n7944), .Z(n8287) );
  OAI21_X1 U10580 ( .B1(n8289), .B2(n8288), .A(n8287), .ZN(n8291) );
  NAND2_X1 U10581 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  INV_X1 U10582 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8296) );
  NOR2_X1 U10583 ( .A1(n8310), .A2(n7756), .ZN(n14298) );
  NAND2_X1 U10584 ( .A1(n14298), .A2(n8293), .ZN(n8295) );
  AOI22_X1 U10585 ( .A1(n8461), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n7929), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n8294) );
  OAI211_X1 U10586 ( .C1(n8465), .C2(n8296), .A(n8295), .B(n8294), .ZN(n14573)
         );
  INV_X1 U10587 ( .A(n14573), .ZN(n14546) );
  INV_X1 U10588 ( .A(n8297), .ZN(n8301) );
  NOR2_X1 U10589 ( .A1(n8298), .A2(n11085), .ZN(n8299) );
  XNOR2_X1 U10590 ( .A(n8302), .B(SI_21_), .ZN(n8303) );
  XNOR2_X1 U10591 ( .A(n8304), .B(n8303), .ZN(n12016) );
  NAND2_X1 U10592 ( .A1(n12016), .A2(n8484), .ZN(n8306) );
  OR2_X1 U10593 ( .A1(n8458), .A2(n7203), .ZN(n8305) );
  INV_X1 U10594 ( .A(n14877), .ZN(n14303) );
  MUX2_X1 U10595 ( .A(n14546), .B(n14303), .S(n7944), .Z(n8309) );
  INV_X1 U10596 ( .A(n8309), .ZN(n8307) );
  MUX2_X1 U10597 ( .A(n14573), .B(n14877), .S(n6677), .Z(n8308) );
  NOR2_X1 U10598 ( .A1(n8310), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8311) );
  OR2_X1 U10599 ( .A1(n8312), .A2(n8311), .ZN(n14690) );
  INV_X1 U10600 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10601 ( .A1(n8461), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10602 ( .A1(n7929), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8313) );
  OAI211_X1 U10603 ( .C1(n8315), .C2(n8465), .A(n8314), .B(n8313), .ZN(n8316)
         );
  INV_X1 U10604 ( .A(n8316), .ZN(n8317) );
  OAI21_X1 U10605 ( .B1(n14690), .B2(n6972), .A(n8317), .ZN(n14548) );
  INV_X1 U10606 ( .A(n14692), .ZN(n14872) );
  MUX2_X1 U10607 ( .A(n14548), .B(n14872), .S(n6677), .Z(n8320) );
  INV_X1 U10608 ( .A(n14548), .ZN(n14575) );
  MUX2_X1 U10609 ( .A(n14575), .B(n14692), .S(n7944), .Z(n8319) );
  MUX2_X1 U10610 ( .A(n14395), .B(n14866), .S(n6677), .Z(n8321) );
  NAND2_X1 U10611 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  OAI21_X1 U10612 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(n8347) );
  NAND2_X1 U10613 ( .A1(n7929), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8333) );
  INV_X1 U10614 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8326) );
  OR2_X1 U10615 ( .A1(n8465), .A2(n8326), .ZN(n8332) );
  OAI21_X1 U10616 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8328), .A(n8353), .ZN(
        n14663) );
  OR2_X1 U10617 ( .A1(n6972), .A2(n14663), .ZN(n8331) );
  INV_X1 U10618 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8329) );
  OR2_X1 U10619 ( .A1(n6970), .A2(n8329), .ZN(n8330) );
  NAND4_X1 U10620 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .ZN(n14577) );
  INV_X1 U10621 ( .A(n9003), .ZN(n8337) );
  INV_X1 U10622 ( .A(n8339), .ZN(n8334) );
  AOI22_X1 U10623 ( .A1(n11185), .A2(n8337), .B1(n8334), .B2(n11511), .ZN(
        n8335) );
  OAI21_X1 U10624 ( .B1(n8337), .B2(n11185), .A(n11511), .ZN(n8340) );
  AND2_X1 U10625 ( .A1(SI_23_), .A2(SI_22_), .ZN(n8338) );
  AOI22_X1 U10626 ( .A1(n8340), .A2(n8339), .B1(n9003), .B2(n8338), .ZN(n8341)
         );
  MUX2_X1 U10627 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n10497), .Z(n8361) );
  XNOR2_X1 U10628 ( .A(n8360), .B(n8361), .ZN(n12206) );
  NAND2_X1 U10629 ( .A1(n12206), .A2(n8484), .ZN(n8344) );
  INV_X1 U10630 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12209) );
  OR2_X1 U10631 ( .A1(n8458), .A2(n12209), .ZN(n8343) );
  MUX2_X1 U10632 ( .A(n14577), .B(n14857), .S(n6677), .Z(n8348) );
  NAND2_X1 U10633 ( .A1(n8347), .A2(n8348), .ZN(n8346) );
  MUX2_X1 U10634 ( .A(n14577), .B(n14857), .S(n7944), .Z(n8345) );
  NAND2_X1 U10635 ( .A1(n8346), .A2(n8345), .ZN(n8352) );
  INV_X1 U10636 ( .A(n8347), .ZN(n8350) );
  INV_X1 U10637 ( .A(n8348), .ZN(n8349) );
  NAND2_X1 U10638 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  NAND2_X1 U10639 ( .A1(n8461), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8359) );
  INV_X1 U10640 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14645) );
  OR2_X1 U10641 ( .A1(n6973), .A2(n14645), .ZN(n8358) );
  NAND2_X1 U10642 ( .A1(n8354), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8373) );
  OAI21_X1 U10643 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8354), .A(n8373), .ZN(
        n14644) );
  OR2_X1 U10644 ( .A1(n6972), .A2(n14644), .ZN(n8357) );
  INV_X1 U10645 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8355) );
  OR2_X1 U10646 ( .A1(n8465), .A2(n8355), .ZN(n8356) );
  INV_X1 U10647 ( .A(n14579), .ZN(n14394) );
  NAND2_X1 U10648 ( .A1(n8363), .A2(SI_24_), .ZN(n8364) );
  MUX2_X1 U10649 ( .A(n12332), .B(n12329), .S(n10497), .Z(n8365) );
  NAND2_X1 U10650 ( .A1(n8365), .A2(n12277), .ZN(n8382) );
  INV_X1 U10651 ( .A(n8365), .ZN(n8366) );
  NAND2_X1 U10652 ( .A1(n8366), .A2(SI_25_), .ZN(n8367) );
  NAND2_X1 U10653 ( .A1(n8382), .A2(n8367), .ZN(n8380) );
  XNOR2_X1 U10654 ( .A(n8381), .B(n8380), .ZN(n12327) );
  NAND2_X1 U10655 ( .A1(n12327), .A2(n8484), .ZN(n8369) );
  OR2_X1 U10656 ( .A1(n8458), .A2(n12329), .ZN(n8368) );
  MUX2_X1 U10657 ( .A(n14394), .B(n14647), .S(n7944), .Z(n8371) );
  MUX2_X1 U10658 ( .A(n14394), .B(n14647), .S(n6677), .Z(n8370) );
  NAND2_X1 U10659 ( .A1(n7929), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8379) );
  INV_X1 U10660 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8372) );
  OR2_X1 U10661 ( .A1(n8465), .A2(n8372), .ZN(n8378) );
  INV_X1 U10662 ( .A(n8373), .ZN(n8374) );
  NAND2_X1 U10663 ( .A1(n8374), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8388) );
  OAI21_X1 U10664 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n8374), .A(n8388), .ZN(
        n14633) );
  OR2_X1 U10665 ( .A1(n6972), .A2(n14633), .ZN(n8377) );
  INV_X1 U10666 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8375) );
  OR2_X1 U10667 ( .A1(n6970), .A2(n8375), .ZN(n8376) );
  INV_X1 U10668 ( .A(n14309), .ZN(n14580) );
  MUX2_X1 U10669 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n10497), .Z(n8395) );
  INV_X1 U10670 ( .A(SI_26_), .ZN(n13670) );
  XNOR2_X1 U10671 ( .A(n8395), .B(n13670), .ZN(n8383) );
  NAND2_X1 U10672 ( .A1(n14251), .A2(n8484), .ZN(n8385) );
  INV_X1 U10673 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14950) );
  OR2_X1 U10674 ( .A1(n8458), .A2(n14950), .ZN(n8384) );
  MUX2_X1 U10675 ( .A(n14580), .B(n14843), .S(n6677), .Z(n8387) );
  MUX2_X1 U10676 ( .A(n14580), .B(n14843), .S(n7944), .Z(n8386) );
  NAND2_X1 U10677 ( .A1(n8461), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8394) );
  INV_X1 U10678 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14621) );
  OR2_X1 U10679 ( .A1(n6973), .A2(n14621), .ZN(n8393) );
  INV_X1 U10680 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U10681 ( .A1(n8389), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8406) );
  OAI21_X1 U10682 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n8389), .A(n8406), .ZN(
        n14620) );
  OR2_X1 U10683 ( .A1(n6972), .A2(n14620), .ZN(n8392) );
  INV_X1 U10684 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10685 ( .A1(n8465), .A2(n8390), .ZN(n8391) );
  INV_X1 U10686 ( .A(n14550), .ZN(n14582) );
  INV_X1 U10687 ( .A(n8395), .ZN(n8396) );
  MUX2_X1 U10688 ( .A(n14250), .B(n7617), .S(n10502), .Z(n8413) );
  XNOR2_X1 U10689 ( .A(n8413), .B(SI_27_), .ZN(n8400) );
  NAND2_X1 U10690 ( .A1(n14945), .A2(n8484), .ZN(n8402) );
  OR2_X1 U10691 ( .A1(n8458), .A2(n7617), .ZN(n8401) );
  MUX2_X1 U10692 ( .A(n14582), .B(n14837), .S(n7944), .Z(n8404) );
  MUX2_X1 U10693 ( .A(n14582), .B(n14837), .S(n6677), .Z(n8403) );
  NAND2_X1 U10694 ( .A1(n8461), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8412) );
  INV_X1 U10695 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8405) );
  OR2_X1 U10696 ( .A1(n6973), .A2(n8405), .ZN(n8411) );
  INV_X1 U10697 ( .A(n8406), .ZN(n8407) );
  NAND2_X1 U10698 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n8407), .ZN(n14588) );
  OAI21_X1 U10699 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n8407), .A(n14588), .ZN(
        n14606) );
  OR2_X1 U10700 ( .A1(n6972), .A2(n14606), .ZN(n8410) );
  INV_X1 U10701 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8408) );
  OR2_X1 U10702 ( .A1(n8465), .A2(n8408), .ZN(n8409) );
  NAND4_X1 U10703 ( .A1(n8412), .A2(n8411), .A3(n8410), .A4(n8409), .ZN(n14557) );
  INV_X1 U10704 ( .A(n8413), .ZN(n8416) );
  NOR2_X1 U10705 ( .A1(n8416), .A2(SI_27_), .ZN(n8414) );
  NAND2_X1 U10706 ( .A1(n8416), .A2(SI_27_), .ZN(n8417) );
  INV_X1 U10707 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14245) );
  INV_X1 U10708 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12605) );
  MUX2_X1 U10709 ( .A(n14245), .B(n12605), .S(n10497), .Z(n8418) );
  INV_X1 U10710 ( .A(SI_28_), .ZN(n12560) );
  NAND2_X1 U10711 ( .A1(n8418), .A2(n12560), .ZN(n8438) );
  INV_X1 U10712 ( .A(n8418), .ZN(n8419) );
  NAND2_X1 U10713 ( .A1(n8419), .A2(SI_28_), .ZN(n8420) );
  NAND2_X1 U10714 ( .A1(n8438), .A2(n8420), .ZN(n8436) );
  NAND2_X1 U10715 ( .A1(n14242), .A2(n8484), .ZN(n8422) );
  OR2_X1 U10716 ( .A1(n8458), .A2(n12605), .ZN(n8421) );
  NAND2_X2 U10717 ( .A1(n8422), .A2(n8421), .ZN(n14830) );
  MUX2_X1 U10718 ( .A(n14557), .B(n14830), .S(n6677), .Z(n8425) );
  INV_X1 U10719 ( .A(n14557), .ZN(n14551) );
  MUX2_X1 U10720 ( .A(n14551), .B(n14610), .S(n7944), .Z(n8423) );
  INV_X1 U10721 ( .A(n8423), .ZN(n8428) );
  INV_X1 U10722 ( .A(n8424), .ZN(n8427) );
  INV_X1 U10723 ( .A(n8425), .ZN(n8426) );
  NAND2_X1 U10724 ( .A1(n8461), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10725 ( .A1(n7929), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8434) );
  OR2_X1 U10726 ( .A1(n6972), .A2(n14588), .ZN(n8433) );
  INV_X1 U10727 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8431) );
  OR2_X1 U10728 ( .A1(n8465), .A2(n8431), .ZN(n8432) );
  NAND4_X1 U10729 ( .A1(n8435), .A2(n8434), .A3(n8433), .A4(n8432), .ZN(n14393) );
  MUX2_X1 U10730 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n10502), .Z(n8449) );
  INV_X1 U10731 ( .A(SI_29_), .ZN(n12643) );
  XNOR2_X1 U10732 ( .A(n8449), .B(n12643), .ZN(n8447) );
  NAND2_X1 U10733 ( .A1(n14239), .A2(n8484), .ZN(n8441) );
  INV_X1 U10734 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14944) );
  OR2_X1 U10735 ( .A1(n8458), .A2(n14944), .ZN(n8440) );
  MUX2_X1 U10736 ( .A(n14393), .B(n14822), .S(n7944), .Z(n8443) );
  MUX2_X1 U10737 ( .A(n14393), .B(n14822), .S(n6677), .Z(n8446) );
  INV_X1 U10738 ( .A(n8443), .ZN(n8444) );
  INV_X1 U10739 ( .A(n8449), .ZN(n8450) );
  NAND2_X1 U10740 ( .A1(n8450), .A2(n12643), .ZN(n8451) );
  MUX2_X1 U10741 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n10497), .Z(n8453) );
  NAND2_X1 U10742 ( .A1(n8453), .A2(SI_30_), .ZN(n8479) );
  OAI21_X1 U10743 ( .B1(SI_30_), .B2(n8453), .A(n8479), .ZN(n8454) );
  NAND2_X1 U10744 ( .A1(n8455), .A2(n8454), .ZN(n8456) );
  INV_X1 U10745 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12639) );
  OR2_X1 U10746 ( .A1(n8458), .A2(n12639), .ZN(n8459) );
  INV_X1 U10747 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10748 ( .A1(n7929), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10749 ( .A1(n8461), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8462) );
  OAI211_X1 U10750 ( .C1(n8465), .C2(n8464), .A(n8463), .B(n8462), .ZN(n14820)
         );
  NAND2_X1 U10751 ( .A1(n8466), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8472) );
  INV_X1 U10752 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8467) );
  OR2_X1 U10753 ( .A1(n6970), .A2(n8467), .ZN(n8471) );
  INV_X1 U10754 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14526) );
  OR2_X1 U10755 ( .A1(n6973), .A2(n14526), .ZN(n8470) );
  AND3_X1 U10756 ( .A1(n8472), .A2(n8471), .A3(n8470), .ZN(n14525) );
  INV_X1 U10757 ( .A(n8473), .ZN(n8474) );
  OAI22_X1 U10758 ( .A1(n14525), .A2(n6677), .B1(n10703), .B2(n8474), .ZN(
        n8475) );
  AOI22_X1 U10759 ( .A1(n14533), .A2(n6677), .B1(n14820), .B2(n8475), .ZN(
        n8477) );
  INV_X1 U10760 ( .A(n14525), .ZN(n10583) );
  NAND2_X1 U10761 ( .A1(n10703), .A2(n8486), .ZN(n8543) );
  OAI21_X1 U10762 ( .B1(n10583), .B2(n8543), .A(n14820), .ZN(n8476) );
  MUX2_X1 U10763 ( .A(n14818), .B(n8476), .S(n6677), .Z(n8478) );
  MUX2_X1 U10764 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10502), .Z(n8481) );
  XNOR2_X1 U10765 ( .A(n8481), .B(SI_31_), .ZN(n8482) );
  NAND2_X1 U10766 ( .A1(n10583), .A2(n6677), .ZN(n8525) );
  INV_X1 U10767 ( .A(n8525), .ZN(n8488) );
  NAND2_X1 U10768 ( .A1(n6681), .A2(n6679), .ZN(n11202) );
  OR2_X1 U10769 ( .A1(n10560), .A2(n10702), .ZN(n8485) );
  NAND2_X1 U10770 ( .A1(n11202), .A2(n8485), .ZN(n8534) );
  INV_X1 U10771 ( .A(n10703), .ZN(n12018) );
  AND2_X1 U10772 ( .A1(n12018), .A2(n8486), .ZN(n10480) );
  INV_X1 U10773 ( .A(n10480), .ZN(n8487) );
  NAND2_X1 U10774 ( .A1(n8534), .A2(n8487), .ZN(n8523) );
  AOI21_X1 U10775 ( .B1(n14522), .B2(n8488), .A(n8523), .ZN(n8491) );
  OR2_X1 U10776 ( .A1(n10583), .A2(n6677), .ZN(n8521) );
  INV_X1 U10777 ( .A(n8521), .ZN(n8489) );
  NAND2_X1 U10778 ( .A1(n7262), .A2(n8489), .ZN(n8490) );
  XNOR2_X1 U10779 ( .A(n14522), .B(n10583), .ZN(n8535) );
  INV_X1 U10780 ( .A(n8535), .ZN(n8519) );
  XOR2_X1 U10781 ( .A(n14820), .B(n14533), .Z(n8517) );
  NAND2_X1 U10782 ( .A1(n14830), .A2(n14557), .ZN(n14584) );
  OR2_X1 U10783 ( .A1(n14830), .A2(n14557), .ZN(n8492) );
  XNOR2_X1 U10784 ( .A(n14866), .B(n14576), .ZN(n14672) );
  INV_X1 U10785 ( .A(n14672), .ZN(n14549) );
  XNOR2_X1 U10786 ( .A(n14877), .B(n14573), .ZN(n14702) );
  XNOR2_X1 U10787 ( .A(n14905), .B(n14564), .ZN(n14781) );
  NOR2_X1 U10788 ( .A1(n15122), .A2(n14985), .ZN(n12351) );
  NAND2_X1 U10789 ( .A1(n15122), .A2(n14985), .ZN(n12352) );
  INV_X1 U10790 ( .A(n12352), .ZN(n8494) );
  OR2_X1 U10791 ( .A1(n12351), .A2(n8494), .ZN(n15112) );
  XNOR2_X1 U10792 ( .A(n15263), .B(n11518), .ZN(n11285) );
  INV_X1 U10793 ( .A(n11285), .ZN(n8504) );
  NAND2_X1 U10794 ( .A1(n8498), .A2(n8497), .ZN(n14803) );
  NOR2_X1 U10795 ( .A1(n11143), .A2(n14803), .ZN(n8501) );
  NAND2_X1 U10796 ( .A1(n11152), .A2(n8499), .ZN(n11148) );
  INV_X1 U10797 ( .A(n11148), .ZN(n11175) );
  INV_X1 U10798 ( .A(n15200), .ZN(n15202) );
  XNOR2_X1 U10799 ( .A(n14406), .B(n11203), .ZN(n11154) );
  NAND4_X1 U10800 ( .A1(n8501), .A2(n11175), .A3(n15202), .A4(n11154), .ZN(
        n8502) );
  XNOR2_X1 U10801 ( .A(n11276), .B(n14405), .ZN(n11208) );
  NOR2_X1 U10802 ( .A1(n8502), .A2(n11208), .ZN(n8503) );
  XNOR2_X1 U10803 ( .A(n11314), .B(n11279), .ZN(n11300) );
  INV_X1 U10804 ( .A(n11300), .ZN(n11305) );
  NAND3_X1 U10805 ( .A1(n8504), .A2(n8503), .A3(n11305), .ZN(n8505) );
  XNOR2_X1 U10806 ( .A(n11705), .B(n11709), .ZN(n11704) );
  NOR2_X1 U10807 ( .A1(n8505), .A2(n11704), .ZN(n8506) );
  XNOR2_X1 U10808 ( .A(n15284), .B(n15096), .ZN(n12033) );
  INV_X1 U10809 ( .A(n12033), .ZN(n12022) );
  XNOR2_X1 U10810 ( .A(n12030), .B(n12020), .ZN(n11699) );
  INV_X1 U10811 ( .A(n11699), .ZN(n11706) );
  AND4_X1 U10812 ( .A1(n15112), .A2(n8506), .A3(n12022), .A4(n11706), .ZN(
        n8507) );
  XNOR2_X1 U10813 ( .A(n15130), .B(n12412), .ZN(n12401) );
  INV_X1 U10814 ( .A(n12401), .ZN(n12406) );
  XNOR2_X1 U10815 ( .A(n15087), .B(n14399), .ZN(n14983) );
  NAND4_X1 U10816 ( .A1(n14781), .A2(n8507), .A3(n12406), .A4(n14983), .ZN(
        n8508) );
  NOR2_X1 U10817 ( .A1(n8508), .A2(n12410), .ZN(n8509) );
  XNOR2_X1 U10818 ( .A(n14899), .B(n14565), .ZN(n14770) );
  NAND3_X1 U10819 ( .A1(n14787), .A2(n8509), .A3(n14770), .ZN(n8510) );
  NOR2_X1 U10820 ( .A1(n14732), .A2(n8510), .ZN(n8512) );
  XNOR2_X1 U10821 ( .A(n14883), .B(n14571), .ZN(n14726) );
  INV_X1 U10822 ( .A(n14726), .ZN(n14544) );
  XNOR2_X1 U10823 ( .A(n14893), .B(n14542), .ZN(n14754) );
  INV_X1 U10824 ( .A(n14754), .ZN(n8511) );
  NAND4_X1 U10825 ( .A1(n14702), .A2(n8512), .A3(n14544), .A4(n8511), .ZN(
        n8513) );
  NOR2_X1 U10826 ( .A1(n8513), .A2(n14685), .ZN(n8514) );
  XNOR2_X1 U10827 ( .A(n14857), .B(n14577), .ZN(n14661) );
  NAND3_X1 U10828 ( .A1(n14549), .A2(n8514), .A3(n14661), .ZN(n8515) );
  OR4_X1 U10829 ( .A1(n14601), .A2(n14630), .A3(n14643), .A4(n8515), .ZN(n8516) );
  NOR3_X1 U10830 ( .A1(n8517), .A2(n14583), .A3(n8516), .ZN(n8518) );
  XNOR2_X1 U10831 ( .A(n14822), .B(n14393), .ZN(n14585) );
  NAND3_X1 U10832 ( .A1(n8519), .A2(n8518), .A3(n14585), .ZN(n8520) );
  XNOR2_X1 U10833 ( .A(n8520), .B(n6681), .ZN(n8531) );
  INV_X1 U10834 ( .A(n8534), .ZN(n8527) );
  NOR2_X1 U10835 ( .A1(n10583), .A2(n8523), .ZN(n8522) );
  MUX2_X1 U10836 ( .A(n8527), .B(n8522), .S(n8521), .Z(n8529) );
  INV_X1 U10837 ( .A(n8523), .ZN(n8524) );
  AND2_X1 U10838 ( .A1(n10583), .A2(n8524), .ZN(n8526) );
  MUX2_X1 U10839 ( .A(n8527), .B(n8526), .S(n8525), .Z(n8528) );
  MUX2_X1 U10840 ( .A(n8529), .B(n8528), .S(n14522), .Z(n8530) );
  NAND2_X1 U10841 ( .A1(n8533), .A2(n8532), .ZN(n8542) );
  NOR3_X1 U10842 ( .A1(n8536), .A2(n8535), .A3(n8534), .ZN(n8541) );
  OAI21_X1 U10843 ( .B1(n8537), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10844 ( .A(n8539), .B(n8538), .ZN(n10559) );
  INV_X2 U10845 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U10846 ( .A1(n10559), .A2(P1_U3086), .ZN(n12180) );
  INV_X1 U10847 ( .A(n12180), .ZN(n8540) );
  OAI21_X1 U10848 ( .B1(n8542), .B2(n8541), .A(n8540), .ZN(n8558) );
  NAND2_X1 U10849 ( .A1(n6681), .A2(n14953), .ZN(n8544) );
  NAND2_X1 U10850 ( .A1(n15253), .A2(n10560), .ZN(n8554) );
  NAND2_X1 U10851 ( .A1(n8545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10852 ( .A1(n6716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8547) );
  XNOR2_X1 U10853 ( .A(n8547), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10477) );
  INV_X1 U10854 ( .A(n8548), .ZN(n8549) );
  NAND2_X1 U10855 ( .A1(n8549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8550) );
  MUX2_X1 U10856 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8550), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8551) );
  AND2_X1 U10857 ( .A1(n10481), .A2(n10559), .ZN(n8553) );
  NAND2_X1 U10858 ( .A1(n8554), .A2(n8553), .ZN(n10486) );
  INV_X1 U10859 ( .A(n8555), .ZN(n10588) );
  INV_X1 U10860 ( .A(n14986), .ZN(n15095) );
  NOR3_X1 U10861 ( .A1(n11322), .A2(n15095), .A3(n6988), .ZN(n8557) );
  OAI21_X1 U10862 ( .B1(n12180), .B2(n14953), .A(P1_B_REG_SCAN_IN), .ZN(n8556)
         );
  NAND2_X1 U10863 ( .A1(n8558), .A2(n7762), .ZN(P1_U3242) );
  INV_X1 U10864 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8563) );
  INV_X1 U10865 ( .A(n8576), .ZN(n8570) );
  INV_X1 U10866 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10867 ( .A1(n8570), .A2(n8569), .ZN(n8578) );
  INV_X1 U10868 ( .A(n9066), .ZN(n8573) );
  XNOR2_X2 U10869 ( .A(n8574), .B(n8573), .ZN(n8612) );
  NAND2_X1 U10870 ( .A1(n8578), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10871 ( .A1(n8576), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8577) );
  MUX2_X1 U10872 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8577), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8579) );
  NOR2_X1 U10873 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8583) );
  NOR2_X1 U10874 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8582) );
  NOR2_X1 U10875 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8581) );
  INV_X1 U10876 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8587) );
  INV_X1 U10877 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10878 ( .A1(n12882), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8602) );
  INV_X2 U10879 ( .A(n8590), .ZN(n14241) );
  INV_X1 U10880 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8591) );
  OR2_X1 U10881 ( .A1(n12885), .A2(n8591), .ZN(n8601) );
  NAND2_X1 U10882 ( .A1(n8685), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U10883 ( .A1(n8722), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8762) );
  INV_X1 U10884 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8761) );
  INV_X1 U10885 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8901) );
  INV_X1 U10886 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8921) );
  INV_X1 U10887 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8973) );
  INV_X1 U10888 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13708) );
  INV_X1 U10889 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U10890 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n9021), .ZN(n9038) );
  INV_X1 U10891 ( .A(n9038), .ZN(n8593) );
  NAND2_X1 U10892 ( .A1(n8593), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9040) );
  INV_X1 U10893 ( .A(n9040), .ZN(n8594) );
  NAND2_X1 U10894 ( .A1(n8594), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9056) );
  INV_X1 U10895 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10896 ( .A1(n9040), .A2(n8595), .ZN(n8596) );
  NAND2_X1 U10897 ( .A1(n9056), .A2(n8596), .ZN(n13971) );
  OR2_X1 U10898 ( .A1(n8721), .A2(n13971), .ZN(n8600) );
  INV_X1 U10899 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8598) );
  OR2_X1 U10900 ( .A1(n12868), .A2(n8598), .ZN(n8599) );
  NAND4_X1 U10901 ( .A1(n8602), .A2(n8601), .A3(n8600), .A4(n8599), .ZN(n13960) );
  NAND2_X1 U10902 ( .A1(n6678), .A2(n13960), .ZN(n9049) );
  INV_X1 U10903 ( .A(n9049), .ZN(n9051) );
  OAI21_X2 U10904 ( .B1(n8864), .B2(n8603), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8605) );
  XNOR2_X2 U10905 ( .A(n8608), .B(n8607), .ZN(n10752) );
  NAND2_X2 U10906 ( .A1(n10782), .A2(n10752), .ZN(n8916) );
  NAND2_X1 U10907 ( .A1(n8916), .A2(n10501), .ZN(n12857) );
  NAND2_X1 U10908 ( .A1(n14251), .A2(n6675), .ZN(n8610) );
  INV_X1 U10909 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14253) );
  OR2_X1 U10910 ( .A1(n12879), .A2(n14253), .ZN(n8609) );
  INV_X1 U10911 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U10912 ( .A1(n8615), .A2(n8614), .ZN(n8892) );
  INV_X1 U10913 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8617) );
  INV_X1 U10914 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8616) );
  NAND3_X1 U10915 ( .A1(n8618), .A2(n8617), .A3(n8616), .ZN(n8619) );
  OAI21_X1 U10916 ( .B1(n8892), .B2(n8619), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8620) );
  NAND2_X1 U10917 ( .A1(n8621), .A2(n13871), .ZN(n10979) );
  INV_X1 U10918 ( .A(n8613), .ZN(n12651) );
  XNOR2_X1 U10919 ( .A(n14154), .B(n13693), .ZN(n9050) );
  NAND2_X1 U10920 ( .A1(n12882), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8626) );
  INV_X1 U10921 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8622) );
  OR2_X1 U10922 ( .A1(n12885), .A2(n8622), .ZN(n8625) );
  OAI21_X1 U10923 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9021), .A(n9038), .ZN(
        n14008) );
  OR2_X1 U10924 ( .A1(n8721), .A2(n14008), .ZN(n8624) );
  INV_X1 U10925 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14009) );
  OR2_X1 U10926 ( .A1(n12868), .A2(n14009), .ZN(n8623) );
  NAND4_X1 U10927 ( .A1(n8626), .A2(n8625), .A3(n8624), .A4(n8623), .ZN(n13920) );
  NAND2_X1 U10928 ( .A1(n6678), .A2(n13920), .ZN(n9031) );
  INV_X1 U10929 ( .A(n9031), .ZN(n9033) );
  NAND2_X1 U10930 ( .A1(n12206), .A2(n6675), .ZN(n8628) );
  INV_X1 U10931 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12212) );
  OR2_X1 U10932 ( .A1(n12879), .A2(n12212), .ZN(n8627) );
  XNOR2_X1 U10933 ( .A(n14165), .B(n13693), .ZN(n9032) );
  INV_X1 U10934 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U10935 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8629) );
  XNOR2_X1 U10936 ( .A(n8630), .B(n8629), .ZN(n10869) );
  OR2_X1 U10937 ( .A1(n8916), .A2(n10869), .ZN(n8633) );
  INV_X1 U10938 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8634) );
  INV_X1 U10939 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10756) );
  OR2_X1 U10940 ( .A1(n8656), .A2(n10756), .ZN(n8636) );
  NAND2_X1 U10941 ( .A1(n8655), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8635) );
  INV_X1 U10942 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U10943 ( .A1(n14018), .A2(n13800), .ZN(n8637) );
  INV_X1 U10944 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10871) );
  INV_X1 U10945 ( .A(SI_0_), .ZN(n10532) );
  NOR2_X1 U10946 ( .A1(n10502), .A2(n10532), .ZN(n8639) );
  XNOR2_X1 U10947 ( .A(n8639), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14256) );
  MUX2_X1 U10948 ( .A(n10871), .B(n14256), .S(n8916), .Z(n15381) );
  OR2_X1 U10949 ( .A1(n8653), .A2(n12648), .ZN(n8644) );
  INV_X1 U10950 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15383) );
  NAND2_X1 U10951 ( .A1(n8655), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8642) );
  INV_X1 U10952 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8640) );
  OR2_X1 U10953 ( .A1(n8656), .A2(n8640), .ZN(n8641) );
  AND2_X1 U10954 ( .A1(n12648), .A2(n10891), .ZN(n11610) );
  NAND2_X1 U10955 ( .A1(n11610), .A2(n14018), .ZN(n8643) );
  NAND2_X1 U10956 ( .A1(n8644), .A2(n8643), .ZN(n10899) );
  OR2_X2 U10957 ( .A1(n10898), .A2(n10899), .ZN(n10896) );
  NAND2_X1 U10958 ( .A1(n10896), .A2(n8645), .ZN(n10993) );
  INV_X1 U10959 ( .A(n8647), .ZN(n8648) );
  NAND2_X1 U10960 ( .A1(n8648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8649) );
  XNOR2_X1 U10961 ( .A(n8649), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10775) );
  NAND2_X1 U10962 ( .A1(n8650), .A2(n12846), .ZN(n8651) );
  NAND2_X2 U10963 ( .A1(n8652), .A2(n8651), .ZN(n12663) );
  XNOR2_X1 U10964 ( .A(n8653), .B(n12663), .ZN(n8662) );
  INV_X1 U10965 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10995) );
  OR2_X1 U10966 ( .A1(n8721), .A2(n10995), .ZN(n8660) );
  INV_X1 U10967 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10968 ( .A1(n8655), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8658) );
  INV_X1 U10969 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10755) );
  OR2_X1 U10970 ( .A1(n8656), .A2(n10755), .ZN(n8657) );
  AND2_X1 U10971 ( .A1(n14018), .A2(n13799), .ZN(n8661) );
  NAND2_X1 U10972 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  AND2_X1 U10973 ( .A1(n8664), .A2(n8663), .ZN(n10994) );
  NAND2_X1 U10974 ( .A1(n10993), .A2(n10994), .ZN(n10992) );
  INV_X1 U10975 ( .A(n8667), .ZN(n8677) );
  NAND2_X1 U10976 ( .A1(n8677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8668) );
  XNOR2_X1 U10977 ( .A(n8668), .B(P2_IR_REG_3__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U10978 ( .A1(n8666), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10747), 
        .B2(n13805), .ZN(n8669) );
  XNOR2_X1 U10979 ( .A(n15410), .B(n13693), .ZN(n8675) );
  NAND2_X1 U10980 ( .A1(n8655), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8673) );
  INV_X1 U10981 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11419) );
  OR2_X1 U10982 ( .A1(n12868), .A2(n11419), .ZN(n8672) );
  OR2_X1 U10983 ( .A1(n12885), .A2(n15415), .ZN(n8671) );
  OR2_X1 U10984 ( .A1(n8721), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8670) );
  AND2_X1 U10985 ( .A1(n14018), .A2(n13798), .ZN(n8674) );
  XNOR2_X1 U10986 ( .A(n8675), .B(n8674), .ZN(n11019) );
  NAND2_X1 U10987 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  NAND2_X1 U10988 ( .A1(n10537), .A2(n12846), .ZN(n8684) );
  NAND2_X1 U10989 ( .A1(n8679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8678) );
  MUX2_X1 U10990 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8678), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8682) );
  INV_X1 U10991 ( .A(n8679), .ZN(n8681) );
  NAND2_X1 U10992 ( .A1(n8681), .A2(n8680), .ZN(n8716) );
  NAND2_X1 U10993 ( .A1(n8682), .A2(n8716), .ZN(n13819) );
  INV_X1 U10994 ( .A(n13819), .ZN(n13815) );
  AOI22_X1 U10995 ( .A1(n8666), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10747), 
        .B2(n13815), .ZN(n8683) );
  XNOR2_X1 U10996 ( .A(n15417), .B(n9007), .ZN(n8691) );
  NAND2_X1 U10997 ( .A1(n12882), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8690) );
  INV_X1 U10998 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11794) );
  OR2_X1 U10999 ( .A1(n12868), .A2(n11794), .ZN(n8689) );
  INV_X1 U11000 ( .A(n8685), .ZN(n8703) );
  OAI21_X1 U11001 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8703), .ZN(n11798) );
  OR2_X1 U11002 ( .A1(n8721), .A2(n11798), .ZN(n8688) );
  INV_X1 U11003 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8686) );
  OR2_X1 U11004 ( .A1(n12885), .A2(n8686), .ZN(n8687) );
  INV_X1 U11005 ( .A(n12678), .ZN(n13797) );
  NAND2_X1 U11006 ( .A1(n13797), .A2(n6678), .ZN(n8692) );
  NAND2_X1 U11007 ( .A1(n8691), .A2(n8692), .ZN(n8698) );
  INV_X1 U11008 ( .A(n8691), .ZN(n8694) );
  INV_X1 U11009 ( .A(n8692), .ZN(n8693) );
  NAND2_X1 U11010 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  NAND2_X1 U11011 ( .A1(n8698), .A2(n8695), .ZN(n10986) );
  NAND2_X1 U11012 ( .A1(n10984), .A2(n8698), .ZN(n11003) );
  NAND2_X1 U11013 ( .A1(n10541), .A2(n6675), .ZN(n8701) );
  NAND2_X1 U11014 ( .A1(n8716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8699) );
  XNOR2_X1 U11015 ( .A(n8699), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U11016 ( .A1(n8666), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10747), 
        .B2(n10780), .ZN(n8700) );
  NAND2_X1 U11017 ( .A1(n8701), .A2(n8700), .ZN(n15423) );
  XNOR2_X1 U11018 ( .A(n15423), .B(n9007), .ZN(n8710) );
  NAND2_X1 U11019 ( .A1(n12882), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8709) );
  INV_X1 U11020 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11783) );
  OR2_X1 U11021 ( .A1(n12868), .A2(n11783), .ZN(n8708) );
  INV_X1 U11022 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11023 ( .A1(n8703), .A2(n8702), .ZN(n8704) );
  NAND2_X1 U11024 ( .A1(n8724), .A2(n8704), .ZN(n11784) );
  OR2_X1 U11025 ( .A1(n8721), .A2(n11784), .ZN(n8707) );
  INV_X1 U11026 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8705) );
  OR2_X1 U11027 ( .A1(n12885), .A2(n8705), .ZN(n8706) );
  NAND4_X1 U11028 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(n13796) );
  NAND2_X1 U11029 ( .A1(n6678), .A2(n13796), .ZN(n8711) );
  NAND2_X1 U11030 ( .A1(n8710), .A2(n8711), .ZN(n8715) );
  INV_X1 U11031 ( .A(n8710), .ZN(n8713) );
  INV_X1 U11032 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U11033 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  AND2_X1 U11034 ( .A1(n8715), .A2(n8714), .ZN(n11004) );
  NAND2_X1 U11035 ( .A1(n10555), .A2(n6675), .ZN(n8719) );
  NAND2_X1 U11036 ( .A1(n8735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8717) );
  XNOR2_X1 U11037 ( .A(n8717), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U11038 ( .A1(n8666), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10747), 
        .B2(n10811), .ZN(n8718) );
  XNOR2_X1 U11039 ( .A(n15429), .B(n9007), .ZN(n8730) );
  NAND2_X1 U11040 ( .A1(n12883), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8729) );
  INV_X1 U11041 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8720) );
  INV_X1 U11042 ( .A(n8722), .ZN(n8743) );
  NAND2_X1 U11043 ( .A1(n8724), .A2(n8723), .ZN(n8725) );
  NAND2_X1 U11044 ( .A1(n8743), .A2(n8725), .ZN(n11841) );
  OR2_X1 U11045 ( .A1(n8721), .A2(n11841), .ZN(n8728) );
  INV_X1 U11046 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8726) );
  OR2_X1 U11047 ( .A1(n12885), .A2(n8726), .ZN(n8727) );
  NAND2_X1 U11048 ( .A1(n6678), .A2(n13795), .ZN(n8731) );
  XNOR2_X1 U11049 ( .A(n8730), .B(n8731), .ZN(n11008) );
  INV_X1 U11050 ( .A(n8730), .ZN(n8733) );
  INV_X1 U11051 ( .A(n8731), .ZN(n8732) );
  NAND2_X1 U11052 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U11053 ( .A1(n10564), .A2(n6675), .ZN(n8740) );
  INV_X1 U11054 ( .A(n8735), .ZN(n8737) );
  NAND2_X1 U11055 ( .A1(n8737), .A2(n8736), .ZN(n8754) );
  NAND2_X1 U11056 ( .A1(n8754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8738) );
  XNOR2_X1 U11057 ( .A(n8738), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13836) );
  AOI22_X1 U11058 ( .A1(n8666), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10747), 
        .B2(n13836), .ZN(n8739) );
  XNOR2_X1 U11059 ( .A(n15434), .B(n13693), .ZN(n8752) );
  NAND2_X1 U11060 ( .A1(n12883), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8749) );
  INV_X1 U11061 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8741) );
  OR2_X1 U11062 ( .A1(n12866), .A2(n8741), .ZN(n8748) );
  INV_X1 U11063 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11064 ( .A1(n8743), .A2(n8742), .ZN(n8744) );
  NAND2_X1 U11065 ( .A1(n8762), .A2(n8744), .ZN(n11824) );
  OR2_X1 U11066 ( .A1(n8721), .A2(n11824), .ZN(n8747) );
  INV_X1 U11067 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8745) );
  OR2_X1 U11068 ( .A1(n12885), .A2(n8745), .ZN(n8746) );
  NAND4_X1 U11069 ( .A1(n8749), .A2(n8748), .A3(n8747), .A4(n8746), .ZN(n13794) );
  NAND2_X1 U11070 ( .A1(n6678), .A2(n13794), .ZN(n8750) );
  XNOR2_X1 U11071 ( .A(n8752), .B(n8750), .ZN(n11038) );
  INV_X1 U11072 ( .A(n8750), .ZN(n8751) );
  AND2_X1 U11073 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U11074 ( .A1(n10571), .A2(n6675), .ZN(n8759) );
  NAND2_X1 U11075 ( .A1(n8756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8755) );
  MUX2_X1 U11076 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8755), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8757) );
  NAND2_X1 U11077 ( .A1(n8757), .A2(n8794), .ZN(n13850) );
  INV_X1 U11078 ( .A(n13850), .ZN(n10817) );
  AOI22_X1 U11079 ( .A1(n8666), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10817), 
        .B2(n10747), .ZN(n8758) );
  XNOR2_X1 U11080 ( .A(n12717), .B(n9007), .ZN(n8769) );
  NAND2_X1 U11081 ( .A1(n12883), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8768) );
  INV_X1 U11082 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8760) );
  OR2_X1 U11083 ( .A1(n12866), .A2(n8760), .ZN(n8767) );
  NAND2_X1 U11084 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  NAND2_X1 U11085 ( .A1(n8781), .A2(n8763), .ZN(n11812) );
  OR2_X1 U11086 ( .A1(n8721), .A2(n11812), .ZN(n8766) );
  INV_X1 U11087 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8764) );
  OR2_X1 U11088 ( .A1(n12885), .A2(n8764), .ZN(n8765) );
  NAND4_X1 U11089 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n13793) );
  NAND2_X1 U11090 ( .A1(n6678), .A2(n13793), .ZN(n8770) );
  NAND2_X1 U11091 ( .A1(n8769), .A2(n8770), .ZN(n8774) );
  INV_X1 U11092 ( .A(n8769), .ZN(n8772) );
  INV_X1 U11093 ( .A(n8770), .ZN(n8771) );
  NAND2_X1 U11094 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  AND2_X1 U11095 ( .A1(n8774), .A2(n8773), .ZN(n11105) );
  NAND2_X1 U11096 ( .A1(n10575), .A2(n6675), .ZN(n8777) );
  NAND2_X1 U11097 ( .A1(n8794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8775) );
  XNOR2_X1 U11098 ( .A(n8775), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U11099 ( .A1(n8666), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10820), 
        .B2(n10747), .ZN(n8776) );
  XNOR2_X1 U11100 ( .A(n15449), .B(n9007), .ZN(n8788) );
  NAND2_X1 U11101 ( .A1(n12883), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8787) );
  INV_X1 U11102 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8778) );
  OR2_X1 U11103 ( .A1(n12866), .A2(n8778), .ZN(n8786) );
  INV_X1 U11104 ( .A(n8779), .ZN(n8802) );
  NAND2_X1 U11105 ( .A1(n8781), .A2(n8780), .ZN(n8782) );
  NAND2_X1 U11106 ( .A1(n8802), .A2(n8782), .ZN(n11451) );
  OR2_X1 U11107 ( .A1(n8721), .A2(n11451), .ZN(n8785) );
  INV_X1 U11108 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8783) );
  OR2_X1 U11109 ( .A1(n12885), .A2(n8783), .ZN(n8784) );
  NAND4_X1 U11110 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(n13792) );
  NAND2_X1 U11111 ( .A1(n6678), .A2(n13792), .ZN(n8789) );
  NAND2_X1 U11112 ( .A1(n8788), .A2(n8789), .ZN(n8793) );
  INV_X1 U11113 ( .A(n8788), .ZN(n8791) );
  INV_X1 U11114 ( .A(n8789), .ZN(n8790) );
  NAND2_X1 U11115 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  AND2_X1 U11116 ( .A1(n8793), .A2(n8792), .ZN(n11166) );
  NAND2_X1 U11117 ( .A1(n10650), .A2(n6675), .ZN(n8799) );
  INV_X1 U11118 ( .A(n8794), .ZN(n8796) );
  INV_X1 U11119 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11120 ( .A1(n8796), .A2(n8795), .ZN(n8813) );
  NAND2_X1 U11121 ( .A1(n8813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8797) );
  XNOR2_X1 U11122 ( .A(n8797), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U11123 ( .A1(n10854), .A2(n10747), .B1(n8666), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11124 ( .A1(n8799), .A2(n8798), .ZN(n12731) );
  XNOR2_X1 U11125 ( .A(n12731), .B(n9007), .ZN(n8809) );
  NAND2_X1 U11126 ( .A1(n12883), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8808) );
  INV_X1 U11127 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10804) );
  OR2_X1 U11128 ( .A1(n12866), .A2(n10804), .ZN(n8807) );
  INV_X1 U11129 ( .A(n8800), .ZN(n8818) );
  INV_X1 U11130 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U11131 ( .A1(n8802), .A2(n8801), .ZN(n8803) );
  NAND2_X1 U11132 ( .A1(n8818), .A2(n8803), .ZN(n11648) );
  OR2_X1 U11133 ( .A1(n8721), .A2(n11648), .ZN(n8806) );
  INV_X1 U11134 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8804) );
  OR2_X1 U11135 ( .A1(n12885), .A2(n8804), .ZN(n8805) );
  NAND4_X1 U11136 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n13791) );
  NAND2_X1 U11137 ( .A1(n6678), .A2(n13791), .ZN(n8810) );
  XNOR2_X1 U11138 ( .A(n8809), .B(n8810), .ZN(n11268) );
  INV_X1 U11139 ( .A(n8809), .ZN(n8812) );
  INV_X1 U11140 ( .A(n8810), .ZN(n8811) );
  NAND2_X1 U11141 ( .A1(n10688), .A2(n6675), .ZN(n8816) );
  OAI21_X1 U11142 ( .B1(n8813), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U11143 ( .A(n8814), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U11144 ( .A1(n10910), .A2(n10747), .B1(n8666), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U11145 ( .A(n12736), .B(n9007), .ZN(n8825) );
  NAND2_X1 U11146 ( .A1(n12882), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8824) );
  INV_X1 U11147 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11148 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  NAND2_X1 U11149 ( .A1(n8854), .A2(n8819), .ZN(n11661) );
  OR2_X1 U11150 ( .A1(n8721), .A2(n11661), .ZN(n8823) );
  INV_X1 U11151 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8820) );
  OR2_X1 U11152 ( .A1(n12885), .A2(n8820), .ZN(n8822) );
  INV_X1 U11153 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11662) );
  OR2_X1 U11154 ( .A1(n12868), .A2(n11662), .ZN(n8821) );
  NAND4_X1 U11155 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n13790) );
  NAND2_X1 U11156 ( .A1(n6678), .A2(n13790), .ZN(n8826) );
  NAND2_X1 U11157 ( .A1(n8825), .A2(n8826), .ZN(n8830) );
  INV_X1 U11158 ( .A(n8825), .ZN(n8828) );
  INV_X1 U11159 ( .A(n8826), .ZN(n8827) );
  NAND2_X1 U11160 ( .A1(n8828), .A2(n8827), .ZN(n8829) );
  NAND2_X1 U11161 ( .A1(n8830), .A2(n8829), .ZN(n11622) );
  NAND2_X1 U11162 ( .A1(n10720), .A2(n6675), .ZN(n8836) );
  NAND2_X1 U11163 ( .A1(n8831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8832) );
  MUX2_X1 U11164 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8832), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8834) );
  NAND2_X1 U11165 ( .A1(n8834), .A2(n8833), .ZN(n15353) );
  INV_X1 U11166 ( .A(n15353), .ZN(n15359) );
  AOI22_X1 U11167 ( .A1(n8666), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10747), 
        .B2(n15359), .ZN(n8835) );
  XNOR2_X1 U11168 ( .A(n12749), .B(n9007), .ZN(n8843) );
  NAND2_X1 U11169 ( .A1(n12882), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8842) );
  INV_X1 U11170 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8837) );
  OR2_X1 U11171 ( .A1(n12868), .A2(n8837), .ZN(n8841) );
  XNOR2_X1 U11172 ( .A(n8854), .B(n8853), .ZN(n11941) );
  OR2_X1 U11173 ( .A1(n8721), .A2(n11941), .ZN(n8840) );
  INV_X1 U11174 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8838) );
  OR2_X1 U11175 ( .A1(n12885), .A2(n8838), .ZN(n8839) );
  NAND4_X1 U11176 ( .A1(n8842), .A2(n8841), .A3(n8840), .A4(n8839), .ZN(n13789) );
  NAND2_X1 U11177 ( .A1(n6678), .A2(n13789), .ZN(n8844) );
  NAND2_X1 U11178 ( .A1(n8843), .A2(n8844), .ZN(n8848) );
  INV_X1 U11179 ( .A(n8843), .ZN(n8846) );
  INV_X1 U11180 ( .A(n8844), .ZN(n8845) );
  NAND2_X1 U11181 ( .A1(n8846), .A2(n8845), .ZN(n8847) );
  AND2_X1 U11182 ( .A1(n8848), .A2(n8847), .ZN(n11939) );
  NAND2_X1 U11183 ( .A1(n10745), .A2(n6675), .ZN(n8851) );
  NAND2_X1 U11184 ( .A1(n8833), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8849) );
  XNOR2_X1 U11185 ( .A(n8849), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U11186 ( .A1(n8666), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10747), 
        .B2(n11077), .ZN(n8850) );
  XNOR2_X1 U11187 ( .A(n12756), .B(n13693), .ZN(n8863) );
  INV_X1 U11188 ( .A(n8721), .ZN(n8944) );
  OAI21_X1 U11189 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8855) );
  AND2_X1 U11190 ( .A1(n8855), .A2(n8871), .ZN(n12234) );
  NAND2_X1 U11191 ( .A1(n8944), .A2(n12234), .ZN(n8860) );
  NAND2_X1 U11192 ( .A1(n12882), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8859) );
  INV_X1 U11193 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11072) );
  OR2_X1 U11194 ( .A1(n12868), .A2(n11072), .ZN(n8858) );
  INV_X1 U11195 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8856) );
  OR2_X1 U11196 ( .A1(n12885), .A2(n8856), .ZN(n8857) );
  NAND4_X1 U11197 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n12755) );
  NAND2_X1 U11198 ( .A1(n6678), .A2(n12755), .ZN(n8861) );
  XNOR2_X1 U11199 ( .A(n8863), .B(n8861), .ZN(n12010) );
  INV_X1 U11200 ( .A(n8861), .ZN(n8862) );
  NAND2_X1 U11201 ( .A1(n8864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U11202 ( .A(n8865), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U11203 ( .A1(n8666), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10747), 
        .B2(n11426), .ZN(n8866) );
  INV_X1 U11204 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11205 ( .A1(n12883), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11206 ( .A1(n12882), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8868) );
  AND2_X1 U11207 ( .A1(n8869), .A2(n8868), .ZN(n8874) );
  INV_X1 U11208 ( .A(n8870), .ZN(n8884) );
  NAND2_X1 U11209 ( .A1(n8871), .A2(n12201), .ZN(n8872) );
  NAND2_X1 U11210 ( .A1(n8884), .A2(n8872), .ZN(n12319) );
  OR2_X1 U11211 ( .A1(n12319), .A2(n8721), .ZN(n8873) );
  OAI211_X1 U11212 ( .C1(n12885), .C2(n8875), .A(n8874), .B(n8873), .ZN(n13788) );
  NAND2_X1 U11213 ( .A1(n6678), .A2(n13788), .ZN(n8877) );
  NAND2_X1 U11214 ( .A1(n8876), .A2(n8877), .ZN(n8879) );
  NAND2_X1 U11215 ( .A1(n11015), .A2(n6675), .ZN(n8882) );
  NAND2_X1 U11216 ( .A1(n8892), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8880) );
  XNOR2_X1 U11217 ( .A(n8880), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U11218 ( .A1(n8666), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10747), 
        .B2(n11906), .ZN(n8881) );
  XNOR2_X1 U11219 ( .A(n12771), .B(n13693), .ZN(n8888) );
  XNOR2_X1 U11220 ( .A(n8890), .B(n8888), .ZN(n12363) );
  INV_X1 U11221 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12294) );
  INV_X1 U11222 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U11223 ( .A1(n8884), .A2(n8883), .ZN(n8885) );
  NAND2_X1 U11224 ( .A1(n8902), .A2(n8885), .ZN(n12364) );
  OR2_X1 U11225 ( .A1(n12364), .A2(n8721), .ZN(n8887) );
  AOI22_X1 U11226 ( .A1(n12882), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n12840), 
        .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n8886) );
  OAI211_X1 U11227 ( .C1(n12868), .C2(n12294), .A(n8887), .B(n8886), .ZN(
        n13787) );
  AND2_X1 U11228 ( .A1(n13787), .A2(n6678), .ZN(n12362) );
  INV_X1 U11229 ( .A(n8888), .ZN(n8889) );
  OR2_X1 U11230 ( .A1(n8890), .A2(n8889), .ZN(n8891) );
  NAND2_X1 U11231 ( .A1(n10880), .A2(n6675), .ZN(n8900) );
  NOR2_X1 U11232 ( .A1(n8892), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8896) );
  INV_X1 U11233 ( .A(n8896), .ZN(n8893) );
  NAND2_X1 U11234 ( .A1(n8893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8894) );
  MUX2_X1 U11235 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8894), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8897) );
  INV_X1 U11236 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11237 ( .A1(n8896), .A2(n8895), .ZN(n8914) );
  NAND2_X1 U11238 ( .A1(n8897), .A2(n8914), .ZN(n12424) );
  OAI22_X1 U11239 ( .A1(n12879), .A2(n10927), .B1(n12424), .B2(n8916), .ZN(
        n8898) );
  INV_X1 U11240 ( .A(n8898), .ZN(n8899) );
  XNOR2_X1 U11241 ( .A(n14207), .B(n9007), .ZN(n8906) );
  NAND2_X1 U11242 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  NAND2_X1 U11243 ( .A1(n8922), .A2(n8903), .ZN(n13723) );
  AOI22_X1 U11244 ( .A1(n12882), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n12883), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U11245 ( .A1(n12840), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8904) );
  OAI211_X1 U11246 ( .C1(n13723), .C2(n8721), .A(n8905), .B(n8904), .ZN(n14125) );
  NAND2_X1 U11247 ( .A1(n14125), .A2(n6678), .ZN(n8907) );
  NAND2_X1 U11248 ( .A1(n8906), .A2(n8907), .ZN(n8912) );
  INV_X1 U11249 ( .A(n8906), .ZN(n8909) );
  INV_X1 U11250 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U11251 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  NAND2_X1 U11252 ( .A1(n8912), .A2(n8910), .ZN(n13722) );
  INV_X1 U11253 ( .A(n13722), .ZN(n8911) );
  NAND2_X1 U11254 ( .A1(n10958), .A2(n6675), .ZN(n8919) );
  NAND2_X1 U11255 ( .A1(n8914), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8913) );
  MUX2_X1 U11256 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8913), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8915) );
  OR2_X1 U11257 ( .A1(n8914), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11258 ( .A1(n8915), .A2(n8935), .ZN(n15378) );
  OAI22_X1 U11259 ( .A1(n15378), .A2(n8916), .B1(n12879), .B2(n10960), .ZN(
        n8917) );
  INV_X1 U11260 ( .A(n8917), .ZN(n8918) );
  XNOR2_X1 U11261 ( .A(n14200), .B(n9007), .ZN(n8929) );
  INV_X1 U11262 ( .A(n8920), .ZN(n8942) );
  NAND2_X1 U11263 ( .A1(n8922), .A2(n8921), .ZN(n8923) );
  NAND2_X1 U11264 ( .A1(n8942), .A2(n8923), .ZN(n14116) );
  OR2_X1 U11265 ( .A1(n14116), .A2(n8721), .ZN(n8928) );
  INV_X1 U11266 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U11267 ( .A1(n12840), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11268 ( .A1(n12882), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8924) );
  OAI211_X1 U11269 ( .C1(n12868), .C2(n12421), .A(n8925), .B(n8924), .ZN(n8926) );
  INV_X1 U11270 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U11271 ( .A1(n8928), .A2(n8927), .ZN(n13889) );
  NAND2_X1 U11272 ( .A1(n13889), .A2(n6678), .ZN(n8930) );
  NAND2_X1 U11273 ( .A1(n8929), .A2(n8930), .ZN(n8934) );
  INV_X1 U11274 ( .A(n8929), .ZN(n8932) );
  INV_X1 U11275 ( .A(n8930), .ZN(n8931) );
  NAND2_X1 U11276 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  AND2_X1 U11277 ( .A1(n8934), .A2(n8933), .ZN(n13731) );
  NAND2_X1 U11278 ( .A1(n11132), .A2(n6675), .ZN(n8939) );
  NAND2_X1 U11279 ( .A1(n8935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8936) );
  XNOR2_X1 U11280 ( .A(n8936), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12426) );
  NOR2_X1 U11281 ( .A1(n12879), .A2(n11135), .ZN(n8937) );
  AOI21_X1 U11282 ( .B1(n12426), .B2(n10747), .A(n8937), .ZN(n8938) );
  XNOR2_X1 U11283 ( .A(n14195), .B(n9007), .ZN(n8951) );
  INV_X1 U11284 ( .A(n8940), .ZN(n8959) );
  INV_X1 U11285 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11286 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  AND2_X1 U11287 ( .A1(n8959), .A2(n8943), .ZN(n14100) );
  NAND2_X1 U11288 ( .A1(n14100), .A2(n8944), .ZN(n8950) );
  INV_X1 U11289 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U11290 ( .A1(n12883), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U11291 ( .A1(n12840), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8945) );
  OAI211_X1 U11292 ( .C1(n12866), .C2(n8947), .A(n8946), .B(n8945), .ZN(n8948)
         );
  INV_X1 U11293 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U11294 ( .A1(n8950), .A2(n8949), .ZN(n14127) );
  NAND2_X1 U11295 ( .A1(n14127), .A2(n6678), .ZN(n8952) );
  XNOR2_X1 U11296 ( .A(n8951), .B(n8952), .ZN(n13764) );
  INV_X1 U11297 ( .A(n8951), .ZN(n8954) );
  INV_X1 U11298 ( .A(n8952), .ZN(n8953) );
  NAND2_X1 U11299 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  NAND2_X1 U11300 ( .A1(n11299), .A2(n6675), .ZN(n8957) );
  AOI22_X1 U11301 ( .A1(n8666), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10747), 
        .B2(n12926), .ZN(n8956) );
  XNOR2_X1 U11302 ( .A(n14191), .B(n9007), .ZN(n8967) );
  INV_X1 U11303 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11304 ( .A1(n8959), .A2(n8958), .ZN(n8960) );
  NAND2_X1 U11305 ( .A1(n8974), .A2(n8960), .ZN(n14081) );
  OR2_X1 U11306 ( .A1(n14081), .A2(n8721), .ZN(n8966) );
  INV_X1 U11307 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11308 ( .A1(n12883), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11309 ( .A1(n12840), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8961) );
  OAI211_X1 U11310 ( .C1(n12866), .C2(n8963), .A(n8962), .B(n8961), .ZN(n8964)
         );
  INV_X1 U11311 ( .A(n8964), .ZN(n8965) );
  NAND2_X1 U11312 ( .A1(n8966), .A2(n8965), .ZN(n13892) );
  NAND2_X1 U11313 ( .A1(n13892), .A2(n6678), .ZN(n8968) );
  NAND2_X1 U11314 ( .A1(n8967), .A2(n8968), .ZN(n13682) );
  INV_X1 U11315 ( .A(n8967), .ZN(n8970) );
  INV_X1 U11316 ( .A(n8968), .ZN(n8969) );
  NAND2_X1 U11317 ( .A1(n8970), .A2(n8969), .ZN(n13681) );
  INV_X1 U11318 ( .A(n13750), .ZN(n8983) );
  NAND2_X1 U11319 ( .A1(n11884), .A2(n6675), .ZN(n8972) );
  OR2_X1 U11320 ( .A1(n12879), .A2(n7635), .ZN(n8971) );
  NAND2_X2 U11321 ( .A1(n8972), .A2(n8971), .ZN(n14185) );
  XNOR2_X1 U11322 ( .A(n14185), .B(n9007), .ZN(n8985) );
  NAND2_X1 U11323 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  NAND2_X1 U11324 ( .A1(n8988), .A2(n8975), .ZN(n14063) );
  OR2_X1 U11325 ( .A1(n14063), .A2(n8721), .ZN(n8981) );
  INV_X1 U11326 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11327 ( .A1(n12883), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11328 ( .A1(n12840), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8976) );
  OAI211_X1 U11329 ( .C1(n12866), .C2(n8978), .A(n8977), .B(n8976), .ZN(n8979)
         );
  INV_X1 U11330 ( .A(n8979), .ZN(n8980) );
  NAND2_X1 U11331 ( .A1(n8981), .A2(n8980), .ZN(n13914) );
  NAND2_X1 U11332 ( .A1(n13914), .A2(n6678), .ZN(n8984) );
  XNOR2_X1 U11333 ( .A(n8985), .B(n8984), .ZN(n13751) );
  NAND2_X1 U11334 ( .A1(n8985), .A2(n8984), .ZN(n8986) );
  OR2_X1 U11335 ( .A1(n12879), .A2(n12017), .ZN(n8987) );
  XNOR2_X1 U11336 ( .A(n14180), .B(n9007), .ZN(n8998) );
  NAND2_X1 U11337 ( .A1(n8988), .A2(n13708), .ZN(n8990) );
  INV_X1 U11338 ( .A(n9008), .ZN(n8989) );
  NAND2_X1 U11339 ( .A1(n8990), .A2(n8989), .ZN(n13706) );
  OR2_X1 U11340 ( .A1(n13706), .A2(n8721), .ZN(n8996) );
  INV_X1 U11341 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U11342 ( .A1(n12883), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U11343 ( .A1(n12840), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8991) );
  OAI211_X1 U11344 ( .C1(n12866), .C2(n8993), .A(n8992), .B(n8991), .ZN(n8994)
         );
  INV_X1 U11345 ( .A(n8994), .ZN(n8995) );
  NAND2_X1 U11346 ( .A1(n8996), .A2(n8995), .ZN(n14031) );
  NAND2_X1 U11347 ( .A1(n14031), .A2(n14018), .ZN(n8999) );
  XNOR2_X1 U11348 ( .A(n8998), .B(n8999), .ZN(n13702) );
  INV_X1 U11349 ( .A(n13702), .ZN(n8997) );
  INV_X1 U11350 ( .A(n8998), .ZN(n9001) );
  INV_X1 U11351 ( .A(n8999), .ZN(n9000) );
  NAND2_X1 U11352 ( .A1(n9001), .A2(n9000), .ZN(n9002) );
  XNOR2_X1 U11353 ( .A(n9004), .B(n9003), .ZN(n12038) );
  NAND2_X1 U11354 ( .A1(n12038), .A2(n6675), .ZN(n9006) );
  OR2_X1 U11355 ( .A1(n12879), .A2(n12040), .ZN(n9005) );
  XNOR2_X1 U11356 ( .A(n14175), .B(n9007), .ZN(n9013) );
  XNOR2_X2 U11357 ( .A(n9015), .B(n9013), .ZN(n13756) );
  NAND2_X1 U11358 ( .A1(n12882), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U11359 ( .A1(n12840), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9011) );
  OAI21_X1 U11360 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n9008), .A(n9020), .ZN(
        n14035) );
  OR2_X1 U11361 ( .A1(n8721), .A2(n14035), .ZN(n9010) );
  INV_X1 U11362 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14036) );
  OR2_X1 U11363 ( .A1(n12868), .A2(n14036), .ZN(n9009) );
  NAND4_X1 U11364 ( .A1(n9012), .A2(n9011), .A3(n9010), .A4(n9009), .ZN(n13915) );
  NAND2_X1 U11365 ( .A1(n6678), .A2(n13915), .ZN(n13757) );
  INV_X1 U11366 ( .A(n9013), .ZN(n9014) );
  NOR2_X1 U11367 ( .A1(n9015), .A2(n9014), .ZN(n9016) );
  AOI21_X2 U11368 ( .B1(n13756), .B2(n13757), .A(n9016), .ZN(n9030) );
  NAND2_X1 U11369 ( .A1(n12179), .A2(n6675), .ZN(n9018) );
  INV_X1 U11370 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12178) );
  OR2_X1 U11371 ( .A1(n12879), .A2(n12178), .ZN(n9017) );
  XNOR2_X1 U11372 ( .A(n14170), .B(n13693), .ZN(n9029) );
  XNOR2_X2 U11373 ( .A(n9030), .B(n9029), .ZN(n13677) );
  NAND2_X1 U11374 ( .A1(n12883), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9028) );
  INV_X1 U11375 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9019) );
  OR2_X1 U11376 ( .A1(n12866), .A2(n9019), .ZN(n9027) );
  INV_X1 U11377 ( .A(n9020), .ZN(n9023) );
  INV_X1 U11378 ( .A(n9021), .ZN(n9022) );
  OAI21_X1 U11379 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n9023), .A(n9022), .ZN(
        n14025) );
  OR2_X1 U11380 ( .A1(n8721), .A2(n14025), .ZN(n9026) );
  INV_X1 U11381 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9024) );
  OR2_X1 U11382 ( .A1(n12885), .A2(n9024), .ZN(n9025) );
  NAND4_X1 U11383 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n14030) );
  NAND2_X1 U11384 ( .A1(n6678), .A2(n14030), .ZN(n13676) );
  NOR2_X2 U11385 ( .A1(n13677), .A2(n13676), .ZN(n13675) );
  NOR2_X2 U11386 ( .A1(n13675), .A2(n7758), .ZN(n13739) );
  XNOR2_X1 U11387 ( .A(n9032), .B(n9031), .ZN(n13738) );
  NAND2_X1 U11388 ( .A1(n12327), .A2(n6675), .ZN(n9035) );
  OR2_X1 U11389 ( .A1(n12879), .A2(n12332), .ZN(n9034) );
  XNOR2_X1 U11390 ( .A(n14159), .B(n13693), .ZN(n9046) );
  NAND2_X1 U11391 ( .A1(n12882), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9044) );
  INV_X1 U11392 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9036) );
  OR2_X1 U11393 ( .A1(n12885), .A2(n9036), .ZN(n9043) );
  INV_X1 U11394 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U11395 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  NAND2_X1 U11396 ( .A1(n9040), .A2(n9039), .ZN(n13988) );
  OR2_X1 U11397 ( .A1(n8721), .A2(n13988), .ZN(n9042) );
  INV_X1 U11398 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13989) );
  OR2_X1 U11399 ( .A1(n12868), .A2(n13989), .ZN(n9041) );
  NAND4_X1 U11400 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n13898) );
  AND2_X1 U11401 ( .A1(n6678), .A2(n13898), .ZN(n9045) );
  NAND2_X1 U11402 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  OAI21_X1 U11403 ( .B1(n9046), .B2(n9045), .A(n9047), .ZN(n13716) );
  INV_X1 U11404 ( .A(n9047), .ZN(n9048) );
  XNOR2_X1 U11405 ( .A(n9050), .B(n9049), .ZN(n13775) );
  NAND2_X1 U11406 ( .A1(n14945), .A2(n6675), .ZN(n9053) );
  OR2_X1 U11407 ( .A1(n12879), .A2(n14250), .ZN(n9052) );
  XNOR2_X1 U11408 ( .A(n14149), .B(n13693), .ZN(n9064) );
  NAND2_X1 U11409 ( .A1(n12882), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9062) );
  INV_X1 U11410 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9054) );
  OR2_X1 U11411 ( .A1(n12885), .A2(n9054), .ZN(n9061) );
  INV_X1 U11412 ( .A(n9056), .ZN(n9055) );
  NAND2_X1 U11413 ( .A1(n9055), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9108) );
  INV_X1 U11414 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U11415 ( .A1(n9056), .A2(n9115), .ZN(n9057) );
  NAND2_X1 U11416 ( .A1(n9108), .A2(n9057), .ZN(n13953) );
  INV_X1 U11417 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9058) );
  OR2_X1 U11418 ( .A1(n12868), .A2(n9058), .ZN(n9059) );
  NAND4_X1 U11419 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n13942) );
  AND2_X1 U11420 ( .A1(n6678), .A2(n13942), .ZN(n9063) );
  NAND2_X1 U11421 ( .A1(n9064), .A2(n9063), .ZN(n13690) );
  NAND2_X1 U11422 ( .A1(n9076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9069) );
  INV_X1 U11423 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9068) );
  NOR2_X1 U11424 ( .A1(n9070), .A2(n8588), .ZN(n9071) );
  MUX2_X1 U11425 ( .A(n8588), .B(n9071), .S(P2_IR_REG_24__SCAN_IN), .Z(n9072)
         );
  INV_X1 U11426 ( .A(P2_B_REG_SCAN_IN), .ZN(n9074) );
  XOR2_X1 U11427 ( .A(n12210), .B(n9074), .Z(n9075) );
  AND2_X1 U11428 ( .A1(n12330), .A2(n9075), .ZN(n9079) );
  INV_X1 U11429 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9077) );
  OR2_X1 U11430 ( .A1(n9095), .A2(P2_D_REG_1__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11431 ( .A1(n14255), .A2(n12330), .ZN(n9080) );
  NAND2_X1 U11432 ( .A1(n9082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11433 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10494), .ZN(n9084) );
  NAND2_X1 U11434 ( .A1(n10964), .A2(n15401), .ZN(n15400) );
  OR2_X1 U11435 ( .A1(n9095), .A2(P2_D_REG_0__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11436 ( .A1(n14255), .A2(n12210), .ZN(n9085) );
  NOR4_X1 U11437 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9090) );
  NOR4_X1 U11438 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9089) );
  NOR4_X1 U11439 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9088) );
  NOR4_X1 U11440 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9087) );
  NAND4_X1 U11441 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9097)
         );
  NOR2_X1 U11442 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9094) );
  NOR4_X1 U11443 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9093) );
  NOR4_X1 U11444 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9092) );
  NOR4_X1 U11445 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9091) );
  NAND4_X1 U11446 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n9096)
         );
  INV_X1 U11447 ( .A(n9095), .ZN(n15395) );
  OAI21_X1 U11448 ( .B1(n9097), .B2(n9096), .A(n15395), .ZN(n10962) );
  NAND2_X1 U11449 ( .A1(n12119), .A2(n10962), .ZN(n9120) );
  INV_X1 U11450 ( .A(n12863), .ZN(n12850) );
  NAND2_X1 U11451 ( .A1(n15380), .A2(n12850), .ZN(n15467) );
  INV_X1 U11452 ( .A(n12862), .ZN(n12925) );
  INV_X1 U11453 ( .A(n10748), .ZN(n9098) );
  AND2_X1 U11454 ( .A1(n15467), .A2(n9098), .ZN(n9099) );
  AND2_X1 U11455 ( .A1(n15380), .A2(n10971), .ZN(n11412) );
  NAND2_X1 U11456 ( .A1(n9105), .A2(n11412), .ZN(n9104) );
  NAND2_X1 U11457 ( .A1(n15380), .A2(n15385), .ZN(n9118) );
  NOR2_X1 U11458 ( .A1(n7344), .A2(n13747), .ZN(n9128) );
  NAND2_X1 U11459 ( .A1(n9105), .A2(n12863), .ZN(n13742) );
  OR2_X1 U11460 ( .A1(n13742), .A2(n15388), .ZN(n13770) );
  NAND2_X1 U11461 ( .A1(n12883), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9114) );
  INV_X1 U11462 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9106) );
  OR2_X1 U11463 ( .A1(n12866), .A2(n9106), .ZN(n9113) );
  INV_X1 U11464 ( .A(n9108), .ZN(n9107) );
  NAND2_X1 U11465 ( .A1(n9107), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13905) );
  INV_X1 U11466 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13697) );
  NAND2_X1 U11467 ( .A1(n9108), .A2(n13697), .ZN(n9109) );
  NAND2_X1 U11468 ( .A1(n13905), .A2(n9109), .ZN(n13947) );
  OR2_X1 U11469 ( .A1(n8721), .A2(n13947), .ZN(n9112) );
  INV_X1 U11470 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9110) );
  OR2_X1 U11471 ( .A1(n12885), .A2(n9110), .ZN(n9111) );
  NAND4_X1 U11472 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9111), .ZN(n13959) );
  INV_X1 U11473 ( .A(n13959), .ZN(n13903) );
  OAI22_X1 U11474 ( .A1(n13770), .A2(n13903), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9115), .ZN(n9116) );
  INV_X1 U11475 ( .A(n9116), .ZN(n9126) );
  INV_X1 U11476 ( .A(n10752), .ZN(n9117) );
  NAND2_X1 U11477 ( .A1(n10748), .A2(n9117), .ZN(n14090) );
  INV_X1 U11478 ( .A(n10964), .ZN(n9119) );
  OAI21_X1 U11479 ( .B1(n9120), .B2(n9119), .A(n9118), .ZN(n9123) );
  NAND2_X1 U11480 ( .A1(n10748), .A2(n12850), .ZN(n10961) );
  INV_X1 U11481 ( .A(n12176), .ZN(n10749) );
  AND2_X1 U11482 ( .A1(n10749), .A2(n10494), .ZN(n9121) );
  NAND2_X1 U11483 ( .A1(n10961), .A2(n9121), .ZN(n12958) );
  INV_X1 U11484 ( .A(n12958), .ZN(n9122) );
  NAND2_X1 U11485 ( .A1(n9123), .A2(n9122), .ZN(n10890) );
  OAI22_X1 U11486 ( .A1(n13759), .A2(n13900), .B1(n13781), .B2(n13953), .ZN(
        n9124) );
  INV_X1 U11487 ( .A(n9124), .ZN(n9125) );
  INV_X1 U11488 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13218) );
  XNOR2_X1 U11489 ( .A(n13218), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n9163) );
  INV_X1 U11490 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9151) );
  INV_X1 U11491 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9149) );
  INV_X1 U11492 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n9317) );
  INV_X1 U11493 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9143) );
  INV_X1 U11494 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9137) );
  NOR2_X1 U11495 ( .A1(n9132), .A2(n9133), .ZN(n9135) );
  INV_X1 U11496 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9290) );
  XOR2_X1 U11497 ( .A(n9290), .B(n9137), .Z(n9183) );
  INV_X1 U11498 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9138) );
  NOR2_X1 U11499 ( .A1(n9139), .A2(n9138), .ZN(n9141) );
  INV_X1 U11500 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15533) );
  XOR2_X1 U11501 ( .A(n15533), .B(n9143), .Z(n9192) );
  XOR2_X1 U11502 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n9195) );
  INV_X1 U11503 ( .A(n9146), .ZN(n9145) );
  NAND2_X1 U11504 ( .A1(n9145), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9147) );
  XOR2_X1 U11505 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n9146), .Z(n9197) );
  XOR2_X1 U11506 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .Z(n9164) );
  XOR2_X1 U11507 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .Z(n9199) );
  AOI21_X2 U11508 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n9151), .A(n9150), .ZN(
        n9202) );
  INV_X1 U11509 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9152) );
  AND2_X1 U11510 ( .A1(n9152), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n9153) );
  INV_X1 U11511 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U11512 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15011), .ZN(n9155) );
  NOR2_X1 U11513 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15011), .ZN(n9159) );
  NAND2_X1 U11514 ( .A1(n9156), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9158) );
  XOR2_X1 U11515 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9156), .Z(n9204) );
  INV_X1 U11516 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13244) );
  NAND2_X1 U11517 ( .A1(n9204), .A2(n13244), .ZN(n9157) );
  NAND2_X1 U11518 ( .A1(n9158), .A2(n9157), .ZN(n9206) );
  XNOR2_X1 U11519 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9206), .ZN(n9207) );
  XNOR2_X1 U11520 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n9207), .ZN(n15006) );
  AOI21_X1 U11521 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15011), .A(n9159), .ZN(
        n9161) );
  XOR2_X1 U11522 ( .A(n9161), .B(n9160), .Z(n15163) );
  XNOR2_X1 U11523 ( .A(n9163), .B(n9162), .ZN(n15159) );
  XOR2_X1 U11524 ( .A(n9165), .B(n9164), .Z(n15146) );
  AND2_X1 U11525 ( .A1(n9177), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9178) );
  INV_X1 U11526 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10877) );
  NOR2_X1 U11527 ( .A1(n9170), .A2(n10877), .ZN(n9171) );
  OAI21_X1 U11528 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9169), .A(n9168), .ZN(
        n15700) );
  NAND2_X1 U11529 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15700), .ZN(n15710) );
  NOR2_X1 U11530 ( .A1(n15710), .A2(n15709), .ZN(n15708) );
  XOR2_X1 U11531 ( .A(n9173), .B(n9172), .Z(n14964) );
  NAND2_X1 U11532 ( .A1(n14965), .A2(n14964), .ZN(n9174) );
  NOR2_X1 U11533 ( .A1(n14965), .A2(n14964), .ZN(n14963) );
  XOR2_X1 U11534 ( .A(n9175), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15705) );
  NOR2_X1 U11535 ( .A1(n15706), .A2(n15705), .ZN(n9176) );
  NAND2_X1 U11536 ( .A1(n15706), .A2(n15705), .ZN(n15704) );
  OAI21_X1 U11537 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n9176), .A(n15704), .ZN(
        n15696) );
  NAND2_X1 U11538 ( .A1(n9180), .A2(n9181), .ZN(n9182) );
  INV_X1 U11539 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15698) );
  INV_X1 U11540 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9185) );
  NOR2_X1 U11541 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  XOR2_X1 U11542 ( .A(n9184), .B(n9183), .Z(n14969) );
  INV_X1 U11543 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9190) );
  NOR2_X1 U11544 ( .A1(n9189), .A2(n9190), .ZN(n9191) );
  XOR2_X1 U11545 ( .A(n9188), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n15703) );
  INV_X1 U11546 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14971) );
  XOR2_X1 U11547 ( .A(n9196), .B(n9195), .Z(n14974) );
  XNOR2_X1 U11548 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n9197), .ZN(n14979) );
  XOR2_X1 U11549 ( .A(n9200), .B(n9199), .Z(n15149) );
  XNOR2_X1 U11550 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n9203) );
  INV_X1 U11551 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15156) );
  NAND2_X1 U11552 ( .A1(n15159), .A2(n15158), .ZN(n15157) );
  XNOR2_X1 U11553 ( .A(n13244), .B(n9204), .ZN(n15167) );
  NAND2_X1 U11554 ( .A1(n15166), .A2(n15167), .ZN(n15165) );
  NAND2_X1 U11555 ( .A1(n15006), .A2(n15005), .ZN(n9205) );
  XNOR2_X1 U11556 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n9210) );
  NOR2_X1 U11557 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9206), .ZN(n9209) );
  INV_X1 U11558 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13275) );
  NOR2_X1 U11559 ( .A1(n13275), .A2(n9207), .ZN(n9208) );
  NOR2_X1 U11560 ( .A1(n9209), .A2(n9208), .ZN(n9213) );
  XNOR2_X1 U11561 ( .A(n9210), .B(n9213), .ZN(n14957) );
  XNOR2_X1 U11562 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9211) );
  INV_X1 U11563 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9214) );
  AND2_X1 U11564 ( .A1(n9214), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n9212) );
  OAI22_X1 U11565 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9214), .B1(n9213), .B2(
        n9212), .ZN(n9215) );
  INV_X1 U11566 ( .A(n9215), .ZN(n9544) );
  OAI22_X1 U11567 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g112), .B1(
        keyinput_g76), .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n9216) );
  AOI221_X1 U11568 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g112), .C1(
        P3_DATAO_REG_20__SCAN_IN), .C2(keyinput_g76), .A(n9216), .ZN(n9223) );
  OAI22_X1 U11569 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        keyinput_g74), .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n9217) );
  AOI221_X1 U11570 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        P3_DATAO_REG_22__SCAN_IN), .C2(keyinput_g74), .A(n9217), .ZN(n9222) );
  OAI22_X1 U11571 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        SI_23_), .B2(keyinput_g9), .ZN(n9218) );
  AOI221_X1 U11572 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        keyinput_g9), .C2(SI_23_), .A(n9218), .ZN(n9221) );
  OAI22_X1 U11573 ( .A1(SI_21_), .A2(keyinput_g11), .B1(SI_19_), .B2(
        keyinput_g13), .ZN(n9219) );
  AOI221_X1 U11574 ( .B1(SI_21_), .B2(keyinput_g11), .C1(keyinput_g13), .C2(
        SI_19_), .A(n9219), .ZN(n9220) );
  NAND4_X1 U11575 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), .ZN(n9252)
         );
  OAI22_X1 U11576 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_g64), .B1(keyinput_g65), .B2(P3_DATAO_REG_31__SCAN_IN), .ZN(n9224) );
  AOI221_X1 U11577 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_g64), .C1(
        P3_DATAO_REG_31__SCAN_IN), .C2(keyinput_g65), .A(n9224), .ZN(n9231) );
  OAI22_X1 U11578 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g72), .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n9225) );
  AOI221_X1 U11579 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P3_DATAO_REG_24__SCAN_IN), .C2(keyinput_g72), .A(n9225), .ZN(n9230) );
  OAI22_X1 U11580 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        keyinput_g101), .B2(P3_ADDR_REG_4__SCAN_IN), .ZN(n9226) );
  AOI221_X1 U11581 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_g101), .A(n9226), .ZN(n9229) );
  OAI22_X1 U11582 ( .A1(SI_16_), .A2(keyinput_g16), .B1(
        P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .ZN(n9227) );
  AOI221_X1 U11583 ( .B1(SI_16_), .B2(keyinput_g16), .C1(keyinput_g69), .C2(
        P3_DATAO_REG_27__SCAN_IN), .A(n9227), .ZN(n9228) );
  NAND4_X1 U11584 ( .A1(n9231), .A2(n9230), .A3(n9229), .A4(n9228), .ZN(n9251)
         );
  OAI22_X1 U11585 ( .A1(SI_15_), .A2(keyinput_g17), .B1(keyinput_g88), .B2(
        P3_DATAO_REG_8__SCAN_IN), .ZN(n9232) );
  AOI221_X1 U11586 ( .B1(SI_15_), .B2(keyinput_g17), .C1(
        P3_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n9232), .ZN(n9239) );
  OAI22_X1 U11587 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g60), .B2(P3_REG3_REG_18__SCAN_IN), .ZN(n9233) );
  AOI221_X1 U11588 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9233), .ZN(n9238) );
  OAI22_X1 U11589 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        keyinput_g113), .B2(P1_IR_REG_6__SCAN_IN), .ZN(n9234) );
  AOI221_X1 U11590 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput_g113), .A(n9234), .ZN(n9237) );
  OAI22_X1 U11591 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        keyinput_g93), .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n9235) );
  AOI221_X1 U11592 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P3_DATAO_REG_3__SCAN_IN), .C2(keyinput_g93), .A(n9235), .ZN(n9236) );
  NAND4_X1 U11593 ( .A1(n9239), .A2(n9238), .A3(n9237), .A4(n9236), .ZN(n9250)
         );
  OAI22_X1 U11594 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_g114), .B1(
        keyinput_g105), .B2(P3_ADDR_REG_8__SCAN_IN), .ZN(n9240) );
  AOI221_X1 U11595 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_g114), .C1(
        P3_ADDR_REG_8__SCAN_IN), .C2(keyinput_g105), .A(n9240), .ZN(n9248) );
  OAI22_X1 U11596 ( .A1(SI_8_), .A2(keyinput_g24), .B1(keyinput_g98), .B2(
        P3_ADDR_REG_1__SCAN_IN), .ZN(n9241) );
  AOI221_X1 U11597 ( .B1(SI_8_), .B2(keyinput_g24), .C1(P3_ADDR_REG_1__SCAN_IN), .C2(keyinput_g98), .A(n9241), .ZN(n9247) );
  OAI22_X1 U11598 ( .A1(SI_13_), .A2(keyinput_g19), .B1(
        P3_DATAO_REG_23__SCAN_IN), .B2(keyinput_g73), .ZN(n9242) );
  AOI221_X1 U11599 ( .B1(SI_13_), .B2(keyinput_g19), .C1(keyinput_g73), .C2(
        P3_DATAO_REG_23__SCAN_IN), .A(n9242), .ZN(n9246) );
  INV_X1 U11600 ( .A(SI_4_), .ZN(n10522) );
  XNOR2_X1 U11601 ( .A(n10522), .B(keyinput_g28), .ZN(n9244) );
  XNOR2_X1 U11602 ( .A(keyinput_g89), .B(P3_DATAO_REG_7__SCAN_IN), .ZN(n9243)
         );
  NOR2_X1 U11603 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  NAND4_X1 U11604 ( .A1(n9248), .A2(n9247), .A3(n9246), .A4(n9245), .ZN(n9249)
         );
  NOR4_X1 U11605 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(n9542)
         );
  OAI22_X1 U11606 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_g111), .ZN(n9253) );
  AOI221_X1 U11607 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g111), .C2(P1_IR_REG_4__SCAN_IN), .A(n9253), .ZN(n9260) );
  OAI22_X1 U11608 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_g110), .ZN(n9254) );
  AOI221_X1 U11609 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        keyinput_g110), .C2(P1_IR_REG_3__SCAN_IN), .A(n9254), .ZN(n9259) );
  OAI22_X1 U11610 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g116), .B2(
        P1_IR_REG_9__SCAN_IN), .ZN(n9255) );
  AOI221_X1 U11611 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P1_IR_REG_9__SCAN_IN), 
        .C2(keyinput_g116), .A(n9255), .ZN(n9258) );
  OAI22_X1 U11612 ( .A1(SI_26_), .A2(keyinput_g6), .B1(P3_ADDR_REG_7__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n9256) );
  AOI221_X1 U11613 ( .B1(SI_26_), .B2(keyinput_g6), .C1(keyinput_g104), .C2(
        P3_ADDR_REG_7__SCAN_IN), .A(n9256), .ZN(n9257) );
  NAND4_X1 U11614 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), .ZN(n9373)
         );
  AOI22_X1 U11615 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n9261) );
  OAI221_X1 U11616 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n9261), .ZN(n9268) );
  AOI22_X1 U11617 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_g92), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9262) );
  OAI221_X1 U11618 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput_g92), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n9262), .ZN(n9267) );
  AOI22_X1 U11619 ( .A1(SI_20_), .A2(keyinput_g12), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n9263) );
  OAI221_X1 U11620 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n9263), .ZN(n9266) );
  AOI22_X1 U11621 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n9264) );
  OAI221_X1 U11622 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        SI_12_), .C2(keyinput_g20), .A(n9264), .ZN(n9265) );
  NOR4_X1 U11623 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .ZN(n9286)
         );
  AOI22_X1 U11624 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n9269) );
  OAI221_X1 U11625 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_24_), .C2(
        keyinput_g8), .A(n9269), .ZN(n9276) );
  AOI22_X1 U11626 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(keyinput_g102), .B1(SI_6_), .B2(keyinput_g26), .ZN(n9270) );
  OAI221_X1 U11627 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_g102), .C1(
        SI_6_), .C2(keyinput_g26), .A(n9270), .ZN(n9275) );
  AOI22_X1 U11628 ( .A1(n14955), .A2(keyinput_g107), .B1(SI_9_), .B2(
        keyinput_g23), .ZN(n9271) );
  OAI221_X1 U11629 ( .B1(n14955), .B2(keyinput_g107), .C1(SI_9_), .C2(
        keyinput_g23), .A(n9271), .ZN(n9274) );
  AOI22_X1 U11630 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P1_IR_REG_20__SCAN_IN), 
        .B2(keyinput_g127), .ZN(n9272) );
  OAI221_X1 U11631 ( .B1(SI_30_), .B2(keyinput_g2), .C1(P1_IR_REG_20__SCAN_IN), 
        .C2(keyinput_g127), .A(n9272), .ZN(n9273) );
  NOR4_X1 U11632 ( .A1(n9276), .A2(n9275), .A3(n9274), .A4(n9273), .ZN(n9285)
         );
  OAI22_X1 U11633 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        keyinput_g32), .B2(SI_0_), .ZN(n9277) );
  AOI221_X1 U11634 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_0_), .C2(keyinput_g32), .A(n9277), .ZN(n9283) );
  OAI22_X1 U11635 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        keyinput_g108), .B2(P1_IR_REG_1__SCAN_IN), .ZN(n9278) );
  AOI221_X1 U11636 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput_g108), .A(n9278), .ZN(n9282) );
  OAI22_X1 U11637 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .ZN(n9279) );
  AOI221_X1 U11638 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        keyinput_g0), .C2(P3_WR_REG_SCAN_IN), .A(n9279), .ZN(n9281) );
  XNOR2_X1 U11639 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g118), .ZN(n9280)
         );
  AND4_X1 U11640 ( .A1(n9283), .A2(n9282), .A3(n9281), .A4(n9280), .ZN(n9284)
         );
  NAND3_X1 U11641 ( .A1(n9286), .A2(n9285), .A3(n9284), .ZN(n9372) );
  INV_X1 U11642 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U11643 ( .A1(n10577), .A2(keyinput_g18), .B1(keyinput_g66), .B2(
        n11296), .ZN(n9287) );
  OAI221_X1 U11644 ( .B1(n10577), .B2(keyinput_g18), .C1(n11296), .C2(
        keyinput_g66), .A(n9287), .ZN(n9295) );
  INV_X1 U11645 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n11253) );
  INV_X1 U11646 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U11647 ( .A1(n11253), .A2(keyinput_g78), .B1(n11248), .B2(
        keyinput_g86), .ZN(n9288) );
  OAI221_X1 U11648 ( .B1(n11253), .B2(keyinput_g78), .C1(n11248), .C2(
        keyinput_g86), .A(n9288), .ZN(n9294) );
  AOI22_X1 U11649 ( .A1(n15590), .A2(keyinput_g59), .B1(keyinput_g103), .B2(
        n9290), .ZN(n9289) );
  OAI221_X1 U11650 ( .B1(n15590), .B2(keyinput_g59), .C1(n9290), .C2(
        keyinput_g103), .A(n9289), .ZN(n9293) );
  INV_X1 U11651 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9474) );
  AOI22_X1 U11652 ( .A1(n9474), .A2(keyinput_g38), .B1(keyinput_g109), .B2(
        n7768), .ZN(n9291) );
  OAI221_X1 U11653 ( .B1(n9474), .B2(keyinput_g38), .C1(n7768), .C2(
        keyinput_g109), .A(n9291), .ZN(n9292) );
  NOR4_X1 U11654 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n9328)
         );
  INV_X1 U11655 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9447) );
  INV_X1 U11656 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U11657 ( .A1(n9447), .A2(keyinput_g41), .B1(keyinput_g70), .B2(
        n11123), .ZN(n9296) );
  OAI221_X1 U11658 ( .B1(n9447), .B2(keyinput_g41), .C1(n11123), .C2(
        keyinput_g70), .A(n9296), .ZN(n9302) );
  INV_X1 U11659 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n10905) );
  INV_X1 U11660 ( .A(SI_27_), .ZN(n12970) );
  AOI22_X1 U11661 ( .A1(n10905), .A2(keyinput_g84), .B1(n12970), .B2(
        keyinput_g5), .ZN(n9297) );
  OAI221_X1 U11662 ( .B1(n10905), .B2(keyinput_g84), .C1(n12970), .C2(
        keyinput_g5), .A(n9297), .ZN(n9301) );
  INV_X1 U11663 ( .A(SI_5_), .ZN(n10529) );
  XNOR2_X1 U11664 ( .A(n10529), .B(keyinput_g27), .ZN(n9300) );
  XNOR2_X1 U11665 ( .A(n9298), .B(keyinput_g121), .ZN(n9299) );
  OR4_X1 U11666 ( .A1(n9302), .A2(n9301), .A3(n9300), .A4(n9299), .ZN(n9305)
         );
  INV_X1 U11667 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14960) );
  XNOR2_X1 U11668 ( .A(n14960), .B(keyinput_g33), .ZN(n9304) );
  INV_X1 U11669 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n11238) );
  XNOR2_X1 U11670 ( .A(n11238), .B(keyinput_g94), .ZN(n9303) );
  NOR3_X1 U11671 ( .A1(n9305), .A2(n9304), .A3(n9303), .ZN(n9327) );
  AOI22_X1 U11672 ( .A1(n9688), .A2(keyinput_g49), .B1(n9749), .B2(
        keyinput_g53), .ZN(n9306) );
  OAI221_X1 U11673 ( .B1(n9688), .B2(keyinput_g49), .C1(n9749), .C2(
        keyinput_g53), .A(n9306), .ZN(n9309) );
  INV_X1 U11674 ( .A(SI_7_), .ZN(n10516) );
  XNOR2_X1 U11675 ( .A(n10516), .B(keyinput_g25), .ZN(n9308) );
  INV_X1 U11676 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n11736) );
  XNOR2_X1 U11677 ( .A(n11736), .B(keyinput_g99), .ZN(n9307) );
  OR3_X1 U11678 ( .A1(n9309), .A2(n9308), .A3(n9307), .ZN(n9314) );
  INV_X1 U11679 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U11680 ( .A1(n11378), .A2(keyinput_g44), .B1(keyinput_g122), .B2(
        n9493), .ZN(n9310) );
  OAI221_X1 U11681 ( .B1(n11378), .B2(keyinput_g44), .C1(n9493), .C2(
        keyinput_g122), .A(n9310), .ZN(n9313) );
  INV_X1 U11682 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n11250) );
  INV_X1 U11683 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U11684 ( .A1(n11250), .A2(keyinput_g80), .B1(keyinput_g87), .B2(
        n11242), .ZN(n9311) );
  OAI221_X1 U11685 ( .B1(n11250), .B2(keyinput_g80), .C1(n11242), .C2(
        keyinput_g87), .A(n9311), .ZN(n9312) );
  NOR3_X1 U11686 ( .A1(n9314), .A2(n9313), .A3(n9312), .ZN(n9326) );
  INV_X1 U11687 ( .A(SI_17_), .ZN(n10696) );
  INV_X1 U11688 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U11689 ( .A1(n10696), .A2(keyinput_g15), .B1(n15505), .B2(
        keyinput_g54), .ZN(n9315) );
  OAI221_X1 U11690 ( .B1(n10696), .B2(keyinput_g15), .C1(n15505), .C2(
        keyinput_g54), .A(n9315), .ZN(n9324) );
  INV_X1 U11691 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U11692 ( .A1(n11263), .A2(keyinput_g96), .B1(n9317), .B2(
        keyinput_g106), .ZN(n9316) );
  OAI221_X1 U11693 ( .B1(n11263), .B2(keyinput_g96), .C1(n9317), .C2(
        keyinput_g106), .A(n9316), .ZN(n9323) );
  INV_X1 U11694 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11919) );
  XOR2_X1 U11695 ( .A(n11919), .B(keyinput_g35), .Z(n9321) );
  XNOR2_X1 U11696 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9320) );
  XNOR2_X1 U11697 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9319) );
  XNOR2_X1 U11698 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g119), .ZN(n9318)
         );
  NAND4_X1 U11699 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(n9322)
         );
  NOR3_X1 U11700 ( .A1(n9324), .A2(n9323), .A3(n9322), .ZN(n9325) );
  NAND4_X1 U11701 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n9371)
         );
  INV_X1 U11702 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n9330) );
  AOI22_X1 U11703 ( .A1(n9330), .A2(keyinput_g39), .B1(keyinput_g4), .B2(
        n12560), .ZN(n9329) );
  OAI221_X1 U11704 ( .B1(n9330), .B2(keyinput_g39), .C1(n12560), .C2(
        keyinput_g4), .A(n9329), .ZN(n9333) );
  INV_X1 U11705 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11298) );
  XNOR2_X1 U11706 ( .A(n11298), .B(keyinput_g67), .ZN(n9332) );
  XOR2_X1 U11707 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g126), .Z(n9331) );
  OR3_X1 U11708 ( .A1(n9333), .A2(n9332), .A3(n9331), .ZN(n9339) );
  INV_X1 U11709 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U11710 ( .A1(n11127), .A2(keyinput_g82), .B1(keyinput_g100), .B2(
        n9335), .ZN(n9334) );
  OAI221_X1 U11711 ( .B1(n11127), .B2(keyinput_g82), .C1(n9335), .C2(
        keyinput_g100), .A(n9334), .ZN(n9338) );
  AOI22_X1 U11712 ( .A1(n8089), .A2(keyinput_g117), .B1(n7771), .B2(
        keyinput_g120), .ZN(n9336) );
  OAI221_X1 U11713 ( .B1(n8089), .B2(keyinput_g117), .C1(n7771), .C2(
        keyinput_g120), .A(n9336), .ZN(n9337) );
  NOR3_X1 U11714 ( .A1(n9339), .A2(n9338), .A3(n9337), .ZN(n9369) );
  INV_X1 U11715 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n11121) );
  INV_X1 U11716 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U11717 ( .A1(n11121), .A2(keyinput_g71), .B1(n11088), .B2(
        keyinput_g75), .ZN(n9340) );
  OAI221_X1 U11718 ( .B1(n11121), .B2(keyinput_g71), .C1(n11088), .C2(
        keyinput_g75), .A(n9340), .ZN(n9343) );
  XOR2_X1 U11719 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_g115), .Z(n9342) );
  INV_X1 U11720 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n11246) );
  XNOR2_X1 U11721 ( .A(n11246), .B(keyinput_g77), .ZN(n9341) );
  OR3_X1 U11722 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(n9348) );
  INV_X1 U11723 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n11232) );
  INV_X1 U11724 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U11725 ( .A1(n11232), .A2(keyinput_g91), .B1(n15506), .B2(
        keyinput_g97), .ZN(n9344) );
  OAI221_X1 U11726 ( .B1(n11232), .B2(keyinput_g91), .C1(n15506), .C2(
        keyinput_g97), .A(n9344), .ZN(n9347) );
  INV_X1 U11727 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U11728 ( .A1(n11244), .A2(keyinput_g81), .B1(n7887), .B2(
        keyinput_g124), .ZN(n9345) );
  OAI221_X1 U11729 ( .B1(n11244), .B2(keyinput_g81), .C1(n7887), .C2(
        keyinput_g124), .A(n9345), .ZN(n9346) );
  NOR3_X1 U11730 ( .A1(n9348), .A2(n9347), .A3(n9346), .ZN(n9368) );
  INV_X1 U11731 ( .A(SI_31_), .ZN(n13668) );
  INV_X1 U11732 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U11733 ( .A1(n13668), .A2(keyinput_g1), .B1(keyinput_g83), .B2(
        n11255), .ZN(n9349) );
  OAI221_X1 U11734 ( .B1(n13668), .B2(keyinput_g1), .C1(n11255), .C2(
        keyinput_g83), .A(n9349), .ZN(n9356) );
  INV_X1 U11735 ( .A(SI_10_), .ZN(n10514) );
  INV_X1 U11736 ( .A(SI_18_), .ZN(n10743) );
  AOI22_X1 U11737 ( .A1(n10514), .A2(keyinput_g22), .B1(n10743), .B2(
        keyinput_g14), .ZN(n9350) );
  OAI221_X1 U11738 ( .B1(n10514), .B2(keyinput_g22), .C1(n10743), .C2(
        keyinput_g14), .A(n9350), .ZN(n9355) );
  INV_X1 U11739 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U11740 ( .A1(n11558), .A2(keyinput_g40), .B1(keyinput_g21), .B2(
        n10519), .ZN(n9351) );
  OAI221_X1 U11741 ( .B1(n11558), .B2(keyinput_g40), .C1(n10519), .C2(
        keyinput_g21), .A(n9351), .ZN(n9354) );
  INV_X1 U11742 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U11743 ( .A1(n11226), .A2(keyinput_g79), .B1(n9880), .B2(
        keyinput_g50), .ZN(n9352) );
  OAI221_X1 U11744 ( .B1(n11226), .B2(keyinput_g79), .C1(n9880), .C2(
        keyinput_g50), .A(n9352), .ZN(n9353) );
  NOR4_X1 U11745 ( .A1(n9356), .A2(n9355), .A3(n9354), .A4(n9353), .ZN(n9367)
         );
  INV_X1 U11746 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U11747 ( .A1(n12643), .A2(keyinput_g3), .B1(keyinput_g95), .B2(
        n11131), .ZN(n9357) );
  OAI221_X1 U11748 ( .B1(n12643), .B2(keyinput_g3), .C1(n11131), .C2(
        keyinput_g95), .A(n9357), .ZN(n9365) );
  INV_X1 U11749 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12264) );
  INV_X1 U11750 ( .A(SI_22_), .ZN(n11185) );
  AOI22_X1 U11751 ( .A1(n12264), .A2(keyinput_g58), .B1(keyinput_g10), .B2(
        n11185), .ZN(n9358) );
  OAI221_X1 U11752 ( .B1(n12264), .B2(keyinput_g58), .C1(n11185), .C2(
        keyinput_g10), .A(n9358), .ZN(n9364) );
  INV_X1 U11753 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n11230) );
  INV_X1 U11754 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11755 ( .A1(n11230), .A2(keyinput_g90), .B1(n9971), .B2(
        keyinput_g47), .ZN(n9359) );
  OAI221_X1 U11756 ( .B1(n11230), .B2(keyinput_g90), .C1(n9971), .C2(
        keyinput_g47), .A(n9359), .ZN(n9363) );
  XNOR2_X1 U11757 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g123), .ZN(n9361)
         );
  XNOR2_X1 U11758 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_g43), .ZN(n9360)
         );
  NAND2_X1 U11759 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  NOR4_X1 U11760 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n9366)
         );
  NAND4_X1 U11761 ( .A1(n9369), .A2(n9368), .A3(n9367), .A4(n9366), .ZN(n9370)
         );
  NOR4_X1 U11762 ( .A1(n9373), .A2(n9372), .A3(n9371), .A4(n9370), .ZN(n9541)
         );
  AOI22_X1 U11763 ( .A1(keyinput_f76), .A2(P3_DATAO_REG_20__SCAN_IN), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n9374) );
  OAI221_X1 U11764 ( .B1(keyinput_f76), .B2(P3_DATAO_REG_20__SCAN_IN), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n9374), .ZN(n9381) );
  AOI22_X1 U11765 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f89), .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n9375) );
  OAI221_X1 U11766 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        keyinput_f89), .C2(P3_DATAO_REG_7__SCAN_IN), .A(n9375), .ZN(n9380) );
  AOI22_X1 U11767 ( .A1(P3_DATAO_REG_19__SCAN_IN), .A2(keyinput_f77), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n9376) );
  OAI221_X1 U11768 ( .B1(P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n9376), .ZN(n9379) );
  AOI22_X1 U11769 ( .A1(keyinput_f92), .A2(P3_DATAO_REG_4__SCAN_IN), .B1(
        keyinput_f80), .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n9377) );
  OAI221_X1 U11770 ( .B1(keyinput_f92), .B2(P3_DATAO_REG_4__SCAN_IN), .C1(
        keyinput_f80), .C2(P3_DATAO_REG_16__SCAN_IN), .A(n9377), .ZN(n9378) );
  NOR4_X1 U11771 ( .A1(n9381), .A2(n9380), .A3(n9379), .A4(n9378), .ZN(n9535)
         );
  OAI22_X1 U11772 ( .A1(SI_13_), .A2(keyinput_f19), .B1(keyinput_f67), .B2(
        P3_DATAO_REG_29__SCAN_IN), .ZN(n9382) );
  AOI221_X1 U11773 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P3_DATAO_REG_29__SCAN_IN), .C2(keyinput_f67), .A(n9382), .ZN(n9389) );
  OAI22_X1 U11774 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput_f98), .B1(
        P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .ZN(n9383) );
  AOI221_X1 U11775 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_f98), .C1(
        keyinput_f87), .C2(P3_DATAO_REG_9__SCAN_IN), .A(n9383), .ZN(n9388) );
  OAI22_X1 U11776 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P1_IR_REG_2__SCAN_IN), 
        .B2(keyinput_f109), .ZN(n9384) );
  AOI221_X1 U11777 ( .B1(SI_3_), .B2(keyinput_f29), .C1(keyinput_f109), .C2(
        P1_IR_REG_2__SCAN_IN), .A(n9384), .ZN(n9387) );
  OAI22_X1 U11778 ( .A1(n14955), .A2(keyinput_f107), .B1(keyinput_f33), .B2(
        P3_RD_REG_SCAN_IN), .ZN(n9385) );
  AOI221_X1 U11779 ( .B1(n14955), .B2(keyinput_f107), .C1(P3_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n9385), .ZN(n9386) );
  NAND4_X1 U11780 ( .A1(n9389), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n9396)
         );
  AOI22_X1 U11781 ( .A1(keyinput_f88), .A2(P3_DATAO_REG_8__SCAN_IN), .B1(
        keyinput_f83), .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n9390) );
  OAI221_X1 U11782 ( .B1(keyinput_f88), .B2(P3_DATAO_REG_8__SCAN_IN), .C1(
        keyinput_f83), .C2(P3_DATAO_REG_13__SCAN_IN), .A(n9390), .ZN(n9395) );
  AOI22_X1 U11783 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_29_), .B2(
        keyinput_f3), .ZN(n9391) );
  OAI221_X1 U11784 ( .B1(SI_10_), .B2(keyinput_f22), .C1(SI_29_), .C2(
        keyinput_f3), .A(n9391), .ZN(n9394) );
  XNOR2_X1 U11785 ( .A(n9392), .B(keyinput_f110), .ZN(n9393) );
  NOR4_X1 U11786 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(n9408)
         );
  OAI22_X1 U11787 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(SI_26_), .B2(keyinput_f6), .ZN(n9397) );
  AOI221_X1 U11788 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f6), .C2(SI_26_), .A(n9397), .ZN(n9407) );
  OAI22_X1 U11789 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n9398) );
  AOI221_X1 U11790 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f35), .C2(P3_REG3_REG_7__SCAN_IN), .A(n9398), .ZN(n9405) );
  OAI22_X1 U11791 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput_f105), .ZN(n9399) );
  AOI221_X1 U11792 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f105), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n9399), .ZN(n9404) );
  OAI22_X1 U11793 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_f101), .B1(
        P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_f104), .ZN(n9400) );
  AOI221_X1 U11794 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f104), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n9400), .ZN(n9403) );
  OAI22_X1 U11795 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f63), .B2(P3_REG3_REG_15__SCAN_IN), .ZN(n9401) );
  AOI221_X1 U11796 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n9401), .ZN(n9402) );
  AND4_X1 U11797 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(n9406)
         );
  AND3_X1 U11798 ( .A1(n9408), .A2(n9407), .A3(n9406), .ZN(n9534) );
  OAI22_X1 U11799 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        keyinput_f123), .B2(P1_IR_REG_16__SCAN_IN), .ZN(n9409) );
  AOI221_X1 U11800 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f123), .A(n9409), .ZN(n9416) );
  OAI22_X1 U11801 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        keyinput_f12), .B2(SI_20_), .ZN(n9410) );
  AOI221_X1 U11802 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        SI_20_), .C2(keyinput_f12), .A(n9410), .ZN(n9415) );
  OAI22_X1 U11803 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_f113), .ZN(n9411) );
  AOI221_X1 U11804 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        keyinput_f113), .C2(P1_IR_REG_6__SCAN_IN), .A(n9411), .ZN(n9414) );
  OAI22_X1 U11805 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f120), .B1(
        P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .ZN(n9412) );
  AOI221_X1 U11806 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f120), .C1(
        keyinput_f86), .C2(P3_DATAO_REG_10__SCAN_IN), .A(n9412), .ZN(n9413) );
  NAND4_X1 U11807 ( .A1(n9416), .A2(n9415), .A3(n9414), .A4(n9413), .ZN(n9444)
         );
  OAI22_X1 U11808 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        keyinput_f75), .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n9417) );
  AOI221_X1 U11809 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        P3_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n9417), .ZN(n9424) );
  OAI22_X1 U11810 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_f121), .B1(
        P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .ZN(n9418) );
  AOI221_X1 U11811 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_f121), .C1(
        keyinput_f74), .C2(P3_DATAO_REG_22__SCAN_IN), .A(n9418), .ZN(n9423) );
  OAI22_X1 U11812 ( .A1(SI_0_), .A2(keyinput_f32), .B1(keyinput_f82), .B2(
        P3_DATAO_REG_14__SCAN_IN), .ZN(n9419) );
  AOI221_X1 U11813 ( .B1(SI_0_), .B2(keyinput_f32), .C1(
        P3_DATAO_REG_14__SCAN_IN), .C2(keyinput_f82), .A(n9419), .ZN(n9422) );
  OAI22_X1 U11814 ( .A1(SI_6_), .A2(keyinput_f26), .B1(keyinput_f111), .B2(
        P1_IR_REG_4__SCAN_IN), .ZN(n9420) );
  AOI221_X1 U11815 ( .B1(SI_6_), .B2(keyinput_f26), .C1(P1_IR_REG_4__SCAN_IN), 
        .C2(keyinput_f111), .A(n9420), .ZN(n9421) );
  NAND4_X1 U11816 ( .A1(n9424), .A2(n9423), .A3(n9422), .A4(n9421), .ZN(n9443)
         );
  OAI22_X1 U11817 ( .A1(keyinput_f65), .A2(P3_DATAO_REG_31__SCAN_IN), .B1(
        keyinput_f93), .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n9425) );
  AOI221_X1 U11818 ( .B1(keyinput_f65), .B2(P3_DATAO_REG_31__SCAN_IN), .C1(
        P3_DATAO_REG_3__SCAN_IN), .C2(keyinput_f93), .A(n9425), .ZN(n9432) );
  OAI22_X1 U11819 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P3_ADDR_REG_6__SCAN_IN), 
        .B2(keyinput_f103), .ZN(n9426) );
  AOI221_X1 U11820 ( .B1(SI_28_), .B2(keyinput_f4), .C1(keyinput_f103), .C2(
        P3_ADDR_REG_6__SCAN_IN), .A(n9426), .ZN(n9431) );
  OAI22_X1 U11821 ( .A1(SI_19_), .A2(keyinput_f13), .B1(
        P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .ZN(n9427) );
  AOI221_X1 U11822 ( .B1(SI_19_), .B2(keyinput_f13), .C1(keyinput_f79), .C2(
        P3_DATAO_REG_17__SCAN_IN), .A(n9427), .ZN(n9430) );
  OAI22_X1 U11823 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f118), .B1(
        keyinput_f95), .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n9428) );
  AOI221_X1 U11824 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f118), .C1(
        P3_DATAO_REG_1__SCAN_IN), .C2(keyinput_f95), .A(n9428), .ZN(n9429) );
  NAND4_X1 U11825 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(n9442)
         );
  OAI22_X1 U11826 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f100), .B2(P3_ADDR_REG_3__SCAN_IN), .ZN(n9433) );
  AOI221_X1 U11827 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P3_ADDR_REG_3__SCAN_IN), .C2(keyinput_f100), .A(n9433), .ZN(n9440) );
  OAI22_X1 U11828 ( .A1(keyinput_f73), .A2(P3_DATAO_REG_23__SCAN_IN), .B1(
        P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_f102), .ZN(n9434) );
  AOI221_X1 U11829 ( .B1(keyinput_f73), .B2(P3_DATAO_REG_23__SCAN_IN), .C1(
        keyinput_f102), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n9434), .ZN(n9439) );
  OAI22_X1 U11830 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        keyinput_f78), .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n9435) );
  AOI221_X1 U11831 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P3_DATAO_REG_18__SCAN_IN), .C2(keyinput_f78), .A(n9435), .ZN(n9438) );
  OAI22_X1 U11832 ( .A1(n11263), .A2(keyinput_f96), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n9436) );
  AOI221_X1 U11833 ( .B1(n11263), .B2(keyinput_f96), .C1(keyinput_f84), .C2(
        P3_DATAO_REG_12__SCAN_IN), .A(n9436), .ZN(n9437) );
  NAND4_X1 U11834 ( .A1(n9440), .A2(n9439), .A3(n9438), .A4(n9437), .ZN(n9441)
         );
  NOR4_X1 U11835 ( .A1(n9444), .A2(n9443), .A3(n9442), .A4(n9441), .ZN(n9533)
         );
  AOI22_X1 U11836 ( .A1(n11736), .A2(keyinput_f99), .B1(P3_U3151), .B2(
        keyinput_f34), .ZN(n9445) );
  OAI221_X1 U11837 ( .B1(n11736), .B2(keyinput_f99), .C1(P3_U3151), .C2(
        keyinput_f34), .A(n9445), .ZN(n9453) );
  AOI22_X1 U11838 ( .A1(n15590), .A2(keyinput_f59), .B1(n9447), .B2(
        keyinput_f41), .ZN(n9446) );
  OAI221_X1 U11839 ( .B1(n15590), .B2(keyinput_f59), .C1(n9447), .C2(
        keyinput_f41), .A(n9446), .ZN(n9452) );
  INV_X1 U11840 ( .A(SI_21_), .ZN(n11267) );
  AOI22_X1 U11841 ( .A1(n11185), .A2(keyinput_f10), .B1(keyinput_f11), .B2(
        n11267), .ZN(n9448) );
  OAI221_X1 U11842 ( .B1(n11185), .B2(keyinput_f10), .C1(n11267), .C2(
        keyinput_f11), .A(n9448), .ZN(n9451) );
  INV_X1 U11843 ( .A(SI_9_), .ZN(n10512) );
  AOI22_X1 U11844 ( .A1(n11244), .A2(keyinput_f81), .B1(n10512), .B2(
        keyinput_f23), .ZN(n9449) );
  OAI221_X1 U11845 ( .B1(n11244), .B2(keyinput_f81), .C1(n10512), .C2(
        keyinput_f23), .A(n9449), .ZN(n9450) );
  NOR4_X1 U11846 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n9472)
         );
  INV_X1 U11847 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U11848 ( .A1(n10519), .A2(keyinput_f21), .B1(n13003), .B2(
        keyinput_f37), .ZN(n9454) );
  OAI221_X1 U11849 ( .B1(n10519), .B2(keyinput_f21), .C1(n13003), .C2(
        keyinput_f37), .A(n9454), .ZN(n9463) );
  AOI22_X1 U11850 ( .A1(n12970), .A2(keyinput_f5), .B1(n11558), .B2(
        keyinput_f40), .ZN(n9455) );
  OAI221_X1 U11851 ( .B1(n12970), .B2(keyinput_f5), .C1(n11558), .C2(
        keyinput_f40), .A(n9455), .ZN(n9462) );
  INV_X1 U11852 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9458) );
  INV_X1 U11853 ( .A(P3_B_REG_SCAN_IN), .ZN(n9457) );
  AOI22_X1 U11854 ( .A1(n9458), .A2(keyinput_f60), .B1(n9457), .B2(
        keyinput_f64), .ZN(n9456) );
  OAI221_X1 U11855 ( .B1(n9458), .B2(keyinput_f60), .C1(n9457), .C2(
        keyinput_f64), .A(n9456), .ZN(n9461) );
  AOI22_X1 U11856 ( .A1(n10577), .A2(keyinput_f18), .B1(n9880), .B2(
        keyinput_f50), .ZN(n9459) );
  OAI221_X1 U11857 ( .B1(n10577), .B2(keyinput_f18), .C1(n9880), .C2(
        keyinput_f50), .A(n9459), .ZN(n9460) );
  NOR4_X1 U11858 ( .A1(n9463), .A2(n9462), .A3(n9461), .A4(n9460), .ZN(n9471)
         );
  INV_X1 U11859 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U11860 ( .A1(n15506), .A2(keyinput_f97), .B1(keyinput_f69), .B2(
        n11259), .ZN(n9464) );
  OAI221_X1 U11861 ( .B1(n15506), .B2(keyinput_f97), .C1(n11259), .C2(
        keyinput_f69), .A(n9464), .ZN(n9469) );
  INV_X1 U11862 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U11863 ( .A1(n9863), .A2(keyinput_f48), .B1(keyinput_f15), .B2(
        n10696), .ZN(n9465) );
  OAI221_X1 U11864 ( .B1(n9863), .B2(keyinput_f48), .C1(n10696), .C2(
        keyinput_f15), .A(n9465), .ZN(n9468) );
  AOI22_X1 U11865 ( .A1(n9731), .A2(keyinput_f43), .B1(keyinput_f7), .B2(
        n12277), .ZN(n9466) );
  OAI221_X1 U11866 ( .B1(n9731), .B2(keyinput_f43), .C1(n12277), .C2(
        keyinput_f7), .A(n9466), .ZN(n9467) );
  NOR3_X1 U11867 ( .A1(n9469), .A2(n9468), .A3(n9467), .ZN(n9470) );
  NAND3_X1 U11868 ( .A1(n9472), .A2(n9471), .A3(n9470), .ZN(n9531) );
  OAI22_X1 U11869 ( .A1(n9474), .A2(keyinput_f38), .B1(n8089), .B2(
        keyinput_f117), .ZN(n9473) );
  AOI221_X1 U11870 ( .B1(n9474), .B2(keyinput_f38), .C1(keyinput_f117), .C2(
        n8089), .A(n9473), .ZN(n9479) );
  INV_X1 U11871 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9916) );
  OAI22_X1 U11872 ( .A1(n9916), .A2(keyinput_f55), .B1(n11123), .B2(
        keyinput_f70), .ZN(n9475) );
  AOI221_X1 U11873 ( .B1(n9916), .B2(keyinput_f55), .C1(keyinput_f70), .C2(
        n11123), .A(n9475), .ZN(n9478) );
  XNOR2_X1 U11874 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f108), .ZN(n9477) );
  XNOR2_X1 U11875 ( .A(keyinput_f0), .B(P3_WR_REG_SCAN_IN), .ZN(n9476) );
  NAND4_X1 U11876 ( .A1(n9479), .A2(n9478), .A3(n9477), .A4(n9476), .ZN(n9530)
         );
  INV_X1 U11877 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n11261) );
  INV_X1 U11878 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U11879 ( .A1(n11261), .A2(keyinput_f72), .B1(n11680), .B2(
        keyinput_f52), .ZN(n9480) );
  OAI221_X1 U11880 ( .B1(n11261), .B2(keyinput_f72), .C1(n11680), .C2(
        keyinput_f52), .A(n9480), .ZN(n9484) );
  XOR2_X1 U11881 ( .A(SI_18_), .B(keyinput_f14), .Z(n9483) );
  XNOR2_X1 U11882 ( .A(n10546), .B(keyinput_f20), .ZN(n9482) );
  XNOR2_X1 U11883 ( .A(keyinput_f44), .B(n11378), .ZN(n9481) );
  OR4_X1 U11884 ( .A1(n9484), .A2(n9483), .A3(n9482), .A4(n9481), .ZN(n9490)
         );
  INV_X1 U11885 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U11886 ( .A1(n11391), .A2(keyinput_f68), .B1(keyinput_f71), .B2(
        n11121), .ZN(n9485) );
  OAI221_X1 U11887 ( .B1(n11391), .B2(keyinput_f68), .C1(n11121), .C2(
        keyinput_f71), .A(n9485), .ZN(n9489) );
  AOI22_X1 U11888 ( .A1(n13668), .A2(keyinput_f1), .B1(keyinput_f90), .B2(
        n11230), .ZN(n9486) );
  OAI221_X1 U11889 ( .B1(n13668), .B2(keyinput_f1), .C1(n11230), .C2(
        keyinput_f90), .A(n9486), .ZN(n9488) );
  INV_X1 U11890 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n11257) );
  XNOR2_X1 U11891 ( .A(n11257), .B(keyinput_f85), .ZN(n9487) );
  OR4_X1 U11892 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n9529)
         );
  AOI22_X1 U11893 ( .A1(n11232), .A2(keyinput_f91), .B1(n11511), .B2(
        keyinput_f9), .ZN(n9491) );
  OAI221_X1 U11894 ( .B1(n11232), .B2(keyinput_f91), .C1(n11511), .C2(
        keyinput_f9), .A(n9491), .ZN(n9495) );
  AOI22_X1 U11895 ( .A1(n9493), .A2(keyinput_f122), .B1(n10693), .B2(
        keyinput_f16), .ZN(n9492) );
  OAI221_X1 U11896 ( .B1(n9493), .B2(keyinput_f122), .C1(n10693), .C2(
        keyinput_f16), .A(n9492), .ZN(n9494) );
  NOR2_X1 U11897 ( .A1(n9495), .A2(n9494), .ZN(n9527) );
  XNOR2_X1 U11898 ( .A(SI_2_), .B(keyinput_f30), .ZN(n9499) );
  XNOR2_X1 U11899 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f114), .ZN(n9498) );
  XNOR2_X1 U11900 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f127), .ZN(n9497)
         );
  XNOR2_X1 U11901 ( .A(SI_15_), .B(keyinput_f17), .ZN(n9496) );
  NAND4_X1 U11902 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n9505)
         );
  XNOR2_X1 U11903 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n9503)
         );
  XNOR2_X1 U11904 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f115), .ZN(n9502) );
  XNOR2_X1 U11905 ( .A(SI_5_), .B(keyinput_f27), .ZN(n9501) );
  XNOR2_X1 U11906 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f126), .ZN(n9500)
         );
  NAND4_X1 U11907 ( .A1(n9503), .A2(n9502), .A3(n9501), .A4(n9500), .ZN(n9504)
         );
  NOR2_X1 U11908 ( .A1(n9505), .A2(n9504), .ZN(n9526) );
  XNOR2_X1 U11909 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_f119), .ZN(n9509)
         );
  XNOR2_X1 U11910 ( .A(SI_30_), .B(keyinput_f2), .ZN(n9508) );
  XNOR2_X1 U11911 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9507) );
  XNOR2_X1 U11912 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9506) );
  NAND4_X1 U11913 ( .A1(n9509), .A2(n9508), .A3(n9507), .A4(n9506), .ZN(n9515)
         );
  XNOR2_X1 U11914 ( .A(SI_8_), .B(keyinput_f24), .ZN(n9513) );
  XNOR2_X1 U11915 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_f116), .ZN(n9512) );
  XNOR2_X1 U11916 ( .A(SI_7_), .B(keyinput_f25), .ZN(n9511) );
  XNOR2_X1 U11917 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f112), .ZN(n9510) );
  NAND4_X1 U11918 ( .A1(n9513), .A2(n9512), .A3(n9511), .A4(n9510), .ZN(n9514)
         );
  NOR2_X1 U11919 ( .A1(n9515), .A2(n9514), .ZN(n9525) );
  INV_X1 U11920 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9517) );
  AOI22_X1 U11921 ( .A1(n11238), .A2(keyinput_f94), .B1(n9517), .B2(
        keyinput_f57), .ZN(n9516) );
  OAI221_X1 U11922 ( .B1(n11238), .B2(keyinput_f94), .C1(n9517), .C2(
        keyinput_f57), .A(n9516), .ZN(n9523) );
  XNOR2_X1 U11923 ( .A(keyinput_f124), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9521)
         );
  XNOR2_X1 U11924 ( .A(keyinput_f49), .B(P3_REG3_REG_5__SCAN_IN), .ZN(n9520)
         );
  XNOR2_X1 U11925 ( .A(keyinput_f8), .B(SI_24_), .ZN(n9519) );
  XNOR2_X1 U11926 ( .A(keyinput_f56), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n9518)
         );
  NAND4_X1 U11927 ( .A1(n9521), .A2(n9520), .A3(n9519), .A4(n9518), .ZN(n9522)
         );
  NOR2_X1 U11928 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NAND4_X1 U11929 ( .A1(n9527), .A2(n9526), .A3(n9525), .A4(n9524), .ZN(n9528)
         );
  NOR4_X1 U11930 ( .A1(n9531), .A2(n9530), .A3(n9529), .A4(n9528), .ZN(n9532)
         );
  NAND4_X1 U11931 ( .A1(n9535), .A2(n9534), .A3(n9533), .A4(n9532), .ZN(n9537)
         );
  AOI21_X1 U11932 ( .B1(keyinput_f125), .B2(n9537), .A(keyinput_g125), .ZN(
        n9539) );
  INV_X1 U11933 ( .A(keyinput_f125), .ZN(n9536) );
  AOI21_X1 U11934 ( .B1(n9537), .B2(n9536), .A(P1_IR_REG_18__SCAN_IN), .ZN(
        n9538) );
  AOI22_X1 U11935 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(n9539), .B1(keyinput_g125), 
        .B2(n9538), .ZN(n9540) );
  AOI21_X1 U11936 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9543) );
  NAND2_X1 U11937 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14245), .ZN(n9585) );
  NOR2_X1 U11938 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7617), .ZN(n9584) );
  NOR2_X1 U11939 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14253), .ZN(n9583) );
  AOI22_X1 U11940 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n12332), .B2(n12329), .ZN(n9967) );
  AOI22_X1 U11941 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12017), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n7203), .ZN(n9924) );
  INV_X1 U11942 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U11943 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11135), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n11133), .ZN(n9887) );
  XNOR2_X1 U11944 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n9870) );
  XNOR2_X1 U11945 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9802) );
  INV_X1 U11946 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U11947 ( .A1(n9653), .A2(n9652), .ZN(n9548) );
  NAND2_X1 U11948 ( .A1(n10496), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U11949 ( .A1(n9548), .A2(n9547), .ZN(n9636) );
  XNOR2_X1 U11950 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9634) );
  NAND2_X1 U11951 ( .A1(n9636), .A2(n9634), .ZN(n9550) );
  NAND2_X1 U11952 ( .A1(n10509), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U11953 ( .A1(n9550), .A2(n9549), .ZN(n9663) );
  XNOR2_X1 U11954 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9661) );
  NAND2_X1 U11955 ( .A1(n9663), .A2(n9661), .ZN(n9552) );
  NAND2_X1 U11956 ( .A1(n7026), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U11957 ( .A1(n9552), .A2(n9551), .ZN(n9678) );
  XNOR2_X1 U11958 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9676) );
  NAND2_X1 U11959 ( .A1(n9678), .A2(n9676), .ZN(n9554) );
  NAND2_X1 U11960 ( .A1(n10540), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U11961 ( .A1(n10544), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U11962 ( .A1(n9557), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U11963 ( .A1(n9745), .A2(n9743), .ZN(n9561) );
  NAND2_X1 U11964 ( .A1(n10572), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U11965 ( .A1(n9561), .A2(n9560), .ZN(n9759) );
  NAND2_X1 U11966 ( .A1(n9759), .A2(n9758), .ZN(n9564) );
  NAND2_X1 U11967 ( .A1(n9562), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U11968 ( .A1(n9564), .A2(n9563), .ZN(n9771) );
  NAND2_X1 U11969 ( .A1(n9771), .A2(n9770), .ZN(n9566) );
  NAND2_X1 U11970 ( .A1(n10653), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U11971 ( .A1(n10689), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U11972 ( .A1(n10790), .A2(n9568), .ZN(n9569) );
  XNOR2_X1 U11973 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9824) );
  INV_X1 U11974 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10941) );
  NAND2_X1 U11975 ( .A1(n10941), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9570) );
  XNOR2_X1 U11976 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9837) );
  XNOR2_X1 U11977 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9853) );
  NAND2_X1 U11978 ( .A1(n9855), .A2(n9853), .ZN(n9573) );
  NAND2_X1 U11979 ( .A1(n9571), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U11980 ( .A1(n9887), .A2(n9889), .ZN(n9575) );
  AOI22_X1 U11981 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12967), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n9576), .ZN(n9899) );
  NAND2_X1 U11982 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n9578), .ZN(n9579) );
  INV_X1 U11983 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9580) );
  AOI22_X1 U11984 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12040), .B2(n9580), .ZN(n9935) );
  AOI22_X1 U11985 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n12178), .B2(n12182), .ZN(n9945) );
  INV_X1 U11986 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14240) );
  AOI22_X1 U11987 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n14240), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14944), .ZN(n10017) );
  INV_X1 U11988 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U11989 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12859), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n12639), .ZN(n9618) );
  XNOR2_X1 U11990 ( .A(n9619), .B(n9618), .ZN(n12972) );
  NOR2_X1 U11991 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n9591) );
  NOR2_X1 U11992 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n9590) );
  NOR2_X1 U11993 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n9589) );
  NAND4_X1 U11994 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n9593)
         );
  NAND2_X1 U11995 ( .A1(n12972), .A2(n9805), .ZN(n9601) );
  NAND2_X1 U11996 ( .A1(n9651), .A2(SI_30_), .ZN(n9600) );
  NAND2_X1 U11997 ( .A1(n9689), .A2(n9688), .ZN(n9704) );
  OR2_X2 U11998 ( .A1(n9777), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9792) );
  INV_X1 U11999 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U12000 ( .A1(n9972), .A2(n9971), .ZN(n9983) );
  INV_X1 U12001 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13034) );
  NOR2_X1 U12002 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), 
        .ZN(n9607) );
  INV_X1 U12003 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9603) );
  AND2_X1 U12004 ( .A1(n9607), .A2(n9603), .ZN(n9604) );
  NAND2_X1 U12005 ( .A1(n10217), .A2(n9607), .ZN(n9608) );
  NAND2_X1 U12006 ( .A1(n9608), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U12007 ( .A1(n15030), .A2(n9816), .ZN(n10027) );
  INV_X1 U12008 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9615) );
  AND2_X2 U12009 ( .A1(n9612), .A2(n12641), .ZN(n9646) );
  NAND2_X1 U12010 ( .A1(n9646), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U12011 ( .A1(n9847), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9613) );
  OAI211_X1 U12012 ( .C1(n6994), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9616)
         );
  INV_X1 U12013 ( .A(n9616), .ZN(n9617) );
  NOR2_X1 U12014 ( .A1(n15040), .A2(n12545), .ZN(n10208) );
  OAI21_X1 U12015 ( .B1(n12639), .B2(P1_DATAO_REG_30__SCAN_IN), .A(n9620), 
        .ZN(n9623) );
  INV_X1 U12016 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10585) );
  INV_X1 U12017 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9621) );
  AOI22_X1 U12018 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n10585), .B2(n9621), .ZN(n9622) );
  INV_X1 U12019 ( .A(n15036), .ZN(n15031) );
  INV_X1 U12020 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U12021 ( .A1(n10000), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U12022 ( .A1(n9847), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9624) );
  OAI211_X1 U12023 ( .C1(n6994), .C2(n9626), .A(n9625), .B(n9624), .ZN(n9627)
         );
  INV_X1 U12024 ( .A(n9627), .ZN(n9628) );
  NAND2_X1 U12025 ( .A1(n10027), .A2(n9628), .ZN(n15029) );
  NAND2_X1 U12026 ( .A1(n9951), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12027 ( .A1(n9816), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U12028 ( .A1(n9847), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9629) );
  INV_X1 U12029 ( .A(n9634), .ZN(n9635) );
  XNOR2_X1 U12030 ( .A(n9636), .B(n9635), .ZN(n10521) );
  NAND2_X1 U12031 ( .A1(n9651), .A2(n7242), .ZN(n9637) );
  INV_X1 U12032 ( .A(n11495), .ZN(n9655) );
  NAND2_X1 U12033 ( .A1(n9951), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U12034 ( .A1(n9646), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12035 ( .A1(n9847), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9638) );
  INV_X1 U12036 ( .A(n9652), .ZN(n9644) );
  INV_X1 U12037 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U12038 ( .A1(n9642), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9643) );
  NAND2_X1 U12039 ( .A1(n9644), .A2(n9643), .ZN(n10531) );
  NAND2_X1 U12040 ( .A1(n9651), .A2(SI_0_), .ZN(n9645) );
  INV_X1 U12041 ( .A(n11366), .ZN(n12637) );
  INV_X1 U12042 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11534) );
  INV_X1 U12043 ( .A(n9633), .ZN(n9650) );
  NAND2_X1 U12044 ( .A1(n9651), .A2(SI_1_), .ZN(n9654) );
  XNOR2_X1 U12045 ( .A(n9653), .B(n9652), .ZN(n10503) );
  NAND2_X1 U12046 ( .A1(n11368), .A2(n10078), .ZN(n15587) );
  NAND2_X1 U12047 ( .A1(n9655), .A2(n15587), .ZN(n9656) );
  INV_X1 U12048 ( .A(n15612), .ZN(n12041) );
  NAND2_X1 U12049 ( .A1(n12041), .A2(n11393), .ZN(n10086) );
  NAND2_X1 U12050 ( .A1(n9646), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U12051 ( .A1(n9816), .A2(n11558), .ZN(n9659) );
  NAND2_X1 U12052 ( .A1(n9847), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9658) );
  INV_X1 U12053 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11545) );
  OR2_X1 U12054 ( .A1(n10024), .A2(n11545), .ZN(n9657) );
  INV_X1 U12055 ( .A(SI_3_), .ZN(n10524) );
  NAND2_X1 U12056 ( .A1(n9651), .A2(n10524), .ZN(n9669) );
  INV_X1 U12057 ( .A(n9661), .ZN(n9662) );
  XNOR2_X1 U12058 ( .A(n9663), .B(n9662), .ZN(n10525) );
  NAND2_X1 U12059 ( .A1(n9805), .A2(n10525), .ZN(n9668) );
  NAND2_X1 U12060 ( .A1(n9664), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9665) );
  MUX2_X1 U12061 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9665), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n9666) );
  AND2_X1 U12062 ( .A1(n9666), .A2(n9679), .ZN(n11588) );
  OR2_X1 U12063 ( .A1(n10229), .A2(n11588), .ZN(n9667) );
  NAND2_X1 U12064 ( .A1(n15596), .A2(n12045), .ZN(n10087) );
  INV_X1 U12065 ( .A(n12045), .ZN(n12115) );
  NAND2_X1 U12066 ( .A1(n11478), .A2(n11502), .ZN(n9670) );
  NAND2_X1 U12067 ( .A1(n10000), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9675) );
  OR2_X1 U12068 ( .A1(n7755), .A2(n9689), .ZN(n15582) );
  NAND2_X1 U12069 ( .A1(n9816), .A2(n15582), .ZN(n9674) );
  NAND2_X1 U12070 ( .A1(n9847), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9673) );
  INV_X1 U12071 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9671) );
  OR2_X1 U12072 ( .A1(n10024), .A2(n9671), .ZN(n9672) );
  NAND2_X1 U12073 ( .A1(n9651), .A2(n10522), .ZN(n9686) );
  INV_X1 U12074 ( .A(n9676), .ZN(n9677) );
  XNOR2_X1 U12075 ( .A(n9678), .B(n9677), .ZN(n10523) );
  NAND2_X1 U12076 ( .A1(n9805), .A2(n10523), .ZN(n9685) );
  NAND2_X1 U12077 ( .A1(n9679), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U12078 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9680), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9683) );
  INV_X1 U12079 ( .A(n9681), .ZN(n9682) );
  OR2_X1 U12080 ( .A1(n10229), .A2(n11596), .ZN(n9684) );
  NAND2_X1 U12081 ( .A1(n12094), .A2(n15581), .ZN(n10095) );
  INV_X1 U12082 ( .A(n15581), .ZN(n12102) );
  INV_X1 U12083 ( .A(n15576), .ZN(n10045) );
  NAND2_X1 U12084 ( .A1(n15572), .A2(n10045), .ZN(n9687) );
  NAND2_X1 U12085 ( .A1(n10000), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9695) );
  OR2_X1 U12086 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  NAND2_X1 U12087 ( .A1(n9704), .A2(n9690), .ZN(n15568) );
  NAND2_X1 U12088 ( .A1(n9816), .A2(n15568), .ZN(n9694) );
  NAND2_X1 U12089 ( .A1(n9847), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9693) );
  INV_X1 U12090 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9691) );
  OR2_X1 U12091 ( .A1(n6994), .A2(n9691), .ZN(n9692) );
  NAND2_X1 U12092 ( .A1(n9651), .A2(n10529), .ZN(n9703) );
  XNOR2_X1 U12093 ( .A(n6979), .B(n7218), .ZN(n10530) );
  NAND2_X1 U12094 ( .A1(n9805), .A2(n10530), .ZN(n9702) );
  NOR2_X1 U12095 ( .A1(n9681), .A2(n10225), .ZN(n9698) );
  MUX2_X1 U12096 ( .A(n10225), .B(n9698), .S(P3_IR_REG_5__SCAN_IN), .Z(n9700)
         );
  OR2_X1 U12097 ( .A1(n9700), .A2(n9699), .ZN(n11598) );
  INV_X1 U12098 ( .A(n11598), .ZN(n11606) );
  OR2_X1 U12099 ( .A1(n10229), .A2(n11606), .ZN(n9701) );
  NAND2_X1 U12100 ( .A1(n12051), .A2(n15567), .ZN(n10100) );
  INV_X1 U12101 ( .A(n15567), .ZN(n12090) );
  NAND2_X1 U12102 ( .A1(n15574), .A2(n12090), .ZN(n10096) );
  NAND2_X1 U12103 ( .A1(n9646), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U12104 ( .A1(n9704), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U12105 ( .A1(n9717), .A2(n9705), .ZN(n12067) );
  NAND2_X1 U12106 ( .A1(n9816), .A2(n12067), .ZN(n9709) );
  NAND2_X1 U12107 ( .A1(n9847), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9708) );
  INV_X1 U12108 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9706) );
  OR2_X1 U12109 ( .A1(n6994), .A2(n9706), .ZN(n9707) );
  OR2_X1 U12110 ( .A1(n9699), .A2(n10225), .ZN(n9711) );
  XNOR2_X1 U12111 ( .A(n9711), .B(n9723), .ZN(n11863) );
  NAND2_X1 U12112 ( .A1(n9651), .A2(SI_6_), .ZN(n9715) );
  XNOR2_X1 U12113 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9712) );
  XNOR2_X1 U12114 ( .A(n9713), .B(n9712), .ZN(n10526) );
  NAND2_X1 U12115 ( .A1(n9805), .A2(n10526), .ZN(n9714) );
  OAI211_X1 U12116 ( .C1(n10229), .C2(n11863), .A(n9715), .B(n9714), .ZN(
        n15649) );
  NAND2_X1 U12117 ( .A1(n12054), .A2(n15649), .ZN(n10107) );
  INV_X1 U12118 ( .A(n15649), .ZN(n12072) );
  NAND2_X1 U12119 ( .A1(n15562), .A2(n12072), .ZN(n10101) );
  NAND2_X1 U12120 ( .A1(n10107), .A2(n10101), .ZN(n11724) );
  INV_X1 U12121 ( .A(n11724), .ZN(n10043) );
  NAND2_X1 U12122 ( .A1(n11719), .A2(n10043), .ZN(n9716) );
  INV_X1 U12123 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11860) );
  OR2_X1 U12124 ( .A1(n10024), .A2(n11860), .ZN(n9722) );
  NAND2_X1 U12125 ( .A1(n10000), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9721) );
  AND2_X1 U12126 ( .A1(n9717), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9718) );
  OR2_X1 U12127 ( .A1(n9718), .A2(n9732), .ZN(n12077) );
  NAND2_X1 U12128 ( .A1(n9816), .A2(n12077), .ZN(n9720) );
  NAND2_X1 U12129 ( .A1(n9847), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9719) );
  NAND4_X1 U12130 ( .A1(n9722), .A2(n9721), .A3(n9720), .A4(n9719), .ZN(n12169) );
  NAND2_X1 U12131 ( .A1(n9699), .A2(n9723), .ZN(n9739) );
  NAND2_X1 U12132 ( .A1(n9739), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9725) );
  INV_X1 U12133 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9724) );
  XNOR2_X1 U12134 ( .A(n9725), .B(n9724), .ZN(n11926) );
  INV_X1 U12135 ( .A(n11926), .ZN(n11861) );
  XNOR2_X1 U12136 ( .A(n9727), .B(n9726), .ZN(n10517) );
  NAND2_X1 U12137 ( .A1(n9805), .A2(n10517), .ZN(n9729) );
  NAND2_X1 U12138 ( .A1(n9651), .A2(n10516), .ZN(n9728) );
  OAI211_X1 U12139 ( .C1(n11861), .C2(n10229), .A(n9729), .B(n9728), .ZN(
        n12083) );
  INV_X1 U12140 ( .A(n12057), .ZN(n11957) );
  INV_X1 U12141 ( .A(n12169), .ZN(n10111) );
  INV_X1 U12142 ( .A(n12083), .ZN(n12161) );
  NAND2_X1 U12143 ( .A1(n10111), .A2(n12161), .ZN(n9730) );
  NAND2_X1 U12144 ( .A1(n10000), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9738) );
  NOR2_X1 U12145 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  OR2_X1 U12146 ( .A1(n9750), .A2(n9733), .ZN(n12173) );
  NAND2_X1 U12147 ( .A1(n9816), .A2(n12173), .ZN(n9737) );
  NAND2_X1 U12148 ( .A1(n9847), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9736) );
  INV_X1 U12149 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9734) );
  OR2_X1 U12150 ( .A1(n6994), .A2(n9734), .ZN(n9735) );
  NAND2_X1 U12151 ( .A1(n9741), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9740) );
  MUX2_X1 U12152 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9740), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n9742) );
  NAND2_X1 U12153 ( .A1(n9742), .A2(n9772), .ZN(n15522) );
  NAND2_X1 U12154 ( .A1(n9651), .A2(SI_8_), .ZN(n9747) );
  INV_X1 U12155 ( .A(n9743), .ZN(n9744) );
  XNOR2_X1 U12156 ( .A(n9745), .B(n9744), .ZN(n10534) );
  NAND2_X1 U12157 ( .A1(n9805), .A2(n10534), .ZN(n9746) );
  OAI211_X1 U12158 ( .C1(n10229), .C2(n15522), .A(n9747), .B(n9746), .ZN(n9748) );
  NAND2_X1 U12159 ( .A1(n12215), .A2(n9748), .ZN(n10117) );
  INV_X1 U12160 ( .A(n9748), .ZN(n12214) );
  NAND2_X1 U12161 ( .A1(n12220), .A2(n12214), .ZN(n10116) );
  INV_X1 U12162 ( .A(n12213), .ZN(n9762) );
  NAND2_X1 U12163 ( .A1(n10000), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9756) );
  OR2_X1 U12164 ( .A1(n9750), .A2(n9749), .ZN(n9751) );
  NAND2_X1 U12165 ( .A1(n9764), .A2(n9751), .ZN(n12224) );
  NAND2_X1 U12166 ( .A1(n9816), .A2(n12224), .ZN(n9755) );
  NAND2_X1 U12167 ( .A1(n9847), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9754) );
  INV_X1 U12168 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9752) );
  OR2_X1 U12169 ( .A1(n6994), .A2(n9752), .ZN(n9753) );
  NAND2_X1 U12170 ( .A1(n9772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9757) );
  XNOR2_X1 U12171 ( .A(n9757), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11997) );
  NAND2_X1 U12172 ( .A1(n9651), .A2(n10512), .ZN(n9761) );
  XNOR2_X1 U12173 ( .A(n9759), .B(n9758), .ZN(n10513) );
  NAND2_X1 U12174 ( .A1(n9805), .A2(n10513), .ZN(n9760) );
  OAI211_X1 U12175 ( .C1(n11997), .C2(n10229), .A(n9761), .B(n9760), .ZN(
        n12223) );
  NAND2_X1 U12176 ( .A1(n12305), .A2(n12223), .ZN(n9763) );
  NAND2_X1 U12177 ( .A1(n9646), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9769) );
  NAND2_X1 U12178 ( .A1(n9764), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U12179 ( .A1(n9777), .A2(n9765), .ZN(n12242) );
  NAND2_X1 U12180 ( .A1(n9816), .A2(n12242), .ZN(n9768) );
  NAND2_X1 U12181 ( .A1(n9847), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9767) );
  INV_X1 U12182 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12000) );
  OR2_X1 U12183 ( .A1(n6994), .A2(n12000), .ZN(n9766) );
  XNOR2_X1 U12184 ( .A(n9771), .B(n9770), .ZN(n10515) );
  NAND2_X1 U12185 ( .A1(n9805), .A2(n10515), .ZN(n9776) );
  NAND2_X1 U12186 ( .A1(n9651), .A2(n10514), .ZN(n9775) );
  NOR2_X1 U12187 ( .A1(n9772), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9784) );
  OR2_X1 U12188 ( .A1(n9784), .A2(n10225), .ZN(n9773) );
  XNOR2_X1 U12189 ( .A(n9773), .B(P3_IR_REG_10__SCAN_IN), .ZN(n12007) );
  OR2_X1 U12190 ( .A1(n10229), .A2(n12007), .ZN(n9774) );
  INV_X1 U12191 ( .A(n12442), .ZN(n12252) );
  NAND2_X1 U12192 ( .A1(n12563), .A2(n12252), .ZN(n10124) );
  NAND2_X1 U12193 ( .A1(n13116), .A2(n12442), .ZN(n12456) );
  NAND2_X1 U12194 ( .A1(n9847), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U12195 ( .A1(n9777), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U12196 ( .A1(n9792), .A2(n9778), .ZN(n12462) );
  NAND2_X1 U12197 ( .A1(n9816), .A2(n12462), .ZN(n9781) );
  NAND2_X1 U12198 ( .A1(n10000), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9780) );
  INV_X1 U12199 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12259) );
  OR2_X1 U12200 ( .A1(n6994), .A2(n12259), .ZN(n9779) );
  NAND2_X1 U12201 ( .A1(n9784), .A2(n9783), .ZN(n9785) );
  NAND2_X1 U12202 ( .A1(n9785), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9786) );
  XNOR2_X1 U12203 ( .A(n9786), .B(P3_IR_REG_11__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U12204 ( .A1(n9651), .A2(n10519), .ZN(n9790) );
  XNOR2_X1 U12205 ( .A(n9788), .B(n9787), .ZN(n10520) );
  NAND2_X1 U12206 ( .A1(n9805), .A2(n10520), .ZN(n9789) );
  OAI211_X1 U12207 ( .C1(n13190), .C2(n10229), .A(n9790), .B(n9789), .ZN(
        n15056) );
  INV_X1 U12208 ( .A(n15056), .ZN(n13118) );
  NAND2_X1 U12209 ( .A1(n13055), .A2(n13118), .ZN(n10128) );
  AND2_X1 U12210 ( .A1(n12456), .A2(n10128), .ZN(n9791) );
  NAND2_X1 U12211 ( .A1(n12457), .A2(n9791), .ZN(n12449) );
  NAND2_X1 U12212 ( .A1(n9646), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9797) );
  AND2_X1 U12213 ( .A1(n9792), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9793) );
  OR2_X1 U12214 ( .A1(n9793), .A2(n9817), .ZN(n13050) );
  NAND2_X1 U12215 ( .A1(n9816), .A2(n13050), .ZN(n9796) );
  NAND2_X1 U12216 ( .A1(n9847), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9795) );
  OR2_X1 U12217 ( .A1(n6994), .A2(n15055), .ZN(n9794) );
  NAND2_X1 U12218 ( .A1(n9798), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9799) );
  MUX2_X1 U12219 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9799), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9801) );
  INV_X1 U12220 ( .A(n9800), .ZN(n9811) );
  NAND2_X1 U12221 ( .A1(n9801), .A2(n9811), .ZN(n15534) );
  INV_X1 U12222 ( .A(n9802), .ZN(n9803) );
  XNOR2_X1 U12223 ( .A(n9804), .B(n9803), .ZN(n10545) );
  NAND2_X1 U12224 ( .A1(n9805), .A2(n10545), .ZN(n9807) );
  NAND2_X1 U12225 ( .A1(n9651), .A2(SI_12_), .ZN(n9806) );
  OAI211_X1 U12226 ( .C1(n10229), .C2(n15534), .A(n9807), .B(n9806), .ZN(
        n13057) );
  NAND2_X1 U12227 ( .A1(n13531), .A2(n13057), .ZN(n10132) );
  INV_X1 U12228 ( .A(n13057), .ZN(n12571) );
  NAND2_X1 U12229 ( .A1(n13114), .A2(n12571), .ZN(n10131) );
  NAND2_X1 U12230 ( .A1(n10132), .A2(n10131), .ZN(n12473) );
  NAND2_X1 U12231 ( .A1(n13111), .A2(n15056), .ZN(n12448) );
  AND2_X1 U12232 ( .A1(n12450), .A2(n12448), .ZN(n9808) );
  NAND2_X1 U12233 ( .A1(n12449), .A2(n9808), .ZN(n9809) );
  XNOR2_X1 U12234 ( .A(n9810), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U12235 ( .A1(n10570), .A2(n9805), .ZN(n9814) );
  NAND2_X1 U12236 ( .A1(n9811), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9812) );
  XNOR2_X1 U12237 ( .A(n9812), .B(P3_IR_REG_13__SCAN_IN), .ZN(n13204) );
  INV_X1 U12238 ( .A(n13204), .ZN(n13209) );
  AOI22_X1 U12239 ( .A1(n9651), .A2(n10569), .B1(n11530), .B2(n13209), .ZN(
        n9813) );
  NAND2_X1 U12240 ( .A1(n9814), .A2(n9813), .ZN(n15046) );
  INV_X1 U12241 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9815) );
  OR2_X1 U12242 ( .A1(n6994), .A2(n9815), .ZN(n9822) );
  NAND2_X1 U12243 ( .A1(n9847), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9821) );
  OR2_X1 U12244 ( .A1(n9817), .A2(n13096), .ZN(n9818) );
  NAND2_X1 U12245 ( .A1(n9829), .A2(n9818), .ZN(n13533) );
  NAND2_X1 U12246 ( .A1(n9816), .A2(n13533), .ZN(n9820) );
  NAND2_X1 U12247 ( .A1(n10000), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9819) );
  NAND4_X1 U12248 ( .A1(n9822), .A2(n9821), .A3(n9820), .A4(n9819), .ZN(n13052) );
  OR2_X1 U12249 ( .A1(n15046), .A2(n13052), .ZN(n10138) );
  INV_X1 U12250 ( .A(n10138), .ZN(n9823) );
  NAND2_X1 U12251 ( .A1(n15046), .A2(n13052), .ZN(n10137) );
  XNOR2_X1 U12252 ( .A(n9825), .B(n9824), .ZN(n10578) );
  NAND2_X1 U12253 ( .A1(n10578), .A2(n9805), .ZN(n9828) );
  NAND2_X1 U12254 ( .A1(n9840), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9826) );
  XNOR2_X1 U12255 ( .A(n9826), .B(n7396), .ZN(n13207) );
  AOI22_X1 U12256 ( .A1(n9651), .A2(n10577), .B1(n11530), .B2(n13207), .ZN(
        n9827) );
  NAND2_X1 U12257 ( .A1(n9828), .A2(n9827), .ZN(n13010) );
  NAND2_X1 U12258 ( .A1(n9951), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U12259 ( .A1(n10000), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U12260 ( .A1(n9829), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12261 ( .A1(n9844), .A2(n9830), .ZN(n13007) );
  NAND2_X1 U12262 ( .A1(n9816), .A2(n13007), .ZN(n9832) );
  NAND2_X1 U12263 ( .A1(n9847), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9831) );
  NAND4_X1 U12264 ( .A1(n9834), .A2(n9833), .A3(n9832), .A4(n9831), .ZN(n13097) );
  NAND2_X1 U12265 ( .A1(n13010), .A2(n13097), .ZN(n10143) );
  OR2_X1 U12266 ( .A1(n13010), .A2(n13097), .ZN(n10142) );
  INV_X1 U12267 ( .A(n9837), .ZN(n9838) );
  XNOR2_X1 U12268 ( .A(n9839), .B(n9838), .ZN(n10646) );
  NAND2_X1 U12269 ( .A1(n10646), .A2(n9805), .ZN(n9843) );
  OR2_X1 U12270 ( .A1(n9857), .A2(n10225), .ZN(n9841) );
  XNOR2_X1 U12271 ( .A(n9841), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U12272 ( .A1(n9651), .A2(SI_15_), .B1(n11530), .B2(n13248), .ZN(
        n9842) );
  NAND2_X1 U12273 ( .A1(n9843), .A2(n9842), .ZN(n13144) );
  INV_X1 U12274 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15015) );
  OR2_X1 U12275 ( .A1(n6994), .A2(n15015), .ZN(n9851) );
  NAND2_X1 U12276 ( .A1(n10000), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9850) );
  INV_X1 U12277 ( .A(n9864), .ZN(n9846) );
  NAND2_X1 U12278 ( .A1(n9844), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U12279 ( .A1(n9846), .A2(n9845), .ZN(n13520) );
  NAND2_X1 U12280 ( .A1(n9816), .A2(n13520), .ZN(n9849) );
  NAND2_X1 U12281 ( .A1(n9847), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9848) );
  NAND4_X1 U12282 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(n13503) );
  INV_X1 U12283 ( .A(n13503), .ZN(n13072) );
  OR2_X1 U12284 ( .A1(n13144), .A2(n13072), .ZN(n10146) );
  NAND2_X1 U12285 ( .A1(n13144), .A2(n13072), .ZN(n10150) );
  NAND2_X1 U12286 ( .A1(n13519), .A2(n13518), .ZN(n9852) );
  INV_X1 U12287 ( .A(n9853), .ZN(n9854) );
  XNOR2_X1 U12288 ( .A(n9855), .B(n9854), .ZN(n10692) );
  NAND2_X1 U12289 ( .A1(n10692), .A2(n9805), .ZN(n9862) );
  NAND2_X1 U12290 ( .A1(n9859), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9858) );
  MUX2_X1 U12291 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9858), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9860) );
  AND2_X1 U12292 ( .A1(n9860), .A2(n9873), .ZN(n13251) );
  AOI22_X1 U12293 ( .A1(n9651), .A2(SI_16_), .B1(n11530), .B2(n13251), .ZN(
        n9861) );
  NAND2_X1 U12294 ( .A1(n9862), .A2(n9861), .ZN(n13067) );
  NAND2_X1 U12295 ( .A1(n10000), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9869) );
  NOR2_X1 U12296 ( .A1(n9864), .A2(n9863), .ZN(n9865) );
  OR2_X1 U12297 ( .A1(n9881), .A2(n9865), .ZN(n13510) );
  NAND2_X1 U12298 ( .A1(n9816), .A2(n13510), .ZN(n9868) );
  NAND2_X1 U12299 ( .A1(n9847), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9867) );
  INV_X1 U12300 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13599) );
  OR2_X1 U12301 ( .A1(n6994), .A2(n13599), .ZN(n9866) );
  OR2_X1 U12302 ( .A1(n13067), .A2(n13517), .ZN(n10145) );
  NAND2_X1 U12303 ( .A1(n13067), .A2(n13517), .ZN(n13492) );
  INV_X1 U12304 ( .A(n9870), .ZN(n9871) );
  XNOR2_X1 U12305 ( .A(n9872), .B(n9871), .ZN(n10695) );
  NAND2_X1 U12306 ( .A1(n10695), .A2(n9805), .ZN(n9879) );
  NAND2_X1 U12307 ( .A1(n9873), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U12308 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9874), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9877) );
  NAND2_X1 U12309 ( .A1(n9877), .A2(n9901), .ZN(n13288) );
  INV_X1 U12310 ( .A(n13288), .ZN(n13299) );
  AOI22_X1 U12311 ( .A1(n9651), .A2(SI_17_), .B1(n11530), .B2(n13299), .ZN(
        n9878) );
  NAND2_X1 U12312 ( .A1(n9879), .A2(n9878), .ZN(n13076) );
  NAND2_X1 U12313 ( .A1(n10000), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9886) );
  OR2_X1 U12314 ( .A1(n9881), .A2(n9880), .ZN(n9882) );
  NAND2_X1 U12315 ( .A1(n9893), .A2(n9882), .ZN(n13494) );
  NAND2_X1 U12316 ( .A1(n9816), .A2(n13494), .ZN(n9885) );
  NAND2_X1 U12317 ( .A1(n9847), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9884) );
  INV_X1 U12318 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13595) );
  OR2_X1 U12319 ( .A1(n6994), .A2(n13595), .ZN(n9883) );
  NAND2_X1 U12320 ( .A1(n13076), .A2(n13128), .ZN(n10157) );
  OR2_X1 U12321 ( .A1(n13076), .A2(n13128), .ZN(n10162) );
  INV_X1 U12322 ( .A(n9887), .ZN(n9888) );
  XNOR2_X1 U12323 ( .A(n9889), .B(n9888), .ZN(n10742) );
  NAND2_X1 U12324 ( .A1(n10742), .A2(n9805), .ZN(n9892) );
  NAND2_X1 U12325 ( .A1(n9901), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9890) );
  XNOR2_X1 U12326 ( .A(n9890), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U12327 ( .A1(n9651), .A2(SI_18_), .B1(n11530), .B2(n13316), .ZN(
        n9891) );
  NAND2_X1 U12328 ( .A1(n9892), .A2(n9891), .ZN(n13589) );
  NAND2_X1 U12329 ( .A1(n9646), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U12330 ( .A1(n9893), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U12331 ( .A1(n9906), .A2(n9894), .ZN(n13478) );
  NAND2_X1 U12332 ( .A1(n9816), .A2(n13478), .ZN(n9897) );
  NAND2_X1 U12333 ( .A1(n9847), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9896) );
  INV_X1 U12334 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13292) );
  OR2_X1 U12335 ( .A1(n6994), .A2(n13292), .ZN(n9895) );
  OR2_X1 U12336 ( .A1(n13589), .A2(n13491), .ZN(n13459) );
  NAND2_X1 U12337 ( .A1(n13589), .A2(n13491), .ZN(n10161) );
  XNOR2_X1 U12338 ( .A(n9900), .B(n9899), .ZN(n10830) );
  NAND2_X1 U12339 ( .A1(n10830), .A2(n9805), .ZN(n9904) );
  AOI22_X1 U12340 ( .A1(n9651), .A2(n10831), .B1(n11530), .B2(n13314), .ZN(
        n9903) );
  INV_X1 U12341 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n9905) );
  OR2_X1 U12342 ( .A1(n6994), .A2(n9905), .ZN(n9911) );
  NAND2_X1 U12343 ( .A1(n9646), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9910) );
  AND2_X1 U12344 ( .A1(n9906), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9907) );
  OR2_X1 U12345 ( .A1(n9907), .A2(n9917), .ZN(n13463) );
  NAND2_X1 U12346 ( .A1(n9816), .A2(n13463), .ZN(n9909) );
  NAND2_X1 U12347 ( .A1(n9847), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9908) );
  NAND4_X1 U12348 ( .A1(n9911), .A2(n9910), .A3(n9909), .A4(n9908), .ZN(n13472) );
  NAND2_X1 U12349 ( .A1(n13644), .A2(n13472), .ZN(n10167) );
  OR2_X1 U12350 ( .A1(n13644), .A2(n13472), .ZN(n10166) );
  NAND2_X1 U12351 ( .A1(n9912), .A2(n10166), .ZN(n13444) );
  XNOR2_X1 U12352 ( .A(n9913), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U12353 ( .A1(n11084), .A2(n9805), .ZN(n9915) );
  NAND2_X1 U12354 ( .A1(n9651), .A2(SI_20_), .ZN(n9914) );
  NAND2_X1 U12355 ( .A1(n9951), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12356 ( .A1(n10000), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U12357 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  OR2_X1 U12358 ( .A1(n9930), .A2(n9918), .ZN(n13445) );
  NAND2_X1 U12359 ( .A1(n13445), .A2(n9816), .ZN(n9920) );
  NAND2_X1 U12360 ( .A1(n9847), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9919) );
  NAND4_X1 U12361 ( .A1(n9922), .A2(n9921), .A3(n9920), .A4(n9919), .ZN(n13454) );
  XNOR2_X1 U12362 ( .A(n13638), .B(n13454), .ZN(n13443) );
  INV_X1 U12363 ( .A(n13638), .ZN(n13447) );
  NAND2_X1 U12364 ( .A1(n13447), .A2(n13454), .ZN(n9923) );
  INV_X1 U12365 ( .A(n9924), .ZN(n9925) );
  XNOR2_X1 U12366 ( .A(n9926), .B(n9925), .ZN(n11265) );
  NAND2_X1 U12367 ( .A1(n11265), .A2(n9805), .ZN(n9928) );
  NAND2_X1 U12368 ( .A1(n9651), .A2(SI_21_), .ZN(n9927) );
  OR2_X1 U12369 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  NAND2_X1 U12370 ( .A1(n9939), .A2(n9931), .ZN(n13431) );
  AOI22_X1 U12371 ( .A1(n13431), .A2(n9816), .B1(n9847), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U12372 ( .A1(n9951), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n9646), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U12373 ( .A1(n13430), .A2(n13439), .ZN(n10175) );
  NAND2_X1 U12374 ( .A1(n13428), .A2(n10175), .ZN(n9934) );
  NAND2_X1 U12375 ( .A1(n9934), .A2(n10176), .ZN(n13416) );
  XNOR2_X1 U12376 ( .A(n9936), .B(n9935), .ZN(n11188) );
  NAND2_X1 U12377 ( .A1(n11188), .A2(n9805), .ZN(n9938) );
  NAND2_X1 U12378 ( .A1(n9651), .A2(SI_22_), .ZN(n9937) );
  INV_X1 U12379 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U12380 ( .A1(n9939), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U12381 ( .A1(n9949), .A2(n9940), .ZN(n13417) );
  NAND2_X1 U12382 ( .A1(n13417), .A2(n9816), .ZN(n9942) );
  AOI22_X1 U12383 ( .A1(n9951), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n10000), 
        .B2(P3_REG2_REG_22__SCAN_IN), .ZN(n9941) );
  OAI211_X1 U12384 ( .C1(n9943), .C2(n13629), .A(n9942), .B(n9941), .ZN(n13423) );
  NAND2_X1 U12385 ( .A1(n13107), .A2(n13403), .ZN(n10071) );
  NAND2_X1 U12386 ( .A1(n13416), .A2(n10071), .ZN(n9944) );
  OR2_X1 U12387 ( .A1(n13107), .A2(n13403), .ZN(n10070) );
  XNOR2_X1 U12388 ( .A(n9946), .B(n9945), .ZN(n11509) );
  NAND2_X1 U12389 ( .A1(n11509), .A2(n9805), .ZN(n9948) );
  NAND2_X1 U12390 ( .A1(n9651), .A2(SI_23_), .ZN(n9947) );
  NAND2_X1 U12391 ( .A1(n9949), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12392 ( .A1(n9959), .A2(n9950), .ZN(n13406) );
  NAND2_X1 U12393 ( .A1(n13406), .A2(n9816), .ZN(n9954) );
  AOI22_X1 U12394 ( .A1(n9951), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n10000), 
        .B2(P3_REG2_REG_23__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U12395 ( .A1(n9847), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9952) );
  XNOR2_X1 U12396 ( .A(n13015), .B(n13412), .ZN(n13404) );
  INV_X1 U12397 ( .A(n13404), .ZN(n10181) );
  NAND2_X1 U12398 ( .A1(n13627), .A2(n13390), .ZN(n10185) );
  XNOR2_X1 U12399 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9956), .ZN(n12230) );
  NAND2_X1 U12400 ( .A1(n12230), .A2(n9805), .ZN(n9958) );
  NAND2_X1 U12401 ( .A1(n9651), .A2(SI_24_), .ZN(n9957) );
  INV_X1 U12402 ( .A(n9972), .ZN(n9961) );
  NAND2_X1 U12403 ( .A1(n9959), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U12404 ( .A1(n9961), .A2(n9960), .ZN(n13395) );
  NAND2_X1 U12405 ( .A1(n13395), .A2(n9816), .ZN(n9966) );
  INV_X1 U12406 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U12407 ( .A1(n9646), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12408 ( .A1(n9847), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9962) );
  OAI211_X1 U12409 ( .C1(n6994), .C2(n13562), .A(n9963), .B(n9962), .ZN(n9964)
         );
  INV_X1 U12410 ( .A(n9964), .ZN(n9965) );
  NAND2_X1 U12411 ( .A1(n12602), .A2(n13402), .ZN(n10189) );
  NAND2_X1 U12412 ( .A1(n10187), .A2(n10189), .ZN(n13387) );
  XNOR2_X1 U12413 ( .A(n9968), .B(n9967), .ZN(n12276) );
  NAND2_X1 U12414 ( .A1(n12276), .A2(n9805), .ZN(n9970) );
  NAND2_X1 U12415 ( .A1(n9651), .A2(SI_25_), .ZN(n9969) );
  OR2_X1 U12416 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  NAND2_X1 U12417 ( .A1(n9983), .A2(n9973), .ZN(n13379) );
  NAND2_X1 U12418 ( .A1(n13379), .A2(n9816), .ZN(n9978) );
  INV_X1 U12419 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U12420 ( .A1(n10000), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U12421 ( .A1(n9847), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9974) );
  OAI211_X1 U12422 ( .C1(n6994), .C2(n13558), .A(n9975), .B(n9974), .ZN(n9976)
         );
  INV_X1 U12423 ( .A(n9976), .ZN(n9977) );
  NAND2_X1 U12424 ( .A1(n13378), .A2(n12992), .ZN(n10195) );
  AOI22_X1 U12425 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n14253), .B2(n14950), .ZN(n9979) );
  XNOR2_X1 U12426 ( .A(n9980), .B(n9979), .ZN(n13669) );
  NAND2_X1 U12427 ( .A1(n13669), .A2(n9805), .ZN(n9982) );
  NAND2_X1 U12428 ( .A1(n9651), .A2(SI_26_), .ZN(n9981) );
  NAND2_X1 U12429 ( .A1(n9983), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U12430 ( .A1(n9997), .A2(n9984), .ZN(n13363) );
  NAND2_X1 U12431 ( .A1(n13363), .A2(n9816), .ZN(n9990) );
  INV_X1 U12432 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U12433 ( .A1(n9847), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12434 ( .A1(n10000), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9985) );
  OAI211_X1 U12435 ( .C1(n6994), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9988)
         );
  INV_X1 U12436 ( .A(n9988), .ZN(n9989) );
  INV_X1 U12437 ( .A(n13372), .ZN(n9991) );
  NAND2_X1 U12438 ( .A1(n13552), .A2(n9991), .ZN(n10067) );
  AOI22_X1 U12439 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n14250), .B2(n7617), .ZN(n9992) );
  INV_X1 U12440 ( .A(n9992), .ZN(n9993) );
  XNOR2_X1 U12441 ( .A(n9994), .B(n9993), .ZN(n12968) );
  NAND2_X1 U12442 ( .A1(n12968), .A2(n9805), .ZN(n9996) );
  NAND2_X1 U12443 ( .A1(n9651), .A2(SI_27_), .ZN(n9995) );
  INV_X1 U12444 ( .A(n10012), .ZN(n9999) );
  NAND2_X1 U12445 ( .A1(n9997), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U12446 ( .A1(n9999), .A2(n9998), .ZN(n13353) );
  NAND2_X1 U12447 ( .A1(n13353), .A2(n9816), .ZN(n10005) );
  INV_X1 U12448 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13550) );
  NAND2_X1 U12449 ( .A1(n10000), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U12450 ( .A1(n9847), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10001) );
  OAI211_X1 U12451 ( .C1(n6994), .C2(n13550), .A(n10002), .B(n10001), .ZN(
        n10003) );
  INV_X1 U12452 ( .A(n10003), .ZN(n10004) );
  NAND2_X1 U12453 ( .A1(n13347), .A2(n13346), .ZN(n10006) );
  NAND2_X1 U12454 ( .A1(n13352), .A2(n13139), .ZN(n10063) );
  AOI22_X1 U12455 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14245), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n12605), .ZN(n10007) );
  INV_X1 U12456 ( .A(n10007), .ZN(n10008) );
  XNOR2_X1 U12457 ( .A(n10009), .B(n10008), .ZN(n12558) );
  NAND2_X1 U12458 ( .A1(n12558), .A2(n9805), .ZN(n10011) );
  NAND2_X1 U12459 ( .A1(n9651), .A2(SI_28_), .ZN(n10010) );
  NOR2_X1 U12460 ( .A1(n10012), .A2(n13034), .ZN(n10013) );
  INV_X1 U12461 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13546) );
  NAND2_X1 U12462 ( .A1(n9646), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U12463 ( .A1(n9847), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10014) );
  OAI211_X1 U12464 ( .C1(n6994), .C2(n13546), .A(n10015), .B(n10014), .ZN(
        n10016) );
  AOI21_X1 U12465 ( .B1(n13337), .B2(n9816), .A(n10016), .ZN(n12996) );
  NAND2_X1 U12466 ( .A1(n12515), .A2(n12996), .ZN(n10064) );
  NAND2_X1 U12467 ( .A1(n9651), .A2(SI_29_), .ZN(n10019) );
  INV_X1 U12468 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12469 ( .A1(n10000), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U12470 ( .A1(n9847), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10021) );
  OAI211_X1 U12471 ( .C1(n6994), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10025) );
  INV_X1 U12472 ( .A(n10025), .ZN(n10026) );
  OR2_X2 U12473 ( .A1(n13606), .A2(n13033), .ZN(n10204) );
  NAND2_X1 U12474 ( .A1(n15036), .A2(n15029), .ZN(n10210) );
  NAND2_X1 U12475 ( .A1(n13606), .A2(n13033), .ZN(n10203) );
  INV_X1 U12476 ( .A(n15029), .ZN(n10028) );
  OAI21_X1 U12477 ( .B1(n10028), .B2(n12545), .A(n15040), .ZN(n10029) );
  XNOR2_X1 U12478 ( .A(n10030), .B(n13325), .ZN(n10060) );
  INV_X1 U12479 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12480 ( .A1(n10040), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U12481 ( .A1(n10038), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U12482 ( .A1(n11487), .A2(n12621), .ZN(n11498) );
  NAND2_X1 U12483 ( .A1(n10070), .A2(n10071), .ZN(n13415) );
  NAND2_X1 U12484 ( .A1(n13376), .A2(n7651), .ZN(n10069) );
  NAND2_X1 U12485 ( .A1(n10162), .A2(n10157), .ZN(n12522) );
  NAND2_X1 U12486 ( .A1(n10142), .A2(n10143), .ZN(n12516) );
  NAND2_X1 U12487 ( .A1(n10138), .A2(n10137), .ZN(n13528) );
  NAND2_X1 U12488 ( .A1(n15614), .A2(n12637), .ZN(n10073) );
  INV_X1 U12489 ( .A(n10073), .ZN(n10042) );
  OR2_X1 U12490 ( .A1(n11369), .A2(n10042), .ZN(n15493) );
  INV_X1 U12491 ( .A(n15493), .ZN(n12555) );
  NAND2_X1 U12492 ( .A1(n10078), .A2(n10080), .ZN(n11492) );
  INV_X1 U12493 ( .A(n11492), .ZN(n15611) );
  NAND4_X1 U12494 ( .A1(n12555), .A2(n11502), .A3(n10043), .A4(n15611), .ZN(
        n10047) );
  NAND2_X1 U12495 ( .A1(n12243), .A2(n12223), .ZN(n10044) );
  INV_X1 U12496 ( .A(n12223), .ZN(n12183) );
  NAND2_X1 U12497 ( .A1(n12305), .A2(n12183), .ZN(n12301) );
  INV_X1 U12498 ( .A(n12218), .ZN(n10119) );
  NAND4_X1 U12499 ( .A1(n10045), .A2(n15561), .A3(n10119), .A4(n12165), .ZN(
        n10046) );
  NOR3_X1 U12500 ( .A1(n10047), .A2(n10046), .A3(n15593), .ZN(n10049) );
  AND2_X1 U12501 ( .A1(n10128), .A2(n12448), .ZN(n10125) );
  NAND2_X1 U12502 ( .A1(n12456), .A2(n10124), .ZN(n12303) );
  NOR2_X1 U12503 ( .A1(n12303), .A2(n12057), .ZN(n10048) );
  NAND4_X1 U12504 ( .A1(n10049), .A2(n10125), .A3(n12450), .A4(n10048), .ZN(
        n10050) );
  NOR3_X1 U12505 ( .A1(n12516), .A2(n13528), .A3(n10050), .ZN(n10051) );
  NAND3_X1 U12506 ( .A1(n13508), .A2(n13518), .A3(n10051), .ZN(n10052) );
  NOR3_X1 U12507 ( .A1(n13477), .A2(n12522), .A3(n10052), .ZN(n10053) );
  NAND4_X1 U12508 ( .A1(n12530), .A2(n13460), .A3(n13443), .A4(n10053), .ZN(
        n10054) );
  NOR4_X1 U12509 ( .A1(n13415), .A2(n13404), .A3(n10069), .A4(n10054), .ZN(
        n10056) );
  NOR2_X1 U12510 ( .A1(n12548), .A2(n13328), .ZN(n10055) );
  XNOR2_X1 U12511 ( .A(n10058), .B(n13325), .ZN(n10059) );
  INV_X1 U12512 ( .A(n12548), .ZN(n10207) );
  NAND2_X1 U12513 ( .A1(n10213), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10062) );
  AOI21_X1 U12514 ( .B1(n10064), .B2(n10063), .A(n12624), .ZN(n10066) );
  MUX2_X1 U12515 ( .A(n12624), .B(n10066), .S(n10065), .Z(n10206) );
  INV_X1 U12516 ( .A(n13328), .ZN(n13330) );
  NAND2_X1 U12517 ( .A1(n13359), .A2(n12624), .ZN(n10201) );
  MUX2_X1 U12518 ( .A(n10068), .B(n10067), .S(n12624), .Z(n10199) );
  INV_X1 U12519 ( .A(n10069), .ZN(n10194) );
  MUX2_X1 U12520 ( .A(n10071), .B(n10070), .S(n11532), .Z(n10182) );
  INV_X1 U12521 ( .A(n13415), .ZN(n10179) );
  NAND2_X1 U12522 ( .A1(n10073), .A2(n11487), .ZN(n10072) );
  NAND2_X1 U12523 ( .A1(n10072), .A2(n12624), .ZN(n10075) );
  NAND3_X1 U12524 ( .A1(n10073), .A2(n10080), .A3(n11485), .ZN(n10074) );
  NAND2_X1 U12525 ( .A1(n10075), .A2(n10074), .ZN(n10077) );
  NAND2_X1 U12526 ( .A1(n11369), .A2(n11362), .ZN(n10076) );
  NAND2_X1 U12527 ( .A1(n10077), .A2(n10076), .ZN(n10079) );
  MUX2_X1 U12528 ( .A(n12624), .B(n10079), .S(n10078), .Z(n10085) );
  NOR2_X1 U12529 ( .A1(n10080), .A2(n11532), .ZN(n10081) );
  NOR2_X1 U12530 ( .A1(n15593), .A2(n10081), .ZN(n10084) );
  NAND2_X1 U12531 ( .A1(n15612), .A2(n15588), .ZN(n10082) );
  AOI21_X1 U12532 ( .B1(n10091), .B2(n10082), .A(n12624), .ZN(n10083) );
  AOI21_X1 U12533 ( .B1(n10085), .B2(n10084), .A(n10083), .ZN(n10090) );
  INV_X1 U12534 ( .A(n10087), .ZN(n10089) );
  AND2_X1 U12535 ( .A1(n10087), .A2(n10086), .ZN(n10088) );
  OAI22_X1 U12536 ( .A1(n10090), .A2(n10089), .B1(n11532), .B2(n10088), .ZN(
        n10094) );
  NOR2_X1 U12537 ( .A1(n10091), .A2(n11532), .ZN(n10092) );
  NOR2_X1 U12538 ( .A1(n15576), .A2(n10092), .ZN(n10093) );
  NAND2_X1 U12539 ( .A1(n10094), .A2(n10093), .ZN(n10099) );
  NAND3_X1 U12540 ( .A1(n10099), .A2(n15561), .A3(n10095), .ZN(n10097) );
  NAND3_X1 U12541 ( .A1(n10097), .A2(n10096), .A3(n10101), .ZN(n10106) );
  NAND3_X1 U12542 ( .A1(n10099), .A2(n15561), .A3(n10098), .ZN(n10104) );
  AND2_X1 U12543 ( .A1(n10107), .A2(n10100), .ZN(n10103) );
  INV_X1 U12544 ( .A(n10101), .ZN(n10102) );
  AOI21_X1 U12545 ( .B1(n10104), .B2(n10103), .A(n10102), .ZN(n10105) );
  MUX2_X1 U12546 ( .A(n10106), .B(n10105), .S(n11532), .Z(n10110) );
  INV_X1 U12547 ( .A(n10107), .ZN(n10108) );
  AOI21_X1 U12548 ( .B1(n10108), .B2(n12624), .A(n12057), .ZN(n10109) );
  NAND2_X1 U12549 ( .A1(n10110), .A2(n10109), .ZN(n10115) );
  NAND2_X1 U12550 ( .A1(n10111), .A2(n11532), .ZN(n10113) );
  NAND2_X1 U12551 ( .A1(n12169), .A2(n12624), .ZN(n10112) );
  MUX2_X1 U12552 ( .A(n10113), .B(n10112), .S(n12083), .Z(n10114) );
  NAND3_X1 U12553 ( .A1(n10115), .A2(n12165), .A3(n10114), .ZN(n10120) );
  MUX2_X1 U12554 ( .A(n10117), .B(n10116), .S(n11532), .Z(n10118) );
  NAND3_X1 U12555 ( .A1(n10120), .A2(n10119), .A3(n10118), .ZN(n10123) );
  MUX2_X1 U12556 ( .A(n12305), .B(n12183), .S(n11532), .Z(n10121) );
  AOI21_X1 U12557 ( .B1(n10121), .B2(n12301), .A(n12303), .ZN(n10122) );
  NAND2_X1 U12558 ( .A1(n10123), .A2(n10122), .ZN(n10127) );
  MUX2_X1 U12559 ( .A(n12456), .B(n10124), .S(n11532), .Z(n10126) );
  INV_X1 U12560 ( .A(n10125), .ZN(n12459) );
  AOI21_X1 U12561 ( .B1(n10127), .B2(n10126), .A(n12459), .ZN(n10136) );
  NAND2_X1 U12562 ( .A1(n10132), .A2(n10128), .ZN(n10130) );
  NAND2_X1 U12563 ( .A1(n10131), .A2(n12448), .ZN(n10129) );
  MUX2_X1 U12564 ( .A(n10130), .B(n10129), .S(n11532), .Z(n10135) );
  INV_X1 U12565 ( .A(n13528), .ZN(n10134) );
  MUX2_X1 U12566 ( .A(n10132), .B(n10131), .S(n12624), .Z(n10133) );
  OAI211_X1 U12567 ( .C1(n10136), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10140) );
  INV_X1 U12568 ( .A(n12516), .ZN(n12482) );
  MUX2_X1 U12569 ( .A(n10138), .B(n10137), .S(n11532), .Z(n10139) );
  NAND3_X1 U12570 ( .A1(n10140), .A2(n12482), .A3(n10139), .ZN(n10141) );
  OAI21_X1 U12571 ( .B1(n10142), .B2(n12624), .A(n10141), .ZN(n10149) );
  INV_X1 U12572 ( .A(n10143), .ZN(n10144) );
  NAND2_X1 U12573 ( .A1(n13518), .A2(n10144), .ZN(n10147) );
  NAND3_X1 U12574 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10148) );
  AOI22_X1 U12575 ( .A1(n10149), .A2(n13518), .B1(n12624), .B2(n10148), .ZN(
        n10153) );
  INV_X1 U12576 ( .A(n13492), .ZN(n10152) );
  AND2_X1 U12577 ( .A1(n13492), .A2(n10150), .ZN(n10151) );
  OAI22_X1 U12578 ( .A1(n10153), .A2(n10152), .B1(n10151), .B2(n12624), .ZN(
        n10156) );
  OR3_X1 U12579 ( .A1(n13067), .A2(n13517), .A3(n12624), .ZN(n10155) );
  NAND2_X1 U12580 ( .A1(n10159), .A2(n12523), .ZN(n10154) );
  AOI21_X1 U12581 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(n10170) );
  INV_X1 U12582 ( .A(n10157), .ZN(n10158) );
  NAND2_X1 U12583 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  NAND3_X1 U12584 ( .A1(n10166), .A2(n10160), .A3(n10161), .ZN(n10165) );
  INV_X1 U12585 ( .A(n10161), .ZN(n10163) );
  OAI211_X1 U12586 ( .C1(n10163), .C2(n10162), .A(n10167), .B(n13459), .ZN(
        n10164) );
  MUX2_X1 U12587 ( .A(n10165), .B(n10164), .S(n11532), .Z(n10169) );
  MUX2_X1 U12588 ( .A(n10167), .B(n10166), .S(n11532), .Z(n10168) );
  OAI211_X1 U12589 ( .C1(n10170), .C2(n10169), .A(n13443), .B(n10168), .ZN(
        n10174) );
  NAND2_X1 U12590 ( .A1(n13638), .A2(n12624), .ZN(n10172) );
  NAND2_X1 U12591 ( .A1(n13447), .A2(n11532), .ZN(n10171) );
  MUX2_X1 U12592 ( .A(n10172), .B(n10171), .S(n13454), .Z(n10173) );
  NAND3_X1 U12593 ( .A1(n10174), .A2(n12530), .A3(n10173), .ZN(n10178) );
  MUX2_X1 U12594 ( .A(n10176), .B(n10175), .S(n11532), .Z(n10177) );
  NAND3_X1 U12595 ( .A1(n10179), .A2(n10178), .A3(n10177), .ZN(n10180) );
  NAND3_X1 U12596 ( .A1(n10182), .A2(n10181), .A3(n10180), .ZN(n10184) );
  NAND3_X1 U12597 ( .A1(n13015), .A2(n13412), .A3(n11532), .ZN(n10183) );
  NAND2_X1 U12598 ( .A1(n10184), .A2(n10183), .ZN(n10193) );
  INV_X1 U12599 ( .A(n10185), .ZN(n10186) );
  NAND2_X1 U12600 ( .A1(n10189), .A2(n10186), .ZN(n10188) );
  NAND2_X1 U12601 ( .A1(n10188), .A2(n10187), .ZN(n10191) );
  INV_X1 U12602 ( .A(n10189), .ZN(n10190) );
  MUX2_X1 U12603 ( .A(n10191), .B(n10190), .S(n11532), .Z(n10192) );
  MUX2_X1 U12604 ( .A(n10196), .B(n10195), .S(n11532), .Z(n10197) );
  NAND3_X1 U12605 ( .A1(n13346), .A2(n10199), .A3(n10198), .ZN(n10200) );
  OAI21_X1 U12606 ( .B1(n13352), .B2(n10201), .A(n10200), .ZN(n10202) );
  MUX2_X1 U12607 ( .A(n10204), .B(n10203), .S(n11532), .Z(n10205) );
  NAND2_X1 U12608 ( .A1(n11483), .A2(n13314), .ZN(n12622) );
  INV_X1 U12609 ( .A(n12622), .ZN(n11488) );
  INV_X1 U12610 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n10214) );
  OR2_X1 U12611 ( .A1(n11531), .A2(P3_U3151), .ZN(n11528) );
  INV_X1 U12612 ( .A(n11528), .ZN(n10216) );
  NOR2_X1 U12613 ( .A1(n10226), .A2(n10225), .ZN(n10219) );
  INV_X1 U12614 ( .A(n10220), .ZN(n10221) );
  NOR2_X1 U12615 ( .A1(n10223), .A2(n10225), .ZN(n10224) );
  NOR2_X1 U12616 ( .A1(n12280), .A2(n12233), .ZN(n10228) );
  OR2_X1 U12617 ( .A1(n11529), .A2(n12622), .ZN(n11356) );
  INV_X1 U12618 ( .A(n12561), .ZN(n12543) );
  NAND2_X1 U12619 ( .A1(n12543), .A2(n6997), .ZN(n11559) );
  NAND2_X1 U12620 ( .A1(n11559), .A2(n10229), .ZN(n11354) );
  INV_X1 U12621 ( .A(n11354), .ZN(n10230) );
  NOR2_X1 U12622 ( .A1(n11356), .A2(n15594), .ZN(n11353) );
  OAI21_X1 U12623 ( .B1(n11528), .B2(n11485), .A(P3_B_REG_SCAN_IN), .ZN(n10231) );
  AOI21_X1 U12624 ( .B1(n11353), .B2(n12543), .A(n10231), .ZN(n10232) );
  INV_X1 U12625 ( .A(n10232), .ZN(n10233) );
  NAND2_X1 U12626 ( .A1(n10234), .A2(n10233), .ZN(P3_U3296) );
  NOR2_X1 U12627 ( .A1(n14570), .A2(n10458), .ZN(n10235) );
  AOI21_X1 U12628 ( .B1(n14888), .B2(n10437), .A(n10235), .ZN(n10381) );
  OAI22_X1 U12629 ( .A1(n14742), .A2(n10457), .B1(n14570), .B2(n10445), .ZN(
        n10236) );
  XNOR2_X1 U12630 ( .A(n10236), .B(n10701), .ZN(n10376) );
  INV_X1 U12631 ( .A(n10376), .ZN(n10380) );
  AOI22_X1 U12632 ( .A1(n14905), .A2(n10437), .B1(n6967), .B2(n14564), .ZN(
        n10367) );
  AOI22_X1 U12633 ( .A1(n14905), .A2(n10444), .B1(n10451), .B2(n14564), .ZN(
        n10237) );
  XNOR2_X1 U12634 ( .A(n10237), .B(n10701), .ZN(n10366) );
  NAND2_X1 U12635 ( .A1(n10241), .A2(n10288), .ZN(n10239) );
  OR2_X1 U12636 ( .A1(n11047), .A2(n10457), .ZN(n10238) );
  NAND2_X1 U12637 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  XNOR2_X1 U12638 ( .A(n10240), .B(n10701), .ZN(n10249) );
  AOI22_X1 U12639 ( .A1(n14806), .A2(n10437), .B1(n14955), .B2(n7586), .ZN(
        n10242) );
  AND2_X1 U12640 ( .A1(n10243), .A2(n10242), .ZN(n10714) );
  NAND2_X1 U12641 ( .A1(n14411), .A2(n10288), .ZN(n10247) );
  NOR2_X1 U12642 ( .A1(n10481), .A2(n10244), .ZN(n10245) );
  AOI21_X1 U12643 ( .B1(n14806), .B2(n10444), .A(n10245), .ZN(n10246) );
  NAND2_X1 U12644 ( .A1(n10247), .A2(n10246), .ZN(n10713) );
  NAND2_X1 U12645 ( .A1(n10714), .A2(n10713), .ZN(n10712) );
  OR2_X1 U12646 ( .A1(n10713), .A2(n10448), .ZN(n10248) );
  NAND2_X1 U12647 ( .A1(n10712), .A2(n10248), .ZN(n10791) );
  INV_X1 U12648 ( .A(n10249), .ZN(n10251) );
  NAND2_X1 U12649 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NAND2_X1 U12650 ( .A1(n10253), .A2(n10252), .ZN(n10883) );
  NAND2_X1 U12651 ( .A1(n14408), .A2(n10288), .ZN(n10255) );
  OR2_X1 U12652 ( .A1(n15232), .A2(n10457), .ZN(n10254) );
  NAND2_X1 U12653 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  XNOR2_X1 U12654 ( .A(n10256), .B(n10701), .ZN(n10257) );
  INV_X1 U12655 ( .A(n15232), .ZN(n15206) );
  AOI22_X1 U12656 ( .A1(n14408), .A2(n10417), .B1(n15206), .B2(n10288), .ZN(
        n10258) );
  XNOR2_X1 U12657 ( .A(n10257), .B(n10258), .ZN(n10882) );
  INV_X1 U12658 ( .A(n10257), .ZN(n10259) );
  NAND2_X1 U12659 ( .A1(n10259), .A2(n10258), .ZN(n10260) );
  NAND2_X1 U12660 ( .A1(n14407), .A2(n10288), .ZN(n10262) );
  NAND2_X1 U12661 ( .A1(n6976), .A2(n10444), .ZN(n10261) );
  NAND2_X1 U12662 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  XNOR2_X1 U12663 ( .A(n10263), .B(n10448), .ZN(n10266) );
  AOI22_X1 U12664 ( .A1(n14407), .A2(n10417), .B1(n6976), .B2(n10288), .ZN(
        n10265) );
  XNOR2_X1 U12665 ( .A(n10266), .B(n10265), .ZN(n10929) );
  OR2_X1 U12666 ( .A1(n10266), .A2(n10265), .ZN(n11026) );
  NAND2_X1 U12667 ( .A1(n14406), .A2(n10288), .ZN(n10268) );
  NAND2_X1 U12668 ( .A1(n11203), .A2(n10444), .ZN(n10267) );
  NAND2_X1 U12669 ( .A1(n10268), .A2(n10267), .ZN(n10269) );
  XNOR2_X1 U12670 ( .A(n10269), .B(n10701), .ZN(n11029) );
  NAND2_X1 U12671 ( .A1(n14406), .A2(n10417), .ZN(n10271) );
  NAND2_X1 U12672 ( .A1(n11203), .A2(n10451), .ZN(n10270) );
  NAND2_X1 U12673 ( .A1(n10271), .A2(n10270), .ZN(n10274) );
  NAND2_X1 U12674 ( .A1(n11029), .A2(n10274), .ZN(n10272) );
  AND2_X1 U12675 ( .A1(n11026), .A2(n10272), .ZN(n10273) );
  NAND2_X1 U12676 ( .A1(n11027), .A2(n10273), .ZN(n10277) );
  INV_X1 U12677 ( .A(n11029), .ZN(n10275) );
  INV_X1 U12678 ( .A(n10274), .ZN(n11028) );
  NAND2_X1 U12679 ( .A1(n10275), .A2(n11028), .ZN(n10276) );
  INV_X1 U12680 ( .A(n10368), .ZN(n10296) );
  OR2_X1 U12681 ( .A1(n11276), .A2(n10296), .ZN(n10279) );
  NAND2_X1 U12682 ( .A1(n14405), .A2(n6967), .ZN(n10278) );
  AND2_X1 U12683 ( .A1(n10279), .A2(n10278), .ZN(n11059) );
  NAND2_X1 U12684 ( .A1(n11061), .A2(n11059), .ZN(n10282) );
  NAND2_X1 U12685 ( .A1(n14405), .A2(n10451), .ZN(n10280) );
  OAI21_X1 U12686 ( .B1(n11276), .B2(n10457), .A(n10280), .ZN(n10281) );
  XNOR2_X1 U12687 ( .A(n10281), .B(n10701), .ZN(n11058) );
  NAND2_X1 U12688 ( .A1(n10282), .A2(n11058), .ZN(n10284) );
  NAND2_X1 U12689 ( .A1(n11314), .A2(n10444), .ZN(n10286) );
  OR2_X1 U12690 ( .A1(n11279), .A2(n10296), .ZN(n10285) );
  NAND2_X1 U12691 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  XNOR2_X1 U12692 ( .A(n10287), .B(n10448), .ZN(n10291) );
  NAND2_X1 U12693 ( .A1(n11314), .A2(n10288), .ZN(n10290) );
  OR2_X1 U12694 ( .A1(n11279), .A2(n10458), .ZN(n10289) );
  NAND2_X1 U12695 ( .A1(n10290), .A2(n10289), .ZN(n10292) );
  XNOR2_X1 U12696 ( .A(n10291), .B(n10292), .ZN(n11111) );
  NAND2_X1 U12697 ( .A1(n11112), .A2(n11111), .ZN(n10295) );
  INV_X1 U12698 ( .A(n10291), .ZN(n10293) );
  NAND2_X1 U12699 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  NAND2_X1 U12700 ( .A1(n10295), .A2(n10294), .ZN(n11191) );
  NAND2_X1 U12701 ( .A1(n15263), .A2(n10444), .ZN(n10298) );
  OR2_X1 U12702 ( .A1(n11518), .A2(n10296), .ZN(n10297) );
  NAND2_X1 U12703 ( .A1(n10298), .A2(n10297), .ZN(n10299) );
  XNOR2_X1 U12704 ( .A(n10299), .B(n10701), .ZN(n10300) );
  AOI22_X1 U12705 ( .A1(n15263), .A2(n10437), .B1(n6967), .B2(n14403), .ZN(
        n10301) );
  XNOR2_X1 U12706 ( .A(n10300), .B(n10301), .ZN(n11190) );
  NAND2_X1 U12707 ( .A1(n11191), .A2(n11190), .ZN(n10304) );
  INV_X1 U12708 ( .A(n10300), .ZN(n10302) );
  OR2_X1 U12709 ( .A1(n10302), .A2(n10301), .ZN(n10303) );
  NAND2_X1 U12710 ( .A1(n11705), .A2(n10444), .ZN(n10306) );
  OR2_X1 U12711 ( .A1(n11709), .A2(n10445), .ZN(n10305) );
  NAND2_X1 U12712 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  XNOR2_X1 U12713 ( .A(n10307), .B(n10448), .ZN(n10310) );
  NOR2_X1 U12714 ( .A1(n11709), .A2(n10458), .ZN(n10308) );
  AOI21_X1 U12715 ( .B1(n11705), .B2(n10451), .A(n10308), .ZN(n10309) );
  XNOR2_X1 U12716 ( .A(n10310), .B(n10309), .ZN(n11472) );
  NAND2_X1 U12717 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  NOR2_X1 U12718 ( .A1(n12020), .A2(n10458), .ZN(n10312) );
  AOI21_X1 U12719 ( .B1(n12030), .B2(n10451), .A(n10312), .ZN(n10316) );
  NAND2_X1 U12720 ( .A1(n10317), .A2(n10316), .ZN(n11946) );
  NAND2_X1 U12721 ( .A1(n12030), .A2(n10444), .ZN(n10314) );
  OR2_X1 U12722 ( .A1(n12020), .A2(n10445), .ZN(n10313) );
  NAND2_X1 U12723 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  XNOR2_X1 U12724 ( .A(n10315), .B(n10701), .ZN(n11949) );
  NAND2_X1 U12725 ( .A1(n11946), .A2(n11949), .ZN(n10318) );
  NAND2_X1 U12726 ( .A1(n10318), .A2(n11947), .ZN(n11972) );
  NAND2_X1 U12727 ( .A1(n15284), .A2(n10444), .ZN(n10320) );
  OR2_X1 U12728 ( .A1(n15096), .A2(n10445), .ZN(n10319) );
  NAND2_X1 U12729 ( .A1(n10320), .A2(n10319), .ZN(n10321) );
  XNOR2_X1 U12730 ( .A(n10321), .B(n10448), .ZN(n10323) );
  NOR2_X1 U12731 ( .A1(n15096), .A2(n10458), .ZN(n10322) );
  AOI21_X1 U12732 ( .B1(n15284), .B2(n10451), .A(n10322), .ZN(n10324) );
  NAND2_X1 U12733 ( .A1(n10323), .A2(n10324), .ZN(n11971) );
  NAND2_X1 U12734 ( .A1(n11972), .A2(n11971), .ZN(n10327) );
  INV_X1 U12735 ( .A(n10323), .ZN(n10326) );
  INV_X1 U12736 ( .A(n10324), .ZN(n10325) );
  NAND2_X1 U12737 ( .A1(n10326), .A2(n10325), .ZN(n11970) );
  NAND2_X1 U12738 ( .A1(n10327), .A2(n11970), .ZN(n15100) );
  INV_X1 U12739 ( .A(n15100), .ZN(n10333) );
  NAND2_X1 U12740 ( .A1(n15122), .A2(n10444), .ZN(n10329) );
  NAND2_X1 U12741 ( .A1(n14985), .A2(n10451), .ZN(n10328) );
  NAND2_X1 U12742 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  XNOR2_X1 U12743 ( .A(n10330), .B(n10448), .ZN(n10335) );
  AND2_X1 U12744 ( .A1(n14985), .A2(n6967), .ZN(n10331) );
  AOI21_X1 U12745 ( .B1(n15122), .B2(n10451), .A(n10331), .ZN(n10334) );
  XNOR2_X1 U12746 ( .A(n10335), .B(n10334), .ZN(n15099) );
  INV_X1 U12747 ( .A(n15099), .ZN(n10332) );
  NAND2_X1 U12748 ( .A1(n10335), .A2(n10334), .ZN(n10336) );
  NAND2_X1 U12749 ( .A1(n15087), .A2(n10444), .ZN(n10338) );
  NAND2_X1 U12750 ( .A1(n14399), .A2(n10451), .ZN(n10337) );
  NAND2_X1 U12751 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  XNOR2_X1 U12752 ( .A(n10339), .B(n10701), .ZN(n10343) );
  AND2_X1 U12753 ( .A1(n14399), .A2(n6967), .ZN(n10340) );
  AOI21_X1 U12754 ( .B1(n15087), .B2(n10451), .A(n10340), .ZN(n10341) );
  XNOR2_X1 U12755 ( .A(n10343), .B(n10341), .ZN(n15083) );
  INV_X1 U12756 ( .A(n10341), .ZN(n10342) );
  NAND2_X1 U12757 ( .A1(n15130), .A2(n10444), .ZN(n10345) );
  OR2_X1 U12758 ( .A1(n12412), .A2(n10445), .ZN(n10344) );
  NAND2_X1 U12759 ( .A1(n10345), .A2(n10344), .ZN(n10346) );
  XNOR2_X1 U12760 ( .A(n10346), .B(n10701), .ZN(n10348) );
  NOR2_X1 U12761 ( .A1(n12412), .A2(n10458), .ZN(n10347) );
  AOI21_X1 U12762 ( .B1(n15130), .B2(n10437), .A(n10347), .ZN(n10349) );
  XNOR2_X1 U12763 ( .A(n10348), .B(n10349), .ZN(n12393) );
  NAND2_X1 U12764 ( .A1(n12394), .A2(n12393), .ZN(n12392) );
  INV_X1 U12765 ( .A(n10348), .ZN(n10350) );
  OR2_X1 U12766 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  NAND2_X1 U12767 ( .A1(n14921), .A2(n10444), .ZN(n10353) );
  OR2_X1 U12768 ( .A1(n14560), .A2(n10445), .ZN(n10352) );
  NAND2_X1 U12769 ( .A1(n10353), .A2(n10352), .ZN(n10354) );
  XNOR2_X1 U12770 ( .A(n10354), .B(n10448), .ZN(n10357) );
  NOR2_X1 U12771 ( .A1(n14560), .A2(n10458), .ZN(n10355) );
  AOI21_X1 U12772 ( .B1(n14921), .B2(n10437), .A(n10355), .ZN(n10356) );
  XNOR2_X1 U12773 ( .A(n10357), .B(n10356), .ZN(n14269) );
  NAND2_X1 U12774 ( .A1(n10357), .A2(n10356), .ZN(n10358) );
  NAND2_X1 U12775 ( .A1(n14911), .A2(n10444), .ZN(n10360) );
  INV_X1 U12776 ( .A(n10368), .ZN(n10445) );
  OR2_X1 U12777 ( .A1(n14562), .A2(n10445), .ZN(n10359) );
  NAND2_X1 U12778 ( .A1(n10360), .A2(n10359), .ZN(n10361) );
  XNOR2_X1 U12779 ( .A(n10361), .B(n10448), .ZN(n10363) );
  INV_X1 U12780 ( .A(n14911), .ZN(n14563) );
  OAI22_X1 U12781 ( .A1(n14563), .A2(n10445), .B1(n14562), .B2(n10458), .ZN(
        n14382) );
  INV_X1 U12782 ( .A(n10362), .ZN(n10365) );
  INV_X1 U12783 ( .A(n10363), .ZN(n10364) );
  NAND2_X1 U12784 ( .A1(n10365), .A2(n10364), .ZN(n14380) );
  XNOR2_X1 U12785 ( .A(n10366), .B(n10367), .ZN(n14318) );
  OAI22_X1 U12786 ( .A1(n8244), .A2(n10457), .B1(n14566), .B2(n10445), .ZN(
        n10369) );
  XOR2_X1 U12787 ( .A(n10701), .B(n10369), .Z(n14325) );
  AOI22_X1 U12788 ( .A1(n14899), .A2(n10437), .B1(n6967), .B2(n14565), .ZN(
        n14324) );
  INV_X1 U12789 ( .A(n14325), .ZN(n10371) );
  INV_X1 U12790 ( .A(n14324), .ZN(n10370) );
  NAND2_X1 U12791 ( .A1(n14893), .A2(n10444), .ZN(n10373) );
  NAND2_X1 U12792 ( .A1(n14398), .A2(n10437), .ZN(n10372) );
  NAND2_X1 U12793 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  XNOR2_X1 U12794 ( .A(n10374), .B(n10701), .ZN(n10377) );
  AND2_X1 U12795 ( .A1(n14398), .A2(n6967), .ZN(n10375) );
  AOI21_X1 U12796 ( .B1(n14893), .B2(n10451), .A(n10375), .ZN(n10378) );
  XNOR2_X1 U12797 ( .A(n10377), .B(n10378), .ZN(n14361) );
  XNOR2_X1 U12798 ( .A(n10376), .B(n10381), .ZN(n14288) );
  INV_X1 U12799 ( .A(n10377), .ZN(n10379) );
  NAND2_X1 U12800 ( .A1(n10379), .A2(n10378), .ZN(n14286) );
  NAND3_X1 U12801 ( .A1(n14359), .A2(n14288), .A3(n14286), .ZN(n14287) );
  OAI22_X1 U12802 ( .A1(n10382), .A2(n10445), .B1(n14571), .B2(n10458), .ZN(
        n10387) );
  NAND2_X1 U12803 ( .A1(n14883), .A2(n10444), .ZN(n10384) );
  NAND2_X1 U12804 ( .A1(n14396), .A2(n10451), .ZN(n10383) );
  NAND2_X1 U12805 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  XNOR2_X1 U12806 ( .A(n10385), .B(n10701), .ZN(n10386) );
  XOR2_X1 U12807 ( .A(n10387), .B(n10386), .Z(n14342) );
  NAND2_X1 U12808 ( .A1(n14877), .A2(n10444), .ZN(n10389) );
  NAND2_X1 U12809 ( .A1(n14573), .A2(n10451), .ZN(n10388) );
  NAND2_X1 U12810 ( .A1(n10389), .A2(n10388), .ZN(n10390) );
  XNOR2_X1 U12811 ( .A(n10390), .B(n10701), .ZN(n10394) );
  NAND2_X1 U12812 ( .A1(n14877), .A2(n10451), .ZN(n10392) );
  NAND2_X1 U12813 ( .A1(n14573), .A2(n6967), .ZN(n10391) );
  NAND2_X1 U12814 ( .A1(n10392), .A2(n10391), .ZN(n10393) );
  NOR2_X1 U12815 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  AOI21_X1 U12816 ( .B1(n10394), .B2(n10393), .A(n10395), .ZN(n14293) );
  INV_X1 U12817 ( .A(n10395), .ZN(n14351) );
  OAI22_X1 U12818 ( .A1(n14692), .A2(n10457), .B1(n14575), .B2(n10445), .ZN(
        n10396) );
  XNOR2_X1 U12819 ( .A(n10396), .B(n10448), .ZN(n10399) );
  OR2_X1 U12820 ( .A1(n14692), .A2(n10445), .ZN(n10398) );
  NAND2_X1 U12821 ( .A1(n14548), .A2(n6967), .ZN(n10397) );
  AND2_X1 U12822 ( .A1(n10398), .A2(n10397), .ZN(n10400) );
  NAND2_X1 U12823 ( .A1(n10399), .A2(n10400), .ZN(n10404) );
  INV_X1 U12824 ( .A(n10399), .ZN(n10402) );
  INV_X1 U12825 ( .A(n10400), .ZN(n10401) );
  NAND2_X1 U12826 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  NAND2_X1 U12827 ( .A1(n10404), .A2(n10403), .ZN(n14350) );
  INV_X1 U12828 ( .A(n10404), .ZN(n14276) );
  NAND2_X1 U12829 ( .A1(n14866), .A2(n10444), .ZN(n10406) );
  NAND2_X1 U12830 ( .A1(n14395), .A2(n10451), .ZN(n10405) );
  NAND2_X1 U12831 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  XNOR2_X1 U12832 ( .A(n10407), .B(n10448), .ZN(n10409) );
  NOR2_X1 U12833 ( .A1(n14576), .A2(n10458), .ZN(n10408) );
  AOI21_X1 U12834 ( .B1(n14866), .B2(n10451), .A(n10408), .ZN(n10410) );
  NAND2_X1 U12835 ( .A1(n10409), .A2(n10410), .ZN(n14333) );
  INV_X1 U12836 ( .A(n10409), .ZN(n10412) );
  INV_X1 U12837 ( .A(n10410), .ZN(n10411) );
  NAND2_X1 U12838 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  AND2_X1 U12839 ( .A1(n14333), .A2(n10413), .ZN(n14275) );
  NAND2_X1 U12840 ( .A1(n14857), .A2(n10444), .ZN(n10415) );
  NAND2_X1 U12841 ( .A1(n14577), .A2(n10451), .ZN(n10414) );
  NAND2_X1 U12842 ( .A1(n10415), .A2(n10414), .ZN(n10416) );
  XNOR2_X1 U12843 ( .A(n10416), .B(n10448), .ZN(n10419) );
  AND2_X1 U12844 ( .A1(n14577), .A2(n6967), .ZN(n10418) );
  AOI21_X1 U12845 ( .B1(n14857), .B2(n10451), .A(n10418), .ZN(n10420) );
  NAND2_X1 U12846 ( .A1(n10419), .A2(n10420), .ZN(n10424) );
  INV_X1 U12847 ( .A(n10419), .ZN(n10422) );
  INV_X1 U12848 ( .A(n10420), .ZN(n10421) );
  NAND2_X1 U12849 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  NAND2_X1 U12850 ( .A1(n10424), .A2(n10423), .ZN(n14332) );
  INV_X1 U12851 ( .A(n10424), .ZN(n14306) );
  NAND2_X1 U12852 ( .A1(n14647), .A2(n10444), .ZN(n10426) );
  OR2_X1 U12853 ( .A1(n14579), .A2(n10445), .ZN(n10425) );
  NAND2_X1 U12854 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  XNOR2_X1 U12855 ( .A(n10427), .B(n10448), .ZN(n10430) );
  NOR2_X1 U12856 ( .A1(n14579), .A2(n10458), .ZN(n10428) );
  AOI21_X1 U12857 ( .B1(n14647), .B2(n10451), .A(n10428), .ZN(n10429) );
  NAND2_X1 U12858 ( .A1(n10430), .A2(n10429), .ZN(n10432) );
  OR2_X1 U12859 ( .A1(n10430), .A2(n10429), .ZN(n10431) );
  AND2_X1 U12860 ( .A1(n10432), .A2(n10431), .ZN(n14305) );
  NAND2_X1 U12861 ( .A1(n14843), .A2(n10444), .ZN(n10434) );
  OR2_X1 U12862 ( .A1(n14309), .A2(n10445), .ZN(n10433) );
  NAND2_X1 U12863 ( .A1(n10434), .A2(n10433), .ZN(n10435) );
  XNOR2_X1 U12864 ( .A(n10435), .B(n10448), .ZN(n10439) );
  INV_X1 U12865 ( .A(n10439), .ZN(n10441) );
  NOR2_X1 U12866 ( .A1(n14309), .A2(n10458), .ZN(n10436) );
  AOI21_X1 U12867 ( .B1(n14843), .B2(n10437), .A(n10436), .ZN(n10438) );
  INV_X1 U12868 ( .A(n10438), .ZN(n10440) );
  AND2_X1 U12869 ( .A1(n10439), .A2(n10438), .ZN(n10442) );
  AOI21_X1 U12870 ( .B1(n10441), .B2(n10440), .A(n10442), .ZN(n14370) );
  NAND2_X1 U12871 ( .A1(n14369), .A2(n14370), .ZN(n14368) );
  INV_X1 U12872 ( .A(n10442), .ZN(n10443) );
  NAND2_X1 U12873 ( .A1(n14368), .A2(n10443), .ZN(n14259) );
  NAND2_X1 U12874 ( .A1(n14837), .A2(n10444), .ZN(n10447) );
  OR2_X1 U12875 ( .A1(n14550), .A2(n10445), .ZN(n10446) );
  NAND2_X1 U12876 ( .A1(n10447), .A2(n10446), .ZN(n10449) );
  XNOR2_X1 U12877 ( .A(n10449), .B(n10448), .ZN(n10453) );
  INV_X1 U12878 ( .A(n10453), .ZN(n10455) );
  NOR2_X1 U12879 ( .A1(n14550), .A2(n10458), .ZN(n10450) );
  AOI21_X1 U12880 ( .B1(n14837), .B2(n10451), .A(n10450), .ZN(n10452) );
  INV_X1 U12881 ( .A(n10452), .ZN(n10454) );
  AND2_X1 U12882 ( .A1(n10453), .A2(n10452), .ZN(n10456) );
  AOI21_X1 U12883 ( .B1(n10455), .B2(n10454), .A(n10456), .ZN(n14260) );
  OAI22_X1 U12884 ( .A1(n14610), .A2(n10457), .B1(n14551), .B2(n10445), .ZN(
        n10461) );
  OAI22_X1 U12885 ( .A1(n14610), .A2(n10445), .B1(n14551), .B2(n10458), .ZN(
        n10459) );
  XNOR2_X1 U12886 ( .A(n10459), .B(n10701), .ZN(n10460) );
  XOR2_X1 U12887 ( .A(n10461), .B(n10460), .Z(n10462) );
  NAND2_X1 U12888 ( .A1(n12207), .A2(P1_B_REG_SCAN_IN), .ZN(n10464) );
  OAI22_X1 U12889 ( .A1(n10477), .A2(n10464), .B1(P1_B_REG_SCAN_IN), .B2(
        n12207), .ZN(n10466) );
  NAND2_X1 U12890 ( .A1(n14952), .A2(n12207), .ZN(n10551) );
  OAI21_X1 U12891 ( .B1(n10708), .B2(P1_D_REG_0__SCAN_IN), .A(n10551), .ZN(
        n11318) );
  NOR4_X1 U12892 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10470) );
  NOR4_X1 U12893 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10469) );
  NOR4_X1 U12894 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10468) );
  NOR4_X1 U12895 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10467) );
  NAND4_X1 U12896 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10476) );
  NOR2_X1 U12897 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n10474) );
  NOR4_X1 U12898 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10473) );
  NOR4_X1 U12899 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10472) );
  NOR4_X1 U12900 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10471) );
  NAND4_X1 U12901 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  NOR2_X1 U12902 ( .A1(n10476), .A2(n10475), .ZN(n10709) );
  AND2_X1 U12903 ( .A1(n10709), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10478) );
  INV_X1 U12904 ( .A(n10477), .ZN(n12328) );
  NAND2_X1 U12905 ( .A1(n14952), .A2(n12328), .ZN(n10706) );
  OAI21_X1 U12906 ( .B1(n10708), .B2(n10478), .A(n10706), .ZN(n11136) );
  OR2_X1 U12907 ( .A1(n11318), .A2(n11136), .ZN(n10485) );
  NAND2_X1 U12908 ( .A1(n10480), .A2(n10479), .ZN(n11156) );
  NAND2_X2 U12909 ( .A1(n11140), .A2(n11156), .ZN(n15283) );
  NAND2_X1 U12910 ( .A1(n10481), .A2(n10552), .ZN(n11139) );
  NOR2_X2 U12911 ( .A1(n10485), .A2(n10482), .ZN(n15081) );
  NAND2_X1 U12912 ( .A1(n10485), .A2(n11140), .ZN(n10715) );
  INV_X1 U12913 ( .A(n11139), .ZN(n10548) );
  NAND2_X1 U12914 ( .A1(n10715), .A2(n10548), .ZN(n15093) );
  OR2_X1 U12915 ( .A1(n14550), .A2(n15095), .ZN(n10484) );
  AND2_X1 U12916 ( .A1(n8555), .A2(n10560), .ZN(n14987) );
  NAND2_X1 U12917 ( .A1(n14393), .A2(n14987), .ZN(n10483) );
  NAND2_X1 U12918 ( .A1(n10484), .A2(n10483), .ZN(n14829) );
  OR2_X1 U12919 ( .A1(n11322), .A2(n10485), .ZN(n15079) );
  INV_X2 U12920 ( .A(n15079), .ZN(n15105) );
  INV_X1 U12921 ( .A(n10486), .ZN(n10487) );
  NAND2_X1 U12922 ( .A1(n10715), .A2(n10487), .ZN(n10488) );
  INV_X1 U12923 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10489) );
  OAI22_X1 U12924 ( .A1(n15090), .A2(n14606), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10489), .ZN(n10490) );
  AOI21_X1 U12925 ( .B1(n14829), .B2(n15105), .A(n10490), .ZN(n10491) );
  INV_X1 U12926 ( .A(n10492), .ZN(n10493) );
  AND2_X2 U12927 ( .A1(n7586), .A2(n10552), .ZN(P1_U4016) );
  NOR2_X1 U12928 ( .A1(n12176), .A2(n10494), .ZN(n10750) );
  INV_X1 U12929 ( .A(n10495), .ZN(n11348) );
  NAND2_X1 U12930 ( .A1(n10497), .A2(P2_U3088), .ZN(n14252) );
  NOR2_X1 U12931 ( .A1(n10497), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14246) );
  INV_X2 U12932 ( .A(n14246), .ZN(n14254) );
  OAI222_X1 U12933 ( .A1(n14252), .A2(n10496), .B1(n14254), .B2(n10499), .C1(
        n10869), .C2(P2_U3088), .ZN(P2_U3326) );
  AND2_X1 U12934 ( .A1(n10502), .A2(P1_U3086), .ZN(n12509) );
  INV_X2 U12935 ( .A(n12509), .ZN(n12208) );
  NOR2_X1 U12936 ( .A1(n10497), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12510) );
  INV_X1 U12937 ( .A(n12510), .ZN(n14949) );
  OAI222_X1 U12938 ( .A1(P1_U3086), .A2(n10598), .B1(n12208), .B2(n10499), 
        .C1(n10498), .C2(n14949), .ZN(P1_U3354) );
  OAI222_X1 U12939 ( .A1(n14949), .A2(n10500), .B1(n12208), .B2(n10508), .C1(
        P1_U3086), .C2(n14429), .ZN(P1_U3353) );
  AND2_X1 U12940 ( .A1(n10501), .A2(P3_U3151), .ZN(n11186) );
  INV_X2 U12941 ( .A(n11186), .ZN(n12971) );
  INV_X1 U12942 ( .A(SI_1_), .ZN(n10505) );
  NAND2_X1 U12943 ( .A1(n10497), .A2(P3_U3151), .ZN(n13672) );
  INV_X1 U12944 ( .A(n10503), .ZN(n10504) );
  OAI222_X1 U12945 ( .A1(P3_U3151), .A2(n11569), .B1(n12971), .B2(n10505), 
        .C1(n13672), .C2(n10504), .ZN(P3_U3294) );
  INV_X1 U12946 ( .A(n14252), .ZN(n10507) );
  AOI22_X1 U12947 ( .A1(n10507), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n13805), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10506) );
  OAI21_X1 U12948 ( .B1(n10510), .B2(n14254), .A(n10506), .ZN(P2_U3324) );
  INV_X1 U12949 ( .A(n10507), .ZN(n14249) );
  INV_X1 U12950 ( .A(n10775), .ZN(n15303) );
  OAI222_X1 U12951 ( .A1(n14249), .A2(n10509), .B1(n14254), .B2(n10508), .C1(
        P2_U3088), .C2(n15303), .ZN(P2_U3325) );
  OAI222_X1 U12952 ( .A1(n14949), .A2(n10511), .B1(n12208), .B2(n10510), .C1(
        P1_U3086), .C2(n14446), .ZN(P1_U3352) );
  INV_X1 U12953 ( .A(n13672), .ZN(n13662) );
  INV_X1 U12954 ( .A(n13662), .ZN(n12279) );
  OAI222_X1 U12955 ( .A1(n12279), .A2(n10513), .B1(n12971), .B2(n10512), .C1(
        n7338), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12956 ( .A1(n12279), .A2(n10515), .B1(n12971), .B2(n10514), .C1(
        n11999), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U12957 ( .A1(n12279), .A2(n10517), .B1(n12971), .B2(n10516), .C1(
        n11926), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12958 ( .A(n13190), .ZN(n10518) );
  OAI222_X1 U12959 ( .A1(n12279), .A2(n10520), .B1(n12971), .B2(n10519), .C1(
        n10518), .C2(P3_U3151), .ZN(P3_U3284) );
  OAI222_X1 U12960 ( .A1(n7564), .A2(P3_U3151), .B1(n12279), .B2(n10521), .C1(
        n7242), .C2(n12971), .ZN(P3_U3293) );
  OAI222_X1 U12961 ( .A1(n11696), .A2(P3_U3151), .B1(n12279), .B2(n10523), 
        .C1(n10522), .C2(n12971), .ZN(P3_U3291) );
  OAI222_X1 U12962 ( .A1(n11577), .A2(P3_U3151), .B1(n12279), .B2(n10525), 
        .C1(n10524), .C2(n12971), .ZN(P3_U3292) );
  INV_X1 U12963 ( .A(n10526), .ZN(n10528) );
  INV_X1 U12964 ( .A(SI_6_), .ZN(n10527) );
  OAI222_X1 U12965 ( .A1(n11863), .A2(P3_U3151), .B1(n12279), .B2(n10528), 
        .C1(n10527), .C2(n12971), .ZN(P3_U3289) );
  OAI222_X1 U12966 ( .A1(n11598), .A2(P3_U3151), .B1(n12279), .B2(n10530), 
        .C1(n10529), .C2(n12971), .ZN(P3_U3290) );
  INV_X1 U12967 ( .A(n10531), .ZN(n10533) );
  OAI222_X1 U12968 ( .A1(n6887), .A2(P3_U3151), .B1(n12279), .B2(n10533), .C1(
        n10532), .C2(n12971), .ZN(P3_U3295) );
  INV_X1 U12969 ( .A(SI_8_), .ZN(n10536) );
  INV_X1 U12970 ( .A(n10534), .ZN(n10535) );
  OAI222_X1 U12971 ( .A1(P3_U3151), .A2(n15522), .B1(n12971), .B2(n10536), 
        .C1(n12279), .C2(n10535), .ZN(P3_U3287) );
  INV_X1 U12972 ( .A(n10537), .ZN(n10539) );
  OAI222_X1 U12973 ( .A1(n14949), .A2(n10538), .B1(n12208), .B2(n10539), .C1(
        P1_U3086), .C2(n14456), .ZN(P1_U3351) );
  OAI222_X1 U12974 ( .A1(n14249), .A2(n10540), .B1(n14254), .B2(n10539), .C1(
        P2_U3088), .C2(n13819), .ZN(P2_U3323) );
  INV_X1 U12975 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10542) );
  INV_X1 U12976 ( .A(n10541), .ZN(n10543) );
  INV_X1 U12977 ( .A(n10619), .ZN(n10613) );
  OAI222_X1 U12978 ( .A1(n14949), .A2(n10542), .B1(n12208), .B2(n10543), .C1(
        P1_U3086), .C2(n10613), .ZN(P1_U3350) );
  INV_X1 U12979 ( .A(n10780), .ZN(n15323) );
  OAI222_X1 U12980 ( .A1(n14249), .A2(n10544), .B1(n14254), .B2(n10543), .C1(
        P2_U3088), .C2(n15323), .ZN(P2_U3322) );
  INV_X1 U12981 ( .A(n10545), .ZN(n10547) );
  OAI222_X1 U12982 ( .A1(n12279), .A2(n10547), .B1(n12971), .B2(n10546), .C1(
        n15534), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U12983 ( .A1(n10548), .A2(n10708), .ZN(n15226) );
  INV_X1 U12984 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10550) );
  INV_X1 U12985 ( .A(n10706), .ZN(n10549) );
  AOI22_X1 U12986 ( .A1(n15226), .A2(n10550), .B1(n10549), .B2(n10552), .ZN(
        P1_U3446) );
  INV_X1 U12987 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10554) );
  INV_X1 U12988 ( .A(n10551), .ZN(n10553) );
  AOI22_X1 U12989 ( .A1(n15226), .A2(n10554), .B1(n10553), .B2(n10552), .ZN(
        P1_U3445) );
  INV_X1 U12990 ( .A(n10555), .ZN(n10557) );
  INV_X1 U12991 ( .A(n10620), .ZN(n10663) );
  OAI222_X1 U12992 ( .A1(n14949), .A2(n10556), .B1(n12208), .B2(n10557), .C1(
        P1_U3086), .C2(n10663), .ZN(P1_U3349) );
  INV_X1 U12993 ( .A(n10811), .ZN(n10788) );
  OAI222_X1 U12994 ( .A1(n14249), .A2(n10558), .B1(n14254), .B2(n10557), .C1(
        P2_U3088), .C2(n10788), .ZN(P2_U3321) );
  NAND2_X1 U12995 ( .A1(n10560), .A2(n10559), .ZN(n10561) );
  NAND2_X1 U12996 ( .A1(n10562), .A2(n10561), .ZN(n10587) );
  AND2_X1 U12997 ( .A1(n11139), .A2(n12180), .ZN(n10586) );
  INV_X1 U12998 ( .A(n10586), .ZN(n10563) );
  AND2_X1 U12999 ( .A1(n10587), .A2(n10563), .ZN(n15177) );
  NOR2_X1 U13000 ( .A1(n15177), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13001 ( .A(n10564), .ZN(n10567) );
  AOI22_X1 U13002 ( .A1(n10636), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n12510), .ZN(n10565) );
  OAI21_X1 U13003 ( .B1(n10567), .B2(n12208), .A(n10565), .ZN(P1_U3348) );
  INV_X1 U13004 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10568) );
  INV_X1 U13005 ( .A(n13836), .ZN(n10566) );
  OAI222_X1 U13006 ( .A1(n14249), .A2(n10568), .B1(n14254), .B2(n10567), .C1(
        P2_U3088), .C2(n10566), .ZN(P2_U3320) );
  OAI222_X1 U13007 ( .A1(n13209), .A2(P3_U3151), .B1(n12279), .B2(n10570), 
        .C1(n10569), .C2(n12971), .ZN(P3_U3282) );
  INV_X1 U13008 ( .A(n10571), .ZN(n10573) );
  INV_X1 U13009 ( .A(n10671), .ZN(n10675) );
  OAI222_X1 U13010 ( .A1(n14949), .A2(n10572), .B1(n12208), .B2(n10573), .C1(
        P1_U3086), .C2(n10675), .ZN(P1_U3347) );
  INV_X1 U13011 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10574) );
  OAI222_X1 U13012 ( .A1(n14249), .A2(n10574), .B1(n14254), .B2(n10573), .C1(
        P2_U3088), .C2(n13850), .ZN(P2_U3319) );
  INV_X1 U13013 ( .A(n10575), .ZN(n10581) );
  AOI22_X1 U13014 ( .A1(n10731), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n12510), .ZN(n10576) );
  OAI21_X1 U13015 ( .B1(n10581), .B2(n12208), .A(n10576), .ZN(P1_U3346) );
  OAI222_X1 U13016 ( .A1(n12279), .A2(n10578), .B1(n12971), .B2(n10577), .C1(
        n13207), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U13017 ( .A(P1_U4016), .ZN(n14409) );
  NAND2_X1 U13018 ( .A1(n14409), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n10579) );
  OAI21_X1 U13019 ( .B1(n14562), .B2(n14409), .A(n10579), .ZN(P1_U3575) );
  NAND2_X1 U13020 ( .A1(n14409), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n10580) );
  OAI21_X1 U13021 ( .B1(n14560), .B2(n14409), .A(n10580), .ZN(P1_U3574) );
  INV_X1 U13022 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10582) );
  INV_X1 U13023 ( .A(n10820), .ZN(n15342) );
  OAI222_X1 U13024 ( .A1(n14249), .A2(n10582), .B1(n14254), .B2(n10581), .C1(
        P2_U3088), .C2(n15342), .ZN(P2_U3318) );
  NAND2_X1 U13025 ( .A1(n10583), .A2(P1_U4016), .ZN(n10584) );
  OAI21_X1 U13026 ( .B1(P1_U4016), .B2(n10585), .A(n10584), .ZN(P1_U3591) );
  OR2_X1 U13027 ( .A1(n10587), .A2(n10586), .ZN(n15180) );
  INV_X1 U13028 ( .A(n6988), .ZN(n15169) );
  INV_X1 U13029 ( .A(n14456), .ZN(n10592) );
  MUX2_X1 U13030 ( .A(n10590), .B(P1_REG1_REG_2__SCAN_IN), .S(n14429), .Z(
        n14436) );
  XNOR2_X1 U13031 ( .A(n10598), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n14414) );
  AND2_X1 U13032 ( .A1(n14955), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U13033 ( .A1(n14414), .A2(n14413), .ZN(n14412) );
  INV_X1 U13034 ( .A(n10598), .ZN(n14417) );
  NAND2_X1 U13035 ( .A1(n14417), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13036 ( .A1(n14412), .A2(n10589), .ZN(n14435) );
  NAND2_X1 U13037 ( .A1(n14436), .A2(n14435), .ZN(n14434) );
  OAI21_X1 U13038 ( .B1(n10590), .B2(n14429), .A(n14434), .ZN(n14443) );
  MUX2_X1 U13039 ( .A(n10591), .B(P1_REG1_REG_3__SCAN_IN), .S(n14446), .Z(
        n14444) );
  NAND2_X1 U13040 ( .A1(n14443), .A2(n14444), .ZN(n14442) );
  OAI21_X1 U13041 ( .B1(n10591), .B2(n14446), .A(n14442), .ZN(n14460) );
  INV_X1 U13042 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15294) );
  MUX2_X1 U13043 ( .A(n15294), .B(P1_REG1_REG_4__SCAN_IN), .S(n14456), .Z(
        n14461) );
  AND2_X1 U13044 ( .A1(n14460), .A2(n14461), .ZN(n14458) );
  MUX2_X1 U13045 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10593), .S(n10619), .Z(
        n10594) );
  NAND2_X1 U13046 ( .A1(n10595), .A2(n10594), .ZN(n10614) );
  OAI21_X1 U13047 ( .B1(n10595), .B2(n10594), .A(n10614), .ZN(n10609) );
  OR2_X1 U13048 ( .A1(n8555), .A2(n6988), .ZN(n10596) );
  INV_X1 U13049 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10597) );
  MUX2_X1 U13050 ( .A(n10597), .B(P1_REG2_REG_2__SCAN_IN), .S(n14429), .Z(
        n14433) );
  MUX2_X1 U13051 ( .A(n10599), .B(P1_REG2_REG_1__SCAN_IN), .S(n10598), .Z(
        n14416) );
  AND2_X1 U13052 ( .A1(n14955), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U13053 ( .A1(n14416), .A2(n10600), .ZN(n14415) );
  NAND2_X1 U13054 ( .A1(n14417), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13055 ( .A1(n14415), .A2(n10601), .ZN(n14432) );
  AND2_X1 U13056 ( .A1(n14433), .A2(n14432), .ZN(n14431) );
  NOR2_X1 U13057 ( .A1(n14429), .A2(n10597), .ZN(n14445) );
  INV_X1 U13058 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11179) );
  MUX2_X1 U13059 ( .A(n11179), .B(P1_REG2_REG_3__SCAN_IN), .S(n14446), .Z(
        n10602) );
  OAI21_X1 U13060 ( .B1(n14431), .B2(n14445), .A(n10602), .ZN(n14465) );
  INV_X1 U13061 ( .A(n14446), .ZN(n10603) );
  NAND2_X1 U13062 ( .A1(n10603), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14464) );
  MUX2_X1 U13063 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7953), .S(n14456), .Z(
        n14463) );
  AOI21_X1 U13064 ( .B1(n14465), .B2(n14464), .A(n14463), .ZN(n14462) );
  NOR2_X1 U13065 ( .A1(n14456), .A2(n7953), .ZN(n10605) );
  MUX2_X1 U13066 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11215), .S(n10619), .Z(
        n10604) );
  OAI21_X1 U13067 ( .B1(n14462), .B2(n10605), .A(n10604), .ZN(n10657) );
  INV_X1 U13068 ( .A(n10657), .ZN(n10607) );
  NOR3_X1 U13069 ( .A1(n14462), .A2(n10605), .A3(n10604), .ZN(n10606) );
  NOR3_X1 U13070 ( .A1(n15183), .A2(n10607), .A3(n10606), .ZN(n10608) );
  AOI21_X1 U13071 ( .B1(n15188), .B2(n10609), .A(n10608), .ZN(n10612) );
  NAND2_X1 U13072 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11064) );
  INV_X1 U13073 ( .A(n11064), .ZN(n10610) );
  AOI21_X1 U13074 ( .B1(n15177), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10610), .ZN(
        n10611) );
  OAI211_X1 U13075 ( .C1(n10613), .C2(n15193), .A(n10612), .B(n10611), .ZN(
        P1_U3248) );
  OAI21_X1 U13076 ( .B1(n10619), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10614), .ZN(
        n10665) );
  INV_X1 U13077 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10615) );
  MUX2_X1 U13078 ( .A(n10615), .B(P1_REG1_REG_6__SCAN_IN), .S(n10620), .Z(
        n10666) );
  NOR2_X1 U13079 ( .A1(n10665), .A2(n10666), .ZN(n10664) );
  INV_X1 U13080 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10616) );
  MUX2_X1 U13081 ( .A(n10616), .B(P1_REG1_REG_7__SCAN_IN), .S(n10636), .Z(
        n10617) );
  NOR2_X1 U13082 ( .A1(n10618), .A2(n10617), .ZN(n10635) );
  AOI211_X1 U13083 ( .C1(n10618), .C2(n10617), .A(n12377), .B(n10635), .ZN(
        n10630) );
  NAND2_X1 U13084 ( .A1(n10619), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10656) );
  MUX2_X1 U13085 ( .A(n8000), .B(P1_REG2_REG_6__SCAN_IN), .S(n10620), .Z(
        n10655) );
  AOI21_X1 U13086 ( .B1(n10657), .B2(n10656), .A(n10655), .ZN(n10654) );
  NOR2_X1 U13087 ( .A1(n10663), .A2(n8000), .ZN(n10623) );
  MUX2_X1 U13088 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10621), .S(n10636), .Z(
        n10622) );
  OAI21_X1 U13089 ( .B1(n10654), .B2(n10623), .A(n10622), .ZN(n10633) );
  INV_X1 U13090 ( .A(n10633), .ZN(n10625) );
  NOR3_X1 U13091 ( .A1(n10654), .A2(n10623), .A3(n10622), .ZN(n10624) );
  NOR3_X1 U13092 ( .A1(n10625), .A2(n10624), .A3(n15183), .ZN(n10629) );
  INV_X1 U13093 ( .A(n10636), .ZN(n10627) );
  NAND2_X1 U13094 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11194) );
  NAND2_X1 U13095 ( .A1(n15177), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10626) );
  OAI211_X1 U13096 ( .C1(n15193), .C2(n10627), .A(n11194), .B(n10626), .ZN(
        n10628) );
  OR3_X1 U13097 ( .A1(n10630), .A2(n10629), .A3(n10628), .ZN(P1_U3250) );
  NAND2_X1 U13098 ( .A1(n10636), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10632) );
  INV_X1 U13099 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10674) );
  MUX2_X1 U13100 ( .A(n10674), .B(P1_REG2_REG_8__SCAN_IN), .S(n10671), .Z(
        n10631) );
  AOI21_X1 U13101 ( .B1(n10633), .B2(n10632), .A(n10631), .ZN(n10678) );
  NAND3_X1 U13102 ( .A1(n10633), .A2(n10632), .A3(n10631), .ZN(n10634) );
  INV_X1 U13103 ( .A(n15183), .ZN(n14515) );
  NAND2_X1 U13104 ( .A1(n10634), .A2(n14515), .ZN(n10645) );
  MUX2_X1 U13105 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10637), .S(n10671), .Z(
        n10638) );
  NAND2_X1 U13106 ( .A1(n10639), .A2(n10638), .ZN(n10670) );
  OAI21_X1 U13107 ( .B1(n10639), .B2(n10638), .A(n10670), .ZN(n10640) );
  NAND2_X1 U13108 ( .A1(n10640), .A2(n15188), .ZN(n10644) );
  NAND2_X1 U13109 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11473) );
  INV_X1 U13110 ( .A(n11473), .ZN(n10642) );
  NOR2_X1 U13111 ( .A1(n15193), .A2(n10675), .ZN(n10641) );
  AOI211_X1 U13112 ( .C1(n15177), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10642), .B(
        n10641), .ZN(n10643) );
  OAI211_X1 U13113 ( .C1(n10678), .C2(n10645), .A(n10644), .B(n10643), .ZN(
        P1_U3251) );
  INV_X1 U13114 ( .A(n10646), .ZN(n10648) );
  INV_X1 U13115 ( .A(n13248), .ZN(n15012) );
  OAI222_X1 U13116 ( .A1(n12279), .A2(n10648), .B1(n12971), .B2(n10647), .C1(
        n15012), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U13117 ( .A1(n12755), .A2(P2_U3947), .ZN(n10649) );
  OAI21_X1 U13118 ( .B1(n10790), .B2(P2_U3947), .A(n10649), .ZN(P2_U3544) );
  INV_X1 U13119 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10651) );
  INV_X1 U13120 ( .A(n10650), .ZN(n10652) );
  INV_X1 U13121 ( .A(n10854), .ZN(n10826) );
  OAI222_X1 U13122 ( .A1(n14249), .A2(n10651), .B1(n14254), .B2(n10652), .C1(
        P2_U3088), .C2(n10826), .ZN(P2_U3317) );
  INV_X1 U13123 ( .A(n10833), .ZN(n10837) );
  OAI222_X1 U13124 ( .A1(n14949), .A2(n10653), .B1(n12208), .B2(n10652), .C1(
        P1_U3086), .C2(n10837), .ZN(P1_U3345) );
  INV_X1 U13125 ( .A(n10654), .ZN(n10659) );
  NAND3_X1 U13126 ( .A1(n10657), .A2(n10656), .A3(n10655), .ZN(n10658) );
  NAND3_X1 U13127 ( .A1(n14515), .A2(n10659), .A3(n10658), .ZN(n10662) );
  INV_X1 U13128 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11115) );
  NOR2_X1 U13129 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11115), .ZN(n10660) );
  AOI21_X1 U13130 ( .B1(n15177), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10660), .ZN(
        n10661) );
  OAI211_X1 U13131 ( .C1(n15193), .C2(n10663), .A(n10662), .B(n10661), .ZN(
        n10668) );
  AOI211_X1 U13132 ( .C1(n10666), .C2(n10665), .A(n12377), .B(n10664), .ZN(
        n10667) );
  OR2_X1 U13133 ( .A1(n10668), .A2(n10667), .ZN(P1_U3249) );
  MUX2_X1 U13134 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10669), .S(n10731), .Z(
        n10673) );
  OAI21_X1 U13135 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10671), .A(n10670), .ZN(
        n10672) );
  NAND2_X1 U13136 ( .A1(n10672), .A2(n10673), .ZN(n10728) );
  OAI21_X1 U13137 ( .B1(n10673), .B2(n10672), .A(n10728), .ZN(n10686) );
  NOR2_X1 U13138 ( .A1(n10675), .A2(n10674), .ZN(n10677) );
  MUX2_X1 U13139 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11701), .S(n10731), .Z(
        n10676) );
  OAI21_X1 U13140 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10734) );
  INV_X1 U13141 ( .A(n10734), .ZN(n10680) );
  NOR3_X1 U13142 ( .A1(n10678), .A2(n10677), .A3(n10676), .ZN(n10679) );
  NOR3_X1 U13143 ( .A1(n10680), .A2(n10679), .A3(n15183), .ZN(n10685) );
  INV_X1 U13144 ( .A(n10731), .ZN(n10683) );
  NOR2_X1 U13145 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11950), .ZN(n10681) );
  AOI21_X1 U13146 ( .B1(n15177), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10681), .ZN(
        n10682) );
  OAI21_X1 U13147 ( .B1(n15193), .B2(n10683), .A(n10682), .ZN(n10684) );
  AOI211_X1 U13148 ( .C1(n10686), .C2(n15188), .A(n10685), .B(n10684), .ZN(
        n10687) );
  INV_X1 U13149 ( .A(n10687), .ZN(P1_U3252) );
  INV_X1 U13150 ( .A(n10688), .ZN(n10690) );
  INV_X1 U13151 ( .A(n10949), .ZN(n10943) );
  OAI222_X1 U13152 ( .A1(n14949), .A2(n10689), .B1(n12208), .B2(n10690), .C1(
        P1_U3086), .C2(n10943), .ZN(P1_U3344) );
  INV_X1 U13153 ( .A(n10910), .ZN(n10915) );
  OAI222_X1 U13154 ( .A1(n14249), .A2(n10691), .B1(n14254), .B2(n10690), .C1(
        P2_U3088), .C2(n10915), .ZN(P2_U3316) );
  INV_X1 U13155 ( .A(n10692), .ZN(n10694) );
  INV_X1 U13156 ( .A(n13251), .ZN(n13250) );
  OAI222_X1 U13157 ( .A1(n12279), .A2(n10694), .B1(n13250), .B2(P3_U3151), 
        .C1(n10693), .C2(n12971), .ZN(P3_U3279) );
  INV_X1 U13158 ( .A(n10695), .ZN(n10697) );
  OAI222_X1 U13159 ( .A1(n12279), .A2(n10697), .B1(n12971), .B2(n10696), .C1(
        n13288), .C2(P3_U3151), .ZN(P3_U3278) );
  OR2_X1 U13160 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  NAND2_X1 U13161 ( .A1(n10701), .A2(n10700), .ZN(n11141) );
  OR2_X1 U13162 ( .A1(n11141), .A2(n6681), .ZN(n15274) );
  NAND2_X1 U13163 ( .A1(n6681), .A2(n10702), .ZN(n15266) );
  INV_X1 U13164 ( .A(n15253), .ZN(n15260) );
  NAND2_X1 U13165 ( .A1(n15248), .A2(n15260), .ZN(n10705) );
  NOR3_X1 U13166 ( .A1(n11046), .A2(n10703), .A3(n14953), .ZN(n10704) );
  AND2_X1 U13167 ( .A1(n14410), .A2(n14987), .ZN(n14808) );
  AOI211_X1 U13168 ( .C1(n14803), .C2(n10705), .A(n10704), .B(n14808), .ZN(
        n15228) );
  OAI21_X1 U13169 ( .B1(n10708), .B2(P1_D_REG_1__SCAN_IN), .A(n10706), .ZN(
        n10707) );
  OAI211_X1 U13170 ( .C1(n10709), .C2(n10708), .A(n10707), .B(n11140), .ZN(
        n11319) );
  OR2_X1 U13171 ( .A1(n11319), .A2(n11318), .ZN(n10710) );
  NOR2_X2 U13172 ( .A1(n11322), .A2(n10710), .ZN(n15296) );
  NAND2_X1 U13173 ( .A1(n15300), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10711) );
  OAI21_X1 U13174 ( .B1(n15228), .B2(n15300), .A(n10711), .ZN(P1_U3528) );
  INV_X1 U13175 ( .A(n14808), .ZN(n10719) );
  OAI21_X1 U13176 ( .B1(n10714), .B2(n10713), .A(n10712), .ZN(n14422) );
  NAND2_X1 U13177 ( .A1(n14422), .A2(n15081), .ZN(n10718) );
  INV_X1 U13178 ( .A(n11322), .ZN(n10716) );
  NAND2_X1 U13179 ( .A1(n10716), .A2(n10715), .ZN(n10887) );
  AOI22_X1 U13180 ( .A1(n15088), .A2(n14806), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10887), .ZN(n10717) );
  OAI211_X1 U13181 ( .C1(n10719), .C2(n15079), .A(n10718), .B(n10717), .ZN(
        P1_U3232) );
  INV_X1 U13182 ( .A(n10720), .ZN(n10722) );
  OAI222_X1 U13183 ( .A1(P2_U3088), .A2(n15353), .B1(n14254), .B2(n10722), 
        .C1(n10721), .C2(n14249), .ZN(P2_U3315) );
  INV_X1 U13184 ( .A(n11093), .ZN(n10944) );
  OAI222_X1 U13185 ( .A1(P1_U3086), .A2(n10944), .B1(n12208), .B2(n10722), 
        .C1(n7613), .C2(n14949), .ZN(P1_U3343) );
  INV_X1 U13186 ( .A(n13660), .ZN(n10725) );
  XNOR2_X1 U13187 ( .A(n12233), .B(P3_B_REG_SCAN_IN), .ZN(n10723) );
  NAND2_X1 U13188 ( .A1(n10723), .A2(n12280), .ZN(n10724) );
  AND2_X1 U13189 ( .A1(n10726), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13190 ( .A1(n10726), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13191 ( .A1(n10726), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13192 ( .A1(n10726), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13193 ( .A1(n10726), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13194 ( .A1(n10726), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13195 ( .A1(n10726), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13196 ( .A1(n10726), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13197 ( .A1(n10726), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13198 ( .A1(n10726), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13199 ( .A1(n10726), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13200 ( .A1(n10726), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13201 ( .A1(n10726), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13202 ( .A1(n10726), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13203 ( .A1(n10726), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13204 ( .A1(n10726), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13205 ( .A1(n10726), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13206 ( .A1(n10726), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13207 ( .A1(n10726), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13208 ( .A1(n10726), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13209 ( .A1(n10726), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13210 ( .A1(n10726), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13211 ( .A1(n10726), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13212 ( .A1(n10726), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13213 ( .A1(n10726), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13214 ( .A1(n10726), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13215 ( .A1(n10726), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13216 ( .A1(n10726), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13217 ( .A1(n10726), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13218 ( .A1(n10726), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  INV_X1 U13219 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U13220 ( .A(n10727), .B(P1_REG1_REG_10__SCAN_IN), .S(n10833), .Z(
        n10730) );
  OAI21_X1 U13221 ( .B1(n10731), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10728), .ZN(
        n10729) );
  NOR2_X1 U13222 ( .A1(n10729), .A2(n10730), .ZN(n10832) );
  AOI211_X1 U13223 ( .C1(n10730), .C2(n10729), .A(n12377), .B(n10832), .ZN(
        n10741) );
  NAND2_X1 U13224 ( .A1(n10731), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10733) );
  MUX2_X1 U13225 ( .A(n8077), .B(P1_REG2_REG_10__SCAN_IN), .S(n10833), .Z(
        n10732) );
  AOI21_X1 U13226 ( .B1(n10734), .B2(n10733), .A(n10732), .ZN(n10840) );
  INV_X1 U13227 ( .A(n10840), .ZN(n10736) );
  NAND3_X1 U13228 ( .A1(n10734), .A2(n10733), .A3(n10732), .ZN(n10735) );
  NAND3_X1 U13229 ( .A1(n10736), .A2(n14515), .A3(n10735), .ZN(n10739) );
  NAND2_X1 U13230 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11974)
         );
  INV_X1 U13231 ( .A(n11974), .ZN(n10737) );
  AOI21_X1 U13232 ( .B1(n15177), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10737), 
        .ZN(n10738) );
  OAI211_X1 U13233 ( .C1(n15193), .C2(n10837), .A(n10739), .B(n10738), .ZN(
        n10740) );
  OR2_X1 U13234 ( .A1(n10741), .A2(n10740), .ZN(P1_U3253) );
  INV_X1 U13235 ( .A(n10742), .ZN(n10744) );
  INV_X1 U13236 ( .A(n13316), .ZN(n13302) );
  OAI222_X1 U13237 ( .A1(n12279), .A2(n10744), .B1(n12971), .B2(n10743), .C1(
        n13302), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13238 ( .A(n11077), .ZN(n11071) );
  INV_X1 U13239 ( .A(n10745), .ZN(n10789) );
  OAI222_X1 U13240 ( .A1(P2_U3088), .A2(n11071), .B1(n14254), .B2(n10789), 
        .C1(n7215), .C2(n14252), .ZN(P2_U3314) );
  AOI21_X1 U13241 ( .B1(n10749), .B2(n10748), .A(n10747), .ZN(n10751) );
  OR2_X1 U13242 ( .A1(n10751), .A2(n10750), .ZN(n10754) );
  AND2_X1 U13243 ( .A1(n10754), .A2(n10752), .ZN(n15302) );
  NOR2_X2 U13244 ( .A1(n10754), .A2(P2_U3088), .ZN(n15371) );
  NAND2_X1 U13245 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n11010) );
  INV_X1 U13246 ( .A(n11010), .ZN(n10771) );
  OR2_X1 U13247 ( .A1(n10752), .A2(P2_U3088), .ZN(n14243) );
  INV_X1 U13248 ( .A(n14243), .ZN(n10753) );
  AND2_X1 U13249 ( .A1(n10754), .A2(n10753), .ZN(n10783) );
  INV_X1 U13250 ( .A(n10782), .ZN(n13878) );
  NAND2_X1 U13251 ( .A1(n10783), .A2(n13878), .ZN(n13867) );
  INV_X1 U13252 ( .A(n13867), .ZN(n15372) );
  MUX2_X1 U13253 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10755), .S(n10775), .Z(
        n15312) );
  MUX2_X1 U13254 ( .A(n10756), .B(P2_REG2_REG_1__SCAN_IN), .S(n10869), .Z(
        n10758) );
  AND2_X1 U13255 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10757) );
  NAND2_X1 U13256 ( .A1(n10758), .A2(n10757), .ZN(n10873) );
  INV_X1 U13257 ( .A(n10869), .ZN(n10868) );
  NAND2_X1 U13258 ( .A1(n10868), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U13259 ( .A1(n10873), .A2(n10759), .ZN(n15313) );
  NAND2_X1 U13260 ( .A1(n15312), .A2(n15313), .ZN(n15311) );
  NAND2_X1 U13261 ( .A1(n10775), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13807) );
  NAND2_X1 U13262 ( .A1(n15311), .A2(n13807), .ZN(n10761) );
  MUX2_X1 U13263 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11419), .S(n13805), .Z(
        n10760) );
  NAND2_X1 U13264 ( .A1(n10761), .A2(n10760), .ZN(n13821) );
  NAND2_X1 U13265 ( .A1(n13805), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U13266 ( .A1(n13821), .A2(n13820), .ZN(n10763) );
  MUX2_X1 U13267 ( .A(n11794), .B(P2_REG2_REG_4__SCAN_IN), .S(n13819), .Z(
        n10762) );
  NAND2_X1 U13268 ( .A1(n10763), .A2(n10762), .ZN(n13824) );
  NAND2_X1 U13269 ( .A1(n13815), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U13270 ( .A1(n13824), .A2(n10764), .ZN(n15327) );
  MUX2_X1 U13271 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11783), .S(n10780), .Z(
        n15326) );
  NAND2_X1 U13272 ( .A1(n15327), .A2(n15326), .ZN(n15325) );
  NAND2_X1 U13273 ( .A1(n10780), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10768) );
  NAND2_X1 U13274 ( .A1(n15325), .A2(n10768), .ZN(n10766) );
  INV_X1 U13275 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11836) );
  MUX2_X1 U13276 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11836), .S(n10811), .Z(
        n10765) );
  NAND2_X1 U13277 ( .A1(n10766), .A2(n10765), .ZN(n13840) );
  MUX2_X1 U13278 ( .A(n11836), .B(P2_REG2_REG_6__SCAN_IN), .S(n10811), .Z(
        n10767) );
  NAND3_X1 U13279 ( .A1(n15325), .A2(n10768), .A3(n10767), .ZN(n10769) );
  AND3_X1 U13280 ( .A1(n15372), .A2(n13840), .A3(n10769), .ZN(n10770) );
  AOI211_X1 U13281 ( .C1(n15371), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n10771), .B(
        n10770), .ZN(n10787) );
  MUX2_X1 U13282 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n8720), .S(n10811), .Z(
        n10785) );
  XNOR2_X1 U13283 ( .A(n10869), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13284 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10866) );
  INV_X1 U13285 ( .A(n10866), .ZN(n10772) );
  NAND2_X1 U13286 ( .A1(n10862), .A2(n10772), .ZN(n10863) );
  NAND2_X1 U13287 ( .A1(n10868), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U13288 ( .A1(n10863), .A2(n10773), .ZN(n15307) );
  INV_X1 U13289 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10774) );
  XNOR2_X1 U13290 ( .A(n10775), .B(n10774), .ZN(n15308) );
  NAND2_X1 U13291 ( .A1(n15307), .A2(n15308), .ZN(n15306) );
  NAND2_X1 U13292 ( .A1(n10775), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13293 ( .A1(n15306), .A2(n10776), .ZN(n13803) );
  INV_X1 U13294 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10777) );
  XNOR2_X1 U13295 ( .A(n13805), .B(n10777), .ZN(n13804) );
  NAND2_X1 U13296 ( .A1(n13803), .A2(n13804), .ZN(n13802) );
  NAND2_X1 U13297 ( .A1(n13805), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U13298 ( .A1(n13802), .A2(n10778), .ZN(n13817) );
  XNOR2_X1 U13299 ( .A(n13819), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n13818) );
  NAND2_X1 U13300 ( .A1(n13817), .A2(n13818), .ZN(n13816) );
  NAND2_X1 U13301 ( .A1(n13815), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10779) );
  NAND2_X1 U13302 ( .A1(n13816), .A2(n10779), .ZN(n15318) );
  INV_X1 U13303 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15480) );
  MUX2_X1 U13304 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n15480), .S(n10780), .Z(
        n15319) );
  NAND2_X1 U13305 ( .A1(n15318), .A2(n15319), .ZN(n15317) );
  NAND2_X1 U13306 ( .A1(n10780), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13307 ( .A1(n15317), .A2(n10781), .ZN(n10784) );
  NAND2_X1 U13308 ( .A1(n10784), .A2(n10785), .ZN(n10806) );
  OAI211_X1 U13309 ( .C1(n10785), .C2(n10784), .A(n15364), .B(n10806), .ZN(
        n10786) );
  OAI211_X1 U13310 ( .C1(n15379), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        P2_U3220) );
  INV_X1 U13311 ( .A(n12141), .ZN(n12149) );
  OAI222_X1 U13312 ( .A1(P1_U3086), .A2(n12149), .B1(n14949), .B2(n10790), 
        .C1(n10789), .C2(n12208), .ZN(P1_U3342) );
  INV_X1 U13313 ( .A(n14408), .ZN(n10932) );
  NOR2_X1 U13314 ( .A1(n10932), .A2(n15097), .ZN(n11054) );
  AOI21_X1 U13315 ( .B1(n14986), .B2(n14411), .A(n11054), .ZN(n10796) );
  XNOR2_X1 U13316 ( .A(n10792), .B(n10791), .ZN(n10793) );
  NAND2_X1 U13317 ( .A1(n10793), .A2(n15081), .ZN(n10795) );
  AOI22_X1 U13318 ( .A1(n15216), .A2(n15088), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10887), .ZN(n10794) );
  OAI211_X1 U13319 ( .C1(n10796), .C2(n15079), .A(n10795), .B(n10794), .ZN(
        P1_U3222) );
  INV_X1 U13320 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10797) );
  NAND2_X1 U13321 ( .A1(n15364), .A2(n10797), .ZN(n10798) );
  OAI211_X1 U13322 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n13867), .A(n10798), .B(
        n15379), .ZN(n10799) );
  INV_X1 U13323 ( .A(n10799), .ZN(n10801) );
  AOI22_X1 U13324 ( .A1(n15372), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n15364), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10800) );
  MUX2_X1 U13325 ( .A(n10801), .B(n10800), .S(n10871), .Z(n10803) );
  AOI22_X1 U13326 ( .A1(n15371), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10802) );
  NAND2_X1 U13327 ( .A1(n10803), .A2(n10802), .ZN(P2_U3214) );
  MUX2_X1 U13328 ( .A(n10804), .B(P2_REG1_REG_10__SCAN_IN), .S(n10854), .Z(
        n10810) );
  NAND2_X1 U13329 ( .A1(n10811), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13330 ( .A1(n10806), .A2(n10805), .ZN(n13834) );
  MUX2_X1 U13331 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8741), .S(n13836), .Z(
        n13835) );
  NAND2_X1 U13332 ( .A1(n13834), .A2(n13835), .ZN(n13833) );
  NAND2_X1 U13333 ( .A1(n13836), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U13334 ( .A1(n13833), .A2(n10807), .ZN(n13848) );
  MUX2_X1 U13335 ( .A(n8760), .B(P2_REG1_REG_8__SCAN_IN), .S(n13850), .Z(
        n13849) );
  NAND2_X1 U13336 ( .A1(n13848), .A2(n13849), .ZN(n13847) );
  NAND2_X1 U13337 ( .A1(n10817), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13338 ( .A1(n13847), .A2(n10808), .ZN(n15336) );
  MUX2_X1 U13339 ( .A(n8778), .B(P2_REG1_REG_9__SCAN_IN), .S(n10820), .Z(
        n15335) );
  OR2_X1 U13340 ( .A1(n15336), .A2(n15335), .ZN(n15338) );
  OAI21_X1 U13341 ( .B1(n10820), .B2(P2_REG1_REG_9__SCAN_IN), .A(n15338), .ZN(
        n10809) );
  NOR2_X1 U13342 ( .A1(n10809), .A2(n10810), .ZN(n10853) );
  AOI211_X1 U13343 ( .C1(n10810), .C2(n10809), .A(n11902), .B(n10853), .ZN(
        n10829) );
  NAND2_X1 U13344 ( .A1(n10811), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13839) );
  NAND2_X1 U13345 ( .A1(n13840), .A2(n13839), .ZN(n10813) );
  MUX2_X1 U13346 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n13837), .S(n13836), .Z(
        n10812) );
  NAND2_X1 U13347 ( .A1(n10813), .A2(n10812), .ZN(n13853) );
  NAND2_X1 U13348 ( .A1(n13836), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U13349 ( .A1(n13853), .A2(n13852), .ZN(n10816) );
  INV_X1 U13350 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10814) );
  MUX2_X1 U13351 ( .A(n10814), .B(P2_REG2_REG_8__SCAN_IN), .S(n13850), .Z(
        n10815) );
  NAND2_X1 U13352 ( .A1(n10816), .A2(n10815), .ZN(n13855) );
  NAND2_X1 U13353 ( .A1(n10817), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13354 ( .A1(n13855), .A2(n10818), .ZN(n15331) );
  INV_X1 U13355 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10819) );
  MUX2_X1 U13356 ( .A(n10819), .B(P2_REG2_REG_9__SCAN_IN), .S(n10820), .Z(
        n15330) );
  OR2_X1 U13357 ( .A1(n15331), .A2(n15330), .ZN(n15333) );
  OAI21_X1 U13358 ( .B1(n10820), .B2(P2_REG2_REG_9__SCAN_IN), .A(n15333), .ZN(
        n10823) );
  INV_X1 U13359 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10821) );
  MUX2_X1 U13360 ( .A(n10821), .B(P2_REG2_REG_10__SCAN_IN), .S(n10854), .Z(
        n10822) );
  NOR2_X1 U13361 ( .A1(n10823), .A2(n10822), .ZN(n10848) );
  AOI211_X1 U13362 ( .C1(n10823), .C2(n10822), .A(n13867), .B(n10848), .ZN(
        n10828) );
  NAND2_X1 U13363 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11271)
         );
  INV_X1 U13364 ( .A(n11271), .ZN(n10824) );
  AOI21_X1 U13365 ( .B1(n15371), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10824), 
        .ZN(n10825) );
  OAI21_X1 U13366 ( .B1(n10826), .B2(n15379), .A(n10825), .ZN(n10827) );
  OR3_X1 U13367 ( .A1(n10829), .A2(n10828), .A3(n10827), .ZN(P2_U3224) );
  OAI222_X1 U13368 ( .A1(P3_U3151), .A2(n13314), .B1(n12971), .B2(n10831), 
        .C1(n12279), .C2(n10830), .ZN(P3_U3276) );
  MUX2_X1 U13369 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10834), .S(n10949), .Z(
        n10835) );
  NAND2_X1 U13370 ( .A1(n10836), .A2(n10835), .ZN(n10948) );
  OAI21_X1 U13371 ( .B1(n10836), .B2(n10835), .A(n10948), .ZN(n10846) );
  NOR2_X1 U13372 ( .A1(n10837), .A2(n8077), .ZN(n10839) );
  MUX2_X1 U13373 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n15119), .S(n10949), .Z(
        n10838) );
  OAI21_X1 U13374 ( .B1(n10840), .B2(n10839), .A(n10838), .ZN(n10942) );
  OR3_X1 U13375 ( .A1(n10840), .A2(n10839), .A3(n10838), .ZN(n10841) );
  NAND3_X1 U13376 ( .A1(n10942), .A2(n14515), .A3(n10841), .ZN(n10844) );
  NOR2_X1 U13377 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15092), .ZN(n10842) );
  AOI21_X1 U13378 ( .B1(n15177), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n10842), 
        .ZN(n10843) );
  OAI211_X1 U13379 ( .C1(n15193), .C2(n10943), .A(n10844), .B(n10843), .ZN(
        n10845) );
  AOI21_X1 U13380 ( .B1(n10846), .B2(n15188), .A(n10845), .ZN(n10847) );
  INV_X1 U13381 ( .A(n10847), .ZN(P1_U3254) );
  AOI21_X1 U13382 ( .B1(n10854), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10848), 
        .ZN(n10850) );
  MUX2_X1 U13383 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11662), .S(n10910), .Z(
        n10849) );
  NAND2_X1 U13384 ( .A1(n10850), .A2(n10849), .ZN(n15349) );
  OAI21_X1 U13385 ( .B1(n10850), .B2(n10849), .A(n15349), .ZN(n10860) );
  NAND2_X1 U13386 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11625)
         );
  INV_X1 U13387 ( .A(n11625), .ZN(n10851) );
  AOI21_X1 U13388 ( .B1(n15371), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10851), 
        .ZN(n10852) );
  OAI21_X1 U13389 ( .B1(n10915), .B2(n15379), .A(n10852), .ZN(n10859) );
  AOI21_X1 U13390 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n10854), .A(n10853), 
        .ZN(n10857) );
  INV_X1 U13391 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10855) );
  MUX2_X1 U13392 ( .A(n10855), .B(P2_REG1_REG_11__SCAN_IN), .S(n10910), .Z(
        n10856) );
  NOR2_X1 U13393 ( .A1(n10857), .A2(n10856), .ZN(n10909) );
  AOI211_X1 U13394 ( .C1(n10857), .C2(n10856), .A(n11902), .B(n10909), .ZN(
        n10858) );
  AOI211_X1 U13395 ( .C1(n15372), .C2(n10860), .A(n10859), .B(n10858), .ZN(
        n10861) );
  INV_X1 U13396 ( .A(n10861), .ZN(P2_U3225) );
  INV_X1 U13397 ( .A(n15379), .ZN(n15358) );
  INV_X1 U13398 ( .A(n10862), .ZN(n10865) );
  INV_X1 U13399 ( .A(n10863), .ZN(n10864) );
  AOI211_X1 U13400 ( .C1(n10866), .C2(n10865), .A(n10864), .B(n11902), .ZN(
        n10867) );
  AOI21_X1 U13401 ( .B1(n15358), .B2(n10868), .A(n10867), .ZN(n10875) );
  MUX2_X1 U13402 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10756), .S(n10869), .Z(
        n10870) );
  OAI21_X1 U13403 ( .B1(n8640), .B2(n10871), .A(n10870), .ZN(n10872) );
  NAND3_X1 U13404 ( .A1(n15372), .A2(n10873), .A3(n10872), .ZN(n10874) );
  OAI211_X1 U13405 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10876), .A(n10875), .B(
        n10874), .ZN(n10879) );
  NOR2_X1 U13406 ( .A1(n10877), .A2(n15363), .ZN(n10878) );
  OR2_X1 U13407 ( .A1(n10879), .A2(n10878), .ZN(P2_U3215) );
  INV_X1 U13408 ( .A(n10880), .ZN(n10928) );
  AOI22_X1 U13409 ( .A1(n12376), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n12510), .ZN(n10881) );
  OAI21_X1 U13410 ( .B1(n10928), .B2(n12208), .A(n10881), .ZN(P1_U3339) );
  XNOR2_X1 U13411 ( .A(n10883), .B(n10882), .ZN(n10884) );
  NAND2_X1 U13412 ( .A1(n10884), .A2(n15081), .ZN(n10889) );
  NAND2_X1 U13413 ( .A1(n14410), .A2(n14986), .ZN(n10886) );
  NAND2_X1 U13414 ( .A1(n14407), .A2(n14987), .ZN(n10885) );
  NAND2_X1 U13415 ( .A1(n10886), .A2(n10885), .ZN(n15205) );
  AOI22_X1 U13416 ( .A1(n15205), .A2(n15105), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10887), .ZN(n10888) );
  OAI211_X1 U13417 ( .C1(n15232), .C2(n14388), .A(n10889), .B(n10888), .ZN(
        P1_U3237) );
  NOR2_X1 U13418 ( .A1(n10890), .A2(P2_U3088), .ZN(n10996) );
  INV_X1 U13419 ( .A(n13770), .ZN(n13734) );
  INV_X1 U13420 ( .A(n12647), .ZN(n12895) );
  NOR3_X1 U13421 ( .A1(n13785), .A2(n8580), .A3(n12895), .ZN(n10892) );
  AOI21_X1 U13422 ( .B1(n13734), .B2(n13800), .A(n10892), .ZN(n10895) );
  AOI21_X1 U13423 ( .B1(n6678), .B2(n10891), .A(n13785), .ZN(n10893) );
  OAI21_X1 U13424 ( .B1(n10893), .B2(n13783), .A(n12648), .ZN(n10894) );
  OAI211_X1 U13425 ( .C1(n10996), .C2(n15383), .A(n10895), .B(n10894), .ZN(
        P2_U3204) );
  INV_X1 U13426 ( .A(n10896), .ZN(n10897) );
  AOI21_X1 U13427 ( .B1(n10899), .B2(n10898), .A(n10897), .ZN(n10903) );
  INV_X1 U13428 ( .A(n10996), .ZN(n10900) );
  INV_X1 U13429 ( .A(n13759), .ZN(n13767) );
  AOI22_X1 U13430 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n10900), .B1(n13767), 
        .B2(n10891), .ZN(n10902) );
  AOI22_X1 U13431 ( .A1(n13734), .A2(n13799), .B1(n12654), .B2(n13783), .ZN(
        n10901) );
  OAI211_X1 U13432 ( .C1(n10903), .C2(n13785), .A(n10902), .B(n10901), .ZN(
        P2_U3194) );
  NAND2_X1 U13433 ( .A1(P3_U3897), .A2(n13114), .ZN(n10904) );
  OAI21_X1 U13434 ( .B1(P3_U3897), .B2(n10905), .A(n10904), .ZN(P3_U3503) );
  INV_X1 U13435 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U13436 ( .A1(n11077), .A2(n10907), .ZN(n10906) );
  OAI21_X1 U13437 ( .B1(n11077), .B2(n10907), .A(n10906), .ZN(n10908) );
  INV_X1 U13438 ( .A(n10908), .ZN(n10914) );
  INV_X1 U13439 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10912) );
  AOI21_X1 U13440 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10910), .A(n10909), 
        .ZN(n15356) );
  NAND2_X1 U13441 ( .A1(n15353), .A2(n10912), .ZN(n10911) );
  OAI211_X1 U13442 ( .C1(n10912), .C2(n15353), .A(n15356), .B(n10911), .ZN(
        n15354) );
  OAI21_X1 U13443 ( .B1(n15359), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15354), 
        .ZN(n10913) );
  NOR2_X1 U13444 ( .A1(n10913), .A2(n10914), .ZN(n11076) );
  AOI211_X1 U13445 ( .C1(n10914), .C2(n10913), .A(n11902), .B(n11076), .ZN(
        n10926) );
  NAND2_X1 U13446 ( .A1(n10915), .A2(n11662), .ZN(n15347) );
  NAND2_X1 U13447 ( .A1(n15359), .A2(n8837), .ZN(n10917) );
  NAND2_X1 U13448 ( .A1(n15353), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10916) );
  AND2_X1 U13449 ( .A1(n10917), .A2(n10916), .ZN(n15348) );
  AOI21_X1 U13450 ( .B1(n15349), .B2(n15347), .A(n15348), .ZN(n15346) );
  AOI21_X1 U13451 ( .B1(n8837), .B2(n15353), .A(n15346), .ZN(n10921) );
  NAND2_X1 U13452 ( .A1(n11077), .A2(n11072), .ZN(n10918) );
  OAI21_X1 U13453 ( .B1(n11077), .B2(n11072), .A(n10918), .ZN(n10920) );
  NAND2_X1 U13454 ( .A1(n11071), .A2(n11072), .ZN(n10919) );
  OAI211_X1 U13455 ( .C1(n11072), .C2(n11071), .A(n10921), .B(n10919), .ZN(
        n11070) );
  OAI211_X1 U13456 ( .C1(n10921), .C2(n10920), .A(n11070), .B(n15372), .ZN(
        n10924) );
  NOR2_X1 U13457 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8852), .ZN(n10922) );
  AOI21_X1 U13458 ( .B1(n15371), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10922), 
        .ZN(n10923) );
  OAI211_X1 U13459 ( .C1(n15379), .C2(n11071), .A(n10924), .B(n10923), .ZN(
        n10925) );
  OR2_X1 U13460 ( .A1(n10926), .A2(n10925), .ZN(P2_U3227) );
  OAI222_X1 U13461 ( .A1(P2_U3088), .A2(n12424), .B1(n14254), .B2(n10928), 
        .C1(n10927), .C2(n14249), .ZN(P2_U3311) );
  INV_X1 U13462 ( .A(n15081), .ZN(n15101) );
  AOI21_X1 U13463 ( .B1(n10930), .B2(n10929), .A(n15101), .ZN(n10931) );
  NAND2_X1 U13464 ( .A1(n10931), .A2(n11027), .ZN(n10937) );
  INV_X1 U13465 ( .A(n14406), .ZN(n10933) );
  OAI22_X1 U13466 ( .A1(n10933), .A2(n15097), .B1(n10932), .B2(n15095), .ZN(
        n11177) );
  INV_X1 U13467 ( .A(n15090), .ZN(n10934) );
  MUX2_X1 U13468 ( .A(n10934), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10935) );
  AOI21_X1 U13469 ( .B1(n11177), .B2(n15105), .A(n10935), .ZN(n10936) );
  OAI211_X1 U13470 ( .C1(n15239), .C2(n14388), .A(n10937), .B(n10936), .ZN(
        P1_U3218) );
  INV_X1 U13471 ( .A(n11426), .ZN(n11075) );
  INV_X1 U13472 ( .A(n10938), .ZN(n10940) );
  INV_X1 U13473 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10939) );
  OAI222_X1 U13474 ( .A1(P2_U3088), .A2(n11075), .B1(n14254), .B2(n10940), 
        .C1(n10939), .C2(n14249), .ZN(P2_U3313) );
  INV_X1 U13475 ( .A(n14475), .ZN(n12150) );
  OAI222_X1 U13476 ( .A1(n14949), .A2(n10941), .B1(n12208), .B2(n10940), .C1(
        n12150), .C2(P1_U3086), .ZN(P1_U3341) );
  OAI21_X1 U13477 ( .B1(n15119), .B2(n10943), .A(n10942), .ZN(n10946) );
  AOI22_X1 U13478 ( .A1(n11093), .A2(n14981), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10944), .ZN(n10945) );
  NOR2_X1 U13479 ( .A1(n10945), .A2(n10946), .ZN(n11094) );
  AOI21_X1 U13480 ( .B1(n10946), .B2(n10945), .A(n11094), .ZN(n10957) );
  MUX2_X1 U13481 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10947), .S(n11093), .Z(
        n10951) );
  OAI21_X1 U13482 ( .B1(n10949), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10948), 
        .ZN(n10950) );
  NAND2_X1 U13483 ( .A1(n10950), .A2(n10951), .ZN(n11089) );
  OAI21_X1 U13484 ( .B1(n10951), .B2(n10950), .A(n11089), .ZN(n10952) );
  NAND2_X1 U13485 ( .A1(n10952), .A2(n15188), .ZN(n10956) );
  OAI22_X1 U13486 ( .A1(n15197), .A2(n9151), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10953), .ZN(n10954) );
  AOI21_X1 U13487 ( .B1(n11093), .B2(n14489), .A(n10954), .ZN(n10955) );
  OAI211_X1 U13488 ( .C1(n10957), .C2(n15183), .A(n10956), .B(n10955), .ZN(
        P1_U3255) );
  INV_X1 U13489 ( .A(n10958), .ZN(n10959) );
  INV_X1 U13490 ( .A(n14494), .ZN(n14491) );
  OAI222_X1 U13491 ( .A1(n14949), .A2(n7016), .B1(n12208), .B2(n10959), .C1(
        n14491), .C2(P1_U3086), .ZN(P1_U3338) );
  OAI222_X1 U13492 ( .A1(n14249), .A2(n10960), .B1(n14254), .B2(n10959), .C1(
        n15378), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13493 ( .A1(n12119), .A2(n15401), .ZN(n15398) );
  INV_X1 U13494 ( .A(n15398), .ZN(n10965) );
  NAND2_X1 U13495 ( .A1(n14213), .A2(n13800), .ZN(n10967) );
  INV_X1 U13496 ( .A(n10891), .ZN(n10968) );
  NAND2_X1 U13497 ( .A1(n10968), .A2(n12648), .ZN(n12896) );
  INV_X1 U13498 ( .A(n12896), .ZN(n11612) );
  NAND2_X1 U13499 ( .A1(n12899), .A2(n11612), .ZN(n11611) );
  NAND2_X1 U13500 ( .A1(n11611), .A2(n10969), .ZN(n10970) );
  OAI21_X1 U13501 ( .B1(n12900), .B2(n10970), .A(n11416), .ZN(n10974) );
  OR2_X1 U13502 ( .A1(n8612), .A2(n13871), .ZN(n10972) );
  NAND2_X1 U13503 ( .A1(n12925), .A2(n10971), .ZN(n12930) );
  OAI22_X1 U13504 ( .A1(n15389), .A2(n14090), .B1(n15388), .B2(n11404), .ZN(
        n10973) );
  AOI21_X1 U13505 ( .B1(n10974), .B2(n14129), .A(n10973), .ZN(n11630) );
  OR2_X1 U13506 ( .A1(n12648), .A2(n12654), .ZN(n11609) );
  NAND2_X1 U13507 ( .A1(n12663), .A2(n11609), .ZN(n10975) );
  NAND2_X1 U13508 ( .A1(n10975), .A2(n8580), .ZN(n10976) );
  NOR2_X1 U13509 ( .A1(n11410), .A2(n10976), .ZN(n11634) );
  AND2_X1 U13510 ( .A1(n12663), .A2(n15450), .ZN(n10977) );
  NOR2_X1 U13511 ( .A1(n11634), .A2(n10977), .ZN(n10982) );
  NAND2_X1 U13512 ( .A1(n7001), .A2(n15389), .ZN(n10978) );
  XNOR2_X1 U13513 ( .A(n11402), .B(n12900), .ZN(n11636) );
  INV_X1 U13514 ( .A(n11636), .ZN(n10980) );
  NAND2_X1 U13515 ( .A1(n8612), .A2(n15385), .ZN(n15470) );
  INV_X1 U13516 ( .A(n15454), .ZN(n15077) );
  NAND2_X1 U13517 ( .A1(n10980), .A2(n15077), .ZN(n10981) );
  AND3_X1 U13518 ( .A1(n11630), .A2(n10982), .A3(n10981), .ZN(n15408) );
  NAND2_X1 U13519 ( .A1(n15487), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10983) );
  OAI21_X1 U13520 ( .B1(n15487), .B2(n15408), .A(n10983), .ZN(P2_U3501) );
  INV_X1 U13521 ( .A(n10984), .ZN(n10985) );
  AOI21_X1 U13522 ( .B1(n10987), .B2(n10986), .A(n10985), .ZN(n10991) );
  NAND2_X1 U13523 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n13825) );
  OAI21_X1 U13524 ( .B1(n13770), .B2(n12692), .A(n13825), .ZN(n10989) );
  OAI22_X1 U13525 ( .A1(n13759), .A2(n11404), .B1(n13781), .B2(n11798), .ZN(
        n10988) );
  AOI211_X1 U13526 ( .C1(n15417), .C2(n13783), .A(n10989), .B(n10988), .ZN(
        n10990) );
  OAI21_X1 U13527 ( .B1(n10991), .B2(n13785), .A(n10990), .ZN(P2_U3202) );
  OAI21_X1 U13528 ( .B1(n10994), .B2(n10993), .A(n10992), .ZN(n10999) );
  OAI22_X1 U13529 ( .A1(n13747), .A2(n6951), .B1(n13770), .B2(n11404), .ZN(
        n10998) );
  OAI22_X1 U13530 ( .A1(n10996), .A2(n10995), .B1(n13759), .B2(n15389), .ZN(
        n10997) );
  AOI211_X1 U13531 ( .C1(n9100), .C2(n10999), .A(n10998), .B(n10997), .ZN(
        n11000) );
  INV_X1 U13532 ( .A(n11000), .ZN(P2_U3209) );
  INV_X1 U13533 ( .A(n15423), .ZN(n11785) );
  AND2_X1 U13534 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15320) );
  OAI22_X1 U13535 ( .A1(n13759), .A2(n12678), .B1(n13781), .B2(n11784), .ZN(
        n11001) );
  AOI211_X1 U13536 ( .C1(n13734), .C2(n13795), .A(n15320), .B(n11001), .ZN(
        n11007) );
  OAI21_X1 U13537 ( .B1(n11004), .B2(n11003), .A(n11002), .ZN(n11005) );
  NAND2_X1 U13538 ( .A1(n11005), .A2(n9100), .ZN(n11006) );
  OAI211_X1 U13539 ( .C1(n11785), .C2(n13747), .A(n11007), .B(n11006), .ZN(
        P2_U3199) );
  XNOR2_X1 U13540 ( .A(n11009), .B(n11008), .ZN(n11014) );
  OAI21_X1 U13541 ( .B1(n13770), .B2(n12706), .A(n11010), .ZN(n11012) );
  OAI22_X1 U13542 ( .A1(n13759), .A2(n12692), .B1(n13781), .B2(n11841), .ZN(
        n11011) );
  AOI211_X1 U13543 ( .C1(n15429), .C2(n13783), .A(n11012), .B(n11011), .ZN(
        n11013) );
  OAI21_X1 U13544 ( .B1(n11014), .B2(n13785), .A(n11013), .ZN(P2_U3211) );
  INV_X1 U13545 ( .A(n12153), .ZN(n15192) );
  INV_X1 U13546 ( .A(n11015), .ZN(n11018) );
  OAI222_X1 U13547 ( .A1(P1_U3086), .A2(n15192), .B1(n12208), .B2(n11018), 
        .C1(n11016), .C2(n14949), .ZN(P1_U3340) );
  INV_X1 U13548 ( .A(n11906), .ZN(n11896) );
  OAI222_X1 U13549 ( .A1(P2_U3088), .A2(n11896), .B1(n14254), .B2(n11018), 
        .C1(n11017), .C2(n14252), .ZN(P2_U3312) );
  XNOR2_X1 U13550 ( .A(n6673), .B(n11019), .ZN(n11025) );
  INV_X1 U13551 ( .A(n13781), .ZN(n13766) );
  INV_X1 U13552 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13809) );
  OAI22_X1 U13553 ( .A1(n13770), .A2(n12678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13809), .ZN(n11023) );
  INV_X1 U13554 ( .A(n15410), .ZN(n11413) );
  OAI22_X1 U13555 ( .A1(n13747), .A2(n11413), .B1(n13759), .B2(n11021), .ZN(
        n11022) );
  AOI211_X1 U13556 ( .C1(n13766), .C2(n13809), .A(n11023), .B(n11022), .ZN(
        n11024) );
  OAI21_X1 U13557 ( .B1(n11025), .B2(n13785), .A(n11024), .ZN(P2_U3190) );
  NAND2_X1 U13558 ( .A1(n11027), .A2(n11026), .ZN(n11031) );
  XNOR2_X1 U13559 ( .A(n11029), .B(n11028), .ZN(n11030) );
  XNOR2_X1 U13560 ( .A(n11031), .B(n11030), .ZN(n11037) );
  NAND2_X1 U13561 ( .A1(n14407), .A2(n14986), .ZN(n11033) );
  NAND2_X1 U13562 ( .A1(n14405), .A2(n14987), .ZN(n11032) );
  NAND2_X1 U13563 ( .A1(n11033), .A2(n11032), .ZN(n15243) );
  NAND2_X1 U13564 ( .A1(n15243), .A2(n15105), .ZN(n11034) );
  NAND2_X1 U13565 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14455) );
  OAI211_X1 U13566 ( .C1(n15090), .C2(n11158), .A(n11034), .B(n14455), .ZN(
        n11035) );
  AOI21_X1 U13567 ( .B1(n15088), .B2(n11203), .A(n11035), .ZN(n11036) );
  OAI21_X1 U13568 ( .B1(n11037), .B2(n15101), .A(n11036), .ZN(P1_U3230) );
  XNOR2_X1 U13569 ( .A(n11039), .B(n11038), .ZN(n11045) );
  NAND2_X1 U13570 ( .A1(n14126), .A2(n13793), .ZN(n11041) );
  NAND2_X1 U13571 ( .A1(n14124), .A2(n13795), .ZN(n11040) );
  AND2_X1 U13572 ( .A1(n11041), .A2(n11040), .ZN(n11819) );
  NAND2_X1 U13573 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13831) );
  OAI21_X1 U13574 ( .B1(n13742), .B2(n11819), .A(n13831), .ZN(n11043) );
  NOR2_X1 U13575 ( .A1(n13781), .A2(n11824), .ZN(n11042) );
  AOI211_X1 U13576 ( .C1(n15434), .C2(n13783), .A(n11043), .B(n11042), .ZN(
        n11044) );
  OAI21_X1 U13577 ( .B1(n11045), .B2(n13785), .A(n11044), .ZN(P2_U3185) );
  INV_X1 U13578 ( .A(n15266), .ZN(n15279) );
  NAND2_X1 U13579 ( .A1(n14411), .A2(n14806), .ZN(n11142) );
  XNOR2_X1 U13580 ( .A(n11143), .B(n11142), .ZN(n15222) );
  OAI21_X1 U13581 ( .B1(n11046), .B2(n11047), .A(n15207), .ZN(n11049) );
  OR2_X1 U13582 ( .A1(n11049), .A2(n14862), .ZN(n15218) );
  OAI21_X1 U13583 ( .B1(n11047), .B2(n15246), .A(n15218), .ZN(n11056) );
  INV_X1 U13584 ( .A(n15274), .ZN(n15271) );
  INV_X1 U13585 ( .A(n14411), .ZN(n11048) );
  OAI21_X1 U13586 ( .B1(n11143), .B2(n11048), .A(n15253), .ZN(n11052) );
  XNOR2_X1 U13587 ( .A(n11049), .B(n14410), .ZN(n11050) );
  AOI21_X1 U13588 ( .B1(n11050), .B2(n15253), .A(n14411), .ZN(n11051) );
  AOI21_X1 U13589 ( .B1(n15095), .B2(n11052), .A(n11051), .ZN(n11053) );
  AOI211_X1 U13590 ( .C1(n15271), .C2(n15222), .A(n11054), .B(n11053), .ZN(
        n15225) );
  INV_X1 U13591 ( .A(n15225), .ZN(n11055) );
  AOI211_X1 U13592 ( .C1(n15279), .C2(n15222), .A(n11056), .B(n11055), .ZN(
        n15230) );
  NAND2_X1 U13593 ( .A1(n15300), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11057) );
  OAI21_X1 U13594 ( .B1(n15230), .B2(n15300), .A(n11057), .ZN(P1_U3529) );
  XOR2_X1 U13595 ( .A(n11059), .B(n11058), .Z(n11060) );
  XNOR2_X1 U13596 ( .A(n11061), .B(n11060), .ZN(n11069) );
  INV_X1 U13597 ( .A(n15093), .ZN(n11067) );
  NOR2_X1 U13598 ( .A1(n11276), .A2(n15246), .ZN(n15255) );
  OR2_X1 U13599 ( .A1(n11279), .A2(n15097), .ZN(n11063) );
  NAND2_X1 U13600 ( .A1(n14406), .A2(n14986), .ZN(n11062) );
  NAND2_X1 U13601 ( .A1(n11063), .A2(n11062), .ZN(n11211) );
  NAND2_X1 U13602 ( .A1(n11211), .A2(n15105), .ZN(n11065) );
  OAI211_X1 U13603 ( .C1(n15090), .C2(n11218), .A(n11065), .B(n11064), .ZN(
        n11066) );
  AOI21_X1 U13604 ( .B1(n11067), .B2(n15255), .A(n11066), .ZN(n11068) );
  OAI21_X1 U13605 ( .B1(n11069), .B2(n15101), .A(n11068), .ZN(P1_U3227) );
  OAI21_X1 U13606 ( .B1(n11072), .B2(n11071), .A(n11070), .ZN(n11425) );
  XNOR2_X1 U13607 ( .A(n11425), .B(n11426), .ZN(n11427) );
  XNOR2_X1 U13608 ( .A(n11427), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11082) );
  NOR2_X1 U13609 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12201), .ZN(n11073) );
  AOI21_X1 U13610 ( .B1(n15371), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n11073), 
        .ZN(n11074) );
  OAI21_X1 U13611 ( .B1(n11075), .B2(n15379), .A(n11074), .ZN(n11081) );
  AOI21_X1 U13612 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11077), .A(n11076), 
        .ZN(n11079) );
  XNOR2_X1 U13613 ( .A(n11426), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11078) );
  NOR2_X1 U13614 ( .A1(n11079), .A2(n11078), .ZN(n11422) );
  AOI211_X1 U13615 ( .C1(n11079), .C2(n11078), .A(n11902), .B(n11422), .ZN(
        n11080) );
  AOI211_X1 U13616 ( .C1(n15372), .C2(n11082), .A(n11081), .B(n11080), .ZN(
        n11083) );
  INV_X1 U13617 ( .A(n11083), .ZN(P2_U3228) );
  INV_X1 U13618 ( .A(n11084), .ZN(n11086) );
  OAI222_X1 U13619 ( .A1(n11483), .A2(P3_U3151), .B1(n12279), .B2(n11086), 
        .C1(n11085), .C2(n12971), .ZN(P3_U3275) );
  INV_X1 U13620 ( .A(n13439), .ZN(n13087) );
  NAND2_X1 U13621 ( .A1(n13087), .A2(P3_U3897), .ZN(n11087) );
  OAI21_X1 U13622 ( .B1(P3_U3897), .B2(n11088), .A(n11087), .ZN(P3_U3512) );
  OAI21_X1 U13623 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n11093), .A(n11089), 
        .ZN(n11092) );
  INV_X1 U13624 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11090) );
  MUX2_X1 U13625 ( .A(n11090), .B(P1_REG1_REG_13__SCAN_IN), .S(n12141), .Z(
        n11091) );
  NOR2_X1 U13626 ( .A1(n11092), .A2(n11091), .ZN(n12140) );
  AOI211_X1 U13627 ( .C1(n11092), .C2(n11091), .A(n12140), .B(n12377), .ZN(
        n11103) );
  OR2_X1 U13628 ( .A1(n11093), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11096) );
  INV_X1 U13629 ( .A(n11094), .ZN(n11095) );
  MUX2_X1 U13630 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n12353), .S(n12141), .Z(
        n11097) );
  NAND2_X1 U13631 ( .A1(n11097), .A2(n11098), .ZN(n12148) );
  OAI211_X1 U13632 ( .C1(n11098), .C2(n11097), .A(n14515), .B(n12148), .ZN(
        n11101) );
  NAND2_X1 U13633 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12395)
         );
  INV_X1 U13634 ( .A(n12395), .ZN(n11099) );
  AOI21_X1 U13635 ( .B1(n15177), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11099), 
        .ZN(n11100) );
  OAI211_X1 U13636 ( .C1(n15193), .C2(n12149), .A(n11101), .B(n11100), .ZN(
        n11102) );
  OR2_X1 U13637 ( .A1(n11103), .A2(n11102), .ZN(P1_U3256) );
  OAI21_X1 U13638 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n11107) );
  NAND2_X1 U13639 ( .A1(n11107), .A2(n9100), .ZN(n11110) );
  AND2_X1 U13640 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n13846) );
  OAI22_X1 U13641 ( .A1(n13759), .A2(n12706), .B1(n13781), .B2(n11812), .ZN(
        n11108) );
  AOI211_X1 U13642 ( .C1(n13734), .C2(n13792), .A(n13846), .B(n11108), .ZN(
        n11109) );
  OAI211_X1 U13643 ( .C1(n7347), .C2(n13747), .A(n11110), .B(n11109), .ZN(
        P2_U3193) );
  XNOR2_X1 U13644 ( .A(n11112), .B(n11111), .ZN(n11119) );
  OR2_X1 U13645 ( .A1(n11518), .A2(n15097), .ZN(n11114) );
  NAND2_X1 U13646 ( .A1(n14405), .A2(n14986), .ZN(n11113) );
  NAND2_X1 U13647 ( .A1(n11114), .A2(n11113), .ZN(n11307) );
  OAI22_X1 U13648 ( .A1(n15090), .A2(n11381), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11115), .ZN(n11117) );
  INV_X1 U13649 ( .A(n11314), .ZN(n11382) );
  NOR2_X1 U13650 ( .A1(n11382), .A2(n14388), .ZN(n11116) );
  AOI211_X1 U13651 ( .C1(n15105), .C2(n11307), .A(n11117), .B(n11116), .ZN(
        n11118) );
  OAI21_X1 U13652 ( .B1(n11119), .B2(n15101), .A(n11118), .ZN(P1_U3239) );
  NAND2_X1 U13653 ( .A1(n13391), .A2(P3_U3897), .ZN(n11120) );
  OAI21_X1 U13654 ( .B1(P3_U3897), .B2(n11121), .A(n11120), .ZN(P3_U3516) );
  NAND2_X1 U13655 ( .A1(n13372), .A2(P3_U3897), .ZN(n11122) );
  OAI21_X1 U13656 ( .B1(P3_U3897), .B2(n11123), .A(n11122), .ZN(P3_U3517) );
  INV_X1 U13657 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U13658 ( .A1(n13390), .A2(P3_U3897), .ZN(n11124) );
  OAI21_X1 U13659 ( .B1(P3_U3897), .B2(n11125), .A(n11124), .ZN(P3_U3514) );
  NAND2_X1 U13660 ( .A1(P3_U3897), .A2(n13097), .ZN(n11126) );
  OAI21_X1 U13661 ( .B1(P3_U3897), .B2(n11127), .A(n11126), .ZN(P3_U3505) );
  INV_X1 U13662 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U13663 ( .A1(P3_U3897), .A2(n12220), .ZN(n11128) );
  OAI21_X1 U13664 ( .B1(P3_U3897), .B2(n11129), .A(n11128), .ZN(P3_U3499) );
  NAND2_X1 U13665 ( .A1(P3_U3897), .A2(n15491), .ZN(n11130) );
  OAI21_X1 U13666 ( .B1(P3_U3897), .B2(n11131), .A(n11130), .ZN(P3_U3492) );
  INV_X1 U13667 ( .A(n11132), .ZN(n11134) );
  INV_X1 U13668 ( .A(n14508), .ZN(n14502) );
  OAI222_X1 U13669 ( .A1(n14949), .A2(n11133), .B1(n12208), .B2(n11134), .C1(
        P1_U3086), .C2(n14502), .ZN(P1_U3337) );
  INV_X1 U13670 ( .A(n12426), .ZN(n12437) );
  OAI222_X1 U13671 ( .A1(n14252), .A2(n11135), .B1(n14254), .B2(n11134), .C1(
        P2_U3088), .C2(n12437), .ZN(P2_U3309) );
  INV_X1 U13672 ( .A(n11136), .ZN(n11137) );
  NAND2_X1 U13673 ( .A1(n11137), .A2(n11318), .ZN(n11138) );
  NAND2_X1 U13674 ( .A1(n11143), .A2(n11142), .ZN(n11145) );
  OR2_X1 U13675 ( .A1(n14410), .A2(n15216), .ZN(n11144) );
  NAND2_X1 U13676 ( .A1(n11145), .A2(n11144), .ZN(n15199) );
  NAND2_X1 U13677 ( .A1(n15199), .A2(n15200), .ZN(n11147) );
  OR2_X1 U13678 ( .A1(n14408), .A2(n15206), .ZN(n11146) );
  NAND2_X1 U13679 ( .A1(n11147), .A2(n11146), .ZN(n11174) );
  NAND2_X1 U13680 ( .A1(n11174), .A2(n11148), .ZN(n11150) );
  OR2_X1 U13681 ( .A1(n14407), .A2(n6976), .ZN(n11149) );
  XNOR2_X1 U13682 ( .A(n11199), .B(n11154), .ZN(n15249) );
  NAND2_X1 U13683 ( .A1(n11176), .A2(n11175), .ZN(n11153) );
  NAND2_X1 U13684 ( .A1(n11153), .A2(n11152), .ZN(n11205) );
  XNOR2_X1 U13685 ( .A(n11205), .B(n11154), .ZN(n15252) );
  NAND2_X1 U13686 ( .A1(n15120), .A2(n15253), .ZN(n14697) );
  INV_X1 U13687 ( .A(n14697), .ZN(n14804) );
  NOR2_X2 U13688 ( .A1(n14590), .A2(n6681), .ZN(n15220) );
  INV_X1 U13689 ( .A(n15220), .ZN(n15124) );
  NAND2_X1 U13690 ( .A1(n15208), .A2(n15239), .ZN(n11180) );
  AOI21_X1 U13691 ( .B1(n11180), .B2(n11203), .A(n14862), .ZN(n11155) );
  OR2_X1 U13692 ( .A1(n11180), .A2(n11203), .ZN(n11217) );
  NAND2_X1 U13693 ( .A1(n11155), .A2(n11217), .ZN(n15245) );
  INV_X1 U13694 ( .A(n11156), .ZN(n11157) );
  NOR2_X1 U13695 ( .A1(n15117), .A2(n11158), .ZN(n11160) );
  MUX2_X1 U13696 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n15243), .S(n15120), .Z(
        n11159) );
  AOI211_X1 U13697 ( .C1(n15215), .C2(n11203), .A(n11160), .B(n11159), .ZN(
        n11161) );
  OAI21_X1 U13698 ( .B1(n15124), .B2(n15245), .A(n11161), .ZN(n11162) );
  AOI21_X1 U13699 ( .B1(n15252), .B2(n14804), .A(n11162), .ZN(n11163) );
  OAI21_X1 U13700 ( .B1(n14802), .B2(n15249), .A(n11163), .ZN(P1_U3289) );
  OAI21_X1 U13701 ( .B1(n11166), .B2(n11165), .A(n11164), .ZN(n11172) );
  INV_X1 U13702 ( .A(n13742), .ZN(n13779) );
  INV_X1 U13703 ( .A(n13791), .ZN(n11658) );
  NAND2_X1 U13704 ( .A1(n14124), .A2(n13793), .ZN(n11167) );
  OAI21_X1 U13705 ( .B1(n11658), .B2(n15388), .A(n11167), .ZN(n11449) );
  NAND2_X1 U13706 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15344) );
  INV_X1 U13707 ( .A(n15344), .ZN(n11168) );
  AOI21_X1 U13708 ( .B1(n13779), .B2(n11449), .A(n11168), .ZN(n11170) );
  NAND2_X1 U13709 ( .A1(n15449), .A2(n13783), .ZN(n11169) );
  OAI211_X1 U13710 ( .C1(n13781), .C2(n11451), .A(n11170), .B(n11169), .ZN(
        n11171) );
  AOI21_X1 U13711 ( .B1(n11172), .B2(n9100), .A(n11171), .ZN(n11173) );
  INV_X1 U13712 ( .A(n11173), .ZN(P2_U3203) );
  XNOR2_X1 U13713 ( .A(n11174), .B(n11175), .ZN(n15240) );
  XNOR2_X1 U13714 ( .A(n11176), .B(n11175), .ZN(n11178) );
  AOI21_X1 U13715 ( .B1(n11178), .B2(n15253), .A(n11177), .ZN(n15238) );
  MUX2_X1 U13716 ( .A(n11179), .B(n15238), .S(n15120), .Z(n11184) );
  OAI211_X1 U13717 ( .C1(n15208), .C2(n15239), .A(n15209), .B(n11180), .ZN(
        n15237) );
  INV_X1 U13718 ( .A(n15237), .ZN(n11182) );
  OAI22_X1 U13719 ( .A1(n14780), .A2(n15239), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15117), .ZN(n11181) );
  AOI21_X1 U13720 ( .B1(n11182), .B2(n15220), .A(n11181), .ZN(n11183) );
  OAI211_X1 U13721 ( .C1(n14802), .C2(n15240), .A(n11184), .B(n11183), .ZN(
        P1_U3290) );
  AOI22_X1 U13722 ( .A1(n13540), .A2(P3_STATE_REG_SCAN_IN), .B1(n11186), .B2(
        n11185), .ZN(n11187) );
  OAI21_X1 U13723 ( .B1(n11188), .B2(n12279), .A(n11187), .ZN(n11189) );
  INV_X1 U13724 ( .A(n11189), .ZN(P3_U3273) );
  XNOR2_X1 U13725 ( .A(n11191), .B(n11190), .ZN(n11198) );
  OR2_X1 U13726 ( .A1(n11279), .A2(n15095), .ZN(n11193) );
  OR2_X1 U13727 ( .A1(n11709), .A2(n15097), .ZN(n11192) );
  NAND2_X1 U13728 ( .A1(n11193), .A2(n11192), .ZN(n15262) );
  NAND2_X1 U13729 ( .A1(n15262), .A2(n15105), .ZN(n11195) );
  OAI211_X1 U13730 ( .C1(n15090), .C2(n11288), .A(n11195), .B(n11194), .ZN(
        n11196) );
  AOI21_X1 U13731 ( .B1(n15088), .B2(n15263), .A(n11196), .ZN(n11197) );
  OAI21_X1 U13732 ( .B1(n11198), .B2(n15101), .A(n11197), .ZN(P1_U3213) );
  NAND2_X1 U13733 ( .A1(n14406), .A2(n11203), .ZN(n11200) );
  OAI21_X1 U13734 ( .B1(n11201), .B2(n11208), .A(n11283), .ZN(n15256) );
  INV_X1 U13735 ( .A(n15256), .ZN(n11222) );
  NOR2_X1 U13736 ( .A1(n6676), .A2(n11202), .ZN(n15221) );
  INV_X1 U13737 ( .A(n15221), .ZN(n11387) );
  NAND2_X1 U13738 ( .A1(n15256), .A2(n15271), .ZN(n11214) );
  INV_X1 U13739 ( .A(n11203), .ZN(n15247) );
  NOR2_X1 U13740 ( .A1(n14406), .A2(n15247), .ZN(n11204) );
  NAND2_X1 U13741 ( .A1(n14406), .A2(n15247), .ZN(n11206) );
  NAND2_X1 U13742 ( .A1(n11209), .A2(n11208), .ZN(n11210) );
  NAND2_X1 U13743 ( .A1(n11278), .A2(n11210), .ZN(n11212) );
  AOI21_X1 U13744 ( .B1(n11212), .B2(n15253), .A(n11211), .ZN(n11213) );
  AND2_X1 U13745 ( .A1(n11214), .A2(n11213), .ZN(n15257) );
  MUX2_X1 U13746 ( .A(n15257), .B(n11215), .S(n6676), .Z(n11221) );
  INV_X1 U13747 ( .A(n11313), .ZN(n11216) );
  AOI211_X1 U13748 ( .C1(n11281), .C2(n11217), .A(n14862), .B(n11216), .ZN(
        n15254) );
  OAI22_X1 U13749 ( .A1(n14780), .A2(n11276), .B1(n15117), .B2(n11218), .ZN(
        n11219) );
  AOI21_X1 U13750 ( .B1(n15254), .B2(n15220), .A(n11219), .ZN(n11220) );
  OAI211_X1 U13751 ( .C1(n11222), .C2(n11387), .A(n11221), .B(n11220), .ZN(
        P1_U3288) );
  INV_X1 U13752 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U13753 ( .A1(P3_U3897), .A2(n15573), .ZN(n11223) );
  OAI21_X1 U13754 ( .B1(P3_U3897), .B2(n11224), .A(n11223), .ZN(P3_U3494) );
  NAND2_X1 U13755 ( .A1(P3_U3897), .A2(n13504), .ZN(n11225) );
  OAI21_X1 U13756 ( .B1(P3_U3897), .B2(n11226), .A(n11225), .ZN(P3_U3508) );
  INV_X1 U13757 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U13758 ( .A1(P3_U3897), .A2(n12169), .ZN(n11227) );
  OAI21_X1 U13759 ( .B1(P3_U3897), .B2(n11228), .A(n11227), .ZN(P3_U3498) );
  NAND2_X1 U13760 ( .A1(P3_U3897), .A2(n15562), .ZN(n11229) );
  OAI21_X1 U13761 ( .B1(P3_U3897), .B2(n11230), .A(n11229), .ZN(P3_U3497) );
  NAND2_X1 U13762 ( .A1(P3_U3897), .A2(n15574), .ZN(n11231) );
  OAI21_X1 U13763 ( .B1(P3_U3897), .B2(n11232), .A(n11231), .ZN(P3_U3496) );
  INV_X1 U13764 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n11234) );
  NAND2_X1 U13765 ( .A1(P3_U3897), .A2(n15563), .ZN(n11233) );
  OAI21_X1 U13766 ( .B1(P3_U3897), .B2(n11234), .A(n11233), .ZN(P3_U3495) );
  INV_X1 U13767 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n11236) );
  NAND2_X1 U13768 ( .A1(P3_U3897), .A2(n13454), .ZN(n11235) );
  OAI21_X1 U13769 ( .B1(P3_U3897), .B2(n11236), .A(n11235), .ZN(P3_U3511) );
  NAND2_X1 U13770 ( .A1(P3_U3897), .A2(n15612), .ZN(n11237) );
  OAI21_X1 U13771 ( .B1(P3_U3897), .B2(n11238), .A(n11237), .ZN(P3_U3493) );
  INV_X1 U13772 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U13773 ( .A1(P3_U3897), .A2(n13423), .ZN(n11239) );
  OAI21_X1 U13774 ( .B1(P3_U3897), .B2(n11240), .A(n11239), .ZN(P3_U3513) );
  NAND2_X1 U13775 ( .A1(P3_U3897), .A2(n12305), .ZN(n11241) );
  OAI21_X1 U13776 ( .B1(P3_U3897), .B2(n11242), .A(n11241), .ZN(P3_U3500) );
  NAND2_X1 U13777 ( .A1(P3_U3897), .A2(n13503), .ZN(n11243) );
  OAI21_X1 U13778 ( .B1(P3_U3897), .B2(n11244), .A(n11243), .ZN(P3_U3506) );
  NAND2_X1 U13779 ( .A1(P3_U3897), .A2(n13472), .ZN(n11245) );
  OAI21_X1 U13780 ( .B1(P3_U3897), .B2(n11246), .A(n11245), .ZN(P3_U3510) );
  NAND2_X1 U13781 ( .A1(P3_U3897), .A2(n12563), .ZN(n11247) );
  OAI21_X1 U13782 ( .B1(P3_U3897), .B2(n11248), .A(n11247), .ZN(P3_U3501) );
  NAND2_X1 U13783 ( .A1(P3_U3897), .A2(n13488), .ZN(n11249) );
  OAI21_X1 U13784 ( .B1(P3_U3897), .B2(n11250), .A(n11249), .ZN(P3_U3507) );
  INV_X1 U13785 ( .A(n13491), .ZN(n11251) );
  NAND2_X1 U13786 ( .A1(P3_U3897), .A2(n11251), .ZN(n11252) );
  OAI21_X1 U13787 ( .B1(P3_U3897), .B2(n11253), .A(n11252), .ZN(P3_U3509) );
  NAND2_X1 U13788 ( .A1(P3_U3897), .A2(n13052), .ZN(n11254) );
  OAI21_X1 U13789 ( .B1(P3_U3897), .B2(n11255), .A(n11254), .ZN(P3_U3504) );
  NAND2_X1 U13790 ( .A1(P3_U3897), .A2(n13111), .ZN(n11256) );
  OAI21_X1 U13791 ( .B1(P3_U3897), .B2(n11257), .A(n11256), .ZN(P3_U3502) );
  NAND2_X1 U13792 ( .A1(n13359), .A2(P3_U3897), .ZN(n11258) );
  OAI21_X1 U13793 ( .B1(P3_U3897), .B2(n11259), .A(n11258), .ZN(P3_U3518) );
  NAND2_X1 U13794 ( .A1(n13371), .A2(P3_U3897), .ZN(n11260) );
  OAI21_X1 U13795 ( .B1(P3_U3897), .B2(n11261), .A(n11260), .ZN(P3_U3515) );
  NAND2_X1 U13796 ( .A1(P3_U3897), .A2(n15614), .ZN(n11262) );
  OAI21_X1 U13797 ( .B1(P3_U3897), .B2(n11263), .A(n11262), .ZN(P3_U3491) );
  INV_X1 U13798 ( .A(n11265), .ZN(n11266) );
  OAI222_X1 U13799 ( .A1(P3_U3151), .A2(n11362), .B1(n12971), .B2(n11267), 
        .C1(n12279), .C2(n11266), .ZN(P3_U3274) );
  XNOR2_X1 U13800 ( .A(n11269), .B(n11268), .ZN(n11275) );
  INV_X1 U13801 ( .A(n13790), .ZN(n12738) );
  NAND2_X1 U13802 ( .A1(n14124), .A2(n13792), .ZN(n11270) );
  OAI21_X1 U13803 ( .B1(n12738), .B2(n15388), .A(n11270), .ZN(n11641) );
  NAND2_X1 U13804 ( .A1(n13779), .A2(n11641), .ZN(n11272) );
  OAI211_X1 U13805 ( .C1(n13781), .C2(n11648), .A(n11272), .B(n11271), .ZN(
        n11273) );
  AOI21_X1 U13806 ( .B1(n12731), .B2(n13783), .A(n11273), .ZN(n11274) );
  OAI21_X1 U13807 ( .B1(n11275), .B2(n13785), .A(n11274), .ZN(P2_U3189) );
  OR2_X1 U13808 ( .A1(n11276), .A2(n14405), .ZN(n11277) );
  NAND2_X1 U13809 ( .A1(n11314), .A2(n11279), .ZN(n11280) );
  NAND2_X1 U13810 ( .A1(n11304), .A2(n11280), .ZN(n11517) );
  XNOR2_X1 U13811 ( .A(n11517), .B(n11285), .ZN(n15261) );
  OR2_X1 U13812 ( .A1(n14405), .A2(n11281), .ZN(n11282) );
  NAND2_X1 U13813 ( .A1(n11283), .A2(n11282), .ZN(n11301) );
  NAND2_X1 U13814 ( .A1(n11301), .A2(n11300), .ZN(n11303) );
  NAND2_X1 U13815 ( .A1(n11279), .A2(n11382), .ZN(n11284) );
  NAND2_X1 U13816 ( .A1(n11303), .A2(n11284), .ZN(n11286) );
  NAND2_X1 U13817 ( .A1(n11286), .A2(n11285), .ZN(n11513) );
  OAI21_X1 U13818 ( .B1(n11286), .B2(n11285), .A(n11513), .ZN(n15270) );
  NOR2_X1 U13819 ( .A1(n11313), .A2(n11314), .ZN(n11312) );
  INV_X1 U13820 ( .A(n15263), .ZN(n11287) );
  NAND2_X1 U13821 ( .A1(n11312), .A2(n11287), .ZN(n11522) );
  OAI211_X1 U13822 ( .C1(n11312), .C2(n11287), .A(n15209), .B(n11522), .ZN(
        n15264) );
  NOR2_X1 U13823 ( .A1(n15117), .A2(n11288), .ZN(n11290) );
  MUX2_X1 U13824 ( .A(n15262), .B(P1_REG2_REG_7__SCAN_IN), .S(n6676), .Z(
        n11289) );
  AOI211_X1 U13825 ( .C1(n15215), .C2(n15263), .A(n11290), .B(n11289), .ZN(
        n11291) );
  OAI21_X1 U13826 ( .B1(n15264), .B2(n15124), .A(n11291), .ZN(n11292) );
  AOI21_X1 U13827 ( .B1(n15270), .B2(n15126), .A(n11292), .ZN(n11293) );
  OAI21_X1 U13828 ( .B1(n15261), .B2(n14697), .A(n11293), .ZN(P1_U3286) );
  INV_X1 U13829 ( .A(n12545), .ZN(n11294) );
  NAND2_X1 U13830 ( .A1(n11294), .A2(P3_U3897), .ZN(n11295) );
  OAI21_X1 U13831 ( .B1(P3_U3897), .B2(n11296), .A(n11295), .ZN(P3_U3521) );
  INV_X1 U13832 ( .A(n13033), .ZN(n13335) );
  NAND2_X1 U13833 ( .A1(n13335), .A2(P3_U3897), .ZN(n11297) );
  OAI21_X1 U13834 ( .B1(P3_U3897), .B2(n11298), .A(n11297), .ZN(P3_U3520) );
  INV_X1 U13835 ( .A(n11299), .ZN(n12966) );
  OAI222_X1 U13836 ( .A1(n14949), .A2(n9576), .B1(n12208), .B2(n12966), .C1(
        P1_U3086), .C2(n6966), .ZN(P1_U3336) );
  OR2_X1 U13837 ( .A1(n11301), .A2(n11300), .ZN(n11302) );
  NAND2_X1 U13838 ( .A1(n11303), .A2(n11302), .ZN(n11309) );
  INV_X1 U13839 ( .A(n11309), .ZN(n11388) );
  OAI21_X1 U13840 ( .B1(n11306), .B2(n11305), .A(n11304), .ZN(n11308) );
  AOI21_X1 U13841 ( .B1(n11308), .B2(n15253), .A(n11307), .ZN(n11311) );
  NAND2_X1 U13842 ( .A1(n11309), .A2(n15271), .ZN(n11310) );
  NAND2_X1 U13843 ( .A1(n11311), .A2(n11310), .ZN(n11379) );
  INV_X1 U13844 ( .A(n11379), .ZN(n11316) );
  AOI211_X1 U13845 ( .C1(n11314), .C2(n11313), .A(n14862), .B(n11312), .ZN(
        n11384) );
  AOI21_X1 U13846 ( .B1(n11314), .B2(n15283), .A(n11384), .ZN(n11315) );
  OAI211_X1 U13847 ( .C1(n11388), .C2(n15266), .A(n11316), .B(n11315), .ZN(
        n11323) );
  NAND2_X1 U13848 ( .A1(n11323), .A2(n15140), .ZN(n11317) );
  OAI21_X1 U13849 ( .B1(n15140), .B2(n10615), .A(n11317), .ZN(P1_U3534) );
  INV_X1 U13850 ( .A(n11318), .ZN(n11320) );
  OR2_X1 U13851 ( .A1(n11320), .A2(n11319), .ZN(n11321) );
  NAND2_X1 U13852 ( .A1(n11323), .A2(n15291), .ZN(n11324) );
  OAI21_X1 U13853 ( .B1(n15291), .B2(n8003), .A(n11324), .ZN(P1_U3477) );
  OAI21_X1 U13854 ( .B1(n13540), .B2(n12621), .A(n13325), .ZN(n11325) );
  NAND2_X1 U13855 ( .A1(n11325), .A2(n11362), .ZN(n11328) );
  NAND2_X1 U13856 ( .A1(n11362), .A2(n11483), .ZN(n11326) );
  NAND2_X1 U13857 ( .A1(n13540), .A2(n11326), .ZN(n11327) );
  NAND2_X1 U13858 ( .A1(n11328), .A2(n11327), .ZN(n12609) );
  INV_X1 U13859 ( .A(n11329), .ZN(n13673) );
  NAND2_X1 U13860 ( .A1(n13673), .A2(n12280), .ZN(n11330) );
  NAND2_X1 U13861 ( .A1(n13673), .A2(n12233), .ZN(n11332) );
  NAND2_X1 U13862 ( .A1(n13659), .A2(n13661), .ZN(n11481) );
  NOR2_X1 U13863 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n11336) );
  NOR4_X1 U13864 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n11335) );
  NOR4_X1 U13865 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n11334) );
  NOR4_X1 U13866 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n11333) );
  NAND4_X1 U13867 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11342) );
  NOR4_X1 U13868 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n11340) );
  NOR4_X1 U13869 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n11339) );
  NOR4_X1 U13870 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n11338) );
  NOR4_X1 U13871 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U13872 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11341) );
  NOR2_X1 U13873 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  INV_X1 U13874 ( .A(n11480), .ZN(n11346) );
  INV_X1 U13875 ( .A(n12610), .ZN(n11345) );
  NAND2_X1 U13876 ( .A1(n12609), .A2(n11345), .ZN(n11349) );
  NAND2_X1 U13877 ( .A1(n11485), .A2(n13325), .ZN(n11499) );
  NOR2_X1 U13878 ( .A1(n11499), .A2(n11361), .ZN(n12611) );
  NAND2_X1 U13879 ( .A1(n12626), .A2(n7033), .ZN(n11479) );
  INV_X1 U13880 ( .A(n12608), .ZN(n11350) );
  NAND2_X1 U13881 ( .A1(n12611), .A2(n11350), .ZN(n11347) );
  NAND2_X1 U13882 ( .A1(n11532), .A2(n12622), .ZN(n12629) );
  AND4_X1 U13883 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n12629), .ZN(
        n11352) );
  NOR2_X1 U13884 ( .A1(n11356), .A2(n12624), .ZN(n12607) );
  NAND2_X1 U13885 ( .A1(n12607), .A2(n11350), .ZN(n11351) );
  NOR2_X1 U13886 ( .A1(n13151), .A2(P3_U3151), .ZN(n15498) );
  NAND2_X1 U13887 ( .A1(n15613), .A2(n12608), .ZN(n11355) );
  NAND2_X1 U13888 ( .A1(n15650), .A2(n15609), .ZN(n11357) );
  NAND2_X1 U13889 ( .A1(n12610), .A2(n15650), .ZN(n11358) );
  OR2_X1 U13890 ( .A1(n11529), .A2(n11358), .ZN(n11359) );
  OAI22_X1 U13891 ( .A1(n13138), .A2(n12041), .B1(n15608), .B2(n13154), .ZN(
        n11360) );
  AOI21_X1 U13892 ( .B1(n13134), .B2(n15614), .A(n11360), .ZN(n11377) );
  XNOR2_X1 U13893 ( .A(n11394), .B(n11364), .ZN(n11363) );
  NAND3_X1 U13894 ( .A1(n15491), .A2(n13030), .A3(n11364), .ZN(n11365) );
  NAND2_X1 U13895 ( .A1(n15614), .A2(n11366), .ZN(n15610) );
  NAND2_X1 U13896 ( .A1(n15610), .A2(n13030), .ZN(n11367) );
  INV_X1 U13897 ( .A(n11369), .ZN(n15616) );
  NAND3_X1 U13898 ( .A1(n15616), .A2(n12598), .A3(n11492), .ZN(n11370) );
  OAI211_X1 U13899 ( .C1(n11371), .C2(n15610), .A(n11396), .B(n11370), .ZN(
        n11375) );
  NAND3_X1 U13900 ( .A1(n12609), .A2(n12610), .A3(n15607), .ZN(n11373) );
  NAND2_X1 U13901 ( .A1(n12611), .A2(n12608), .ZN(n11372) );
  NAND2_X1 U13902 ( .A1(n11373), .A2(n11372), .ZN(n11374) );
  INV_X1 U13903 ( .A(n11529), .ZN(n12614) );
  NAND2_X1 U13904 ( .A1(n11375), .A2(n15494), .ZN(n11376) );
  OAI211_X1 U13905 ( .C1(n15498), .C2(n11378), .A(n11377), .B(n11376), .ZN(
        P3_U3162) );
  MUX2_X1 U13906 ( .A(n11379), .B(P1_REG2_REG_6__SCAN_IN), .S(n6676), .Z(
        n11380) );
  INV_X1 U13907 ( .A(n11380), .ZN(n11386) );
  OAI22_X1 U13908 ( .A1(n11382), .A2(n14780), .B1(n11381), .B2(n15117), .ZN(
        n11383) );
  AOI21_X1 U13909 ( .B1(n11384), .B2(n15220), .A(n11383), .ZN(n11385) );
  OAI211_X1 U13910 ( .C1(n11388), .C2(n11387), .A(n11386), .B(n11385), .ZN(
        P1_U3287) );
  INV_X1 U13911 ( .A(n12996), .ZN(n13345) );
  NAND2_X1 U13912 ( .A1(n13345), .A2(P3_U3897), .ZN(n11390) );
  OAI21_X1 U13913 ( .B1(P3_U3897), .B2(n11391), .A(n11390), .ZN(P3_U3519) );
  OAI22_X1 U13914 ( .A1(n13138), .A2(n15596), .B1(n13154), .B2(n15588), .ZN(
        n11392) );
  AOI21_X1 U13915 ( .B1(n13134), .B2(n15491), .A(n11392), .ZN(n11401) );
  XNOR2_X1 U13916 ( .A(n12042), .B(n15612), .ZN(n11398) );
  OAI21_X1 U13917 ( .B1(n11398), .B2(n11397), .A(n12044), .ZN(n11399) );
  NAND2_X1 U13918 ( .A1(n11399), .A2(n15494), .ZN(n11400) );
  OAI211_X1 U13919 ( .C1(n15498), .C2(n15590), .A(n11401), .B(n11400), .ZN(
        P3_U3177) );
  OR2_X1 U13920 ( .A1(n12663), .A2(n13799), .ZN(n11403) );
  OR2_X1 U13921 ( .A1(n15410), .A2(n11404), .ZN(n11405) );
  XNOR2_X1 U13922 ( .A(n11455), .B(n12901), .ZN(n15413) );
  INV_X1 U13923 ( .A(n15400), .ZN(n11407) );
  INV_X1 U13924 ( .A(n12119), .ZN(n11406) );
  NAND3_X1 U13925 ( .A1(n11407), .A2(n12121), .A3(n11406), .ZN(n11408) );
  NAND2_X1 U13926 ( .A1(n8613), .A2(n12926), .ZN(n11776) );
  NAND2_X1 U13927 ( .A1(n15471), .A2(n11776), .ZN(n11409) );
  INV_X1 U13928 ( .A(n11410), .ZN(n11411) );
  AOI211_X1 U13929 ( .C1(n15410), .C2(n11411), .A(n6678), .B(n7346), .ZN(
        n15409) );
  OAI22_X1 U13930 ( .A1(n14102), .A2(n11413), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15384), .ZN(n11414) );
  AOI21_X1 U13931 ( .B1(n14108), .B2(n15409), .A(n11414), .ZN(n11421) );
  INV_X2 U13932 ( .A(n14095), .ZN(n14129) );
  OAI21_X1 U13933 ( .B1(n12901), .B2(n11417), .A(n11438), .ZN(n11418) );
  AOI222_X1 U13934 ( .A1(n14129), .A2(n11418), .B1(n13797), .B2(n14126), .C1(
        n13799), .C2(n14124), .ZN(n15412) );
  MUX2_X1 U13935 ( .A(n11419), .B(n15412), .S(n15392), .Z(n11420) );
  OAI211_X1 U13936 ( .C1(n15413), .C2(n14133), .A(n11421), .B(n11420), .ZN(
        P2_U3262) );
  AOI21_X1 U13937 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n11426), .A(n11422), 
        .ZN(n11897) );
  XNOR2_X1 U13938 ( .A(n11897), .B(n11896), .ZN(n11424) );
  INV_X1 U13939 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11423) );
  NOR2_X1 U13940 ( .A1(n11423), .A2(n11424), .ZN(n11898) );
  AOI211_X1 U13941 ( .C1(n11424), .C2(n11423), .A(n11898), .B(n11902), .ZN(
        n11436) );
  NAND2_X1 U13942 ( .A1(n11426), .A2(n11425), .ZN(n11430) );
  INV_X1 U13943 ( .A(n11427), .ZN(n11428) );
  NAND2_X1 U13944 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n11428), .ZN(n11429) );
  NAND2_X1 U13945 ( .A1(n11430), .A2(n11429), .ZN(n11905) );
  XNOR2_X1 U13946 ( .A(n11896), .B(n11905), .ZN(n11431) );
  NAND2_X1 U13947 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11431), .ZN(n11907) );
  OAI211_X1 U13948 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n11431), .A(n15372), 
        .B(n11907), .ZN(n11434) );
  NOR2_X1 U13949 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8883), .ZN(n11432) );
  AOI21_X1 U13950 ( .B1(n15371), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n11432), 
        .ZN(n11433) );
  OAI211_X1 U13951 ( .C1(n15379), .C2(n11896), .A(n11434), .B(n11433), .ZN(
        n11435) );
  OR2_X1 U13952 ( .A1(n11436), .A2(n11435), .ZN(P2_U3229) );
  INV_X2 U13953 ( .A(n15392), .ZN(n15394) );
  NAND2_X1 U13954 ( .A1(n15417), .A2(n12678), .ZN(n11440) );
  OR2_X1 U13955 ( .A1(n15417), .A2(n12678), .ZN(n11439) );
  NAND2_X1 U13956 ( .A1(n11440), .A2(n11439), .ZN(n12903) );
  INV_X1 U13957 ( .A(n12903), .ZN(n11792) );
  NAND2_X1 U13958 ( .A1(n15423), .A2(n12692), .ZN(n11442) );
  OR2_X1 U13959 ( .A1(n15423), .A2(n12692), .ZN(n11441) );
  AND2_X1 U13960 ( .A1(n11442), .A2(n11441), .ZN(n12906) );
  XNOR2_X1 U13961 ( .A(n15429), .B(n13795), .ZN(n12904) );
  NAND2_X1 U13962 ( .A1(n15429), .A2(n11779), .ZN(n11443) );
  OR2_X1 U13963 ( .A1(n15434), .A2(n12706), .ZN(n11444) );
  NAND2_X1 U13964 ( .A1(n15434), .A2(n12706), .ZN(n11445) );
  INV_X1 U13965 ( .A(n13793), .ZN(n11446) );
  XNOR2_X1 U13966 ( .A(n12717), .B(n11446), .ZN(n12909) );
  INV_X1 U13967 ( .A(n12909), .ZN(n11804) );
  NAND2_X1 U13968 ( .A1(n11805), .A2(n11804), .ZN(n11448) );
  NAND2_X1 U13969 ( .A1(n12717), .A2(n11446), .ZN(n11447) );
  NAND2_X1 U13970 ( .A1(n11448), .A2(n11447), .ZN(n11638) );
  INV_X1 U13971 ( .A(n13792), .ZN(n12726) );
  XNOR2_X1 U13972 ( .A(n15449), .B(n12726), .ZN(n12910) );
  INV_X1 U13973 ( .A(n12910), .ZN(n11637) );
  XNOR2_X1 U13974 ( .A(n11638), .B(n11637), .ZN(n11450) );
  AOI21_X1 U13975 ( .B1(n11450), .B2(n14129), .A(n11449), .ZN(n15451) );
  INV_X1 U13976 ( .A(n15429), .ZN(n11842) );
  NAND2_X1 U13977 ( .A1(n11842), .A2(n11837), .ZN(n11838) );
  AOI211_X1 U13978 ( .C1(n15449), .C2(n11810), .A(n6678), .B(n11647), .ZN(
        n15448) );
  INV_X1 U13979 ( .A(n15449), .ZN(n11454) );
  INV_X1 U13980 ( .A(n11451), .ZN(n11452) );
  INV_X1 U13981 ( .A(n15384), .ZN(n14117) );
  AOI22_X1 U13982 ( .A1(n15394), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11452), 
        .B2(n14117), .ZN(n11453) );
  OAI21_X1 U13983 ( .B1(n11454), .B2(n14102), .A(n11453), .ZN(n11469) );
  NAND2_X1 U13984 ( .A1(n11455), .A2(n7489), .ZN(n11457) );
  OR2_X1 U13985 ( .A1(n15410), .A2(n13798), .ZN(n11456) );
  OR2_X1 U13986 ( .A1(n15417), .A2(n13797), .ZN(n11458) );
  NOR2_X1 U13987 ( .A1(n15423), .A2(n13796), .ZN(n11459) );
  NAND2_X1 U13988 ( .A1(n15423), .A2(n13796), .ZN(n11460) );
  INV_X1 U13989 ( .A(n12904), .ZN(n11829) );
  NAND2_X1 U13990 ( .A1(n11830), .A2(n11829), .ZN(n11462) );
  NAND2_X1 U13991 ( .A1(n15429), .A2(n13795), .ZN(n11461) );
  NAND2_X1 U13992 ( .A1(n11462), .A2(n11461), .ZN(n11817) );
  AND2_X1 U13993 ( .A1(n15434), .A2(n13794), .ZN(n11463) );
  OR2_X1 U13994 ( .A1(n15434), .A2(n13794), .ZN(n11464) );
  NAND2_X1 U13995 ( .A1(n12717), .A2(n13793), .ZN(n11466) );
  OAI21_X1 U13996 ( .B1(n11467), .B2(n12910), .A(n11644), .ZN(n15453) );
  NOR2_X1 U13997 ( .A1(n15453), .A2(n14133), .ZN(n11468) );
  AOI211_X1 U13998 ( .C1(n14108), .C2(n15448), .A(n11469), .B(n11468), .ZN(
        n11470) );
  OAI21_X1 U13999 ( .B1(n15394), .B2(n15451), .A(n11470), .ZN(P2_U3256) );
  XOR2_X1 U14000 ( .A(n11471), .B(n11472), .Z(n11477) );
  OAI22_X1 U14001 ( .A1(n12020), .A2(n15097), .B1(n11518), .B2(n15095), .ZN(
        n11520) );
  NAND2_X1 U14002 ( .A1(n11520), .A2(n15105), .ZN(n11474) );
  OAI211_X1 U14003 ( .C1(n15090), .C2(n11523), .A(n11474), .B(n11473), .ZN(
        n11475) );
  AOI21_X1 U14004 ( .B1(n15088), .B2(n11705), .A(n11475), .ZN(n11476) );
  OAI21_X1 U14005 ( .B1(n11477), .B2(n15101), .A(n11476), .ZN(P1_U3221) );
  XNOR2_X1 U14006 ( .A(n11478), .B(n11502), .ZN(n15639) );
  INV_X1 U14007 ( .A(n15639), .ZN(n11508) );
  NAND3_X1 U14008 ( .A1(n11481), .A2(n11480), .A3(n11479), .ZN(n11482) );
  NOR2_X1 U14009 ( .A1(n11483), .A2(n13325), .ZN(n11484) );
  NAND2_X1 U14010 ( .A1(n11485), .A2(n11484), .ZN(n11490) );
  NAND2_X1 U14011 ( .A1(n12624), .A2(n11490), .ZN(n12628) );
  XNOR2_X1 U14012 ( .A(n12628), .B(n12626), .ZN(n11486) );
  NAND3_X1 U14013 ( .A1(n12633), .A2(n12629), .A3(n11486), .ZN(n11505) );
  AND2_X1 U14014 ( .A1(n11487), .A2(n15609), .ZN(n15605) );
  NAND2_X1 U14015 ( .A1(n15625), .A2(n15605), .ZN(n13351) );
  INV_X1 U14016 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11546) );
  AND2_X1 U14017 ( .A1(n15607), .A2(n11488), .ZN(n11489) );
  NAND2_X1 U14018 ( .A1(n12609), .A2(n11489), .ZN(n11491) );
  OAI22_X1 U14019 ( .A1(n15597), .A2(n12094), .B1(n12041), .B2(n15594), .ZN(
        n11504) );
  NAND2_X1 U14020 ( .A1(n11492), .A2(n15610), .ZN(n11494) );
  NAND2_X1 U14021 ( .A1(n15595), .A2(n15608), .ZN(n11493) );
  NAND2_X1 U14022 ( .A1(n11494), .A2(n11493), .ZN(n15592) );
  NAND2_X1 U14023 ( .A1(n15592), .A2(n15593), .ZN(n11497) );
  NAND2_X1 U14024 ( .A1(n12041), .A2(n15588), .ZN(n11496) );
  INV_X1 U14025 ( .A(n11721), .ZN(n11500) );
  AOI211_X1 U14026 ( .C1(n11502), .C2(n11501), .A(n15619), .B(n11500), .ZN(
        n11503) );
  AOI211_X1 U14027 ( .C1(n15639), .C2(n15656), .A(n11504), .B(n11503), .ZN(
        n15636) );
  MUX2_X1 U14028 ( .A(n11546), .B(n15636), .S(n15625), .Z(n11507) );
  OR2_X1 U14029 ( .A1(n11505), .A2(n15609), .ZN(n12488) );
  INV_X1 U14030 ( .A(n12488), .ZN(n15583) );
  AND2_X1 U14031 ( .A1(n15650), .A2(n12045), .ZN(n15638) );
  AOI22_X1 U14032 ( .A1(n15583), .A2(n15638), .B1(n15622), .B2(n11558), .ZN(
        n11506) );
  OAI211_X1 U14033 ( .C1(n11508), .C2(n13351), .A(n11507), .B(n11506), .ZN(
        P3_U3230) );
  NAND2_X1 U14034 ( .A1(n11509), .A2(n13662), .ZN(n11510) );
  OAI211_X1 U14035 ( .C1(n11511), .C2(n12971), .A(n11510), .B(n11528), .ZN(
        P3_U3272) );
  OAI21_X1 U14036 ( .B1(n11514), .B2(n11704), .A(n11698), .ZN(n11515) );
  INV_X1 U14037 ( .A(n11515), .ZN(n11671) );
  OR2_X1 U14038 ( .A1(n15263), .A2(n11518), .ZN(n11516) );
  NAND2_X1 U14039 ( .A1(n15263), .A2(n11518), .ZN(n11519) );
  XOR2_X1 U14040 ( .A(n11703), .B(n11704), .Z(n11521) );
  AOI21_X1 U14041 ( .B1(n11521), .B2(n15253), .A(n11520), .ZN(n11670) );
  MUX2_X1 U14042 ( .A(n11670), .B(n10674), .S(n6676), .Z(n11527) );
  AOI211_X1 U14043 ( .C1(n11705), .C2(n11522), .A(n14862), .B(n7260), .ZN(
        n11668) );
  INV_X1 U14044 ( .A(n11705), .ZN(n11524) );
  OAI22_X1 U14045 ( .A1(n11524), .A2(n14780), .B1(n11523), .B2(n15117), .ZN(
        n11525) );
  AOI21_X1 U14046 ( .B1(n11668), .B2(n15220), .A(n11525), .ZN(n11526) );
  OAI211_X1 U14047 ( .C1(n11671), .C2(n14802), .A(n11527), .B(n11526), .ZN(
        P1_U3285) );
  NAND2_X1 U14048 ( .A1(n11529), .A2(n11528), .ZN(n11556) );
  AOI21_X1 U14049 ( .B1(n11532), .B2(n11531), .A(n11530), .ZN(n11555) );
  MUX2_X1 U14050 ( .A(P3_U3897), .B(n11568), .S(n12561), .Z(n15503) );
  INV_X1 U14051 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11535) );
  INV_X2 U14052 ( .A(n6997), .ZN(n13268) );
  MUX2_X1 U14053 ( .A(n11535), .B(n11534), .S(n13268), .Z(n11536) );
  INV_X1 U14054 ( .A(n11569), .ZN(n13156) );
  NAND2_X1 U14055 ( .A1(n11536), .A2(n13156), .ZN(n11732) );
  INV_X1 U14056 ( .A(n11536), .ZN(n11537) );
  NAND2_X1 U14057 ( .A1(n11537), .A2(n11569), .ZN(n11538) );
  NAND2_X1 U14058 ( .A1(n11732), .A2(n11538), .ZN(n13157) );
  INV_X1 U14059 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11540) );
  INV_X1 U14060 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11539) );
  MUX2_X1 U14061 ( .A(n11540), .B(n11539), .S(n13268), .Z(n15502) );
  NAND2_X1 U14062 ( .A1(n15502), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15511) );
  OR2_X1 U14063 ( .A1(n13157), .A2(n15511), .ZN(n13159) );
  NAND2_X1 U14064 ( .A1(n13159), .A2(n11732), .ZN(n11544) );
  INV_X1 U14065 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11562) );
  INV_X1 U14066 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11574) );
  MUX2_X1 U14067 ( .A(n11562), .B(n11574), .S(n13268), .Z(n11541) );
  NAND2_X1 U14068 ( .A1(n11541), .A2(n11575), .ZN(n11553) );
  INV_X1 U14069 ( .A(n11541), .ZN(n11542) );
  NAND2_X1 U14070 ( .A1(n11542), .A2(n7564), .ZN(n11543) );
  AND2_X1 U14071 ( .A1(n11553), .A2(n11543), .ZN(n11731) );
  NAND2_X1 U14072 ( .A1(n11544), .A2(n11731), .ZN(n11735) );
  NAND2_X1 U14073 ( .A1(n11735), .A2(n11553), .ZN(n11550) );
  MUX2_X1 U14074 ( .A(n11546), .B(n11545), .S(n13268), .Z(n11547) );
  NAND2_X1 U14075 ( .A1(n11547), .A2(n11588), .ZN(n11690) );
  INV_X1 U14076 ( .A(n11547), .ZN(n11548) );
  NAND2_X1 U14077 ( .A1(n11548), .A2(n11577), .ZN(n11549) );
  AND2_X1 U14078 ( .A1(n11690), .A2(n11549), .ZN(n11551) );
  INV_X1 U14079 ( .A(n11551), .ZN(n11552) );
  NAND3_X1 U14080 ( .A1(n11735), .A2(n11553), .A3(n11552), .ZN(n11554) );
  AOI21_X1 U14081 ( .B1(n11691), .B2(n11554), .A(n15520), .ZN(n11587) );
  INV_X1 U14082 ( .A(n11555), .ZN(n11557) );
  NOR2_X1 U14083 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11558), .ZN(n12113) );
  AOI21_X1 U14084 ( .B1(n15538), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n12113), .ZN(
        n11585) );
  INV_X1 U14085 ( .A(n11559), .ZN(n11560) );
  NOR2_X1 U14086 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11540), .ZN(n15501) );
  NAND2_X1 U14087 ( .A1(n9633), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14088 ( .A1(n11740), .A2(n11739), .ZN(n11738) );
  OR2_X1 U14089 ( .A1(n11575), .A2(n11562), .ZN(n11563) );
  NAND2_X1 U14090 ( .A1(n11738), .A2(n11563), .ZN(n11564) );
  NAND2_X1 U14091 ( .A1(n11564), .A2(n11577), .ZN(n11675) );
  OAI21_X1 U14092 ( .B1(n11566), .B2(P3_REG2_REG_3__SCAN_IN), .A(n11677), .ZN(
        n11567) );
  NAND2_X1 U14093 ( .A1(n15539), .A2(n11567), .ZN(n11584) );
  NAND2_X1 U14094 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n6887), .ZN(n11572) );
  NAND2_X1 U14095 ( .A1(n11569), .A2(n11572), .ZN(n11571) );
  INV_X1 U14096 ( .A(n11572), .ZN(n15499) );
  NAND2_X1 U14097 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n15499), .ZN(n11570) );
  NAND2_X1 U14098 ( .A1(n11571), .A2(n11570), .ZN(n13167) );
  NAND2_X1 U14099 ( .A1(n13167), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n13166) );
  OR2_X1 U14100 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11572), .ZN(n11573) );
  NAND2_X1 U14101 ( .A1(n13166), .A2(n11573), .ZN(n11742) );
  NAND2_X1 U14102 ( .A1(n11743), .A2(n11742), .ZN(n11741) );
  OR2_X1 U14103 ( .A1(n11575), .A2(n11574), .ZN(n11576) );
  NAND2_X1 U14104 ( .A1(n11741), .A2(n11576), .ZN(n11578) );
  OR2_X1 U14105 ( .A1(n11578), .A2(n11577), .ZN(n11579) );
  NAND2_X1 U14106 ( .A1(n11580), .A2(n11545), .ZN(n11581) );
  NAND2_X1 U14107 ( .A1(n11682), .A2(n11581), .ZN(n11582) );
  NAND2_X1 U14108 ( .A1(n15500), .A2(n11582), .ZN(n11583) );
  NAND3_X1 U14109 ( .A1(n11585), .A2(n11584), .A3(n11583), .ZN(n11586) );
  AOI211_X1 U14110 ( .C1(n15503), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        n11589) );
  INV_X1 U14111 ( .A(n11589), .ZN(P3_U3185) );
  INV_X1 U14112 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15585) );
  MUX2_X1 U14113 ( .A(n15585), .B(n9671), .S(n13268), .Z(n11590) );
  XNOR2_X1 U14114 ( .A(n11590), .B(n11596), .ZN(n11689) );
  MUX2_X1 U14115 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13268), .Z(n11591) );
  OR2_X1 U14116 ( .A1(n11591), .A2(n11598), .ZN(n11752) );
  INV_X1 U14117 ( .A(n11752), .ZN(n11592) );
  AND2_X1 U14118 ( .A1(n11591), .A2(n11598), .ZN(n11753) );
  NOR2_X1 U14119 ( .A1(n11592), .A2(n11753), .ZN(n11593) );
  XNOR2_X1 U14120 ( .A(n6835), .B(n11593), .ZN(n11608) );
  XNOR2_X1 U14121 ( .A(n11596), .B(n15585), .ZN(n11676) );
  INV_X1 U14122 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15570) );
  AOI21_X1 U14123 ( .B1(n11595), .B2(n15570), .A(n11759), .ZN(n11604) );
  NOR2_X1 U14124 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9688), .ZN(n12092) );
  NAND2_X1 U14125 ( .A1(n11696), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14126 ( .A1(n11684), .A2(n11597), .ZN(n11599) );
  AOI21_X1 U14127 ( .B1(n11600), .B2(n9691), .A(n11764), .ZN(n11601) );
  NOR2_X1 U14128 ( .A1(n15547), .A2(n11601), .ZN(n11602) );
  AOI211_X1 U14129 ( .C1(n15538), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n12092), .B(
        n11602), .ZN(n11603) );
  OAI21_X1 U14130 ( .B1(n11604), .B2(n15515), .A(n11603), .ZN(n11605) );
  AOI21_X1 U14131 ( .B1(n11606), .B2(n15503), .A(n11605), .ZN(n11607) );
  OAI21_X1 U14132 ( .B1(n15520), .B2(n11608), .A(n11607), .ZN(P3_U3187) );
  INV_X1 U14133 ( .A(n14108), .ZN(n13886) );
  OAI211_X1 U14134 ( .C1(n7001), .C2(n15381), .A(n8580), .B(n11609), .ZN(
        n14212) );
  OAI22_X1 U14135 ( .A1(n13886), .A2(n14212), .B1(n7001), .B2(n14102), .ZN(
        n11619) );
  INV_X1 U14136 ( .A(n14133), .ZN(n12324) );
  XNOR2_X1 U14137 ( .A(n12899), .B(n11610), .ZN(n14211) );
  NAND2_X1 U14138 ( .A1(n12324), .A2(n14211), .ZN(n11617) );
  OAI21_X1 U14139 ( .B1(n12899), .B2(n11612), .A(n11611), .ZN(n11613) );
  NAND2_X1 U14140 ( .A1(n11613), .A2(n14129), .ZN(n11615) );
  AOI22_X1 U14141 ( .A1(n14124), .A2(n10891), .B1(n14126), .B2(n13799), .ZN(
        n11614) );
  NAND2_X1 U14142 ( .A1(n11615), .A2(n11614), .ZN(n14215) );
  AOI22_X1 U14143 ( .A1(n15392), .A2(n14215), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14117), .ZN(n11616) );
  OAI211_X1 U14144 ( .C1(n10756), .C2(n15392), .A(n11617), .B(n11616), .ZN(
        n11618) );
  OR2_X1 U14145 ( .A1(n11619), .A2(n11618), .ZN(P2_U3264) );
  INV_X1 U14146 ( .A(n11620), .ZN(n11621) );
  AOI21_X1 U14147 ( .B1(n11623), .B2(n11622), .A(n11621), .ZN(n11629) );
  INV_X1 U14148 ( .A(n13789), .ZN(n12127) );
  NAND2_X1 U14149 ( .A1(n14124), .A2(n13791), .ZN(n11624) );
  OAI21_X1 U14150 ( .B1(n12127), .B2(n15388), .A(n11624), .ZN(n11655) );
  NAND2_X1 U14151 ( .A1(n13779), .A2(n11655), .ZN(n11626) );
  OAI211_X1 U14152 ( .C1(n13781), .C2(n11661), .A(n11626), .B(n11625), .ZN(
        n11627) );
  AOI21_X1 U14153 ( .B1(n12736), .B2(n13783), .A(n11627), .ZN(n11628) );
  OAI21_X1 U14154 ( .B1(n11629), .B2(n13785), .A(n11628), .ZN(P2_U3208) );
  NOR2_X1 U14155 ( .A1(n15394), .A2(n11630), .ZN(n11633) );
  AOI22_X1 U14156 ( .A1(n15394), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14117), .ZN(n11631) );
  OAI21_X1 U14157 ( .B1(n6951), .B2(n14102), .A(n11631), .ZN(n11632) );
  AOI211_X1 U14158 ( .C1(n11634), .C2(n14108), .A(n11633), .B(n11632), .ZN(
        n11635) );
  OAI21_X1 U14159 ( .B1(n11636), .B2(n14133), .A(n11635), .ZN(P2_U3263) );
  NAND2_X1 U14160 ( .A1(n11638), .A2(n11637), .ZN(n11640) );
  NAND2_X1 U14161 ( .A1(n15449), .A2(n12726), .ZN(n11639) );
  XNOR2_X1 U14162 ( .A(n12731), .B(n11658), .ZN(n12911) );
  INV_X1 U14163 ( .A(n12911), .ZN(n11653) );
  XNOR2_X1 U14164 ( .A(n11654), .B(n11653), .ZN(n11642) );
  AOI21_X1 U14165 ( .B1(n11642), .B2(n14129), .A(n11641), .ZN(n15463) );
  NAND2_X1 U14166 ( .A1(n15449), .A2(n13792), .ZN(n11643) );
  NAND2_X1 U14167 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  OR2_X1 U14168 ( .A1(n11645), .A2(n12911), .ZN(n11646) );
  NAND2_X1 U14169 ( .A1(n11645), .A2(n12911), .ZN(n11657) );
  AND2_X1 U14170 ( .A1(n11657), .A2(n11646), .ZN(n15461) );
  INV_X1 U14171 ( .A(n12731), .ZN(n15457) );
  OAI211_X1 U14172 ( .C1(n15457), .C2(n11647), .A(n8580), .B(n11659), .ZN(
        n15456) );
  INV_X1 U14173 ( .A(n14102), .ZN(n14038) );
  OAI22_X1 U14174 ( .A1(n15392), .A2(n10821), .B1(n11648), .B2(n15384), .ZN(
        n11649) );
  AOI21_X1 U14175 ( .B1(n12731), .B2(n14038), .A(n11649), .ZN(n11650) );
  OAI21_X1 U14176 ( .B1(n15456), .B2(n13886), .A(n11650), .ZN(n11651) );
  AOI21_X1 U14177 ( .B1(n15461), .B2(n12324), .A(n11651), .ZN(n11652) );
  OAI21_X1 U14178 ( .B1(n15463), .B2(n15394), .A(n11652), .ZN(P2_U3255) );
  XNOR2_X1 U14179 ( .A(n12736), .B(n12738), .ZN(n12913) );
  XNOR2_X1 U14180 ( .A(n11887), .B(n12913), .ZN(n11656) );
  AOI21_X1 U14181 ( .B1(n11656), .B2(n14129), .A(n11655), .ZN(n15466) );
  XNOR2_X1 U14182 ( .A(n11889), .B(n12913), .ZN(n15469) );
  INV_X1 U14183 ( .A(n15469), .ZN(n11666) );
  INV_X1 U14184 ( .A(n11659), .ZN(n11660) );
  INV_X1 U14185 ( .A(n12736), .ZN(n15468) );
  OR2_X2 U14186 ( .A1(n11659), .A2(n12736), .ZN(n11890) );
  OAI211_X1 U14187 ( .C1(n11660), .C2(n15468), .A(n8580), .B(n11890), .ZN(
        n15465) );
  OAI22_X1 U14188 ( .A1(n15392), .A2(n11662), .B1(n11661), .B2(n15384), .ZN(
        n11663) );
  AOI21_X1 U14189 ( .B1(n12736), .B2(n14038), .A(n11663), .ZN(n11664) );
  OAI21_X1 U14190 ( .B1(n15465), .B2(n13886), .A(n11664), .ZN(n11665) );
  AOI21_X1 U14191 ( .B1(n11666), .B2(n12324), .A(n11665), .ZN(n11667) );
  OAI21_X1 U14192 ( .B1(n15394), .B2(n15466), .A(n11667), .ZN(P2_U3254) );
  AOI21_X1 U14193 ( .B1(n11705), .B2(n15283), .A(n11668), .ZN(n11669) );
  OAI211_X1 U14194 ( .C1(n11671), .C2(n15248), .A(n11670), .B(n11669), .ZN(
        n11673) );
  NAND2_X1 U14195 ( .A1(n11673), .A2(n15140), .ZN(n11672) );
  OAI21_X1 U14196 ( .B1(n15140), .B2(n10637), .A(n11672), .ZN(P1_U3536) );
  NAND2_X1 U14197 ( .A1(n11673), .A2(n15291), .ZN(n11674) );
  OAI21_X1 U14198 ( .B1(n15291), .B2(n8041), .A(n11674), .ZN(P1_U3483) );
  INV_X1 U14199 ( .A(n15503), .ZN(n15535) );
  AND3_X1 U14200 ( .A1(n11675), .A2(n11676), .A3(n11677), .ZN(n11678) );
  OAI21_X1 U14201 ( .B1(n11679), .B2(n11678), .A(n15539), .ZN(n11688) );
  NOR2_X1 U14202 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11680), .ZN(n12104) );
  AOI21_X1 U14203 ( .B1(n15538), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n12104), .ZN(
        n11687) );
  NAND3_X1 U14204 ( .A1(n11682), .A2(n6714), .A3(n11681), .ZN(n11683) );
  NAND2_X1 U14205 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  NAND2_X1 U14206 ( .A1(n15500), .A2(n11685), .ZN(n11686) );
  AND3_X1 U14207 ( .A1(n11688), .A2(n11687), .A3(n11686), .ZN(n11695) );
  AND3_X1 U14208 ( .A1(n11691), .A2(n11690), .A3(n11689), .ZN(n11692) );
  OAI21_X1 U14209 ( .B1(n11693), .B2(n11692), .A(n15550), .ZN(n11694) );
  OAI211_X1 U14210 ( .C1(n15535), .C2(n11696), .A(n11695), .B(n11694), .ZN(
        P3_U3186) );
  NAND2_X1 U14211 ( .A1(n11524), .A2(n11709), .ZN(n11697) );
  OAI21_X1 U14212 ( .B1(n11700), .B2(n11699), .A(n12032), .ZN(n15278) );
  INV_X1 U14213 ( .A(n15278), .ZN(n15275) );
  OAI22_X1 U14214 ( .A1(n15120), .A2(n11701), .B1(n11951), .B2(n15117), .ZN(
        n11702) );
  AOI21_X1 U14215 ( .B1(n12030), .B2(n15215), .A(n11702), .ZN(n11717) );
  NAND2_X1 U14216 ( .A1(n11707), .A2(n11706), .ZN(n12021) );
  OAI21_X1 U14217 ( .B1(n11707), .B2(n11706), .A(n12021), .ZN(n11708) );
  NAND2_X1 U14218 ( .A1(n11708), .A2(n15253), .ZN(n11713) );
  OR2_X1 U14219 ( .A1(n11709), .A2(n15095), .ZN(n11711) );
  OR2_X1 U14220 ( .A1(n15096), .A2(n15097), .ZN(n11710) );
  NAND2_X1 U14221 ( .A1(n11711), .A2(n11710), .ZN(n11954) );
  INV_X1 U14222 ( .A(n11954), .ZN(n11712) );
  NAND2_X1 U14223 ( .A1(n11713), .A2(n11712), .ZN(n15277) );
  INV_X1 U14224 ( .A(n12030), .ZN(n11714) );
  OAI211_X1 U14225 ( .C1(n11714), .C2(n7260), .A(n6708), .B(n15209), .ZN(
        n15273) );
  NOR2_X1 U14226 ( .A1(n15273), .A2(n6681), .ZN(n11715) );
  OAI21_X1 U14227 ( .B1(n15277), .B2(n11715), .A(n15120), .ZN(n11716) );
  OAI211_X1 U14228 ( .C1(n15275), .C2(n14802), .A(n11717), .B(n11716), .ZN(
        P1_U3284) );
  NAND2_X1 U14229 ( .A1(n15625), .A2(n15656), .ZN(n11718) );
  XNOR2_X1 U14230 ( .A(n11719), .B(n11724), .ZN(n15653) );
  NAND2_X1 U14231 ( .A1(n15573), .A2(n12045), .ZN(n11720) );
  NAND2_X1 U14232 ( .A1(n15563), .A2(n15581), .ZN(n11722) );
  NAND2_X1 U14233 ( .A1(n12051), .A2(n12090), .ZN(n11723) );
  NAND2_X1 U14234 ( .A1(n11725), .A2(n11724), .ZN(n11960) );
  OAI211_X1 U14235 ( .C1(n11725), .C2(n11724), .A(n11960), .B(n15599), .ZN(
        n11727) );
  AOI22_X1 U14236 ( .A1(n15574), .A2(n15615), .B1(n15613), .B2(n12169), .ZN(
        n11726) );
  AND2_X1 U14237 ( .A1(n11727), .A2(n11726), .ZN(n15652) );
  INV_X1 U14238 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11728) );
  MUX2_X1 U14239 ( .A(n15652), .B(n11728), .S(n15627), .Z(n11730) );
  AOI22_X1 U14240 ( .A1(n15033), .A2(n15649), .B1(n15622), .B2(n12067), .ZN(
        n11729) );
  OAI211_X1 U14241 ( .C1(n13539), .C2(n15653), .A(n11730), .B(n11729), .ZN(
        P3_U3227) );
  INV_X1 U14242 ( .A(n11731), .ZN(n11733) );
  NAND3_X1 U14243 ( .A1(n11733), .A2(n11732), .A3(n13159), .ZN(n11734) );
  NAND2_X1 U14244 ( .A1(n11735), .A2(n11734), .ZN(n11749) );
  NAND2_X1 U14245 ( .A1(n15538), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n11737) );
  OAI21_X1 U14246 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15590), .A(n11737), .ZN(
        n11748) );
  OAI21_X1 U14247 ( .B1(n11740), .B2(n11739), .A(n11738), .ZN(n11745) );
  OAI21_X1 U14248 ( .B1(n11743), .B2(n11742), .A(n11741), .ZN(n11744) );
  AOI22_X1 U14249 ( .A1(n15539), .A2(n11745), .B1(n15500), .B2(n11744), .ZN(
        n11746) );
  INV_X1 U14250 ( .A(n11746), .ZN(n11747) );
  AOI211_X1 U14251 ( .C1(n15550), .C2(n11749), .A(n11748), .B(n11747), .ZN(
        n11750) );
  OAI21_X1 U14252 ( .B1(n7564), .B2(n15535), .A(n11750), .ZN(P3_U3184) );
  MUX2_X1 U14253 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13268), .Z(n11864) );
  INV_X1 U14254 ( .A(n11863), .ZN(n11751) );
  XNOR2_X1 U14255 ( .A(n11864), .B(n11751), .ZN(n11755) );
  NAND2_X1 U14256 ( .A1(n11755), .A2(n11754), .ZN(n11865) );
  OAI21_X1 U14257 ( .B1(n11755), .B2(n11754), .A(n11865), .ZN(n11773) );
  NAND2_X1 U14258 ( .A1(n15538), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n11758) );
  INV_X1 U14259 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11756) );
  NOR2_X1 U14260 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11756), .ZN(n12070) );
  INV_X1 U14261 ( .A(n12070), .ZN(n11757) );
  NAND2_X1 U14262 ( .A1(n11758), .A2(n11757), .ZN(n11772) );
  NAND2_X1 U14263 ( .A1(n11863), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11852) );
  OR2_X1 U14264 ( .A1(n11863), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11761) );
  NAND2_X1 U14265 ( .A1(n11852), .A2(n11761), .ZN(n11762) );
  AOI21_X1 U14266 ( .B1(n11763), .B2(n11762), .A(n11854), .ZN(n11770) );
  NAND2_X1 U14267 ( .A1(n11863), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11846) );
  OR2_X1 U14268 ( .A1(n11863), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U14269 ( .A1(n11846), .A2(n11766), .ZN(n11767) );
  AOI21_X1 U14270 ( .B1(n11768), .B2(n11767), .A(n11847), .ZN(n11769) );
  OAI22_X1 U14271 ( .A1(n11770), .A2(n15515), .B1(n15547), .B2(n11769), .ZN(
        n11771) );
  AOI211_X1 U14272 ( .C1(n15550), .C2(n11773), .A(n11772), .B(n11771), .ZN(
        n11774) );
  OAI21_X1 U14273 ( .B1(n11863), .B2(n15535), .A(n11774), .ZN(P3_U3188) );
  XNOR2_X1 U14274 ( .A(n11775), .B(n12906), .ZN(n15426) );
  INV_X1 U14275 ( .A(n11776), .ZN(n15391) );
  NAND2_X1 U14276 ( .A1(n15392), .A2(n15391), .ZN(n14105) );
  OAI21_X1 U14277 ( .B1(n12906), .B2(n11778), .A(n11777), .ZN(n11782) );
  OAI22_X1 U14278 ( .A1(n11779), .A2(n15388), .B1(n14090), .B2(n12678), .ZN(
        n11781) );
  NOR2_X1 U14279 ( .A1(n15426), .A2(n15471), .ZN(n11780) );
  AOI211_X1 U14280 ( .C1(n14129), .C2(n11782), .A(n11781), .B(n11780), .ZN(
        n15425) );
  MUX2_X1 U14281 ( .A(n11783), .B(n15425), .S(n15392), .Z(n11788) );
  AOI211_X1 U14282 ( .C1(n15423), .C2(n11795), .A(n6678), .B(n11837), .ZN(
        n15422) );
  OAI22_X1 U14283 ( .A1(n14102), .A2(n11785), .B1(n15384), .B2(n11784), .ZN(
        n11786) );
  AOI21_X1 U14284 ( .B1(n14108), .B2(n15422), .A(n11786), .ZN(n11787) );
  OAI211_X1 U14285 ( .C1(n15426), .C2(n14105), .A(n11788), .B(n11787), .ZN(
        P2_U3260) );
  XNOR2_X1 U14286 ( .A(n11789), .B(n11792), .ZN(n15420) );
  OAI21_X1 U14287 ( .B1(n11792), .B2(n11791), .A(n11790), .ZN(n11793) );
  AOI222_X1 U14288 ( .A1(n14129), .A2(n11793), .B1(n13796), .B2(n14126), .C1(
        n13798), .C2(n14124), .ZN(n15419) );
  MUX2_X1 U14289 ( .A(n11794), .B(n15419), .S(n15392), .Z(n11801) );
  INV_X1 U14290 ( .A(n11795), .ZN(n11796) );
  AOI211_X1 U14291 ( .C1(n15417), .C2(n11797), .A(n6678), .B(n11796), .ZN(
        n15416) );
  OAI22_X1 U14292 ( .A1(n14102), .A2(n7345), .B1(n15384), .B2(n11798), .ZN(
        n11799) );
  AOI21_X1 U14293 ( .B1(n14108), .B2(n15416), .A(n11799), .ZN(n11800) );
  OAI211_X1 U14294 ( .C1(n14133), .C2(n15420), .A(n11801), .B(n11800), .ZN(
        P2_U3261) );
  OAI21_X1 U14295 ( .B1(n11803), .B2(n12909), .A(n11802), .ZN(n15442) );
  AOI22_X1 U14296 ( .A1(n14124), .A2(n13794), .B1(n14126), .B2(n13792), .ZN(
        n11808) );
  XNOR2_X1 U14297 ( .A(n11805), .B(n11804), .ZN(n11806) );
  NAND2_X1 U14298 ( .A1(n11806), .A2(n14129), .ZN(n11807) );
  OAI211_X1 U14299 ( .C1(n15442), .C2(n15471), .A(n11808), .B(n11807), .ZN(
        n15445) );
  MUX2_X1 U14300 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n15445), .S(n15392), .Z(
        n11809) );
  INV_X1 U14301 ( .A(n11809), .ZN(n11815) );
  AOI21_X1 U14302 ( .B1(n12717), .B2(n11822), .A(n6678), .ZN(n11811) );
  AND2_X1 U14303 ( .A1(n11811), .A2(n11810), .ZN(n15443) );
  OAI22_X1 U14304 ( .A1(n7347), .A2(n14102), .B1(n15384), .B2(n11812), .ZN(
        n11813) );
  AOI21_X1 U14305 ( .B1(n14108), .B2(n15443), .A(n11813), .ZN(n11814) );
  OAI211_X1 U14306 ( .C1(n15442), .C2(n14105), .A(n11815), .B(n11814), .ZN(
        P2_U3257) );
  XNOR2_X1 U14307 ( .A(n15434), .B(n13794), .ZN(n12907) );
  INV_X1 U14308 ( .A(n12907), .ZN(n11816) );
  XNOR2_X1 U14309 ( .A(n11817), .B(n11816), .ZN(n15438) );
  XNOR2_X1 U14310 ( .A(n11818), .B(n12907), .ZN(n11821) );
  INV_X1 U14311 ( .A(n11819), .ZN(n11820) );
  AOI21_X1 U14312 ( .B1(n11821), .B2(n14129), .A(n11820), .ZN(n15440) );
  MUX2_X1 U14313 ( .A(n13837), .B(n15440), .S(n15392), .Z(n11828) );
  AOI21_X1 U14314 ( .B1(n11838), .B2(n15434), .A(n6678), .ZN(n11823) );
  AND2_X1 U14315 ( .A1(n11823), .A2(n11822), .ZN(n15435) );
  INV_X1 U14316 ( .A(n15434), .ZN(n11825) );
  OAI22_X1 U14317 ( .A1(n14102), .A2(n11825), .B1(n15384), .B2(n11824), .ZN(
        n11826) );
  AOI21_X1 U14318 ( .B1(n14108), .B2(n15435), .A(n11826), .ZN(n11827) );
  OAI211_X1 U14319 ( .C1(n15438), .C2(n14133), .A(n11828), .B(n11827), .ZN(
        P2_U3258) );
  XNOR2_X1 U14320 ( .A(n11830), .B(n11829), .ZN(n15432) );
  OAI21_X1 U14321 ( .B1(n11832), .B2(n12904), .A(n11831), .ZN(n11835) );
  OAI22_X1 U14322 ( .A1(n12692), .A2(n14090), .B1(n15388), .B2(n12706), .ZN(
        n11834) );
  NOR2_X1 U14323 ( .A1(n15432), .A2(n15471), .ZN(n11833) );
  AOI211_X1 U14324 ( .C1(n14129), .C2(n11835), .A(n11834), .B(n11833), .ZN(
        n15431) );
  MUX2_X1 U14325 ( .A(n11836), .B(n15431), .S(n15392), .Z(n11845) );
  INV_X1 U14326 ( .A(n11837), .ZN(n11840) );
  INV_X1 U14327 ( .A(n11838), .ZN(n11839) );
  AOI211_X1 U14328 ( .C1(n15429), .C2(n11840), .A(n6678), .B(n11839), .ZN(
        n15428) );
  OAI22_X1 U14329 ( .A1(n14102), .A2(n11842), .B1(n15384), .B2(n11841), .ZN(
        n11843) );
  AOI21_X1 U14330 ( .B1(n15428), .B2(n14108), .A(n11843), .ZN(n11844) );
  OAI211_X1 U14331 ( .C1(n15432), .C2(n14105), .A(n11845), .B(n11844), .ZN(
        P2_U3259) );
  NOR2_X1 U14332 ( .A1(n11861), .A2(n11848), .ZN(n11849) );
  NAND2_X1 U14333 ( .A1(n15522), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11850) );
  OAI21_X1 U14334 ( .B1(n15522), .B2(P3_REG1_REG_8__SCAN_IN), .A(n11850), .ZN(
        n15523) );
  AOI21_X1 U14335 ( .B1(n9752), .B2(n11851), .A(n11998), .ZN(n11883) );
  INV_X1 U14336 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11873) );
  INV_X1 U14337 ( .A(n11852), .ZN(n11853) );
  NOR2_X1 U14338 ( .A1(n11861), .A2(n11855), .ZN(n11856) );
  INV_X1 U14339 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11929) );
  NAND2_X1 U14340 ( .A1(n15522), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11857) );
  OAI21_X1 U14341 ( .B1(n15522), .B2(P3_REG2_REG_8__SCAN_IN), .A(n11857), .ZN(
        n15513) );
  AOI21_X1 U14342 ( .B1(n11873), .B2(n11858), .A(n11980), .ZN(n11859) );
  NOR2_X1 U14343 ( .A1(n11859), .A2(n15515), .ZN(n11881) );
  MUX2_X1 U14344 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13268), .Z(n11868) );
  INV_X1 U14345 ( .A(n15522), .ZN(n11869) );
  XNOR2_X1 U14346 ( .A(n11868), .B(n11869), .ZN(n15518) );
  MUX2_X1 U14347 ( .A(n11929), .B(n11860), .S(n13268), .Z(n11862) );
  NAND2_X1 U14348 ( .A1(n11862), .A2(n11861), .ZN(n11867) );
  XNOR2_X1 U14349 ( .A(n11862), .B(n11926), .ZN(n11922) );
  OR2_X1 U14350 ( .A1(n11864), .A2(n11863), .ZN(n11866) );
  NAND2_X1 U14351 ( .A1(n11866), .A2(n11865), .ZN(n11921) );
  NAND2_X1 U14352 ( .A1(n11922), .A2(n11921), .ZN(n11920) );
  NAND2_X1 U14353 ( .A1(n11867), .A2(n11920), .ZN(n15519) );
  NAND2_X1 U14354 ( .A1(n15518), .A2(n15519), .ZN(n11872) );
  INV_X1 U14355 ( .A(n11868), .ZN(n11870) );
  NAND2_X1 U14356 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  MUX2_X1 U14357 ( .A(n11873), .B(n9752), .S(n13268), .Z(n11874) );
  AND2_X1 U14358 ( .A1(n11874), .A2(n11997), .ZN(n11989) );
  INV_X1 U14359 ( .A(n11989), .ZN(n11875) );
  OR2_X1 U14360 ( .A1(n11874), .A2(n11997), .ZN(n11991) );
  NAND2_X1 U14361 ( .A1(n11875), .A2(n11991), .ZN(n11876) );
  XNOR2_X1 U14362 ( .A(n11990), .B(n11876), .ZN(n11879) );
  NAND2_X1 U14363 ( .A1(n15503), .A2(n11997), .ZN(n11878) );
  NOR2_X1 U14364 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9749), .ZN(n12192) );
  AOI21_X1 U14365 ( .B1(n15538), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12192), .ZN(
        n11877) );
  OAI211_X1 U14366 ( .C1(n11879), .C2(n15520), .A(n11878), .B(n11877), .ZN(
        n11880) );
  NOR2_X1 U14367 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  OAI21_X1 U14368 ( .B1(n11883), .B2(n15547), .A(n11882), .ZN(P3_U3191) );
  INV_X1 U14369 ( .A(n11884), .ZN(n11936) );
  OAI222_X1 U14370 ( .A1(n14949), .A2(n11886), .B1(n12208), .B2(n11936), .C1(
        n11885), .C2(P1_U3086), .ZN(P1_U3335) );
  XNOR2_X1 U14371 ( .A(n12749), .B(n12127), .ZN(n12914) );
  XNOR2_X1 U14372 ( .A(n12128), .B(n12914), .ZN(n11888) );
  AOI222_X1 U14373 ( .A1(n14129), .A2(n11888), .B1(n12755), .B2(n14126), .C1(
        n13790), .C2(n14124), .ZN(n15073) );
  XOR2_X1 U14374 ( .A(n12123), .B(n12914), .Z(n15076) );
  AOI21_X1 U14375 ( .B1(n12749), .B2(n11890), .A(n6678), .ZN(n11891) );
  NAND2_X1 U14376 ( .A1(n11891), .A2(n12133), .ZN(n15072) );
  OAI22_X1 U14377 ( .A1(n15392), .A2(n8837), .B1(n11941), .B2(n15384), .ZN(
        n11892) );
  AOI21_X1 U14378 ( .B1(n12749), .B2(n14038), .A(n11892), .ZN(n11893) );
  OAI21_X1 U14379 ( .B1(n15072), .B2(n13886), .A(n11893), .ZN(n11894) );
  AOI21_X1 U14380 ( .B1(n15076), .B2(n12324), .A(n11894), .ZN(n11895) );
  OAI21_X1 U14381 ( .B1(n15073), .B2(n15394), .A(n11895), .ZN(P2_U3253) );
  NOR2_X1 U14382 ( .A1(n11897), .A2(n11896), .ZN(n11899) );
  NOR2_X1 U14383 ( .A1(n11899), .A2(n11898), .ZN(n11904) );
  INV_X1 U14384 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11900) );
  XNOR2_X1 U14385 ( .A(n12424), .B(n11900), .ZN(n11903) );
  INV_X1 U14386 ( .A(n12431), .ZN(n11901) );
  AOI211_X1 U14387 ( .C1(n11904), .C2(n11903), .A(n11902), .B(n11901), .ZN(
        n11918) );
  NAND2_X1 U14388 ( .A1(n11906), .A2(n11905), .ZN(n11908) );
  NAND2_X1 U14389 ( .A1(n11908), .A2(n11907), .ZN(n11913) );
  INV_X1 U14390 ( .A(n12424), .ZN(n12429) );
  INV_X1 U14391 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U14392 ( .A1(n12429), .A2(n11910), .ZN(n11909) );
  OAI21_X1 U14393 ( .B1(n12429), .B2(n11910), .A(n11909), .ZN(n11912) );
  NAND2_X1 U14394 ( .A1(n12424), .A2(n11910), .ZN(n11911) );
  OAI211_X1 U14395 ( .C1(n11910), .C2(n12424), .A(n11913), .B(n11911), .ZN(
        n12423) );
  OAI211_X1 U14396 ( .C1(n11913), .C2(n11912), .A(n12423), .B(n15372), .ZN(
        n11916) );
  NAND2_X1 U14397 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13724)
         );
  INV_X1 U14398 ( .A(n13724), .ZN(n11914) );
  AOI21_X1 U14399 ( .B1(n15371), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11914), 
        .ZN(n11915) );
  OAI211_X1 U14400 ( .C1(n15379), .C2(n12424), .A(n11916), .B(n11915), .ZN(
        n11917) );
  OR2_X1 U14401 ( .A1(n11918), .A2(n11917), .ZN(P2_U3230) );
  NOR2_X1 U14402 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11919), .ZN(n12081) );
  AOI21_X1 U14403 ( .B1(n15538), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12081), .ZN(
        n11925) );
  OAI21_X1 U14404 ( .B1(n11922), .B2(n11921), .A(n11920), .ZN(n11923) );
  NAND2_X1 U14405 ( .A1(n15550), .A2(n11923), .ZN(n11924) );
  OAI211_X1 U14406 ( .C1(n15535), .C2(n11926), .A(n11925), .B(n11924), .ZN(
        n11935) );
  AOI21_X1 U14407 ( .B1(n11929), .B2(n11928), .A(n11927), .ZN(n11933) );
  AOI21_X1 U14408 ( .B1(n11860), .B2(n11931), .A(n11930), .ZN(n11932) );
  OAI22_X1 U14409 ( .A1(n11933), .A2(n15515), .B1(n15547), .B2(n11932), .ZN(
        n11934) );
  OR2_X1 U14410 ( .A1(n11935), .A2(n11934), .ZN(P3_U3189) );
  OAI222_X1 U14411 ( .A1(n14252), .A2(n7635), .B1(P2_U3088), .B2(n12897), .C1(
        n14254), .C2(n11936), .ZN(P2_U3307) );
  INV_X1 U14412 ( .A(n12749), .ZN(n15074) );
  OAI21_X1 U14413 ( .B1(n11939), .B2(n11938), .A(n11937), .ZN(n11940) );
  NAND2_X1 U14414 ( .A1(n11940), .A2(n9100), .ZN(n11945) );
  NAND2_X1 U14415 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15361)
         );
  INV_X1 U14416 ( .A(n15361), .ZN(n11943) );
  OAI22_X1 U14417 ( .A1(n13759), .A2(n12738), .B1(n13781), .B2(n11941), .ZN(
        n11942) );
  AOI211_X1 U14418 ( .C1(n13734), .C2(n12755), .A(n11943), .B(n11942), .ZN(
        n11944) );
  OAI211_X1 U14419 ( .C1(n15074), .C2(n13747), .A(n11945), .B(n11944), .ZN(
        P2_U3196) );
  NAND2_X1 U14420 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  XOR2_X1 U14421 ( .A(n11949), .B(n11948), .Z(n11956) );
  OAI22_X1 U14422 ( .A1(n15090), .A2(n11951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11950), .ZN(n11953) );
  NAND2_X1 U14423 ( .A1(n12030), .A2(n15283), .ZN(n15272) );
  NOR2_X1 U14424 ( .A1(n15272), .A2(n15093), .ZN(n11952) );
  AOI211_X1 U14425 ( .C1(n15105), .C2(n11954), .A(n11953), .B(n11952), .ZN(
        n11955) );
  OAI21_X1 U14426 ( .B1(n11956), .B2(n15101), .A(n11955), .ZN(P1_U3231) );
  XNOR2_X1 U14427 ( .A(n11958), .B(n11957), .ZN(n15661) );
  INV_X1 U14428 ( .A(n15661), .ZN(n11969) );
  NAND2_X1 U14429 ( .A1(n15562), .A2(n15649), .ZN(n11959) );
  NAND2_X1 U14430 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  NAND2_X1 U14431 ( .A1(n11961), .A2(n12057), .ZN(n12163) );
  OAI211_X1 U14432 ( .C1(n11961), .C2(n12057), .A(n12163), .B(n15599), .ZN(
        n11965) );
  OAI22_X1 U14433 ( .A1(n15597), .A2(n12215), .B1(n12054), .B2(n15594), .ZN(
        n11962) );
  INV_X1 U14434 ( .A(n11962), .ZN(n11964) );
  NAND2_X1 U14435 ( .A1(n15661), .A2(n15656), .ZN(n11963) );
  NAND3_X1 U14436 ( .A1(n11965), .A2(n11964), .A3(n11963), .ZN(n15659) );
  MUX2_X1 U14437 ( .A(n15659), .B(P3_REG2_REG_7__SCAN_IN), .S(n15627), .Z(
        n11966) );
  INV_X1 U14438 ( .A(n11966), .ZN(n11968) );
  NOR2_X1 U14439 ( .A1(n15607), .A2(n12083), .ZN(n15660) );
  AOI22_X1 U14440 ( .A1(n15583), .A2(n15660), .B1(n15622), .B2(n12077), .ZN(
        n11967) );
  OAI211_X1 U14441 ( .C1(n11969), .C2(n13351), .A(n11968), .B(n11967), .ZN(
        P3_U3226) );
  NAND2_X1 U14442 ( .A1(n11971), .A2(n11970), .ZN(n11973) );
  XOR2_X1 U14443 ( .A(n11973), .B(n11972), .Z(n11978) );
  NAND2_X1 U14444 ( .A1(n14401), .A2(n14986), .ZN(n12024) );
  NAND2_X1 U14445 ( .A1(n14985), .A2(n14987), .ZN(n12026) );
  NAND2_X1 U14446 ( .A1(n12024), .A2(n12026), .ZN(n15282) );
  NAND2_X1 U14447 ( .A1(n15282), .A2(n15105), .ZN(n11975) );
  OAI211_X1 U14448 ( .C1(n15090), .C2(n12025), .A(n11975), .B(n11974), .ZN(
        n11976) );
  AOI21_X1 U14449 ( .B1(n15284), .B2(n15088), .A(n11976), .ZN(n11977) );
  OAI21_X1 U14450 ( .B1(n11978), .B2(n15101), .A(n11977), .ZN(P1_U3217) );
  NOR2_X1 U14451 ( .A1(n11997), .A2(n11979), .ZN(n11981) );
  NAND2_X1 U14452 ( .A1(n11999), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n12268) );
  INV_X1 U14453 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U14454 ( .A1(n12007), .A2(n11982), .ZN(n11983) );
  NAND2_X1 U14455 ( .A1(n12268), .A2(n11983), .ZN(n11985) );
  INV_X1 U14456 ( .A(n12269), .ZN(n11984) );
  AOI21_X1 U14457 ( .B1(n11986), .B2(n11985), .A(n11984), .ZN(n12009) );
  MUX2_X1 U14458 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13268), .Z(n11987) );
  NOR2_X1 U14459 ( .A1(n11987), .A2(n11999), .ZN(n12260) );
  AOI21_X1 U14460 ( .B1(n11987), .B2(n11999), .A(n12260), .ZN(n11988) );
  INV_X1 U14461 ( .A(n11988), .ZN(n11993) );
  AOI21_X1 U14462 ( .B1(n11993), .B2(n11992), .A(n6832), .ZN(n11995) );
  NAND2_X1 U14463 ( .A1(n15538), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U14464 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n12250)
         );
  OAI211_X1 U14465 ( .C1(n11995), .C2(n15520), .A(n11994), .B(n12250), .ZN(
        n12006) );
  NAND2_X1 U14466 ( .A1(n11999), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U14467 ( .A1(n12007), .A2(n12000), .ZN(n12001) );
  NAND2_X1 U14468 ( .A1(n12256), .A2(n12001), .ZN(n12002) );
  NAND2_X1 U14469 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  AOI21_X1 U14470 ( .B1(n12257), .B2(n12004), .A(n15547), .ZN(n12005) );
  AOI211_X1 U14471 ( .C1(n15503), .C2(n12007), .A(n12006), .B(n12005), .ZN(
        n12008) );
  OAI21_X1 U14472 ( .B1(n12009), .B2(n15515), .A(n12008), .ZN(P3_U3192) );
  XNOR2_X1 U14473 ( .A(n12011), .B(n12010), .ZN(n12015) );
  AOI22_X1 U14474 ( .A1(n14124), .A2(n13789), .B1(n14126), .B2(n13788), .ZN(
        n12129) );
  OAI22_X1 U14475 ( .A1(n13742), .A2(n12129), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8852), .ZN(n12013) );
  INV_X1 U14476 ( .A(n12756), .ZN(n12284) );
  NOR2_X1 U14477 ( .A1(n12284), .A2(n13747), .ZN(n12012) );
  AOI211_X1 U14478 ( .C1(n13766), .C2(n12234), .A(n12013), .B(n12012), .ZN(
        n12014) );
  OAI21_X1 U14479 ( .B1(n12015), .B2(n13785), .A(n12014), .ZN(P2_U3206) );
  INV_X1 U14480 ( .A(n12016), .ZN(n12019) );
  OAI222_X1 U14481 ( .A1(n14252), .A2(n12017), .B1(n14254), .B2(n12019), .C1(
        n12862), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U14482 ( .A1(n14949), .A2(n7203), .B1(n12208), .B2(n12019), .C1(
        P1_U3086), .C2(n12018), .ZN(P1_U3334) );
  OAI211_X1 U14483 ( .C1(n12023), .C2(n12022), .A(n15253), .B(n12342), .ZN(
        n15286) );
  AND2_X1 U14484 ( .A1(n15286), .A2(n12024), .ZN(n12037) );
  OAI22_X1 U14485 ( .A1(n15120), .A2(n8077), .B1(n12025), .B2(n15117), .ZN(
        n12029) );
  AOI211_X1 U14486 ( .C1(n15284), .C2(n6708), .A(n14862), .B(n15115), .ZN(
        n15281) );
  INV_X1 U14487 ( .A(n15281), .ZN(n12027) );
  AOI21_X1 U14488 ( .B1(n12027), .B2(n12026), .A(n15124), .ZN(n12028) );
  AOI211_X1 U14489 ( .C1(n15215), .C2(n15284), .A(n12029), .B(n12028), .ZN(
        n12036) );
  NAND2_X1 U14490 ( .A1(n11714), .A2(n12020), .ZN(n12031) );
  OAI21_X1 U14491 ( .B1(n12034), .B2(n12033), .A(n12350), .ZN(n15288) );
  NAND2_X1 U14492 ( .A1(n15288), .A2(n15126), .ZN(n12035) );
  OAI211_X1 U14493 ( .C1(n6676), .C2(n12037), .A(n12036), .B(n12035), .ZN(
        P1_U3283) );
  INV_X1 U14494 ( .A(n12038), .ZN(n12039) );
  OAI222_X1 U14495 ( .A1(n14252), .A2(n12040), .B1(n14254), .B2(n12039), .C1(
        n8612), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U14496 ( .A(n12173), .ZN(n12066) );
  NAND2_X1 U14497 ( .A1(n12042), .A2(n12041), .ZN(n12043) );
  XNOR2_X1 U14498 ( .A(n12046), .B(n15596), .ZN(n12109) );
  INV_X1 U14499 ( .A(n12046), .ZN(n12047) );
  XNOR2_X1 U14500 ( .A(n12049), .B(n12094), .ZN(n12101) );
  NAND2_X1 U14501 ( .A1(n12049), .A2(n12094), .ZN(n12050) );
  XNOR2_X1 U14502 ( .A(n12598), .B(n15567), .ZN(n12052) );
  AND2_X1 U14503 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  XNOR2_X1 U14504 ( .A(n12598), .B(n12072), .ZN(n12055) );
  XNOR2_X1 U14505 ( .A(n12055), .B(n12054), .ZN(n12069) );
  NAND2_X1 U14506 ( .A1(n12055), .A2(n15562), .ZN(n12056) );
  XNOR2_X1 U14507 ( .A(n12057), .B(n13030), .ZN(n12079) );
  INV_X1 U14508 ( .A(n12079), .ZN(n12058) );
  NAND2_X1 U14509 ( .A1(n12058), .A2(n12169), .ZN(n12059) );
  XNOR2_X1 U14510 ( .A(n12598), .B(n12214), .ZN(n12184) );
  XNOR2_X1 U14511 ( .A(n12184), .B(n12215), .ZN(n12060) );
  OAI211_X1 U14512 ( .C1(n12061), .C2(n12060), .A(n12186), .B(n15494), .ZN(
        n12065) );
  NAND2_X1 U14513 ( .A1(n15492), .A2(n12305), .ZN(n12062) );
  NAND2_X1 U14514 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15530) );
  OAI211_X1 U14515 ( .C1(n13154), .C2(n12214), .A(n12062), .B(n15530), .ZN(
        n12063) );
  AOI21_X1 U14516 ( .B1(n13134), .B2(n12169), .A(n12063), .ZN(n12064) );
  OAI211_X1 U14517 ( .C1(n12066), .C2(n13121), .A(n12065), .B(n12064), .ZN(
        P3_U3161) );
  INV_X1 U14518 ( .A(n12067), .ZN(n12076) );
  AOI21_X1 U14519 ( .B1(n15492), .B2(n12169), .A(n12070), .ZN(n12071) );
  OAI21_X1 U14520 ( .B1(n12072), .B2(n13154), .A(n12071), .ZN(n12073) );
  AOI21_X1 U14521 ( .B1(n13134), .B2(n15574), .A(n12073), .ZN(n12074) );
  OAI211_X1 U14522 ( .C1(n12076), .C2(n13121), .A(n12075), .B(n12074), .ZN(
        P3_U3179) );
  INV_X1 U14523 ( .A(n12077), .ZN(n12087) );
  OAI211_X1 U14524 ( .C1(n12080), .C2(n12079), .A(n12078), .B(n15494), .ZN(
        n12086) );
  AOI21_X1 U14525 ( .B1(n15492), .B2(n12220), .A(n12081), .ZN(n12082) );
  OAI21_X1 U14526 ( .B1(n13154), .B2(n12083), .A(n12082), .ZN(n12084) );
  AOI21_X1 U14527 ( .B1(n13134), .B2(n15562), .A(n12084), .ZN(n12085) );
  OAI211_X1 U14528 ( .C1(n12087), .C2(n13121), .A(n12086), .B(n12085), .ZN(
        P3_U3153) );
  XOR2_X1 U14529 ( .A(n12089), .B(n12088), .Z(n12097) );
  NOR2_X1 U14530 ( .A1(n13154), .A2(n12090), .ZN(n12091) );
  AOI211_X1 U14531 ( .C1(n15492), .C2(n15562), .A(n12092), .B(n12091), .ZN(
        n12093) );
  OAI21_X1 U14532 ( .B1(n12094), .B2(n13149), .A(n12093), .ZN(n12095) );
  AOI21_X1 U14533 ( .B1(n15568), .B2(n13135), .A(n12095), .ZN(n12096) );
  OAI21_X1 U14534 ( .B1(n12097), .B2(n13142), .A(n12096), .ZN(P3_U3167) );
  INV_X1 U14535 ( .A(n12098), .ZN(n12099) );
  AOI21_X1 U14536 ( .B1(n12101), .B2(n12100), .A(n12099), .ZN(n12108) );
  NOR2_X1 U14537 ( .A1(n13154), .A2(n12102), .ZN(n12103) );
  AOI211_X1 U14538 ( .C1(n15492), .C2(n15574), .A(n12104), .B(n12103), .ZN(
        n12105) );
  OAI21_X1 U14539 ( .B1(n15596), .B2(n13149), .A(n12105), .ZN(n12106) );
  AOI21_X1 U14540 ( .B1(n15582), .B2(n13135), .A(n12106), .ZN(n12107) );
  OAI21_X1 U14541 ( .B1(n12108), .B2(n13142), .A(n12107), .ZN(P3_U3170) );
  AOI21_X1 U14542 ( .B1(n12110), .B2(n12109), .A(n13142), .ZN(n12112) );
  NAND2_X1 U14543 ( .A1(n12112), .A2(n12111), .ZN(n12118) );
  AOI21_X1 U14544 ( .B1(n15492), .B2(n15563), .A(n12113), .ZN(n12114) );
  OAI21_X1 U14545 ( .B1(n13154), .B2(n12115), .A(n12114), .ZN(n12116) );
  AOI21_X1 U14546 ( .B1(n13134), .B2(n15612), .A(n12116), .ZN(n12117) );
  OAI211_X1 U14547 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n13121), .A(n12118), .B(
        n12117), .ZN(P3_U3158) );
  NOR2_X1 U14548 ( .A1(n12119), .A2(n15396), .ZN(n12120) );
  NAND2_X1 U14549 ( .A1(n12749), .A2(n13789), .ZN(n12125) );
  INV_X1 U14550 ( .A(n12755), .ZN(n12283) );
  OR2_X1 U14551 ( .A1(n12756), .A2(n12283), .ZN(n12287) );
  NAND2_X1 U14552 ( .A1(n12756), .A2(n12283), .ZN(n12286) );
  NAND2_X1 U14553 ( .A1(n12287), .A2(n12286), .ZN(n12915) );
  XNOR2_X1 U14554 ( .A(n12281), .B(n12915), .ZN(n12236) );
  XOR2_X1 U14555 ( .A(n12915), .B(n12289), .Z(n12131) );
  INV_X1 U14556 ( .A(n12129), .ZN(n12130) );
  AOI21_X1 U14557 ( .B1(n12131), .B2(n14129), .A(n12130), .ZN(n12241) );
  INV_X1 U14558 ( .A(n12316), .ZN(n12132) );
  AOI211_X1 U14559 ( .C1(n12756), .C2(n12133), .A(n6678), .B(n12132), .ZN(
        n12239) );
  AOI21_X1 U14560 ( .B1(n15450), .B2(n12756), .A(n12239), .ZN(n12134) );
  OAI211_X1 U14561 ( .C1(n15454), .C2(n12236), .A(n12241), .B(n12134), .ZN(
        n12136) );
  NAND2_X1 U14562 ( .A1(n12136), .A2(n15475), .ZN(n12135) );
  OAI21_X1 U14563 ( .B1(n15475), .B2(n8856), .A(n12135), .ZN(P2_U3469) );
  NAND2_X1 U14564 ( .A1(n12136), .A2(n15489), .ZN(n12137) );
  OAI21_X1 U14565 ( .B1(n15489), .B2(n10907), .A(n12137), .ZN(P2_U3512) );
  INV_X1 U14566 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U14567 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14319)
         );
  OAI21_X1 U14568 ( .B1(n15197), .B2(n12138), .A(n14319), .ZN(n12147) );
  XNOR2_X1 U14569 ( .A(n14475), .B(n12139), .ZN(n14480) );
  NAND2_X1 U14570 ( .A1(n14480), .A2(n14481), .ZN(n14479) );
  OAI21_X1 U14571 ( .B1(n14475), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14479), 
        .ZN(n12142) );
  NAND2_X1 U14572 ( .A1(n15192), .A2(n12142), .ZN(n12143) );
  NAND2_X1 U14573 ( .A1(n12143), .A2(n15185), .ZN(n12145) );
  XNOR2_X1 U14574 ( .A(n12376), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12144) );
  NOR2_X1 U14575 ( .A1(n12144), .A2(n12145), .ZN(n12375) );
  AOI211_X1 U14576 ( .C1(n12145), .C2(n12144), .A(n12375), .B(n12377), .ZN(
        n12146) );
  AOI211_X1 U14577 ( .C1(n14489), .C2(n12376), .A(n12147), .B(n12146), .ZN(
        n12159) );
  XNOR2_X1 U14578 ( .A(n12150), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n14478) );
  OAI21_X1 U14579 ( .B1(n12149), .B2(n12353), .A(n12148), .ZN(n14477) );
  NAND2_X1 U14580 ( .A1(n14478), .A2(n14477), .ZN(n14476) );
  OAI21_X1 U14581 ( .B1(n12151), .B2(n12150), .A(n14476), .ZN(n12152) );
  NOR2_X1 U14582 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  XNOR2_X1 U14583 ( .A(n12153), .B(n12152), .ZN(n15182) );
  NOR2_X1 U14584 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15182), .ZN(n15181) );
  NOR2_X1 U14585 ( .A1(n12154), .A2(n15181), .ZN(n12157) );
  MUX2_X1 U14586 ( .A(n8194), .B(P1_REG2_REG_16__SCAN_IN), .S(n12376), .Z(
        n12155) );
  INV_X1 U14587 ( .A(n12155), .ZN(n12156) );
  NAND2_X1 U14588 ( .A1(n12156), .A2(n12157), .ZN(n12369) );
  OAI211_X1 U14589 ( .C1(n12157), .C2(n12156), .A(n14515), .B(n12369), .ZN(
        n12158) );
  NAND2_X1 U14590 ( .A1(n12159), .A2(n12158), .ZN(P1_U3259) );
  XNOR2_X1 U14591 ( .A(n12160), .B(n12164), .ZN(n15663) );
  NAND2_X1 U14592 ( .A1(n12169), .A2(n12161), .ZN(n12162) );
  NAND2_X1 U14593 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  NAND2_X1 U14594 ( .A1(n12217), .A2(n12167), .ZN(n12168) );
  NAND2_X1 U14595 ( .A1(n12168), .A2(n15599), .ZN(n12171) );
  AOI22_X1 U14596 ( .A1(n12305), .A2(n15613), .B1(n15615), .B2(n12169), .ZN(
        n12170) );
  OAI211_X1 U14597 ( .C1(n15602), .C2(n15663), .A(n12171), .B(n12170), .ZN(
        n15664) );
  MUX2_X1 U14598 ( .A(n15664), .B(P3_REG2_REG_8__SCAN_IN), .S(n15627), .Z(
        n12172) );
  INV_X1 U14599 ( .A(n12172), .ZN(n12175) );
  NOR2_X1 U14600 ( .A1(n12214), .A2(n15607), .ZN(n15665) );
  AOI22_X1 U14601 ( .A1(n15583), .A2(n15665), .B1(n15622), .B2(n12173), .ZN(
        n12174) );
  OAI211_X1 U14602 ( .C1(n15663), .C2(n13351), .A(n12175), .B(n12174), .ZN(
        P3_U3225) );
  NAND2_X1 U14603 ( .A1(n12179), .A2(n14246), .ZN(n12177) );
  NAND2_X1 U14604 ( .A1(n12176), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12960) );
  OAI211_X1 U14605 ( .C1(n12178), .C2(n14249), .A(n12177), .B(n12960), .ZN(
        P2_U3304) );
  NAND2_X1 U14606 ( .A1(n12179), .A2(n12509), .ZN(n12181) );
  OAI211_X1 U14607 ( .C1(n12182), .C2(n14949), .A(n12181), .B(n12180), .ZN(
        P1_U3332) );
  XNOR2_X1 U14608 ( .A(n12598), .B(n12183), .ZN(n12244) );
  XNOR2_X1 U14609 ( .A(n12244), .B(n12243), .ZN(n12190) );
  NAND2_X1 U14610 ( .A1(n12184), .A2(n12220), .ZN(n12185) );
  INV_X1 U14611 ( .A(n12190), .ZN(n12187) );
  INV_X1 U14612 ( .A(n12246), .ZN(n12188) );
  AOI21_X1 U14613 ( .B1(n12190), .B2(n12189), .A(n12188), .ZN(n12196) );
  NOR2_X1 U14614 ( .A1(n13154), .A2(n12223), .ZN(n12191) );
  AOI211_X1 U14615 ( .C1(n15492), .C2(n12563), .A(n12192), .B(n12191), .ZN(
        n12193) );
  OAI21_X1 U14616 ( .B1(n12215), .B2(n13149), .A(n12193), .ZN(n12194) );
  AOI21_X1 U14617 ( .B1(n12224), .B2(n13151), .A(n12194), .ZN(n12195) );
  OAI21_X1 U14618 ( .B1(n12196), .B2(n13142), .A(n12195), .ZN(P3_U3171) );
  INV_X1 U14619 ( .A(n12761), .ZN(n12334) );
  OAI21_X1 U14620 ( .B1(n12199), .B2(n12198), .A(n12197), .ZN(n12200) );
  NAND2_X1 U14621 ( .A1(n12200), .A2(n9100), .ZN(n12205) );
  INV_X1 U14622 ( .A(n12319), .ZN(n12203) );
  AOI22_X1 U14623 ( .A1(n14126), .A2(n13787), .B1(n14124), .B2(n12755), .ZN(
        n12313) );
  OAI22_X1 U14624 ( .A1(n13742), .A2(n12313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12201), .ZN(n12202) );
  AOI21_X1 U14625 ( .B1(n12203), .B2(n13766), .A(n12202), .ZN(n12204) );
  OAI211_X1 U14626 ( .C1(n12334), .C2(n13747), .A(n12205), .B(n12204), .ZN(
        P2_U3187) );
  INV_X1 U14627 ( .A(n12206), .ZN(n12211) );
  OAI222_X1 U14628 ( .A1(n14949), .A2(n12209), .B1(n12208), .B2(n12211), .C1(
        n12207), .C2(P1_U3086), .ZN(P1_U3331) );
  OAI222_X1 U14629 ( .A1(n14252), .A2(n12212), .B1(n14254), .B2(n12211), .C1(
        n12210), .C2(P2_U3088), .ZN(P2_U3303) );
  XNOR2_X1 U14630 ( .A(n12213), .B(n12218), .ZN(n15668) );
  NAND2_X1 U14631 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  NAND2_X1 U14632 ( .A1(n12219), .A2(n12218), .ZN(n12302) );
  OAI211_X1 U14633 ( .C1(n12219), .C2(n12218), .A(n12302), .B(n15599), .ZN(
        n12222) );
  AOI22_X1 U14634 ( .A1(n15615), .A2(n12220), .B1(n12563), .B2(n15613), .ZN(
        n12221) );
  OAI211_X1 U14635 ( .C1(n15602), .C2(n15668), .A(n12222), .B(n12221), .ZN(
        n15669) );
  NAND2_X1 U14636 ( .A1(n15669), .A2(n15625), .ZN(n12229) );
  NOR2_X1 U14637 ( .A1(n15607), .A2(n12223), .ZN(n15670) );
  INV_X1 U14638 ( .A(n15670), .ZN(n12226) );
  INV_X1 U14639 ( .A(n12224), .ZN(n12225) );
  OAI22_X1 U14640 ( .A1(n12488), .A2(n12226), .B1(n12225), .B2(n15591), .ZN(
        n12227) );
  AOI21_X1 U14641 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15627), .A(n12227), .ZN(
        n12228) );
  OAI211_X1 U14642 ( .C1(n15668), .C2(n13351), .A(n12229), .B(n12228), .ZN(
        P3_U3224) );
  INV_X1 U14643 ( .A(SI_24_), .ZN(n12232) );
  INV_X1 U14644 ( .A(n12230), .ZN(n12231) );
  OAI222_X1 U14645 ( .A1(n12233), .A2(P3_U3151), .B1(n12971), .B2(n12232), 
        .C1(n13672), .C2(n12231), .ZN(P3_U3271) );
  AOI22_X1 U14646 ( .A1(n15394), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12234), 
        .B2(n14117), .ZN(n12235) );
  OAI21_X1 U14647 ( .B1(n12284), .B2(n14102), .A(n12235), .ZN(n12238) );
  NOR2_X1 U14648 ( .A1(n12236), .A2(n14133), .ZN(n12237) );
  AOI211_X1 U14649 ( .C1(n12239), .C2(n14108), .A(n12238), .B(n12237), .ZN(
        n12240) );
  OAI21_X1 U14650 ( .B1(n15394), .B2(n12241), .A(n12240), .ZN(P2_U3252) );
  INV_X1 U14651 ( .A(n12242), .ZN(n12308) );
  NAND2_X1 U14652 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  XNOR2_X1 U14653 ( .A(n12598), .B(n12442), .ZN(n12562) );
  XNOR2_X1 U14654 ( .A(n12562), .B(n13116), .ZN(n12248) );
  AOI21_X1 U14655 ( .B1(n12247), .B2(n12248), .A(n13142), .ZN(n12249) );
  NAND2_X1 U14656 ( .A1(n12249), .A2(n12566), .ZN(n12255) );
  NAND2_X1 U14657 ( .A1(n15492), .A2(n13111), .ZN(n12251) );
  OAI211_X1 U14658 ( .C1(n13154), .C2(n12252), .A(n12251), .B(n12250), .ZN(
        n12253) );
  AOI21_X1 U14659 ( .B1(n13134), .B2(n12305), .A(n12253), .ZN(n12254) );
  OAI211_X1 U14660 ( .C1(n12308), .C2(n13121), .A(n12255), .B(n12254), .ZN(
        P3_U3157) );
  AND2_X2 U14661 ( .A1(n12257), .A2(n12256), .ZN(n13189) );
  AOI21_X1 U14662 ( .B1(n12259), .B2(n12258), .A(n13191), .ZN(n12275) );
  INV_X1 U14663 ( .A(n15538), .ZN(n15532) );
  INV_X1 U14664 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12267) );
  INV_X1 U14665 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12463) );
  MUX2_X1 U14666 ( .A(n12463), .B(n12259), .S(n13268), .Z(n13182) );
  XNOR2_X1 U14667 ( .A(n13182), .B(n13190), .ZN(n12262) );
  NOR2_X1 U14668 ( .A1(n12261), .A2(n12262), .ZN(n13181) );
  AOI21_X1 U14669 ( .B1(n12262), .B2(n12261), .A(n13181), .ZN(n12263) );
  OR2_X1 U14670 ( .A1(n15520), .A2(n12263), .ZN(n12266) );
  NOR2_X1 U14671 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12264), .ZN(n13113) );
  INV_X1 U14672 ( .A(n13113), .ZN(n12265) );
  OAI211_X1 U14673 ( .C1(n15532), .C2(n12267), .A(n12266), .B(n12265), .ZN(
        n12273) );
  AOI21_X1 U14674 ( .B1(n12463), .B2(n12270), .A(n13174), .ZN(n12271) );
  NOR2_X1 U14675 ( .A1(n12271), .A2(n15515), .ZN(n12272) );
  AOI211_X1 U14676 ( .C1(n15503), .C2(n13190), .A(n12273), .B(n12272), .ZN(
        n12274) );
  OAI21_X1 U14677 ( .B1(n12275), .B2(n15547), .A(n12274), .ZN(P3_U3193) );
  INV_X1 U14678 ( .A(n12276), .ZN(n12278) );
  OAI222_X1 U14679 ( .A1(P3_U3151), .A2(n12280), .B1(n12279), .B2(n12278), 
        .C1(n12277), .C2(n12971), .ZN(P3_U3270) );
  OAI21_X1 U14680 ( .B1(n12756), .B2(n12755), .A(n12281), .ZN(n12282) );
  INV_X1 U14681 ( .A(n13788), .ZN(n12285) );
  XNOR2_X1 U14682 ( .A(n12761), .B(n12285), .ZN(n12917) );
  INV_X1 U14683 ( .A(n13787), .ZN(n12496) );
  XNOR2_X1 U14684 ( .A(n12771), .B(n12496), .ZN(n12920) );
  XNOR2_X1 U14685 ( .A(n12498), .B(n12920), .ZN(n12388) );
  INV_X1 U14686 ( .A(n12388), .ZN(n12299) );
  INV_X1 U14687 ( .A(n12286), .ZN(n12288) );
  XNOR2_X1 U14688 ( .A(n12493), .B(n12920), .ZN(n12290) );
  NOR2_X1 U14689 ( .A1(n12290), .A2(n14095), .ZN(n12386) );
  NAND2_X1 U14690 ( .A1(n14125), .A2(n14126), .ZN(n12292) );
  NAND2_X1 U14691 ( .A1(n14124), .A2(n13788), .ZN(n12291) );
  AND2_X1 U14692 ( .A1(n12292), .A2(n12291), .ZN(n12384) );
  INV_X1 U14693 ( .A(n12384), .ZN(n12293) );
  OAI21_X1 U14694 ( .B1(n12386), .B2(n12293), .A(n15392), .ZN(n12298) );
  OAI22_X1 U14695 ( .A1(n15392), .A2(n12294), .B1(n12364), .B2(n15384), .ZN(
        n12296) );
  INV_X1 U14696 ( .A(n12771), .ZN(n12497) );
  OAI211_X1 U14697 ( .C1(n12497), .C2(n7351), .A(n12500), .B(n8580), .ZN(
        n12385) );
  NOR2_X1 U14698 ( .A1(n12385), .A2(n13886), .ZN(n12295) );
  AOI211_X1 U14699 ( .C1(n14038), .C2(n12771), .A(n12296), .B(n12295), .ZN(
        n12297) );
  OAI211_X1 U14700 ( .C1(n12299), .C2(n14133), .A(n12298), .B(n12297), .ZN(
        P2_U3250) );
  XOR2_X1 U14701 ( .A(n12303), .B(n12300), .Z(n15676) );
  NAND2_X1 U14702 ( .A1(n12302), .A2(n12301), .ZN(n12304) );
  NAND2_X1 U14703 ( .A1(n12304), .A2(n12303), .ZN(n12479) );
  OAI211_X1 U14704 ( .C1(n12304), .C2(n12303), .A(n12479), .B(n15599), .ZN(
        n12307) );
  AOI22_X1 U14705 ( .A1(n15615), .A2(n12305), .B1(n13111), .B2(n15613), .ZN(
        n12306) );
  NAND2_X1 U14706 ( .A1(n12307), .A2(n12306), .ZN(n15678) );
  NAND2_X1 U14707 ( .A1(n15678), .A2(n15625), .ZN(n12311) );
  NAND2_X1 U14708 ( .A1(n15650), .A2(n12442), .ZN(n15674) );
  OAI22_X1 U14709 ( .A1(n12488), .A2(n15674), .B1(n12308), .B2(n15591), .ZN(
        n12309) );
  AOI21_X1 U14710 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15627), .A(n12309), 
        .ZN(n12310) );
  OAI211_X1 U14711 ( .C1(n13539), .C2(n15676), .A(n12311), .B(n12310), .ZN(
        P3_U3223) );
  XOR2_X1 U14712 ( .A(n12917), .B(n12312), .Z(n12314) );
  OAI21_X1 U14713 ( .B1(n12314), .B2(n14095), .A(n12313), .ZN(n12335) );
  INV_X1 U14714 ( .A(n12335), .ZN(n12326) );
  XOR2_X1 U14715 ( .A(n12917), .B(n12315), .Z(n12337) );
  AOI21_X1 U14716 ( .B1(n12761), .B2(n12316), .A(n6678), .ZN(n12318) );
  NAND2_X1 U14717 ( .A1(n12318), .A2(n12317), .ZN(n12333) );
  INV_X1 U14718 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12320) );
  OAI22_X1 U14719 ( .A1(n15392), .A2(n12320), .B1(n12319), .B2(n15384), .ZN(
        n12321) );
  AOI21_X1 U14720 ( .B1(n12761), .B2(n14038), .A(n12321), .ZN(n12322) );
  OAI21_X1 U14721 ( .B1(n12333), .B2(n13886), .A(n12322), .ZN(n12323) );
  AOI21_X1 U14722 ( .B1(n12337), .B2(n12324), .A(n12323), .ZN(n12325) );
  OAI21_X1 U14723 ( .B1(n12326), .B2(n15394), .A(n12325), .ZN(P2_U3251) );
  INV_X1 U14724 ( .A(n12327), .ZN(n12331) );
  OAI222_X1 U14725 ( .A1(n14949), .A2(n12329), .B1(n12208), .B2(n12331), .C1(
        n12328), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U14726 ( .A1(n14252), .A2(n12332), .B1(n14254), .B2(n12331), .C1(
        n12330), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI21_X1 U14727 ( .B1(n12334), .B2(n15467), .A(n12333), .ZN(n12336) );
  AOI211_X1 U14728 ( .C1(n15077), .C2(n12337), .A(n12336), .B(n12335), .ZN(
        n12340) );
  NAND2_X1 U14729 ( .A1(n15487), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12338) );
  OAI21_X1 U14730 ( .B1(n12340), .B2(n15487), .A(n12338), .ZN(P2_U3513) );
  NAND2_X1 U14731 ( .A1(n15474), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n12339) );
  OAI21_X1 U14732 ( .B1(n12340), .B2(n15474), .A(n12339), .ZN(P2_U3472) );
  OR2_X1 U14733 ( .A1(n15284), .A2(n15096), .ZN(n12341) );
  INV_X1 U14734 ( .A(n14985), .ZN(n12344) );
  NAND2_X1 U14735 ( .A1(n15122), .A2(n12344), .ZN(n12343) );
  OR2_X1 U14736 ( .A1(n15122), .A2(n12344), .ZN(n12345) );
  NAND2_X1 U14737 ( .A1(n12346), .A2(n12345), .ZN(n14984) );
  NAND2_X1 U14738 ( .A1(n14984), .A2(n14983), .ZN(n12348) );
  OR2_X1 U14739 ( .A1(n15087), .A2(n15098), .ZN(n12347) );
  NAND2_X1 U14740 ( .A1(n12348), .A2(n12347), .ZN(n12407) );
  XNOR2_X1 U14741 ( .A(n12407), .B(n12406), .ZN(n15132) );
  XNOR2_X1 U14742 ( .A(n12402), .B(n12401), .ZN(n15134) );
  NAND2_X1 U14743 ( .A1(n15134), .A2(n15126), .ZN(n12361) );
  OAI22_X1 U14744 ( .A1(n15120), .A2(n12353), .B1(n12396), .B2(n15117), .ZN(
        n12359) );
  INV_X1 U14745 ( .A(n15122), .ZN(n15116) );
  NAND2_X1 U14746 ( .A1(n15113), .A2(n14998), .ZN(n14993) );
  INV_X1 U14747 ( .A(n12404), .ZN(n12354) );
  AOI211_X1 U14748 ( .C1(n15130), .C2(n14993), .A(n14862), .B(n12354), .ZN(
        n15128) );
  OR2_X1 U14749 ( .A1(n14560), .A2(n15097), .ZN(n12356) );
  NAND2_X1 U14750 ( .A1(n14399), .A2(n14986), .ZN(n12355) );
  NAND2_X1 U14751 ( .A1(n12356), .A2(n12355), .ZN(n15129) );
  AOI21_X1 U14752 ( .B1(n15128), .B2(n6966), .A(n15129), .ZN(n12357) );
  NOR2_X1 U14753 ( .A1(n12357), .A2(n6676), .ZN(n12358) );
  AOI211_X1 U14754 ( .C1(n15215), .C2(n15130), .A(n12359), .B(n12358), .ZN(
        n12360) );
  OAI211_X1 U14755 ( .C1(n15132), .C2(n14697), .A(n12361), .B(n12360), .ZN(
        P1_U3280) );
  XNOR2_X1 U14756 ( .A(n12363), .B(n12362), .ZN(n12368) );
  NOR2_X1 U14757 ( .A1(n13781), .A2(n12364), .ZN(n12366) );
  OAI22_X1 U14758 ( .A1(n13742), .A2(n12384), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8883), .ZN(n12365) );
  AOI211_X1 U14759 ( .C1(n12771), .C2(n13783), .A(n12366), .B(n12365), .ZN(
        n12367) );
  OAI21_X1 U14760 ( .B1(n12368), .B2(n13785), .A(n12367), .ZN(P2_U3213) );
  NAND2_X1 U14761 ( .A1(n12376), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U14762 ( .A1(n12370), .A2(n12369), .ZN(n12373) );
  NOR2_X1 U14763 ( .A1(n14491), .A2(n14767), .ZN(n12371) );
  AOI21_X1 U14764 ( .B1(n14767), .B2(n14491), .A(n12371), .ZN(n12372) );
  NAND2_X1 U14765 ( .A1(n12372), .A2(n12373), .ZN(n14490) );
  OAI211_X1 U14766 ( .C1(n12373), .C2(n12372), .A(n14515), .B(n14490), .ZN(
        n12383) );
  INV_X1 U14767 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n12374) );
  NAND2_X1 U14768 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14328)
         );
  OAI21_X1 U14769 ( .B1(n15197), .B2(n12374), .A(n14328), .ZN(n12381) );
  XNOR2_X1 U14770 ( .A(n14494), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12378) );
  NOR2_X1 U14771 ( .A1(n12379), .A2(n12378), .ZN(n14493) );
  AOI211_X1 U14772 ( .C1(n12379), .C2(n12378), .A(n14493), .B(n12377), .ZN(
        n12380) );
  AOI211_X1 U14773 ( .C1(n14489), .C2(n14494), .A(n12381), .B(n12380), .ZN(
        n12382) );
  NAND2_X1 U14774 ( .A1(n12383), .A2(n12382), .ZN(P1_U3260) );
  OAI211_X1 U14775 ( .C1(n12497), .C2(n15467), .A(n12385), .B(n12384), .ZN(
        n12387) );
  AOI211_X1 U14776 ( .C1(n15077), .C2(n12388), .A(n12387), .B(n12386), .ZN(
        n12391) );
  NAND2_X1 U14777 ( .A1(n15487), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n12389) );
  OAI21_X1 U14778 ( .B1(n12391), .B2(n15487), .A(n12389), .ZN(P2_U3514) );
  NAND2_X1 U14779 ( .A1(n15474), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n12390) );
  OAI21_X1 U14780 ( .B1(n12391), .B2(n15474), .A(n12390), .ZN(P2_U3475) );
  INV_X1 U14781 ( .A(n15130), .ZN(n12400) );
  OAI211_X1 U14782 ( .C1(n12394), .C2(n12393), .A(n12392), .B(n15081), .ZN(
        n12399) );
  OAI21_X1 U14783 ( .B1(n15090), .B2(n12396), .A(n12395), .ZN(n12397) );
  AOI21_X1 U14784 ( .B1(n15129), .B2(n15105), .A(n12397), .ZN(n12398) );
  OAI211_X1 U14785 ( .C1(n12400), .C2(n14388), .A(n12399), .B(n12398), .ZN(
        P1_U3234) );
  AOI22_X1 U14786 ( .A1(n12402), .A2(n12401), .B1(n12400), .B2(n12412), .ZN(
        n12403) );
  NAND2_X1 U14787 ( .A1(n12403), .A2(n12410), .ZN(n14559) );
  OAI21_X1 U14788 ( .B1(n12403), .B2(n12410), .A(n14559), .ZN(n14924) );
  AOI22_X1 U14789 ( .A1(n14921), .A2(n15215), .B1(n6676), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n12420) );
  AOI21_X1 U14790 ( .B1(n14921), .B2(n12404), .A(n14862), .ZN(n12405) );
  OR2_X2 U14791 ( .A1(n14921), .A2(n12404), .ZN(n14788) );
  AND2_X1 U14792 ( .A1(n12405), .A2(n14788), .ZN(n14919) );
  INV_X1 U14793 ( .A(n14919), .ZN(n12417) );
  NAND2_X1 U14794 ( .A1(n12407), .A2(n12406), .ZN(n12409) );
  OR2_X1 U14795 ( .A1(n15130), .A2(n12412), .ZN(n12408) );
  XNOR2_X1 U14796 ( .A(n14538), .B(n12410), .ZN(n12411) );
  NAND2_X1 U14797 ( .A1(n12411), .A2(n15253), .ZN(n14922) );
  INV_X1 U14798 ( .A(n14271), .ZN(n12415) );
  INV_X1 U14799 ( .A(n15117), .ZN(n15217) );
  OR2_X1 U14800 ( .A1(n14562), .A2(n15097), .ZN(n12414) );
  OR2_X1 U14801 ( .A1(n12412), .A2(n15095), .ZN(n12413) );
  NAND2_X1 U14802 ( .A1(n12414), .A2(n12413), .ZN(n14920) );
  AOI21_X1 U14803 ( .B1(n12415), .B2(n15217), .A(n14920), .ZN(n12416) );
  OAI211_X1 U14804 ( .C1(n6681), .C2(n12417), .A(n14922), .B(n12416), .ZN(
        n12418) );
  NAND2_X1 U14805 ( .A1(n12418), .A2(n15120), .ZN(n12419) );
  OAI211_X1 U14806 ( .C1(n14924), .C2(n14802), .A(n12420), .B(n12419), .ZN(
        P1_U3279) );
  NOR2_X1 U14807 ( .A1(n15378), .A2(n12421), .ZN(n12422) );
  AOI21_X1 U14808 ( .B1(n12421), .B2(n15378), .A(n12422), .ZN(n15374) );
  OAI21_X1 U14809 ( .B1(n11910), .B2(n12424), .A(n12423), .ZN(n15375) );
  NAND2_X1 U14810 ( .A1(n15374), .A2(n15375), .ZN(n15373) );
  OAI21_X1 U14811 ( .B1(n15378), .B2(n12421), .A(n15373), .ZN(n12425) );
  NOR2_X1 U14812 ( .A1(n12425), .A2(n12426), .ZN(n13859) );
  AOI21_X1 U14813 ( .B1(n12426), .B2(n12425), .A(n13859), .ZN(n12427) );
  INV_X1 U14814 ( .A(n12427), .ZN(n12428) );
  NOR2_X1 U14815 ( .A1(n12428), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13860) );
  AOI21_X1 U14816 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12428), .A(n13860), 
        .ZN(n12441) );
  INV_X1 U14817 ( .A(n15378), .ZN(n12432) );
  NAND2_X1 U14818 ( .A1(n12429), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12430) );
  NAND2_X1 U14819 ( .A1(n12431), .A2(n12430), .ZN(n15366) );
  XNOR2_X1 U14820 ( .A(n15378), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15365) );
  AOI21_X1 U14821 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n12432), .A(n15367), 
        .ZN(n12433) );
  NOR2_X1 U14822 ( .A1(n12433), .A2(n12437), .ZN(n13862) );
  AOI21_X1 U14823 ( .B1(n12433), .B2(n12437), .A(n13862), .ZN(n12435) );
  AND2_X1 U14824 ( .A1(n12435), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13863) );
  INV_X1 U14825 ( .A(n13863), .ZN(n12434) );
  OAI211_X1 U14826 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n12435), .A(n12434), 
        .B(n15364), .ZN(n12440) );
  NAND2_X1 U14827 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13768)
         );
  NAND2_X1 U14828 ( .A1(n15371), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n12436) );
  OAI211_X1 U14829 ( .C1(n15379), .C2(n12437), .A(n13768), .B(n12436), .ZN(
        n12438) );
  INV_X1 U14830 ( .A(n12438), .ZN(n12439) );
  OAI211_X1 U14831 ( .C1(n12441), .C2(n13867), .A(n12440), .B(n12439), .ZN(
        P2_U3232) );
  NAND2_X1 U14832 ( .A1(n12563), .A2(n12442), .ZN(n12468) );
  NAND2_X1 U14833 ( .A1(n12479), .A2(n12468), .ZN(n12460) );
  NAND2_X1 U14834 ( .A1(n13055), .A2(n15056), .ZN(n12470) );
  NAND2_X1 U14835 ( .A1(n12460), .A2(n12470), .ZN(n12443) );
  NAND2_X1 U14836 ( .A1(n13111), .A2(n13118), .ZN(n12467) );
  NAND2_X1 U14837 ( .A1(n12443), .A2(n12467), .ZN(n12444) );
  XNOR2_X1 U14838 ( .A(n12444), .B(n12450), .ZN(n12447) );
  NAND2_X1 U14839 ( .A1(n15613), .A2(n13052), .ZN(n12445) );
  OAI21_X1 U14840 ( .B1(n13055), .B2(n15594), .A(n12445), .ZN(n12446) );
  AOI21_X1 U14841 ( .B1(n12447), .B2(n15599), .A(n12446), .ZN(n15054) );
  AND2_X1 U14842 ( .A1(n12449), .A2(n12448), .ZN(n12451) );
  XNOR2_X1 U14843 ( .A(n12451), .B(n12450), .ZN(n15052) );
  NOR2_X1 U14844 ( .A1(n12571), .A2(n15607), .ZN(n15050) );
  INV_X1 U14845 ( .A(n15050), .ZN(n12453) );
  AOI22_X1 U14846 ( .A1(n15627), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15622), 
        .B2(n13050), .ZN(n12452) );
  OAI21_X1 U14847 ( .B1(n12488), .B2(n12453), .A(n12452), .ZN(n12454) );
  AOI21_X1 U14848 ( .B1(n15052), .B2(n13524), .A(n12454), .ZN(n12455) );
  OAI21_X1 U14849 ( .B1(n15054), .B2(n15627), .A(n12455), .ZN(P3_U3221) );
  NAND2_X1 U14850 ( .A1(n12457), .A2(n12456), .ZN(n12458) );
  XNOR2_X1 U14851 ( .A(n12458), .B(n12459), .ZN(n15057) );
  XNOR2_X1 U14852 ( .A(n12460), .B(n12459), .ZN(n12461) );
  OAI222_X1 U14853 ( .A1(n15597), .A2(n13531), .B1(n15594), .B2(n13116), .C1(
        n12461), .C2(n15619), .ZN(n15059) );
  NAND2_X1 U14854 ( .A1(n15059), .A2(n15625), .ZN(n12466) );
  INV_X1 U14855 ( .A(n12462), .ZN(n13122) );
  OAI22_X1 U14856 ( .A1(n15625), .A2(n12463), .B1(n13122), .B2(n15591), .ZN(
        n12464) );
  AOI21_X1 U14857 ( .B1(n15033), .B2(n13118), .A(n12464), .ZN(n12465) );
  OAI211_X1 U14858 ( .C1(n13539), .C2(n15057), .A(n12466), .B(n12465), .ZN(
        P3_U3222) );
  NAND2_X1 U14859 ( .A1(n13114), .A2(n13057), .ZN(n12472) );
  AND2_X1 U14860 ( .A1(n12467), .A2(n12472), .ZN(n12469) );
  AND2_X1 U14861 ( .A1(n12468), .A2(n12469), .ZN(n12478) );
  INV_X1 U14862 ( .A(n12469), .ZN(n12471) );
  OR2_X1 U14863 ( .A1(n12471), .A2(n12470), .ZN(n12476) );
  INV_X1 U14864 ( .A(n12472), .ZN(n12474) );
  OR2_X1 U14865 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  AOI21_X2 U14866 ( .B1(n12479), .B2(n12478), .A(n12477), .ZN(n13529) );
  NAND2_X1 U14867 ( .A1(n13529), .A2(n13528), .ZN(n12481) );
  INV_X1 U14868 ( .A(n13052), .ZN(n13005) );
  OR2_X1 U14869 ( .A1(n15046), .A2(n13005), .ZN(n12480) );
  XNOR2_X1 U14870 ( .A(n12517), .B(n12482), .ZN(n12485) );
  NAND2_X1 U14871 ( .A1(n15613), .A2(n13503), .ZN(n12483) );
  OAI21_X1 U14872 ( .B1(n13005), .B2(n15594), .A(n12483), .ZN(n12484) );
  AOI21_X1 U14873 ( .B1(n12485), .B2(n15599), .A(n12484), .ZN(n15044) );
  XNOR2_X1 U14874 ( .A(n12486), .B(n12516), .ZN(n15042) );
  NOR2_X1 U14875 ( .A1(n13010), .A2(n15607), .ZN(n15041) );
  INV_X1 U14876 ( .A(n15041), .ZN(n12489) );
  AOI22_X1 U14877 ( .A1(n15627), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15622), 
        .B2(n13007), .ZN(n12487) );
  OAI21_X1 U14878 ( .B1(n12489), .B2(n12488), .A(n12487), .ZN(n12490) );
  AOI21_X1 U14879 ( .B1(n15042), .B2(n13524), .A(n12490), .ZN(n12491) );
  OAI21_X1 U14880 ( .B1(n15044), .B2(n15627), .A(n12491), .ZN(P3_U3219) );
  NOR2_X1 U14881 ( .A1(n12497), .A2(n13787), .ZN(n12492) );
  INV_X1 U14882 ( .A(n14125), .ZN(n13887) );
  XNOR2_X1 U14883 ( .A(n14207), .B(n13887), .ZN(n13908) );
  XNOR2_X1 U14884 ( .A(n13911), .B(n13908), .ZN(n12494) );
  NAND2_X1 U14885 ( .A1(n12494), .A2(n14129), .ZN(n14208) );
  AND2_X1 U14886 ( .A1(n14124), .A2(n13787), .ZN(n12495) );
  AOI21_X1 U14887 ( .B1(n13889), .B2(n14126), .A(n12495), .ZN(n14204) );
  OAI211_X1 U14888 ( .C1(n15384), .C2(n13723), .A(n14208), .B(n14204), .ZN(
        n12506) );
  NAND2_X1 U14889 ( .A1(n12499), .A2(n13908), .ZN(n13888) );
  OAI21_X1 U14890 ( .B1(n12499), .B2(n13908), .A(n13888), .ZN(n14210) );
  AOI22_X1 U14891 ( .A1(n14207), .A2(n14038), .B1(n15394), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U14892 ( .A1(n12500), .A2(n14207), .ZN(n12501) );
  NAND2_X1 U14893 ( .A1(n12501), .A2(n8580), .ZN(n12502) );
  NOR2_X1 U14894 ( .A1(n14112), .A2(n12502), .ZN(n14205) );
  NAND2_X1 U14895 ( .A1(n14205), .A2(n14108), .ZN(n12503) );
  OAI211_X1 U14896 ( .C1(n14210), .C2(n14133), .A(n12504), .B(n12503), .ZN(
        n12505) );
  AOI21_X1 U14897 ( .B1(n15392), .B2(n12506), .A(n12505), .ZN(n12507) );
  INV_X1 U14898 ( .A(n12507), .ZN(P2_U3249) );
  NAND3_X1 U14899 ( .A1(n12508), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n12513) );
  NAND2_X1 U14900 ( .A1(n14237), .A2(n12509), .ZN(n12512) );
  NAND2_X1 U14901 ( .A1(n12510), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12511) );
  OAI211_X1 U14902 ( .C1(n12514), .C2(n12513), .A(n12512), .B(n12511), .ZN(
        P1_U3324) );
  OR2_X1 U14903 ( .A1(n13010), .A2(n13532), .ZN(n12518) );
  AND2_X1 U14904 ( .A1(n13144), .A2(n13503), .ZN(n12521) );
  OR2_X1 U14905 ( .A1(n13144), .A2(n13503), .ZN(n12520) );
  INV_X1 U14906 ( .A(n12522), .ZN(n12523) );
  OR2_X1 U14907 ( .A1(n13508), .A2(n12523), .ZN(n13467) );
  INV_X1 U14908 ( .A(n13589), .ZN(n13480) );
  AND2_X1 U14909 ( .A1(n13480), .A2(n13491), .ZN(n12525) );
  OR2_X1 U14910 ( .A1(n13467), .A2(n12525), .ZN(n13450) );
  OR2_X1 U14911 ( .A1(n13450), .A2(n13460), .ZN(n12527) );
  NAND2_X1 U14912 ( .A1(n13076), .A2(n13504), .ZN(n12524) );
  NAND2_X1 U14913 ( .A1(n13067), .A2(n13488), .ZN(n13485) );
  OR2_X1 U14914 ( .A1(n12523), .A2(n13485), .ZN(n13483) );
  AND2_X1 U14915 ( .A1(n12524), .A2(n13483), .ZN(n13468) );
  AND2_X1 U14916 ( .A1(n13477), .A2(n13468), .ZN(n13469) );
  OR2_X1 U14917 ( .A1(n12525), .A2(n13469), .ZN(n13451) );
  OR2_X1 U14918 ( .A1(n13460), .A2(n13451), .ZN(n12526) );
  INV_X1 U14919 ( .A(n13472), .ZN(n13438) );
  OR2_X1 U14920 ( .A1(n13644), .A2(n13438), .ZN(n12528) );
  NAND2_X1 U14921 ( .A1(n13638), .A2(n13454), .ZN(n12529) );
  NOR2_X1 U14922 ( .A1(n13107), .A2(n13423), .ZN(n12531) );
  INV_X1 U14923 ( .A(n13107), .ZN(n13631) );
  NAND2_X1 U14924 ( .A1(n13400), .A2(n13404), .ZN(n12533) );
  NAND2_X1 U14925 ( .A1(n13015), .A2(n13390), .ZN(n12532) );
  AND2_X1 U14926 ( .A1(n12602), .A2(n13371), .ZN(n12535) );
  NAND2_X1 U14927 ( .A1(n13623), .A2(n13402), .ZN(n12534) );
  OR2_X1 U14928 ( .A1(n13552), .A2(n13372), .ZN(n12536) );
  NAND2_X1 U14929 ( .A1(n13358), .A2(n12536), .ZN(n12538) );
  NAND2_X1 U14930 ( .A1(n13552), .A2(n13372), .ZN(n12537) );
  OR2_X1 U14931 ( .A1(n13352), .A2(n13359), .ZN(n12541) );
  XNOR2_X1 U14932 ( .A(n12542), .B(n12548), .ZN(n12547) );
  NAND2_X1 U14933 ( .A1(n12543), .A2(P3_B_REG_SCAN_IN), .ZN(n12544) );
  NAND2_X1 U14934 ( .A1(n15613), .A2(n12544), .ZN(n15027) );
  OAI22_X1 U14935 ( .A1(n12996), .A2(n15594), .B1(n12545), .B2(n15027), .ZN(
        n12546) );
  XNOR2_X1 U14936 ( .A(n12549), .B(n12548), .ZN(n13542) );
  AOI22_X1 U14937 ( .A1(n15030), .A2(n15622), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15627), .ZN(n12551) );
  NAND2_X1 U14938 ( .A1(n13606), .A2(n15033), .ZN(n12550) );
  OAI211_X1 U14939 ( .C1(n13542), .C2(n13539), .A(n12551), .B(n12550), .ZN(
        n12552) );
  INV_X1 U14940 ( .A(n12552), .ZN(n12553) );
  OAI21_X1 U14941 ( .B1(n13541), .B2(n15627), .A(n12553), .ZN(P3_U3204) );
  AOI21_X1 U14942 ( .B1(n12609), .B2(n15607), .A(n15599), .ZN(n12554) );
  OAI22_X1 U14943 ( .A1(n12555), .A2(n12554), .B1(n15595), .B2(n15597), .ZN(
        n12635) );
  AOI22_X1 U14944 ( .A1(n12635), .A2(n15625), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15622), .ZN(n12557) );
  NAND2_X1 U14945 ( .A1(n15033), .A2(n11366), .ZN(n12556) );
  OAI211_X1 U14946 ( .C1(n11540), .C2(n15625), .A(n12557), .B(n12556), .ZN(
        P3_U3233) );
  INV_X1 U14947 ( .A(n12558), .ZN(n12559) );
  OAI222_X1 U14948 ( .A1(P3_U3151), .A2(n12561), .B1(n12971), .B2(n12560), 
        .C1(n13672), .C2(n12559), .ZN(P3_U3267) );
  INV_X1 U14949 ( .A(n12562), .ZN(n12564) );
  NAND2_X1 U14950 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  XNOR2_X1 U14951 ( .A(n12598), .B(n13118), .ZN(n12567) );
  INV_X1 U14952 ( .A(n12567), .ZN(n12568) );
  NAND2_X1 U14953 ( .A1(n12569), .A2(n12568), .ZN(n12570) );
  XNOR2_X1 U14954 ( .A(n12598), .B(n12571), .ZN(n13047) );
  NAND2_X1 U14955 ( .A1(n13049), .A2(n13114), .ZN(n12572) );
  XNOR2_X1 U14956 ( .A(n15046), .B(n13030), .ZN(n12573) );
  NAND2_X1 U14957 ( .A1(n12573), .A2(n13005), .ZN(n13092) );
  INV_X1 U14958 ( .A(n12573), .ZN(n12574) );
  NAND2_X1 U14959 ( .A1(n12574), .A2(n13052), .ZN(n13093) );
  XNOR2_X1 U14960 ( .A(n13010), .B(n12598), .ZN(n12575) );
  XNOR2_X1 U14961 ( .A(n12575), .B(n13532), .ZN(n13001) );
  NAND2_X1 U14962 ( .A1(n12575), .A2(n13097), .ZN(n12576) );
  XNOR2_X1 U14963 ( .A(n13144), .B(n12598), .ZN(n12577) );
  XNOR2_X1 U14964 ( .A(n12577), .B(n13503), .ZN(n13146) );
  INV_X1 U14965 ( .A(n12577), .ZN(n12578) );
  NAND2_X1 U14966 ( .A1(n12578), .A2(n13503), .ZN(n12579) );
  XNOR2_X1 U14967 ( .A(n13067), .B(n12598), .ZN(n12580) );
  XNOR2_X1 U14968 ( .A(n12580), .B(n13488), .ZN(n13069) );
  INV_X1 U14969 ( .A(n12580), .ZN(n12581) );
  NAND2_X1 U14970 ( .A1(n12581), .A2(n13488), .ZN(n12582) );
  XNOR2_X1 U14971 ( .A(n13076), .B(n12598), .ZN(n12583) );
  XNOR2_X1 U14972 ( .A(n12583), .B(n13504), .ZN(n13078) );
  INV_X1 U14973 ( .A(n12583), .ZN(n12584) );
  NAND2_X1 U14974 ( .A1(n12584), .A2(n13504), .ZN(n12585) );
  XNOR2_X1 U14975 ( .A(n13589), .B(n12598), .ZN(n12586) );
  XNOR2_X1 U14976 ( .A(n12586), .B(n13491), .ZN(n13126) );
  NAND2_X1 U14977 ( .A1(n12586), .A2(n13491), .ZN(n12587) );
  XNOR2_X1 U14978 ( .A(n13644), .B(n12598), .ZN(n12589) );
  XNOR2_X1 U14979 ( .A(n12589), .B(n13472), .ZN(n13018) );
  NAND2_X1 U14980 ( .A1(n12589), .A2(n13472), .ZN(n12590) );
  XNOR2_X1 U14981 ( .A(n13638), .B(n12598), .ZN(n12591) );
  XNOR2_X1 U14982 ( .A(n12591), .B(n13454), .ZN(n13085) );
  INV_X1 U14983 ( .A(n12591), .ZN(n12592) );
  NAND2_X1 U14984 ( .A1(n12592), .A2(n13454), .ZN(n12593) );
  XNOR2_X1 U14985 ( .A(n13430), .B(n12598), .ZN(n12594) );
  XNOR2_X1 U14986 ( .A(n12594), .B(n13439), .ZN(n13041) );
  XNOR2_X1 U14987 ( .A(n13107), .B(n13030), .ZN(n12982) );
  INV_X1 U14988 ( .A(n12982), .ZN(n12977) );
  AND2_X1 U14989 ( .A1(n12979), .A2(n12977), .ZN(n12595) );
  AOI21_X2 U14990 ( .B1(n13103), .B2(n13403), .A(n12595), .ZN(n12597) );
  XNOR2_X1 U14991 ( .A(n13015), .B(n12598), .ZN(n12596) );
  INV_X1 U14992 ( .A(n12596), .ZN(n12980) );
  XNOR2_X1 U14993 ( .A(n12602), .B(n12598), .ZN(n12987) );
  AOI22_X1 U14994 ( .A1(n13391), .A2(n15492), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12600) );
  NAND2_X1 U14995 ( .A1(n13151), .A2(n13395), .ZN(n12599) );
  OAI211_X1 U14996 ( .C1(n13412), .C2(n13149), .A(n12600), .B(n12599), .ZN(
        n12601) );
  AOI21_X1 U14997 ( .B1(n12602), .B2(n15490), .A(n12601), .ZN(n12603) );
  INV_X1 U14998 ( .A(n14242), .ZN(n12604) );
  OAI222_X1 U14999 ( .A1(n14949), .A2(n12605), .B1(n12208), .B2(n12604), .C1(
        P1_U3086), .C2(n8555), .ZN(P1_U3327) );
  OAI222_X1 U15000 ( .A1(n14254), .A2(n12858), .B1(P2_U3088), .B2(n12606), 
        .C1(n12859), .C2(n14252), .ZN(P2_U3297) );
  NAND2_X1 U15001 ( .A1(n12607), .A2(n12610), .ZN(n12617) );
  NAND2_X1 U15002 ( .A1(n12609), .A2(n12608), .ZN(n12613) );
  NAND2_X1 U15003 ( .A1(n12611), .A2(n12610), .ZN(n12612) );
  NAND2_X1 U15004 ( .A1(n12613), .A2(n12612), .ZN(n12615) );
  NAND2_X1 U15005 ( .A1(n12615), .A2(n12614), .ZN(n12616) );
  INV_X1 U15006 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12618) );
  NOR2_X1 U15007 ( .A1(n15679), .A2(n12618), .ZN(n12619) );
  AOI21_X1 U15008 ( .B1(n15679), .B2(n12635), .A(n12619), .ZN(n12620) );
  OAI21_X1 U15009 ( .B1(n12637), .B2(n13657), .A(n12620), .ZN(P3_U3390) );
  OAI22_X1 U15010 ( .A1(n15607), .A2(n12621), .B1(n13325), .B2(n13540), .ZN(
        n12623) );
  NAND2_X1 U15011 ( .A1(n12623), .A2(n12622), .ZN(n12625) );
  NAND2_X1 U15012 ( .A1(n12625), .A2(n12624), .ZN(n12627) );
  NAND2_X1 U15013 ( .A1(n12627), .A2(n12626), .ZN(n12632) );
  NAND2_X1 U15014 ( .A1(n12629), .A2(n12628), .ZN(n12630) );
  NAND2_X1 U15015 ( .A1(n12630), .A2(n13659), .ZN(n12631) );
  AND2_X1 U15016 ( .A1(n15693), .A2(n15650), .ZN(n13582) );
  NOR2_X1 U15017 ( .A1(n15693), .A2(n11539), .ZN(n12634) );
  AOI21_X1 U15018 ( .B1(n12635), .B2(n15693), .A(n12634), .ZN(n12636) );
  OAI21_X1 U15019 ( .B1(n12637), .B2(n13604), .A(n12636), .ZN(P3_U3459) );
  OAI222_X1 U15020 ( .A1(n14949), .A2(n12639), .B1(P1_U3086), .B2(n12638), 
        .C1(n12208), .C2(n12858), .ZN(P1_U3325) );
  INV_X1 U15021 ( .A(n12640), .ZN(n12642) );
  OAI222_X1 U15022 ( .A1(n12971), .A2(n12643), .B1(n13672), .B2(n12642), .C1(
        P3_U3151), .C2(n12641), .ZN(P3_U3266) );
  OAI21_X1 U15023 ( .B1(n12647), .B2(n12674), .A(n8613), .ZN(n12650) );
  NAND2_X1 U15024 ( .A1(n12674), .A2(n12648), .ZN(n12649) );
  NAND2_X1 U15025 ( .A1(n12650), .A2(n12649), .ZN(n12653) );
  OAI211_X1 U15026 ( .C1(n15381), .C2(n12651), .A(n12674), .B(n10891), .ZN(
        n12652) );
  NAND2_X1 U15027 ( .A1(n12653), .A2(n12652), .ZN(n12660) );
  NAND2_X1 U15028 ( .A1(n12844), .A2(n13800), .ZN(n12656) );
  NAND2_X1 U15029 ( .A1(n12674), .A2(n12654), .ZN(n12655) );
  NAND2_X1 U15030 ( .A1(n12674), .A2(n13800), .ZN(n12657) );
  OAI21_X1 U15031 ( .B1(n7001), .B2(n12674), .A(n12657), .ZN(n12658) );
  NAND2_X1 U15032 ( .A1(n13799), .A2(n12844), .ZN(n12662) );
  NAND2_X1 U15033 ( .A1(n12663), .A2(n12674), .ZN(n12661) );
  NAND2_X1 U15034 ( .A1(n12663), .A2(n12844), .ZN(n12665) );
  NAND2_X1 U15035 ( .A1(n12674), .A2(n13799), .ZN(n12664) );
  NAND2_X1 U15036 ( .A1(n12665), .A2(n12664), .ZN(n12667) );
  NAND2_X1 U15037 ( .A1(n12668), .A2(n12667), .ZN(n12666) );
  INV_X1 U15038 ( .A(n12667), .ZN(n12670) );
  INV_X1 U15039 ( .A(n12668), .ZN(n12669) );
  NAND2_X1 U15040 ( .A1(n12670), .A2(n12669), .ZN(n12671) );
  NAND2_X1 U15041 ( .A1(n15410), .A2(n12787), .ZN(n12673) );
  NAND2_X1 U15042 ( .A1(n12825), .A2(n13798), .ZN(n12672) );
  NAND2_X1 U15043 ( .A1(n12673), .A2(n12672), .ZN(n12676) );
  AOI22_X1 U15044 ( .A1(n15410), .A2(n12825), .B1(n13798), .B2(n12787), .ZN(
        n12675) );
  NOR2_X1 U15045 ( .A1(n12677), .A2(n12676), .ZN(n12683) );
  NOR2_X1 U15046 ( .A1(n12787), .A2(n12678), .ZN(n12679) );
  AOI21_X1 U15047 ( .B1(n15417), .B2(n12787), .A(n12679), .ZN(n12686) );
  NAND2_X1 U15048 ( .A1(n15417), .A2(n12825), .ZN(n12681) );
  NAND2_X1 U15049 ( .A1(n12787), .A2(n13797), .ZN(n12680) );
  NAND2_X1 U15050 ( .A1(n12681), .A2(n12680), .ZN(n12685) );
  AND2_X1 U15051 ( .A1(n12686), .A2(n12685), .ZN(n12682) );
  INV_X1 U15052 ( .A(n12685), .ZN(n12688) );
  INV_X1 U15053 ( .A(n12686), .ZN(n12687) );
  NAND2_X1 U15054 ( .A1(n12688), .A2(n12687), .ZN(n12694) );
  INV_X1 U15055 ( .A(n12844), .ZN(n12702) );
  NAND2_X1 U15056 ( .A1(n15423), .A2(n12702), .ZN(n12690) );
  NAND2_X1 U15057 ( .A1(n12837), .A2(n13796), .ZN(n12689) );
  NAND2_X1 U15058 ( .A1(n15423), .A2(n12825), .ZN(n12691) );
  OAI21_X1 U15059 ( .B1(n12692), .B2(n12844), .A(n12691), .ZN(n12693) );
  NAND2_X1 U15060 ( .A1(n15429), .A2(n12825), .ZN(n12696) );
  NAND2_X1 U15061 ( .A1(n12702), .A2(n13795), .ZN(n12695) );
  NAND2_X1 U15062 ( .A1(n12696), .A2(n12695), .ZN(n12698) );
  AOI22_X1 U15063 ( .A1(n15429), .A2(n12702), .B1(n12837), .B2(n13795), .ZN(
        n12697) );
  AOI21_X1 U15064 ( .B1(n12699), .B2(n12698), .A(n12697), .ZN(n12701) );
  NOR2_X1 U15065 ( .A1(n12699), .A2(n12698), .ZN(n12700) );
  NAND2_X1 U15066 ( .A1(n15434), .A2(n12702), .ZN(n12704) );
  NAND2_X1 U15067 ( .A1(n12837), .A2(n13794), .ZN(n12703) );
  NAND2_X1 U15068 ( .A1(n12704), .A2(n12703), .ZN(n12710) );
  NAND2_X1 U15069 ( .A1(n12709), .A2(n12710), .ZN(n12708) );
  NAND2_X1 U15070 ( .A1(n15434), .A2(n12825), .ZN(n12705) );
  OAI21_X1 U15071 ( .B1(n12706), .B2(n12844), .A(n12705), .ZN(n12707) );
  NAND2_X1 U15072 ( .A1(n12708), .A2(n12707), .ZN(n12714) );
  INV_X1 U15073 ( .A(n12709), .ZN(n12712) );
  INV_X1 U15074 ( .A(n12710), .ZN(n12711) );
  NAND2_X1 U15075 ( .A1(n12712), .A2(n12711), .ZN(n12713) );
  NAND2_X1 U15076 ( .A1(n12714), .A2(n12713), .ZN(n12720) );
  NAND2_X1 U15077 ( .A1(n12717), .A2(n12825), .ZN(n12716) );
  NAND2_X1 U15078 ( .A1(n12702), .A2(n13793), .ZN(n12715) );
  NAND2_X1 U15079 ( .A1(n12716), .A2(n12715), .ZN(n12719) );
  AOI22_X1 U15080 ( .A1(n12717), .A2(n12702), .B1(n12837), .B2(n13793), .ZN(
        n12718) );
  AOI21_X1 U15081 ( .B1(n12720), .B2(n12719), .A(n12718), .ZN(n12722) );
  NOR2_X1 U15082 ( .A1(n12720), .A2(n12719), .ZN(n12721) );
  NAND2_X1 U15083 ( .A1(n15449), .A2(n12702), .ZN(n12724) );
  NAND2_X1 U15084 ( .A1(n12837), .A2(n13792), .ZN(n12723) );
  NAND2_X1 U15085 ( .A1(n15449), .A2(n12825), .ZN(n12725) );
  OAI21_X1 U15086 ( .B1(n12726), .B2(n12844), .A(n12725), .ZN(n12727) );
  NAND2_X1 U15087 ( .A1(n12731), .A2(n12837), .ZN(n12730) );
  NAND2_X1 U15088 ( .A1(n12702), .A2(n13791), .ZN(n12729) );
  NAND2_X1 U15089 ( .A1(n12730), .A2(n12729), .ZN(n12733) );
  AOI22_X1 U15090 ( .A1(n12731), .A2(n12702), .B1(n12837), .B2(n13791), .ZN(
        n12732) );
  NAND2_X1 U15091 ( .A1(n12736), .A2(n12702), .ZN(n12735) );
  NAND2_X1 U15092 ( .A1(n12837), .A2(n13790), .ZN(n12734) );
  NAND2_X1 U15093 ( .A1(n12735), .A2(n12734), .ZN(n12742) );
  NAND2_X1 U15094 ( .A1(n12741), .A2(n12742), .ZN(n12740) );
  NAND2_X1 U15095 ( .A1(n12736), .A2(n12837), .ZN(n12737) );
  OAI21_X1 U15096 ( .B1(n12738), .B2(n12844), .A(n12737), .ZN(n12739) );
  NAND2_X1 U15097 ( .A1(n12740), .A2(n12739), .ZN(n12746) );
  INV_X1 U15098 ( .A(n12741), .ZN(n12744) );
  INV_X1 U15099 ( .A(n12742), .ZN(n12743) );
  NAND2_X1 U15100 ( .A1(n12744), .A2(n12743), .ZN(n12745) );
  NAND2_X1 U15101 ( .A1(n12746), .A2(n12745), .ZN(n12752) );
  NAND2_X1 U15102 ( .A1(n12749), .A2(n12837), .ZN(n12748) );
  NAND2_X1 U15103 ( .A1(n12702), .A2(n13789), .ZN(n12747) );
  NAND2_X1 U15104 ( .A1(n12748), .A2(n12747), .ZN(n12751) );
  AOI22_X1 U15105 ( .A1(n12749), .A2(n12702), .B1(n12837), .B2(n13789), .ZN(
        n12750) );
  NAND2_X1 U15106 ( .A1(n12756), .A2(n12702), .ZN(n12754) );
  NAND2_X1 U15107 ( .A1(n12837), .A2(n12755), .ZN(n12753) );
  AOI22_X1 U15108 ( .A1(n12756), .A2(n12837), .B1(n12755), .B2(n12787), .ZN(
        n12757) );
  NAND2_X1 U15109 ( .A1(n12761), .A2(n12825), .ZN(n12760) );
  NAND2_X1 U15110 ( .A1(n12787), .A2(n13788), .ZN(n12759) );
  NAND2_X1 U15111 ( .A1(n12760), .A2(n12759), .ZN(n12766) );
  NAND2_X1 U15112 ( .A1(n12761), .A2(n12702), .ZN(n12763) );
  NAND2_X1 U15113 ( .A1(n12837), .A2(n13788), .ZN(n12762) );
  NAND2_X1 U15114 ( .A1(n12763), .A2(n12762), .ZN(n12764) );
  INV_X1 U15115 ( .A(n12766), .ZN(n12767) );
  NAND2_X1 U15116 ( .A1(n6773), .A2(n12767), .ZN(n12768) );
  NAND2_X1 U15117 ( .A1(n12771), .A2(n12787), .ZN(n12770) );
  NAND2_X1 U15118 ( .A1(n12837), .A2(n13787), .ZN(n12769) );
  AOI22_X1 U15119 ( .A1(n12771), .A2(n12837), .B1(n13787), .B2(n12702), .ZN(
        n12772) );
  INV_X1 U15120 ( .A(n12772), .ZN(n12773) );
  NAND2_X1 U15121 ( .A1(n14207), .A2(n12825), .ZN(n12775) );
  NAND2_X1 U15122 ( .A1(n14125), .A2(n12702), .ZN(n12774) );
  NAND2_X1 U15123 ( .A1(n12775), .A2(n12774), .ZN(n12777) );
  AOI22_X1 U15124 ( .A1(n14207), .A2(n12702), .B1(n12837), .B2(n14125), .ZN(
        n12776) );
  AND2_X1 U15125 ( .A1(n13889), .A2(n12837), .ZN(n12778) );
  AOI21_X1 U15126 ( .B1(n14200), .B2(n12702), .A(n12778), .ZN(n12781) );
  INV_X1 U15127 ( .A(n13889), .ZN(n14091) );
  NAND2_X1 U15128 ( .A1(n14200), .A2(n12837), .ZN(n12779) );
  OAI21_X1 U15129 ( .B1(n14091), .B2(n12844), .A(n12779), .ZN(n12780) );
  OAI21_X1 U15130 ( .B1(n12782), .B2(n12781), .A(n12780), .ZN(n12784) );
  NAND2_X1 U15131 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  AND2_X1 U15132 ( .A1(n14127), .A2(n12702), .ZN(n12785) );
  AOI21_X1 U15133 ( .B1(n14195), .B2(n12837), .A(n12785), .ZN(n12789) );
  INV_X1 U15134 ( .A(n14127), .ZN(n13913) );
  NAND2_X1 U15135 ( .A1(n14195), .A2(n12702), .ZN(n12786) );
  OAI21_X1 U15136 ( .B1(n13913), .B2(n12787), .A(n12786), .ZN(n12788) );
  NAND2_X1 U15137 ( .A1(n14191), .A2(n12787), .ZN(n12791) );
  NAND2_X1 U15138 ( .A1(n13892), .A2(n12837), .ZN(n12790) );
  AOI22_X1 U15139 ( .A1(n14191), .A2(n12837), .B1(n13892), .B2(n12702), .ZN(
        n12792) );
  NAND2_X1 U15140 ( .A1(n14185), .A2(n12837), .ZN(n12794) );
  NAND2_X1 U15141 ( .A1(n13914), .A2(n12787), .ZN(n12793) );
  NAND2_X1 U15142 ( .A1(n12794), .A2(n12793), .ZN(n12796) );
  AOI22_X1 U15143 ( .A1(n14185), .A2(n12702), .B1(n12837), .B2(n13914), .ZN(
        n12795) );
  AOI21_X1 U15144 ( .B1(n12797), .B2(n12796), .A(n12795), .ZN(n12799) );
  NOR2_X1 U15145 ( .A1(n12797), .A2(n12796), .ZN(n12798) );
  NAND2_X1 U15146 ( .A1(n14180), .A2(n12787), .ZN(n12801) );
  NAND2_X1 U15147 ( .A1(n14031), .A2(n12825), .ZN(n12800) );
  NAND2_X1 U15148 ( .A1(n12801), .A2(n12800), .ZN(n12805) );
  NAND2_X1 U15149 ( .A1(n14180), .A2(n12837), .ZN(n12802) );
  OAI21_X1 U15150 ( .B1(n7047), .B2(n12844), .A(n12802), .ZN(n12803) );
  NAND2_X1 U15151 ( .A1(n14175), .A2(n12837), .ZN(n12807) );
  NAND2_X1 U15152 ( .A1(n12787), .A2(n13915), .ZN(n12806) );
  NAND2_X1 U15153 ( .A1(n12807), .A2(n12806), .ZN(n12809) );
  AOI22_X1 U15154 ( .A1(n14175), .A2(n12702), .B1(n12837), .B2(n13915), .ZN(
        n12808) );
  NAND2_X1 U15155 ( .A1(n14170), .A2(n12702), .ZN(n12811) );
  NAND2_X1 U15156 ( .A1(n12837), .A2(n14030), .ZN(n12810) );
  NAND2_X1 U15157 ( .A1(n12811), .A2(n12810), .ZN(n12814) );
  NAND2_X1 U15158 ( .A1(n14170), .A2(n12837), .ZN(n12813) );
  NAND2_X1 U15159 ( .A1(n12787), .A2(n14030), .ZN(n12812) );
  NAND2_X1 U15160 ( .A1(n14165), .A2(n12825), .ZN(n12816) );
  NAND2_X1 U15161 ( .A1(n12674), .A2(n13920), .ZN(n12815) );
  NAND2_X1 U15162 ( .A1(n12816), .A2(n12815), .ZN(n12819) );
  INV_X1 U15163 ( .A(n13920), .ZN(n13712) );
  NOR2_X1 U15164 ( .A1(n12674), .A2(n13712), .ZN(n12817) );
  AOI21_X1 U15165 ( .B1(n14165), .B2(n12674), .A(n12817), .ZN(n12818) );
  NOR2_X1 U15166 ( .A1(n12820), .A2(n12819), .ZN(n12821) );
  NAND2_X1 U15167 ( .A1(n14159), .A2(n12787), .ZN(n12824) );
  NAND2_X1 U15168 ( .A1(n12837), .A2(n13898), .ZN(n12823) );
  NAND2_X1 U15169 ( .A1(n14159), .A2(n12825), .ZN(n12827) );
  NAND2_X1 U15170 ( .A1(n12787), .A2(n13898), .ZN(n12826) );
  NAND2_X1 U15171 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  INV_X1 U15172 ( .A(n12833), .ZN(n12836) );
  NAND2_X1 U15173 ( .A1(n14154), .A2(n12837), .ZN(n12830) );
  NAND2_X1 U15174 ( .A1(n12674), .A2(n13960), .ZN(n12829) );
  NAND2_X1 U15175 ( .A1(n12830), .A2(n12829), .ZN(n12832) );
  INV_X1 U15176 ( .A(n12832), .ZN(n12835) );
  AOI22_X1 U15177 ( .A1(n14154), .A2(n12674), .B1(n12825), .B2(n13960), .ZN(
        n12831) );
  AOI21_X1 U15178 ( .B1(n12833), .B2(n12832), .A(n12831), .ZN(n12834) );
  AOI22_X1 U15179 ( .A1(n14149), .A2(n12674), .B1(n12837), .B2(n13942), .ZN(
        n12838) );
  AOI22_X1 U15180 ( .A1(n14149), .A2(n12837), .B1(n13942), .B2(n12674), .ZN(
        n12839) );
  INV_X1 U15181 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U15182 ( .A1(n12883), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12842) );
  NAND2_X1 U15183 ( .A1(n12840), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12841) );
  OAI211_X1 U15184 ( .C1(n12866), .C2(n12843), .A(n12842), .B(n12841), .ZN(
        n13879) );
  NAND2_X1 U15185 ( .A1(n12702), .A2(n13879), .ZN(n12874) );
  NAND2_X1 U15186 ( .A1(n12874), .A2(n12674), .ZN(n12848) );
  NAND2_X1 U15187 ( .A1(n12844), .A2(n13879), .ZN(n12847) );
  NOR2_X1 U15188 ( .A1(n12879), .A2(n10585), .ZN(n12845) );
  AOI21_X2 U15189 ( .B1(n14237), .B2(n6675), .A(n12845), .ZN(n14135) );
  MUX2_X1 U15190 ( .A(n12848), .B(n12847), .S(n14135), .Z(n12946) );
  NAND2_X1 U15191 ( .A1(n12925), .A2(n13871), .ZN(n12849) );
  NAND4_X1 U15192 ( .A1(n12644), .A2(n12946), .A3(n12850), .A4(n12849), .ZN(
        n12942) );
  NAND2_X1 U15193 ( .A1(n14242), .A2(n6675), .ZN(n12852) );
  OR2_X1 U15194 ( .A1(n12879), .A2(n14245), .ZN(n12851) );
  AND2_X1 U15195 ( .A1(n12787), .A2(n13959), .ZN(n12853) );
  AOI21_X1 U15196 ( .B1(n14145), .B2(n12837), .A(n12853), .ZN(n12933) );
  NAND2_X1 U15197 ( .A1(n14145), .A2(n12674), .ZN(n12855) );
  NAND2_X1 U15198 ( .A1(n12837), .A2(n13959), .ZN(n12854) );
  NAND2_X1 U15199 ( .A1(n12855), .A2(n12854), .ZN(n12932) );
  INV_X1 U15200 ( .A(n14135), .ZN(n12856) );
  OR2_X1 U15201 ( .A1(n12858), .A2(n12857), .ZN(n12861) );
  OR2_X1 U15202 ( .A1(n12879), .A2(n12859), .ZN(n12860) );
  NOR2_X1 U15203 ( .A1(n12863), .A2(n12862), .ZN(n12864) );
  NAND2_X1 U15204 ( .A1(n12961), .A2(n15385), .ZN(n12929) );
  AND2_X1 U15205 ( .A1(n12864), .A2(n12929), .ZN(n12873) );
  INV_X1 U15206 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n12865) );
  OR2_X1 U15207 ( .A1(n12866), .A2(n12865), .ZN(n12872) );
  INV_X1 U15208 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12867) );
  OR2_X1 U15209 ( .A1(n12868), .A2(n12867), .ZN(n12871) );
  INV_X1 U15210 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n12869) );
  OR2_X1 U15211 ( .A1(n12885), .A2(n12869), .ZN(n12870) );
  AND3_X1 U15212 ( .A1(n12872), .A2(n12871), .A3(n12870), .ZN(n12876) );
  AOI21_X1 U15213 ( .B1(n12874), .B2(n12873), .A(n12876), .ZN(n12875) );
  AOI21_X1 U15214 ( .B1(n13876), .B2(n12825), .A(n12875), .ZN(n12939) );
  NAND2_X1 U15215 ( .A1(n13876), .A2(n12674), .ZN(n12878) );
  INV_X1 U15216 ( .A(n12876), .ZN(n13930) );
  NAND2_X1 U15217 ( .A1(n12837), .A2(n13930), .ZN(n12877) );
  NAND2_X1 U15218 ( .A1(n12878), .A2(n12877), .ZN(n12938) );
  NAND2_X1 U15219 ( .A1(n14239), .A2(n6675), .ZN(n12881) );
  OR2_X1 U15220 ( .A1(n12879), .A2(n14240), .ZN(n12880) );
  NAND2_X1 U15221 ( .A1(n12882), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n12889) );
  NAND2_X1 U15222 ( .A1(n12883), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12888) );
  OR2_X1 U15223 ( .A1(n8721), .A2(n13905), .ZN(n12887) );
  INV_X1 U15224 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n12884) );
  OR2_X1 U15225 ( .A1(n12885), .A2(n12884), .ZN(n12886) );
  NAND4_X1 U15226 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        n13943) );
  AND2_X1 U15227 ( .A1(n12787), .A2(n13943), .ZN(n12890) );
  AOI21_X1 U15228 ( .B1(n14140), .B2(n12837), .A(n12890), .ZN(n12935) );
  NAND2_X1 U15229 ( .A1(n14140), .A2(n12787), .ZN(n12892) );
  NAND2_X1 U15230 ( .A1(n12837), .A2(n13943), .ZN(n12891) );
  NAND2_X1 U15231 ( .A1(n12892), .A2(n12891), .ZN(n12934) );
  OAI22_X1 U15232 ( .A1(n12939), .A2(n12938), .B1(n12935), .B2(n12934), .ZN(
        n12893) );
  OAI21_X1 U15233 ( .B1(n12933), .B2(n12932), .A(n12940), .ZN(n12948) );
  NOR3_X1 U15234 ( .A1(n12941), .A2(n12942), .A3(n12948), .ZN(n12965) );
  XNOR2_X1 U15235 ( .A(n13876), .B(n13930), .ZN(n12924) );
  NAND2_X1 U15236 ( .A1(n14145), .A2(n13903), .ZN(n12894) );
  NAND2_X1 U15237 ( .A1(n13927), .A2(n12894), .ZN(n13902) );
  OR2_X1 U15238 ( .A1(n14154), .A2(n13900), .ZN(n13923) );
  NAND2_X1 U15239 ( .A1(n14154), .A2(n13900), .ZN(n13924) );
  NAND2_X1 U15240 ( .A1(n13923), .A2(n13924), .ZN(n13976) );
  INV_X1 U15241 ( .A(n13898), .ZN(n13922) );
  XNOR2_X1 U15242 ( .A(n14159), .B(n13922), .ZN(n13985) );
  XNOR2_X1 U15243 ( .A(n14165), .B(n13712), .ZN(n13998) );
  OR2_X1 U15244 ( .A1(n14170), .A2(n14030), .ZN(n13896) );
  NAND2_X1 U15245 ( .A1(n14170), .A2(n14030), .ZN(n13895) );
  NAND2_X1 U15246 ( .A1(n13896), .A2(n13895), .ZN(n14022) );
  INV_X1 U15247 ( .A(n13914), .ZN(n13893) );
  XNOR2_X1 U15248 ( .A(n14185), .B(n13893), .ZN(n14068) );
  XNOR2_X1 U15249 ( .A(n14191), .B(n14092), .ZN(n14074) );
  XNOR2_X1 U15250 ( .A(n14195), .B(n13913), .ZN(n14093) );
  NAND2_X1 U15251 ( .A1(n12896), .A2(n12895), .ZN(n15405) );
  NOR2_X1 U15252 ( .A1(n15405), .A2(n12897), .ZN(n12898) );
  NAND4_X1 U15253 ( .A1(n12901), .A2(n12900), .A3(n12899), .A4(n12898), .ZN(
        n12902) );
  NOR2_X1 U15254 ( .A1(n12903), .A2(n12902), .ZN(n12905) );
  NAND4_X1 U15255 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12908) );
  OR4_X1 U15256 ( .A1(n12915), .A2(n12914), .A3(n12913), .A4(n12912), .ZN(
        n12918) );
  NAND2_X1 U15257 ( .A1(n14200), .A2(n14091), .ZN(n13912) );
  OR2_X1 U15258 ( .A1(n14200), .A2(n14091), .ZN(n12916) );
  NAND2_X1 U15259 ( .A1(n13912), .A2(n12916), .ZN(n14110) );
  OR4_X1 U15260 ( .A1(n12918), .A2(n14110), .A3(n12917), .A4(n13908), .ZN(
        n12919) );
  NOR2_X1 U15261 ( .A1(n14068), .A2(n12921), .ZN(n12922) );
  XNOR2_X1 U15262 ( .A(n14180), .B(n14031), .ZN(n14054) );
  XNOR2_X1 U15263 ( .A(n14175), .B(n13915), .ZN(n13917) );
  NAND4_X1 U15264 ( .A1(n14022), .A2(n12922), .A3(n14054), .A4(n13917), .ZN(
        n12923) );
  XNOR2_X1 U15265 ( .A(n14140), .B(n13943), .ZN(n13928) );
  XNOR2_X1 U15266 ( .A(n14149), .B(n13942), .ZN(n13957) );
  AOI21_X1 U15267 ( .B1(n12927), .B2(n12926), .A(n12925), .ZN(n12957) );
  INV_X1 U15268 ( .A(n12927), .ZN(n12928) );
  NAND2_X1 U15269 ( .A1(n12928), .A2(n13871), .ZN(n12954) );
  OAI21_X1 U15270 ( .B1(n12930), .B2(n13871), .A(n12929), .ZN(n12931) );
  AOI21_X1 U15271 ( .B1(n12957), .B2(n12954), .A(n12931), .ZN(n12945) );
  AOI22_X1 U15272 ( .A1(n12935), .A2(n12934), .B1(n12933), .B2(n12932), .ZN(
        n12936) );
  INV_X1 U15273 ( .A(n12942), .ZN(n12944) );
  AOI21_X1 U15274 ( .B1(n12944), .B2(n12943), .A(n12960), .ZN(n12952) );
  INV_X1 U15275 ( .A(n12946), .ZN(n12947) );
  AOI21_X1 U15276 ( .B1(n12949), .B2(n12948), .A(n12947), .ZN(n12950) );
  INV_X1 U15277 ( .A(n12960), .ZN(n12956) );
  INV_X1 U15278 ( .A(n15385), .ZN(n12955) );
  NAND4_X1 U15279 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12963) );
  NAND2_X1 U15280 ( .A1(n13878), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14247) );
  OR3_X1 U15281 ( .A1(n12958), .A2(n14090), .A3(n14247), .ZN(n12959) );
  OAI211_X1 U15282 ( .C1(n12961), .C2(n12960), .A(n12959), .B(P2_B_REG_SCAN_IN), .ZN(n12962) );
  OAI211_X1 U15283 ( .C1(n12965), .C2(n12964), .A(n12963), .B(n12962), .ZN(
        P2_U3328) );
  OAI222_X1 U15284 ( .A1(n14252), .A2(n12967), .B1(n14254), .B2(n12966), .C1(
        n13871), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U15285 ( .A(n12968), .ZN(n12969) );
  INV_X1 U15286 ( .A(n12972), .ZN(n12974) );
  INV_X1 U15287 ( .A(SI_30_), .ZN(n12973) );
  XNOR2_X1 U15288 ( .A(n13352), .B(n13030), .ZN(n13026) );
  XNOR2_X1 U15289 ( .A(n13026), .B(n13139), .ZN(n13028) );
  INV_X1 U15290 ( .A(n12987), .ZN(n12976) );
  AOI22_X1 U15291 ( .A1(n12976), .A2(n13371), .B1(n12980), .B2(n13390), .ZN(
        n12981) );
  OAI21_X1 U15292 ( .B1(n12980), .B2(n13390), .A(n13371), .ZN(n12986) );
  NOR3_X1 U15293 ( .A1(n12980), .A2(n13390), .A3(n13371), .ZN(n12985) );
  INV_X1 U15294 ( .A(n12981), .ZN(n12983) );
  NOR3_X1 U15295 ( .A1(n12983), .A2(n12982), .A3(n13423), .ZN(n12984) );
  AOI211_X1 U15296 ( .C1(n12987), .C2(n12986), .A(n12985), .B(n12984), .ZN(
        n12988) );
  XNOR2_X1 U15297 ( .A(n13378), .B(n13030), .ZN(n12990) );
  XNOR2_X1 U15298 ( .A(n12990), .B(n12992), .ZN(n13061) );
  INV_X1 U15299 ( .A(n12990), .ZN(n12991) );
  XNOR2_X1 U15300 ( .A(n13552), .B(n13030), .ZN(n12993) );
  XNOR2_X1 U15301 ( .A(n12993), .B(n13372), .ZN(n13133) );
  XOR2_X1 U15302 ( .A(n13028), .B(n13029), .Z(n12999) );
  AOI22_X1 U15303 ( .A1(n13372), .A2(n13134), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12995) );
  NAND2_X1 U15304 ( .A1(n13353), .A2(n13135), .ZN(n12994) );
  OAI211_X1 U15305 ( .C1(n12996), .C2(n13138), .A(n12995), .B(n12994), .ZN(
        n12997) );
  AOI21_X1 U15306 ( .B1(n13352), .B2(n15490), .A(n12997), .ZN(n12998) );
  OAI21_X1 U15307 ( .B1(n12999), .B2(n13142), .A(n12998), .ZN(P3_U3154) );
  OAI211_X1 U15308 ( .C1(n13002), .C2(n13001), .A(n13000), .B(n15494), .ZN(
        n13009) );
  NOR2_X1 U15309 ( .A1(n13003), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13208) );
  AOI21_X1 U15310 ( .B1(n15492), .B2(n13503), .A(n13208), .ZN(n13004) );
  OAI21_X1 U15311 ( .B1(n13149), .B2(n13005), .A(n13004), .ZN(n13006) );
  AOI21_X1 U15312 ( .B1(n13007), .B2(n13135), .A(n13006), .ZN(n13008) );
  OAI211_X1 U15313 ( .C1(n13154), .C2(n13010), .A(n13009), .B(n13008), .ZN(
        P3_U3155) );
  XNOR2_X1 U15314 ( .A(n13011), .B(n13412), .ZN(n13017) );
  AOI22_X1 U15315 ( .A1(n13371), .A2(n15492), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13013) );
  NAND2_X1 U15316 ( .A1(n13135), .A2(n13406), .ZN(n13012) );
  OAI211_X1 U15317 ( .C1(n13403), .C2(n13149), .A(n13013), .B(n13012), .ZN(
        n13014) );
  AOI21_X1 U15318 ( .B1(n13015), .B2(n15490), .A(n13014), .ZN(n13016) );
  OAI21_X1 U15319 ( .B1(n13017), .B2(n13142), .A(n13016), .ZN(P3_U3156) );
  AOI21_X1 U15320 ( .B1(n13019), .B2(n13018), .A(n13142), .ZN(n13021) );
  NAND2_X1 U15321 ( .A1(n13021), .A2(n13020), .ZN(n13025) );
  AND2_X1 U15322 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13326) );
  AOI21_X1 U15323 ( .B1(n15492), .B2(n13454), .A(n13326), .ZN(n13022) );
  OAI21_X1 U15324 ( .B1(n13149), .B2(n13491), .A(n13022), .ZN(n13023) );
  AOI21_X1 U15325 ( .B1(n13463), .B2(n13151), .A(n13023), .ZN(n13024) );
  OAI211_X1 U15326 ( .C1(n13154), .C2(n13644), .A(n13025), .B(n13024), .ZN(
        P3_U3159) );
  INV_X1 U15327 ( .A(n13026), .ZN(n13027) );
  XNOR2_X1 U15328 ( .A(n13328), .B(n13030), .ZN(n13031) );
  XNOR2_X1 U15329 ( .A(n13032), .B(n13031), .ZN(n13039) );
  NOR2_X1 U15330 ( .A1(n13033), .A2(n13138), .ZN(n13036) );
  OAI22_X1 U15331 ( .A1(n13139), .A2(n13149), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13034), .ZN(n13035) );
  AOI211_X1 U15332 ( .C1(n13135), .C2(n13337), .A(n13036), .B(n13035), .ZN(
        n13038) );
  NAND2_X1 U15333 ( .A1(n12515), .A2(n15490), .ZN(n13037) );
  AOI21_X1 U15334 ( .B1(n13041), .B2(n13040), .A(n6757), .ZN(n13046) );
  INV_X1 U15335 ( .A(n13454), .ZN(n13425) );
  NAND2_X1 U15336 ( .A1(n13151), .A2(n13431), .ZN(n13043) );
  AOI22_X1 U15337 ( .A1(n15492), .A2(n13423), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13042) );
  OAI211_X1 U15338 ( .C1(n13425), .C2(n13149), .A(n13043), .B(n13042), .ZN(
        n13044) );
  AOI21_X1 U15339 ( .B1(n13430), .B2(n15490), .A(n13044), .ZN(n13045) );
  OAI21_X1 U15340 ( .B1(n13046), .B2(n13142), .A(n13045), .ZN(P3_U3163) );
  XNOR2_X1 U15341 ( .A(n13047), .B(n13531), .ZN(n13048) );
  XNOR2_X1 U15342 ( .A(n13049), .B(n13048), .ZN(n13059) );
  NAND2_X1 U15343 ( .A1(n13151), .A2(n13050), .ZN(n13054) );
  INV_X1 U15344 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13051) );
  NOR2_X1 U15345 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13051), .ZN(n15537) );
  AOI21_X1 U15346 ( .B1(n15492), .B2(n13052), .A(n15537), .ZN(n13053) );
  OAI211_X1 U15347 ( .C1(n13055), .C2(n13149), .A(n13054), .B(n13053), .ZN(
        n13056) );
  AOI21_X1 U15348 ( .B1(n13057), .B2(n15490), .A(n13056), .ZN(n13058) );
  OAI21_X1 U15349 ( .B1(n13059), .B2(n13142), .A(n13058), .ZN(P3_U3164) );
  XOR2_X1 U15350 ( .A(n13061), .B(n13060), .Z(n13066) );
  AOI22_X1 U15351 ( .A1(n13372), .A2(n15492), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13063) );
  NAND2_X1 U15352 ( .A1(n13135), .A2(n13379), .ZN(n13062) );
  OAI211_X1 U15353 ( .C1(n13402), .C2(n13149), .A(n13063), .B(n13062), .ZN(
        n13064) );
  AOI21_X1 U15354 ( .B1(n13378), .B2(n15490), .A(n13064), .ZN(n13065) );
  OAI21_X1 U15355 ( .B1(n13066), .B2(n13142), .A(n13065), .ZN(P3_U3165) );
  INV_X1 U15356 ( .A(n13067), .ZN(n13653) );
  OAI211_X1 U15357 ( .C1(n13070), .C2(n13069), .A(n13068), .B(n15494), .ZN(
        n13075) );
  NAND2_X1 U15358 ( .A1(n15492), .A2(n13504), .ZN(n13071) );
  NAND2_X1 U15359 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13242)
         );
  OAI211_X1 U15360 ( .C1(n13149), .C2(n13072), .A(n13071), .B(n13242), .ZN(
        n13073) );
  AOI21_X1 U15361 ( .B1(n13510), .B2(n13135), .A(n13073), .ZN(n13074) );
  OAI211_X1 U15362 ( .C1(n13653), .C2(n13154), .A(n13075), .B(n13074), .ZN(
        P3_U3166) );
  INV_X1 U15363 ( .A(n13076), .ZN(n13649) );
  OAI211_X1 U15364 ( .C1(n13079), .C2(n13078), .A(n13077), .B(n15494), .ZN(
        n13083) );
  NAND2_X1 U15365 ( .A1(n13134), .A2(n13488), .ZN(n13080) );
  NAND2_X1 U15366 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13274)
         );
  OAI211_X1 U15367 ( .C1(n13491), .C2(n13138), .A(n13080), .B(n13274), .ZN(
        n13081) );
  AOI21_X1 U15368 ( .B1(n13494), .B2(n13135), .A(n13081), .ZN(n13082) );
  OAI211_X1 U15369 ( .C1(n13649), .C2(n13154), .A(n13083), .B(n13082), .ZN(
        P3_U3168) );
  OAI211_X1 U15370 ( .C1(n13086), .C2(n13085), .A(n13084), .B(n15494), .ZN(
        n13091) );
  AOI22_X1 U15371 ( .A1(n15492), .A2(n13087), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13088) );
  OAI21_X1 U15372 ( .B1(n13438), .B2(n13149), .A(n13088), .ZN(n13089) );
  AOI21_X1 U15373 ( .B1(n13445), .B2(n13135), .A(n13089), .ZN(n13090) );
  OAI211_X1 U15374 ( .C1(n13447), .C2(n13154), .A(n13091), .B(n13090), .ZN(
        P3_U3173) );
  NAND2_X1 U15375 ( .A1(n13093), .A2(n13092), .ZN(n13095) );
  XOR2_X1 U15376 ( .A(n13095), .B(n13094), .Z(n13102) );
  INV_X1 U15377 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n13096) );
  NOR2_X1 U15378 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13096), .ZN(n13186) );
  AOI21_X1 U15379 ( .B1(n15492), .B2(n13097), .A(n13186), .ZN(n13098) );
  OAI21_X1 U15380 ( .B1(n13149), .B2(n13531), .A(n13098), .ZN(n13100) );
  NOR2_X1 U15381 ( .A1(n15046), .A2(n13154), .ZN(n13099) );
  AOI211_X1 U15382 ( .C1(n13533), .C2(n13151), .A(n13100), .B(n13099), .ZN(
        n13101) );
  OAI21_X1 U15383 ( .B1(n13102), .B2(n13142), .A(n13101), .ZN(P3_U3174) );
  XNOR2_X1 U15384 ( .A(n13103), .B(n13423), .ZN(n13109) );
  NAND2_X1 U15385 ( .A1(n13135), .A2(n13417), .ZN(n13105) );
  AOI22_X1 U15386 ( .A1(n13390), .A2(n15492), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13104) );
  OAI211_X1 U15387 ( .C1(n13439), .C2(n13149), .A(n13105), .B(n13104), .ZN(
        n13106) );
  AOI21_X1 U15388 ( .B1(n13107), .B2(n15490), .A(n13106), .ZN(n13108) );
  OAI21_X1 U15389 ( .B1(n13109), .B2(n13142), .A(n13108), .ZN(P3_U3175) );
  OAI211_X1 U15390 ( .C1(n13112), .C2(n13111), .A(n13110), .B(n15494), .ZN(
        n13120) );
  AOI21_X1 U15391 ( .B1(n15492), .B2(n13114), .A(n13113), .ZN(n13115) );
  OAI21_X1 U15392 ( .B1(n13149), .B2(n13116), .A(n13115), .ZN(n13117) );
  AOI21_X1 U15393 ( .B1(n13118), .B2(n15490), .A(n13117), .ZN(n13119) );
  OAI211_X1 U15394 ( .C1(n13122), .C2(n13121), .A(n13120), .B(n13119), .ZN(
        P3_U3176) );
  INV_X1 U15395 ( .A(n13123), .ZN(n13124) );
  AOI21_X1 U15396 ( .B1(n13126), .B2(n13125), .A(n13124), .ZN(n13132) );
  NAND2_X1 U15397 ( .A1(n15492), .A2(n13472), .ZN(n13127) );
  NAND2_X1 U15398 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13297)
         );
  OAI211_X1 U15399 ( .C1(n13149), .C2(n13128), .A(n13127), .B(n13297), .ZN(
        n13130) );
  NOR2_X1 U15400 ( .A1(n13480), .A2(n13154), .ZN(n13129) );
  AOI211_X1 U15401 ( .C1(n13478), .C2(n13151), .A(n13130), .B(n13129), .ZN(
        n13131) );
  OAI21_X1 U15402 ( .B1(n13132), .B2(n13142), .A(n13131), .ZN(P3_U3178) );
  AOI22_X1 U15403 ( .A1(n13391), .A2(n13134), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13137) );
  NAND2_X1 U15404 ( .A1(n13135), .A2(n13363), .ZN(n13136) );
  OAI211_X1 U15405 ( .C1(n13139), .C2(n13138), .A(n13137), .B(n13136), .ZN(
        n13140) );
  AOI21_X1 U15406 ( .B1(n13552), .B2(n15490), .A(n13140), .ZN(n13141) );
  OAI21_X1 U15407 ( .B1(n13143), .B2(n13142), .A(n13141), .ZN(P3_U3180) );
  INV_X1 U15408 ( .A(n13144), .ZN(n13658) );
  OAI211_X1 U15409 ( .C1(n13147), .C2(n13146), .A(n13145), .B(n15494), .ZN(
        n13153) );
  AND2_X1 U15410 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n15024) );
  AOI21_X1 U15411 ( .B1(n15492), .B2(n13488), .A(n15024), .ZN(n13148) );
  OAI21_X1 U15412 ( .B1(n13149), .B2(n13532), .A(n13148), .ZN(n13150) );
  AOI21_X1 U15413 ( .B1(n13520), .B2(n13151), .A(n13150), .ZN(n13152) );
  OAI211_X1 U15414 ( .C1(n13658), .C2(n13154), .A(n13153), .B(n13152), .ZN(
        P3_U3181) );
  MUX2_X1 U15415 ( .A(n15029), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13155), .Z(
        P3_U3522) );
  NAND2_X1 U15416 ( .A1(n15503), .A2(n13156), .ZN(n13172) );
  NAND2_X1 U15417 ( .A1(n13157), .A2(n15511), .ZN(n13158) );
  AND2_X1 U15418 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  OAI22_X1 U15419 ( .A1(n15520), .A2(n13160), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11378), .ZN(n13161) );
  AOI21_X1 U15420 ( .B1(n15538), .B2(P3_ADDR_REG_1__SCAN_IN), .A(n13161), .ZN(
        n13171) );
  NAND2_X1 U15421 ( .A1(n13162), .A2(n11535), .ZN(n13163) );
  NAND2_X1 U15422 ( .A1(n13164), .A2(n13163), .ZN(n13165) );
  NAND2_X1 U15423 ( .A1(n15539), .A2(n13165), .ZN(n13170) );
  OAI21_X1 U15424 ( .B1(n13167), .B2(P3_REG1_REG_1__SCAN_IN), .A(n13166), .ZN(
        n13168) );
  NAND2_X1 U15425 ( .A1(n15500), .A2(n13168), .ZN(n13169) );
  NAND4_X1 U15426 ( .A1(n13172), .A2(n13171), .A3(n13170), .A4(n13169), .ZN(
        P3_U3183) );
  INV_X1 U15427 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13177) );
  NOR2_X1 U15428 ( .A1(n13190), .A2(n13173), .ZN(n13175) );
  INV_X1 U15429 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13178) );
  MUX2_X1 U15430 ( .A(n13178), .B(P3_REG2_REG_12__SCAN_IN), .S(n15534), .Z(
        n15540) );
  AOI21_X1 U15431 ( .B1(n13177), .B2(n13176), .A(n13205), .ZN(n13199) );
  MUX2_X1 U15432 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13268), .Z(n13210) );
  XNOR2_X1 U15433 ( .A(n13210), .B(n13209), .ZN(n13185) );
  MUX2_X1 U15434 ( .A(n13178), .B(n15055), .S(n13268), .Z(n13180) );
  INV_X1 U15435 ( .A(n13180), .ZN(n13179) );
  NAND2_X1 U15436 ( .A1(n13179), .A2(n15534), .ZN(n13183) );
  XNOR2_X1 U15437 ( .A(n13180), .B(n15534), .ZN(n15551) );
  AOI21_X1 U15438 ( .B1(n13182), .B2(n13190), .A(n13181), .ZN(n15552) );
  AOI21_X1 U15439 ( .B1(n13185), .B2(n13184), .A(n13213), .ZN(n13188) );
  AOI21_X1 U15440 ( .B1(n15538), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13186), 
        .ZN(n13187) );
  OAI21_X1 U15441 ( .B1(n13188), .B2(n15520), .A(n13187), .ZN(n13197) );
  NOR2_X1 U15442 ( .A1(n13189), .A2(n13190), .ZN(n13192) );
  MUX2_X1 U15443 ( .A(n15055), .B(P3_REG1_REG_12__SCAN_IN), .S(n15534), .Z(
        n15545) );
  NAND2_X1 U15444 ( .A1(n15534), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13193) );
  AOI21_X1 U15445 ( .B1(n9815), .B2(n13194), .A(n13201), .ZN(n13195) );
  NOR2_X1 U15446 ( .A1(n13195), .A2(n15547), .ZN(n13196) );
  AOI211_X1 U15447 ( .C1(n15503), .C2(n13204), .A(n13197), .B(n13196), .ZN(
        n13198) );
  OAI21_X1 U15448 ( .B1(n13199), .B2(n15515), .A(n13198), .ZN(P3_U3195) );
  AND2_X1 U15449 ( .A1(n13207), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13246) );
  INV_X1 U15450 ( .A(n13246), .ZN(n13232) );
  OAI21_X1 U15451 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n13207), .A(n13232), 
        .ZN(n13211) );
  AOI21_X1 U15452 ( .B1(n13202), .B2(n13211), .A(n13245), .ZN(n13223) );
  NOR2_X1 U15453 ( .A1(n13204), .A2(n13203), .ZN(n13206) );
  NAND2_X1 U15454 ( .A1(n13207), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U15455 ( .B1(n13207), .B2(P3_REG2_REG_14__SCAN_IN), .A(n13233), 
        .ZN(n13224) );
  XNOR2_X1 U15456 ( .A(n13225), .B(n13224), .ZN(n13221) );
  NOR2_X1 U15457 ( .A1(n15535), .A2(n13207), .ZN(n13220) );
  INV_X1 U15458 ( .A(n13208), .ZN(n13217) );
  NOR2_X1 U15459 ( .A1(n13210), .A2(n13209), .ZN(n13214) );
  MUX2_X1 U15460 ( .A(n13224), .B(n13211), .S(n13268), .Z(n13212) );
  OAI21_X1 U15461 ( .B1(n13214), .B2(n13213), .A(n13212), .ZN(n13215) );
  NAND3_X1 U15462 ( .A1(n15550), .A2(n13235), .A3(n13215), .ZN(n13216) );
  OAI211_X1 U15463 ( .C1(n15532), .C2(n13218), .A(n13217), .B(n13216), .ZN(
        n13219) );
  AOI211_X1 U15464 ( .C1(n13221), .C2(n15539), .A(n13220), .B(n13219), .ZN(
        n13222) );
  OAI21_X1 U15465 ( .B1(n13223), .B2(n15547), .A(n13222), .ZN(P3_U3196) );
  AND2_X1 U15466 ( .A1(n15012), .A2(n13226), .ZN(n13227) );
  INV_X1 U15467 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15010) );
  NAND2_X1 U15468 ( .A1(n13250), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n13264) );
  INV_X1 U15469 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U15470 ( .A1(n13251), .A2(n13238), .ZN(n13228) );
  NAND2_X1 U15471 ( .A1(n13264), .A2(n13228), .ZN(n13230) );
  OR2_X2 U15472 ( .A1(n13231), .A2(n13230), .ZN(n13265) );
  INV_X1 U15473 ( .A(n13265), .ZN(n13229) );
  AOI21_X1 U15474 ( .B1(n13231), .B2(n13230), .A(n13229), .ZN(n13260) );
  MUX2_X1 U15475 ( .A(n13233), .B(n13232), .S(n13268), .Z(n13234) );
  NAND2_X1 U15476 ( .A1(n13235), .A2(n13234), .ZN(n13236) );
  NOR2_X1 U15477 ( .A1(n13236), .A2(n15012), .ZN(n13237) );
  AOI21_X1 U15478 ( .B1(n15012), .B2(n13236), .A(n13237), .ZN(n15017) );
  MUX2_X1 U15479 ( .A(n15010), .B(n15015), .S(n13268), .Z(n15016) );
  AND2_X1 U15480 ( .A1(n15017), .A2(n15016), .ZN(n15019) );
  MUX2_X1 U15481 ( .A(n13238), .B(n13599), .S(n13268), .Z(n13239) );
  NAND2_X1 U15482 ( .A1(n13239), .A2(n13251), .ZN(n13271) );
  INV_X1 U15483 ( .A(n13239), .ZN(n13240) );
  NAND2_X1 U15484 ( .A1(n13240), .A2(n13250), .ZN(n13270) );
  NAND2_X1 U15485 ( .A1(n13271), .A2(n13270), .ZN(n13241) );
  XNOR2_X1 U15486 ( .A(n13269), .B(n13241), .ZN(n13258) );
  NAND2_X1 U15487 ( .A1(n15503), .A2(n13251), .ZN(n13243) );
  OAI211_X1 U15488 ( .C1(n13244), .C2(n15532), .A(n13243), .B(n13242), .ZN(
        n13257) );
  NOR2_X1 U15489 ( .A1(n13248), .A2(n13247), .ZN(n13249) );
  NAND2_X1 U15490 ( .A1(n13250), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U15491 ( .A1(n13251), .A2(n13599), .ZN(n13252) );
  NAND2_X1 U15492 ( .A1(n13261), .A2(n13252), .ZN(n13253) );
  NAND2_X1 U15493 ( .A1(n13254), .A2(n13253), .ZN(n13255) );
  AOI21_X1 U15494 ( .B1(n13262), .B2(n13255), .A(n15547), .ZN(n13256) );
  AOI211_X1 U15495 ( .C1(n15550), .C2(n13258), .A(n13257), .B(n13256), .ZN(
        n13259) );
  OAI21_X1 U15496 ( .B1(n13260), .B2(n15515), .A(n13259), .ZN(P3_U3198) );
  AOI21_X1 U15497 ( .B1(n13595), .B2(n13263), .A(n13300), .ZN(n13282) );
  INV_X1 U15498 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13266) );
  MUX2_X1 U15499 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13268), .Z(n13289) );
  XNOR2_X1 U15500 ( .A(n13289), .B(n13288), .ZN(n13273) );
  AOI21_X1 U15501 ( .B1(n13273), .B2(n13272), .A(n15520), .ZN(n13277) );
  OAI21_X1 U15502 ( .B1(n15532), .B2(n13275), .A(n13274), .ZN(n13276) );
  AOI21_X1 U15503 ( .B1(n13277), .B2(n13291), .A(n13276), .ZN(n13278) );
  OAI21_X1 U15504 ( .B1(n13279), .B2(n15515), .A(n13278), .ZN(n13280) );
  OAI21_X1 U15505 ( .B1(n13282), .B2(n15547), .A(n13281), .ZN(P3_U3199) );
  NOR2_X1 U15506 ( .A1(n13299), .A2(n13283), .ZN(n13285) );
  NAND2_X1 U15507 ( .A1(n13302), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13309) );
  OAI21_X1 U15508 ( .B1(n13302), .B2(P3_REG2_REG_18__SCAN_IN), .A(n13309), 
        .ZN(n13286) );
  NAND2_X1 U15509 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  NAND2_X1 U15510 ( .A1(n13291), .A2(n13290), .ZN(n13315) );
  XNOR2_X1 U15511 ( .A(n13315), .B(n13316), .ZN(n13295) );
  INV_X1 U15512 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13293) );
  MUX2_X1 U15513 ( .A(n13293), .B(n13292), .S(n13268), .Z(n13294) );
  NAND2_X1 U15514 ( .A1(n13295), .A2(n13294), .ZN(n13319) );
  OAI21_X1 U15515 ( .B1(n13295), .B2(n13294), .A(n13319), .ZN(n13306) );
  NAND2_X1 U15516 ( .A1(n15538), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13296) );
  OAI211_X1 U15517 ( .C1(n15535), .C2(n13302), .A(n13297), .B(n13296), .ZN(
        n13305) );
  NOR2_X1 U15518 ( .A1(n13299), .A2(n13298), .ZN(n13301) );
  NAND2_X1 U15519 ( .A1(n13302), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13311) );
  OAI21_X1 U15520 ( .B1(n13302), .B2(P3_REG1_REG_18__SCAN_IN), .A(n13311), 
        .ZN(n13303) );
  INV_X1 U15521 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13308) );
  MUX2_X1 U15522 ( .A(n13308), .B(P3_REG2_REG_19__SCAN_IN), .S(n13314), .Z(
        n13322) );
  INV_X1 U15523 ( .A(n13309), .ZN(n13310) );
  INV_X1 U15524 ( .A(n13311), .ZN(n13312) );
  XNOR2_X1 U15525 ( .A(n13314), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13321) );
  INV_X1 U15526 ( .A(n13315), .ZN(n13317) );
  NAND2_X1 U15527 ( .A1(n13317), .A2(n13316), .ZN(n13318) );
  NAND2_X1 U15528 ( .A1(n13319), .A2(n13318), .ZN(n13324) );
  MUX2_X1 U15529 ( .A(n13322), .B(n13321), .S(n13268), .Z(n13323) );
  AOI21_X1 U15530 ( .B1(n15538), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n13326), 
        .ZN(n13327) );
  XNOR2_X1 U15531 ( .A(n13329), .B(n13328), .ZN(n13543) );
  NAND2_X1 U15532 ( .A1(n13331), .A2(n13330), .ZN(n13332) );
  NAND2_X1 U15533 ( .A1(n13332), .A2(n15599), .ZN(n13334) );
  AOI22_X1 U15534 ( .A1(n13335), .A2(n15613), .B1(n15615), .B2(n13359), .ZN(
        n13336) );
  NAND2_X1 U15535 ( .A1(n13545), .A2(n15625), .ZN(n13342) );
  INV_X1 U15536 ( .A(n13337), .ZN(n13339) );
  INV_X1 U15537 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13338) );
  OAI22_X1 U15538 ( .A1(n13339), .A2(n15591), .B1(n13338), .B2(n15625), .ZN(
        n13340) );
  AOI21_X1 U15539 ( .B1(n12515), .B2(n15033), .A(n13340), .ZN(n13341) );
  OAI211_X1 U15540 ( .C1(n13539), .C2(n13543), .A(n13342), .B(n13341), .ZN(
        P3_U3205) );
  INV_X1 U15541 ( .A(n13343), .ZN(n13344) );
  AOI21_X1 U15542 ( .B1(n13346), .B2(n7309), .A(n13344), .ZN(n13350) );
  AOI22_X1 U15543 ( .A1(n13345), .A2(n15613), .B1(n15615), .B2(n13372), .ZN(
        n13349) );
  XNOR2_X1 U15544 ( .A(n13347), .B(n13346), .ZN(n13549) );
  NAND2_X1 U15545 ( .A1(n13549), .A2(n15656), .ZN(n13348) );
  OAI211_X1 U15546 ( .C1(n13350), .C2(n15619), .A(n13349), .B(n13348), .ZN(
        n13548) );
  INV_X1 U15547 ( .A(n13548), .ZN(n13357) );
  INV_X1 U15548 ( .A(n13351), .ZN(n15623) );
  INV_X1 U15549 ( .A(n13352), .ZN(n13614) );
  AOI22_X1 U15550 ( .A1(n13353), .A2(n15622), .B1(P3_REG2_REG_27__SCAN_IN), 
        .B2(n15627), .ZN(n13354) );
  OAI21_X1 U15551 ( .B1(n13614), .B2(n13522), .A(n13354), .ZN(n13355) );
  AOI21_X1 U15552 ( .B1(n13549), .B2(n15623), .A(n13355), .ZN(n13356) );
  OAI21_X1 U15553 ( .B1(n13357), .B2(n15627), .A(n13356), .ZN(P3_U3206) );
  XNOR2_X1 U15554 ( .A(n13358), .B(n13362), .ZN(n13360) );
  AOI222_X1 U15555 ( .A1(n13391), .A2(n15615), .B1(n15599), .B2(n13360), .C1(
        n13359), .C2(n15613), .ZN(n13554) );
  XOR2_X1 U15556 ( .A(n13361), .B(n13362), .Z(n13555) );
  INV_X1 U15557 ( .A(n13555), .ZN(n13367) );
  INV_X1 U15558 ( .A(n13552), .ZN(n13365) );
  AOI22_X1 U15559 ( .A1(n15627), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15622), 
        .B2(n13363), .ZN(n13364) );
  OAI21_X1 U15560 ( .B1(n13365), .B2(n13522), .A(n13364), .ZN(n13366) );
  AOI21_X1 U15561 ( .B1(n13367), .B2(n13524), .A(n13366), .ZN(n13368) );
  OAI21_X1 U15562 ( .B1(n13554), .B2(n15627), .A(n13368), .ZN(P3_U3207) );
  INV_X1 U15563 ( .A(n13376), .ZN(n13370) );
  OAI211_X1 U15564 ( .C1(n6766), .C2(n13370), .A(n15599), .B(n13369), .ZN(
        n13374) );
  AOI22_X1 U15565 ( .A1(n13372), .A2(n15613), .B1(n15615), .B2(n13371), .ZN(
        n13373) );
  NAND2_X1 U15566 ( .A1(n13374), .A2(n13373), .ZN(n13556) );
  INV_X1 U15567 ( .A(n13556), .ZN(n13383) );
  OAI21_X1 U15568 ( .B1(n13377), .B2(n13376), .A(n13375), .ZN(n13557) );
  INV_X1 U15569 ( .A(n13378), .ZN(n13619) );
  AOI22_X1 U15570 ( .A1(n15627), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15622), 
        .B2(n13379), .ZN(n13380) );
  OAI21_X1 U15571 ( .B1(n13619), .B2(n13522), .A(n13380), .ZN(n13381) );
  AOI21_X1 U15572 ( .B1(n13557), .B2(n13524), .A(n13381), .ZN(n13382) );
  OAI21_X1 U15573 ( .B1(n13383), .B2(n15627), .A(n13382), .ZN(P3_U3208) );
  INV_X1 U15574 ( .A(n13384), .ZN(n13385) );
  AOI21_X1 U15575 ( .B1(n13387), .B2(n13386), .A(n13385), .ZN(n13394) );
  XNOR2_X1 U15576 ( .A(n13388), .B(n7651), .ZN(n13389) );
  NAND2_X1 U15577 ( .A1(n13389), .A2(n15599), .ZN(n13393) );
  AOI22_X1 U15578 ( .A1(n13391), .A2(n15613), .B1(n15615), .B2(n13390), .ZN(
        n13392) );
  OAI211_X1 U15579 ( .C1(n15602), .C2(n13394), .A(n13393), .B(n13392), .ZN(
        n13560) );
  INV_X1 U15580 ( .A(n13560), .ZN(n13399) );
  INV_X1 U15581 ( .A(n13394), .ZN(n13561) );
  AOI22_X1 U15582 ( .A1(n15627), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15622), 
        .B2(n13395), .ZN(n13396) );
  OAI21_X1 U15583 ( .B1(n13623), .B2(n13522), .A(n13396), .ZN(n13397) );
  AOI21_X1 U15584 ( .B1(n13561), .B2(n15623), .A(n13397), .ZN(n13398) );
  OAI21_X1 U15585 ( .B1(n13399), .B2(n15627), .A(n13398), .ZN(P3_U3209) );
  XNOR2_X1 U15586 ( .A(n13400), .B(n13404), .ZN(n13401) );
  OAI222_X1 U15587 ( .A1(n15594), .A2(n13403), .B1(n15597), .B2(n13402), .C1(
        n15619), .C2(n13401), .ZN(n13564) );
  INV_X1 U15588 ( .A(n13564), .ZN(n13410) );
  XNOR2_X1 U15589 ( .A(n13405), .B(n13404), .ZN(n13565) );
  AOI22_X1 U15590 ( .A1(n15627), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15622), 
        .B2(n13406), .ZN(n13407) );
  OAI21_X1 U15591 ( .B1(n13627), .B2(n13522), .A(n13407), .ZN(n13408) );
  AOI21_X1 U15592 ( .B1(n13565), .B2(n13524), .A(n13408), .ZN(n13409) );
  OAI21_X1 U15593 ( .B1(n13410), .B2(n15627), .A(n13409), .ZN(P3_U3210) );
  XNOR2_X1 U15594 ( .A(n13411), .B(n13415), .ZN(n13414) );
  OAI22_X1 U15595 ( .A1(n13412), .A2(n15597), .B1(n13439), .B2(n15594), .ZN(
        n13413) );
  AOI21_X1 U15596 ( .B1(n13414), .B2(n15599), .A(n13413), .ZN(n13570) );
  XNOR2_X1 U15597 ( .A(n13416), .B(n13415), .ZN(n13568) );
  AOI22_X1 U15598 ( .A1(n15627), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15622), 
        .B2(n13417), .ZN(n13418) );
  OAI21_X1 U15599 ( .B1(n13631), .B2(n13522), .A(n13418), .ZN(n13419) );
  AOI21_X1 U15600 ( .B1(n13568), .B2(n13524), .A(n13419), .ZN(n13420) );
  OAI21_X1 U15601 ( .B1(n13570), .B2(n15627), .A(n13420), .ZN(P3_U3211) );
  OAI21_X1 U15602 ( .B1(n13422), .B2(n13429), .A(n13421), .ZN(n13427) );
  NAND2_X1 U15603 ( .A1(n13423), .A2(n15613), .ZN(n13424) );
  OAI21_X1 U15604 ( .B1(n13425), .B2(n15594), .A(n13424), .ZN(n13426) );
  AOI21_X1 U15605 ( .B1(n13427), .B2(n15599), .A(n13426), .ZN(n13575) );
  XNOR2_X1 U15606 ( .A(n13428), .B(n13429), .ZN(n13573) );
  INV_X1 U15607 ( .A(n13430), .ZN(n13635) );
  AOI22_X1 U15608 ( .A1(n15627), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15622), 
        .B2(n13431), .ZN(n13432) );
  OAI21_X1 U15609 ( .B1(n13635), .B2(n13522), .A(n13432), .ZN(n13433) );
  AOI21_X1 U15610 ( .B1(n13573), .B2(n13524), .A(n13433), .ZN(n13434) );
  OAI21_X1 U15611 ( .B1(n13575), .B2(n15627), .A(n13434), .ZN(P3_U3212) );
  OAI211_X1 U15612 ( .C1(n13437), .C2(n13436), .A(n13435), .B(n15599), .ZN(
        n13442) );
  OAI22_X1 U15613 ( .A1(n13439), .A2(n15597), .B1(n13438), .B2(n15594), .ZN(
        n13440) );
  INV_X1 U15614 ( .A(n13440), .ZN(n13441) );
  XNOR2_X1 U15615 ( .A(n13444), .B(n13443), .ZN(n13578) );
  AOI22_X1 U15616 ( .A1(n15627), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15622), 
        .B2(n13445), .ZN(n13446) );
  OAI21_X1 U15617 ( .B1(n13447), .B2(n13522), .A(n13446), .ZN(n13448) );
  AOI21_X1 U15618 ( .B1(n13578), .B2(n13524), .A(n13448), .ZN(n13449) );
  OAI21_X1 U15619 ( .B1(n13580), .B2(n15627), .A(n13449), .ZN(P3_U3213) );
  OR2_X1 U15620 ( .A1(n13499), .A2(n13450), .ZN(n13452) );
  AND2_X1 U15621 ( .A1(n13452), .A2(n13451), .ZN(n13453) );
  AOI21_X1 U15622 ( .B1(n13453), .B2(n13460), .A(n15619), .ZN(n13458) );
  NAND2_X1 U15623 ( .A1(n15613), .A2(n13454), .ZN(n13455) );
  OAI21_X1 U15624 ( .B1(n13491), .B2(n15594), .A(n13455), .ZN(n13456) );
  AOI21_X1 U15625 ( .B1(n13458), .B2(n13457), .A(n13456), .ZN(n13586) );
  NAND2_X1 U15626 ( .A1(n13474), .A2(n13459), .ZN(n13462) );
  INV_X1 U15627 ( .A(n13460), .ZN(n13461) );
  XNOR2_X1 U15628 ( .A(n13462), .B(n13461), .ZN(n13584) );
  AOI22_X1 U15629 ( .A1(n15627), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15622), 
        .B2(n13463), .ZN(n13464) );
  OAI21_X1 U15630 ( .B1(n13644), .B2(n13522), .A(n13464), .ZN(n13465) );
  AOI21_X1 U15631 ( .B1(n13584), .B2(n13524), .A(n13465), .ZN(n13466) );
  OAI21_X1 U15632 ( .B1(n13586), .B2(n15627), .A(n13466), .ZN(P3_U3214) );
  AND2_X1 U15633 ( .A1(n13484), .A2(n13468), .ZN(n13471) );
  NAND2_X1 U15634 ( .A1(n13484), .A2(n13469), .ZN(n13470) );
  OAI21_X1 U15635 ( .B1(n13471), .B2(n13477), .A(n13470), .ZN(n13473) );
  AOI222_X1 U15636 ( .A1(n15599), .A2(n13473), .B1(n13472), .B2(n15613), .C1(
        n13504), .C2(n15615), .ZN(n13592) );
  INV_X1 U15637 ( .A(n13474), .ZN(n13475) );
  AOI21_X1 U15638 ( .B1(n13477), .B2(n13476), .A(n13475), .ZN(n13590) );
  AOI22_X1 U15639 ( .A1(n15627), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15622), 
        .B2(n13478), .ZN(n13479) );
  OAI21_X1 U15640 ( .B1(n13480), .B2(n13522), .A(n13479), .ZN(n13481) );
  AOI21_X1 U15641 ( .B1(n13590), .B2(n13524), .A(n13481), .ZN(n13482) );
  OAI21_X1 U15642 ( .B1(n13592), .B2(n15627), .A(n13482), .ZN(P3_U3215) );
  AND2_X1 U15643 ( .A1(n13484), .A2(n13483), .ZN(n13487) );
  OR2_X1 U15644 ( .A1(n13499), .A2(n13508), .ZN(n13500) );
  NAND3_X1 U15645 ( .A1(n13500), .A2(n12523), .A3(n13485), .ZN(n13486) );
  NAND3_X1 U15646 ( .A1(n13487), .A2(n15599), .A3(n13486), .ZN(n13490) );
  NAND2_X1 U15647 ( .A1(n13488), .A2(n15615), .ZN(n13489) );
  OAI211_X1 U15648 ( .C1(n13491), .C2(n15597), .A(n13490), .B(n13489), .ZN(
        n13593) );
  INV_X1 U15649 ( .A(n13593), .ZN(n13498) );
  NAND2_X1 U15650 ( .A1(n13507), .A2(n13492), .ZN(n13493) );
  XNOR2_X1 U15651 ( .A(n13493), .B(n12523), .ZN(n13594) );
  AOI22_X1 U15652 ( .A1(n15627), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15622), 
        .B2(n13494), .ZN(n13495) );
  OAI21_X1 U15653 ( .B1(n13649), .B2(n13522), .A(n13495), .ZN(n13496) );
  AOI21_X1 U15654 ( .B1(n13594), .B2(n13524), .A(n13496), .ZN(n13497) );
  OAI21_X1 U15655 ( .B1(n13498), .B2(n15627), .A(n13497), .ZN(P3_U3216) );
  INV_X1 U15656 ( .A(n13499), .ZN(n13502) );
  INV_X1 U15657 ( .A(n13508), .ZN(n13501) );
  OAI211_X1 U15658 ( .C1(n13502), .C2(n13501), .A(n15599), .B(n13500), .ZN(
        n13506) );
  AOI22_X1 U15659 ( .A1(n13504), .A2(n15613), .B1(n15615), .B2(n13503), .ZN(
        n13505) );
  NAND2_X1 U15660 ( .A1(n13506), .A2(n13505), .ZN(n13597) );
  INV_X1 U15661 ( .A(n13597), .ZN(n13514) );
  OAI21_X1 U15662 ( .B1(n13509), .B2(n13508), .A(n13507), .ZN(n13598) );
  AOI22_X1 U15663 ( .A1(n15627), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15622), 
        .B2(n13510), .ZN(n13511) );
  OAI21_X1 U15664 ( .B1(n13653), .B2(n13522), .A(n13511), .ZN(n13512) );
  AOI21_X1 U15665 ( .B1(n13598), .B2(n13524), .A(n13512), .ZN(n13513) );
  OAI21_X1 U15666 ( .B1(n13514), .B2(n15627), .A(n13513), .ZN(P3_U3217) );
  XOR2_X1 U15667 ( .A(n13515), .B(n13518), .Z(n13516) );
  OAI222_X1 U15668 ( .A1(n15597), .A2(n13517), .B1(n15594), .B2(n13532), .C1(
        n13516), .C2(n15619), .ZN(n13601) );
  INV_X1 U15669 ( .A(n13601), .ZN(n13526) );
  XNOR2_X1 U15670 ( .A(n13519), .B(n13518), .ZN(n13602) );
  AOI22_X1 U15671 ( .A1(n15627), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15622), 
        .B2(n13520), .ZN(n13521) );
  OAI21_X1 U15672 ( .B1(n13658), .B2(n13522), .A(n13521), .ZN(n13523) );
  AOI21_X1 U15673 ( .B1(n13602), .B2(n13524), .A(n13523), .ZN(n13525) );
  OAI21_X1 U15674 ( .B1(n13526), .B2(n15627), .A(n13525), .ZN(P3_U3218) );
  XNOR2_X1 U15675 ( .A(n13527), .B(n13528), .ZN(n15047) );
  XNOR2_X1 U15676 ( .A(n13529), .B(n13528), .ZN(n13530) );
  OAI222_X1 U15677 ( .A1(n15597), .A2(n13532), .B1(n15594), .B2(n13531), .C1(
        n13530), .C2(n15619), .ZN(n15049) );
  NAND2_X1 U15678 ( .A1(n15049), .A2(n15625), .ZN(n13538) );
  INV_X1 U15679 ( .A(n15046), .ZN(n13536) );
  INV_X1 U15680 ( .A(n13533), .ZN(n13534) );
  OAI22_X1 U15681 ( .A1(n15625), .A2(n13177), .B1(n13534), .B2(n15591), .ZN(
        n13535) );
  AOI21_X1 U15682 ( .B1(n13536), .B2(n15033), .A(n13535), .ZN(n13537) );
  OAI211_X1 U15683 ( .C1(n13539), .C2(n15047), .A(n13538), .B(n13537), .ZN(
        P3_U3220) );
  NAND2_X1 U15684 ( .A1(n13540), .A2(n15609), .ZN(n15654) );
  INV_X1 U15685 ( .A(n12515), .ZN(n13610) );
  NOR2_X1 U15686 ( .A1(n13543), .A2(n15675), .ZN(n13544) );
  NOR2_X1 U15687 ( .A1(n13545), .A2(n13544), .ZN(n13608) );
  MUX2_X1 U15688 ( .A(n13608), .B(n13546), .S(n15691), .Z(n13547) );
  OAI21_X1 U15689 ( .B1(n13610), .B2(n13604), .A(n13547), .ZN(P3_U3487) );
  AOI21_X1 U15690 ( .B1(n15672), .B2(n13549), .A(n13548), .ZN(n13611) );
  MUX2_X1 U15691 ( .A(n13550), .B(n13611), .S(n15693), .Z(n13551) );
  OAI21_X1 U15692 ( .B1(n13614), .B2(n13604), .A(n13551), .ZN(P3_U3486) );
  NAND2_X1 U15693 ( .A1(n13552), .A2(n15650), .ZN(n13553) );
  OAI211_X1 U15694 ( .C1(n15675), .C2(n13555), .A(n13554), .B(n13553), .ZN(
        n13615) );
  MUX2_X1 U15695 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13615), .S(n15693), .Z(
        P3_U3485) );
  AOI21_X1 U15696 ( .B1(n15051), .B2(n13557), .A(n13556), .ZN(n13616) );
  MUX2_X1 U15697 ( .A(n13558), .B(n13616), .S(n15693), .Z(n13559) );
  OAI21_X1 U15698 ( .B1(n13619), .B2(n13604), .A(n13559), .ZN(P3_U3484) );
  AOI21_X1 U15699 ( .B1(n15672), .B2(n13561), .A(n13560), .ZN(n13620) );
  MUX2_X1 U15700 ( .A(n13562), .B(n13620), .S(n15693), .Z(n13563) );
  OAI21_X1 U15701 ( .B1(n13623), .B2(n13604), .A(n13563), .ZN(P3_U3483) );
  INV_X1 U15702 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13566) );
  AOI21_X1 U15703 ( .B1(n13565), .B2(n15051), .A(n13564), .ZN(n13624) );
  MUX2_X1 U15704 ( .A(n13566), .B(n13624), .S(n15693), .Z(n13567) );
  OAI21_X1 U15705 ( .B1(n13627), .B2(n13604), .A(n13567), .ZN(P3_U3482) );
  INV_X1 U15706 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13571) );
  NAND2_X1 U15707 ( .A1(n13568), .A2(n15051), .ZN(n13569) );
  AND2_X1 U15708 ( .A1(n13570), .A2(n13569), .ZN(n13628) );
  MUX2_X1 U15709 ( .A(n13571), .B(n13628), .S(n15693), .Z(n13572) );
  OAI21_X1 U15710 ( .B1(n13631), .B2(n13604), .A(n13572), .ZN(P3_U3481) );
  INV_X1 U15711 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U15712 ( .A1(n13573), .A2(n15051), .ZN(n13574) );
  AND2_X1 U15713 ( .A1(n13575), .A2(n13574), .ZN(n13632) );
  MUX2_X1 U15714 ( .A(n13576), .B(n13632), .S(n15693), .Z(n13577) );
  OAI21_X1 U15715 ( .B1(n13635), .B2(n13604), .A(n13577), .ZN(P3_U3480) );
  NAND2_X1 U15716 ( .A1(n13578), .A2(n15051), .ZN(n13579) );
  NAND2_X1 U15717 ( .A1(n13580), .A2(n13579), .ZN(n13636) );
  MUX2_X1 U15718 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13636), .S(n15693), .Z(
        n13581) );
  AOI21_X1 U15719 ( .B1(n13582), .B2(n13638), .A(n13581), .ZN(n13583) );
  INV_X1 U15720 ( .A(n13583), .ZN(P3_U3479) );
  NAND2_X1 U15721 ( .A1(n13584), .A2(n15051), .ZN(n13585) );
  NAND2_X1 U15722 ( .A1(n13586), .A2(n13585), .ZN(n13641) );
  MUX2_X1 U15723 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13641), .S(n15693), .Z(
        n13587) );
  INV_X1 U15724 ( .A(n13587), .ZN(n13588) );
  OAI21_X1 U15725 ( .B1(n13604), .B2(n13644), .A(n13588), .ZN(P3_U3478) );
  AOI22_X1 U15726 ( .A1(n13590), .A2(n15051), .B1(n15650), .B2(n13589), .ZN(
        n13591) );
  NAND2_X1 U15727 ( .A1(n13592), .A2(n13591), .ZN(n13645) );
  MUX2_X1 U15728 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13645), .S(n15693), .Z(
        P3_U3477) );
  AOI21_X1 U15729 ( .B1(n13594), .B2(n15051), .A(n13593), .ZN(n13646) );
  MUX2_X1 U15730 ( .A(n13595), .B(n13646), .S(n15693), .Z(n13596) );
  OAI21_X1 U15731 ( .B1(n13649), .B2(n13604), .A(n13596), .ZN(P3_U3476) );
  AOI21_X1 U15732 ( .B1(n15051), .B2(n13598), .A(n13597), .ZN(n13650) );
  MUX2_X1 U15733 ( .A(n13599), .B(n13650), .S(n15693), .Z(n13600) );
  OAI21_X1 U15734 ( .B1(n13653), .B2(n13604), .A(n13600), .ZN(P3_U3475) );
  AOI21_X1 U15735 ( .B1(n13602), .B2(n15051), .A(n13601), .ZN(n13654) );
  MUX2_X1 U15736 ( .A(n15015), .B(n13654), .S(n15693), .Z(n13603) );
  OAI21_X1 U15737 ( .B1(n13658), .B2(n13604), .A(n13603), .ZN(P3_U3474) );
  INV_X1 U15738 ( .A(n13657), .ZN(n13639) );
  INV_X1 U15739 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13607) );
  MUX2_X1 U15740 ( .A(n13608), .B(n13607), .S(n15681), .Z(n13609) );
  OAI21_X1 U15741 ( .B1(n13610), .B2(n13657), .A(n13609), .ZN(P3_U3455) );
  INV_X1 U15742 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13612) );
  MUX2_X1 U15743 ( .A(n13612), .B(n13611), .S(n15679), .Z(n13613) );
  OAI21_X1 U15744 ( .B1(n13614), .B2(n13657), .A(n13613), .ZN(P3_U3454) );
  MUX2_X1 U15745 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13615), .S(n15679), .Z(
        P3_U3453) );
  INV_X1 U15746 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13617) );
  MUX2_X1 U15747 ( .A(n13617), .B(n13616), .S(n15679), .Z(n13618) );
  OAI21_X1 U15748 ( .B1(n13619), .B2(n13657), .A(n13618), .ZN(P3_U3452) );
  INV_X1 U15749 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13621) );
  MUX2_X1 U15750 ( .A(n13621), .B(n13620), .S(n15679), .Z(n13622) );
  OAI21_X1 U15751 ( .B1(n13623), .B2(n13657), .A(n13622), .ZN(P3_U3451) );
  INV_X1 U15752 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13625) );
  MUX2_X1 U15753 ( .A(n13625), .B(n13624), .S(n15679), .Z(n13626) );
  OAI21_X1 U15754 ( .B1(n13627), .B2(n13657), .A(n13626), .ZN(P3_U3450) );
  MUX2_X1 U15755 ( .A(n13629), .B(n13628), .S(n15679), .Z(n13630) );
  OAI21_X1 U15756 ( .B1(n13631), .B2(n13657), .A(n13630), .ZN(P3_U3449) );
  INV_X1 U15757 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13633) );
  MUX2_X1 U15758 ( .A(n13633), .B(n13632), .S(n15679), .Z(n13634) );
  OAI21_X1 U15759 ( .B1(n13635), .B2(n13657), .A(n13634), .ZN(P3_U3448) );
  MUX2_X1 U15760 ( .A(n13636), .B(P3_REG0_REG_20__SCAN_IN), .S(n15681), .Z(
        n13637) );
  AOI21_X1 U15761 ( .B1(n13639), .B2(n13638), .A(n13637), .ZN(n13640) );
  INV_X1 U15762 ( .A(n13640), .ZN(P3_U3447) );
  MUX2_X1 U15763 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13641), .S(n15679), .Z(
        n13642) );
  INV_X1 U15764 ( .A(n13642), .ZN(n13643) );
  OAI21_X1 U15765 ( .B1(n13657), .B2(n13644), .A(n13643), .ZN(P3_U3446) );
  MUX2_X1 U15766 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13645), .S(n15679), .Z(
        P3_U3444) );
  INV_X1 U15767 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13647) );
  MUX2_X1 U15768 ( .A(n13647), .B(n13646), .S(n15679), .Z(n13648) );
  OAI21_X1 U15769 ( .B1(n13649), .B2(n13657), .A(n13648), .ZN(P3_U3441) );
  INV_X1 U15770 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13651) );
  MUX2_X1 U15771 ( .A(n13651), .B(n13650), .S(n15679), .Z(n13652) );
  OAI21_X1 U15772 ( .B1(n13653), .B2(n13657), .A(n13652), .ZN(P3_U3438) );
  INV_X1 U15773 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13655) );
  MUX2_X1 U15774 ( .A(n13655), .B(n13654), .S(n15679), .Z(n13656) );
  OAI21_X1 U15775 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(P3_U3435) );
  MUX2_X1 U15776 ( .A(n13659), .B(P3_D_REG_1__SCAN_IN), .S(n13660), .Z(
        P3_U3377) );
  MUX2_X1 U15777 ( .A(n13661), .B(P3_D_REG_0__SCAN_IN), .S(n13660), .Z(
        P3_U3376) );
  NAND2_X1 U15778 ( .A1(n13663), .A2(n13662), .ZN(n13667) );
  INV_X1 U15779 ( .A(n13664), .ZN(n13665) );
  NAND4_X1 U15780 ( .A1(n13665), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .A4(n9605), .ZN(n13666) );
  OAI211_X1 U15781 ( .C1(n12971), .C2(n13668), .A(n13667), .B(n13666), .ZN(
        P3_U3264) );
  INV_X1 U15782 ( .A(n13669), .ZN(n13671) );
  OAI222_X1 U15783 ( .A1(P3_U3151), .A2(n13673), .B1(n13672), .B2(n13671), 
        .C1(n13670), .C2(n12971), .ZN(P3_U3269) );
  INV_X1 U15784 ( .A(n13915), .ZN(n13894) );
  OAI22_X1 U15785 ( .A1(n13894), .A2(n14090), .B1(n15388), .B2(n13712), .ZN(
        n14023) );
  AOI22_X1 U15786 ( .A1(n13779), .A2(n14023), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13674) );
  OAI21_X1 U15787 ( .B1(n14025), .B2(n13781), .A(n13674), .ZN(n13679) );
  AOI211_X1 U15788 ( .C1(n13677), .C2(n13676), .A(n13785), .B(n13675), .ZN(
        n13678) );
  AOI211_X1 U15789 ( .C1(n14170), .C2(n13783), .A(n13679), .B(n13678), .ZN(
        n13680) );
  INV_X1 U15790 ( .A(n13680), .ZN(P2_U3188) );
  NAND2_X1 U15791 ( .A1(n13682), .A2(n13681), .ZN(n13684) );
  XOR2_X1 U15792 ( .A(n13684), .B(n13683), .Z(n13689) );
  NOR2_X1 U15793 ( .A1(n13781), .A2(n14081), .ZN(n13687) );
  AND2_X1 U15794 ( .A1(n14127), .A2(n14124), .ZN(n13685) );
  AOI21_X1 U15795 ( .B1(n13914), .B2(n14126), .A(n13685), .ZN(n14076) );
  NAND2_X1 U15796 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13874)
         );
  OAI21_X1 U15797 ( .B1(n13742), .B2(n14076), .A(n13874), .ZN(n13686) );
  AOI211_X1 U15798 ( .C1(n14191), .C2(n13783), .A(n13687), .B(n13686), .ZN(
        n13688) );
  OAI21_X1 U15799 ( .B1(n13689), .B2(n13785), .A(n13688), .ZN(P2_U3191) );
  INV_X1 U15800 ( .A(n13690), .ZN(n13691) );
  NAND2_X1 U15801 ( .A1(n6678), .A2(n13959), .ZN(n13694) );
  XOR2_X1 U15802 ( .A(n13694), .B(n13693), .Z(n13695) );
  XNOR2_X1 U15803 ( .A(n14145), .B(n13695), .ZN(n13696) );
  INV_X1 U15804 ( .A(n13942), .ZN(n13926) );
  OAI22_X1 U15805 ( .A1(n13759), .A2(n13926), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13697), .ZN(n13700) );
  INV_X1 U15806 ( .A(n13943), .ZN(n13698) );
  OAI22_X1 U15807 ( .A1(n13770), .A2(n13698), .B1(n13781), .B2(n13947), .ZN(
        n13699) );
  AOI211_X1 U15808 ( .C1(n14145), .C2(n13783), .A(n13700), .B(n13699), .ZN(
        n13701) );
  AOI21_X1 U15809 ( .B1(n13703), .B2(n13702), .A(n13785), .ZN(n13705) );
  NAND2_X1 U15810 ( .A1(n13705), .A2(n13704), .ZN(n13711) );
  INV_X1 U15811 ( .A(n13706), .ZN(n14051) );
  NOR2_X1 U15812 ( .A1(n15388), .A2(n13894), .ZN(n13707) );
  AOI21_X1 U15813 ( .B1(n13914), .B2(n14124), .A(n13707), .ZN(n14046) );
  OAI22_X1 U15814 ( .A1(n13742), .A2(n14046), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13708), .ZN(n13709) );
  AOI21_X1 U15815 ( .B1(n14051), .B2(n13766), .A(n13709), .ZN(n13710) );
  OAI211_X1 U15816 ( .C1(n14053), .C2(n13747), .A(n13711), .B(n13710), .ZN(
        P2_U3195) );
  OAI22_X1 U15817 ( .A1(n13712), .A2(n14090), .B1(n15388), .B2(n13900), .ZN(
        n13982) );
  AOI22_X1 U15818 ( .A1(n13779), .A2(n13982), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13713) );
  OAI21_X1 U15819 ( .B1(n13988), .B2(n13781), .A(n13713), .ZN(n13717) );
  INV_X1 U15820 ( .A(n13718), .ZN(P2_U3197) );
  INV_X1 U15821 ( .A(n13719), .ZN(n13720) );
  AOI21_X1 U15822 ( .B1(n13722), .B2(n13721), .A(n13720), .ZN(n13728) );
  NOR2_X1 U15823 ( .A1(n13781), .A2(n13723), .ZN(n13726) );
  OAI21_X1 U15824 ( .B1(n13742), .B2(n14204), .A(n13724), .ZN(n13725) );
  AOI211_X1 U15825 ( .C1(n14207), .C2(n13783), .A(n13726), .B(n13725), .ZN(
        n13727) );
  OAI21_X1 U15826 ( .B1(n13728), .B2(n13785), .A(n13727), .ZN(P2_U3198) );
  INV_X1 U15827 ( .A(n14200), .ZN(n14120) );
  OAI21_X1 U15828 ( .B1(n13731), .B2(n13730), .A(n6990), .ZN(n13732) );
  NAND2_X1 U15829 ( .A1(n13732), .A2(n9100), .ZN(n13736) );
  AND2_X1 U15830 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15370) );
  OAI22_X1 U15831 ( .A1(n13759), .A2(n13887), .B1(n13781), .B2(n14116), .ZN(
        n13733) );
  AOI211_X1 U15832 ( .C1(n13734), .C2(n14127), .A(n15370), .B(n13733), .ZN(
        n13735) );
  OAI211_X1 U15833 ( .C1(n14120), .C2(n13747), .A(n13736), .B(n13735), .ZN(
        P2_U3200) );
  INV_X1 U15834 ( .A(n14165), .ZN(n13921) );
  OAI21_X1 U15835 ( .B1(n13739), .B2(n13738), .A(n6672), .ZN(n13740) );
  NAND2_X1 U15836 ( .A1(n13740), .A2(n9100), .ZN(n13746) );
  INV_X1 U15837 ( .A(n14008), .ZN(n13744) );
  AOI22_X1 U15838 ( .A1(n14124), .A2(n14030), .B1(n14126), .B2(n13898), .ZN(
        n14000) );
  INV_X1 U15839 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13741) );
  OAI22_X1 U15840 ( .A1(n13742), .A2(n14000), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13741), .ZN(n13743) );
  AOI21_X1 U15841 ( .B1(n13744), .B2(n13766), .A(n13743), .ZN(n13745) );
  OAI211_X1 U15842 ( .C1(n13921), .C2(n13747), .A(n13746), .B(n13745), .ZN(
        P2_U3201) );
  INV_X1 U15843 ( .A(n13748), .ZN(n13749) );
  AOI21_X1 U15844 ( .B1(n13751), .B2(n13750), .A(n13749), .ZN(n13755) );
  OAI22_X1 U15845 ( .A1(n7047), .A2(n15388), .B1(n14092), .B2(n14090), .ZN(
        n14060) );
  AOI22_X1 U15846 ( .A1(n13779), .A2(n14060), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13752) );
  OAI21_X1 U15847 ( .B1(n14063), .B2(n13781), .A(n13752), .ZN(n13753) );
  AOI21_X1 U15848 ( .B1(n14185), .B2(n13783), .A(n13753), .ZN(n13754) );
  OAI21_X1 U15849 ( .B1(n13755), .B2(n13785), .A(n13754), .ZN(P2_U3205) );
  XOR2_X1 U15850 ( .A(n13757), .B(n13756), .Z(n13763) );
  INV_X1 U15851 ( .A(n14030), .ZN(n13918) );
  INV_X1 U15852 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13758) );
  OAI22_X1 U15853 ( .A1(n13770), .A2(n13918), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13758), .ZN(n13761) );
  OAI22_X1 U15854 ( .A1(n13759), .A2(n7047), .B1(n13781), .B2(n14035), .ZN(
        n13760) );
  AOI211_X1 U15855 ( .C1(n14175), .C2(n13783), .A(n13761), .B(n13760), .ZN(
        n13762) );
  OAI21_X1 U15856 ( .B1(n13763), .B2(n13785), .A(n13762), .ZN(P2_U3207) );
  XNOR2_X1 U15857 ( .A(n13765), .B(n13764), .ZN(n13773) );
  AOI22_X1 U15858 ( .A1(n13767), .A2(n13889), .B1(n13766), .B2(n14100), .ZN(
        n13769) );
  OAI211_X1 U15859 ( .C1(n14092), .C2(n13770), .A(n13769), .B(n13768), .ZN(
        n13771) );
  AOI21_X1 U15860 ( .B1(n14195), .B2(n13783), .A(n13771), .ZN(n13772) );
  OAI21_X1 U15861 ( .B1(n13773), .B2(n13785), .A(n13772), .ZN(P2_U3210) );
  OAI21_X1 U15862 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(n13777) );
  INV_X1 U15863 ( .A(n13777), .ZN(n13786) );
  NAND2_X1 U15864 ( .A1(n14124), .A2(n13898), .ZN(n13778) );
  OAI21_X1 U15865 ( .B1(n13926), .B2(n15388), .A(n13778), .ZN(n13966) );
  AOI22_X1 U15866 ( .A1(n13779), .A2(n13966), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13780) );
  OAI21_X1 U15867 ( .B1(n13971), .B2(n13781), .A(n13780), .ZN(n13782) );
  AOI21_X1 U15868 ( .B1(n14154), .B2(n13783), .A(n13782), .ZN(n13784) );
  OAI21_X1 U15869 ( .B1(n13786), .B2(n13785), .A(n13784), .ZN(P2_U3212) );
  MUX2_X1 U15870 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13879), .S(P2_U3947), .Z(
        P2_U3562) );
  INV_X2 U15871 ( .A(P2_U3947), .ZN(n13801) );
  MUX2_X1 U15872 ( .A(n13930), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13801), .Z(
        P2_U3561) );
  MUX2_X1 U15873 ( .A(n13943), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13801), .Z(
        P2_U3560) );
  MUX2_X1 U15874 ( .A(n13959), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13801), .Z(
        P2_U3559) );
  MUX2_X1 U15875 ( .A(n13942), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13801), .Z(
        P2_U3558) );
  MUX2_X1 U15876 ( .A(n13960), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13801), .Z(
        P2_U3557) );
  MUX2_X1 U15877 ( .A(n13898), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13801), .Z(
        P2_U3556) );
  MUX2_X1 U15878 ( .A(n13920), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13801), .Z(
        P2_U3555) );
  MUX2_X1 U15879 ( .A(n14030), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13801), .Z(
        P2_U3554) );
  MUX2_X1 U15880 ( .A(n13915), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13801), .Z(
        P2_U3553) );
  MUX2_X1 U15881 ( .A(n14031), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13801), .Z(
        P2_U3552) );
  MUX2_X1 U15882 ( .A(n13914), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13801), .Z(
        P2_U3551) );
  MUX2_X1 U15883 ( .A(n13892), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13801), .Z(
        P2_U3550) );
  MUX2_X1 U15884 ( .A(n14127), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13801), .Z(
        P2_U3549) );
  MUX2_X1 U15885 ( .A(n13889), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13801), .Z(
        P2_U3548) );
  MUX2_X1 U15886 ( .A(n14125), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13801), .Z(
        P2_U3547) );
  MUX2_X1 U15887 ( .A(n13787), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13801), .Z(
        P2_U3546) );
  MUX2_X1 U15888 ( .A(n13788), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13801), .Z(
        P2_U3545) );
  MUX2_X1 U15889 ( .A(n13789), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13801), .Z(
        P2_U3543) );
  MUX2_X1 U15890 ( .A(n13790), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13801), .Z(
        P2_U3542) );
  MUX2_X1 U15891 ( .A(n13791), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13801), .Z(
        P2_U3541) );
  MUX2_X1 U15892 ( .A(n13792), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13801), .Z(
        P2_U3540) );
  MUX2_X1 U15893 ( .A(n13793), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13801), .Z(
        P2_U3539) );
  MUX2_X1 U15894 ( .A(n13794), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13801), .Z(
        P2_U3538) );
  MUX2_X1 U15895 ( .A(n13795), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13801), .Z(
        P2_U3537) );
  MUX2_X1 U15896 ( .A(n13796), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13801), .Z(
        P2_U3536) );
  MUX2_X1 U15897 ( .A(n13797), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13801), .Z(
        P2_U3535) );
  MUX2_X1 U15898 ( .A(n13798), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13801), .Z(
        P2_U3534) );
  MUX2_X1 U15899 ( .A(n13799), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13801), .Z(
        P2_U3533) );
  MUX2_X1 U15900 ( .A(n13800), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13801), .Z(
        P2_U3532) );
  MUX2_X1 U15901 ( .A(n10891), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13801), .Z(
        P2_U3531) );
  NAND2_X1 U15902 ( .A1(n15358), .A2(n13805), .ZN(n13814) );
  OAI211_X1 U15903 ( .C1(n13804), .C2(n13803), .A(n15364), .B(n13802), .ZN(
        n13813) );
  MUX2_X1 U15904 ( .A(n11419), .B(P2_REG2_REG_3__SCAN_IN), .S(n13805), .Z(
        n13806) );
  NAND3_X1 U15905 ( .A1(n15311), .A2(n13807), .A3(n13806), .ZN(n13808) );
  NAND3_X1 U15906 ( .A1(n15372), .A2(n13821), .A3(n13808), .ZN(n13812) );
  NOR2_X1 U15907 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13809), .ZN(n13810) );
  AOI21_X1 U15908 ( .B1(n15371), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13810), .ZN(
        n13811) );
  NAND4_X1 U15909 ( .A1(n13814), .A2(n13813), .A3(n13812), .A4(n13811), .ZN(
        P2_U3217) );
  NAND2_X1 U15910 ( .A1(n15358), .A2(n13815), .ZN(n13830) );
  OAI211_X1 U15911 ( .C1(n13818), .C2(n13817), .A(n15364), .B(n13816), .ZN(
        n13829) );
  MUX2_X1 U15912 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11794), .S(n13819), .Z(
        n13822) );
  NAND3_X1 U15913 ( .A1(n13822), .A2(n13821), .A3(n13820), .ZN(n13823) );
  NAND3_X1 U15914 ( .A1(n15372), .A2(n13824), .A3(n13823), .ZN(n13828) );
  INV_X1 U15915 ( .A(n13825), .ZN(n13826) );
  AOI21_X1 U15916 ( .B1(n15371), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n13826), .ZN(
        n13827) );
  NAND4_X1 U15917 ( .A1(n13830), .A2(n13829), .A3(n13828), .A4(n13827), .ZN(
        P2_U3218) );
  OAI21_X1 U15918 ( .B1(n15363), .B2(n9190), .A(n13831), .ZN(n13832) );
  AOI21_X1 U15919 ( .B1(n13836), .B2(n15358), .A(n13832), .ZN(n13844) );
  OAI211_X1 U15920 ( .C1(n13835), .C2(n13834), .A(n15364), .B(n13833), .ZN(
        n13843) );
  INV_X1 U15921 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n13837) );
  MUX2_X1 U15922 ( .A(n13837), .B(P2_REG2_REG_7__SCAN_IN), .S(n13836), .Z(
        n13838) );
  NAND3_X1 U15923 ( .A1(n13840), .A2(n13839), .A3(n13838), .ZN(n13841) );
  NAND3_X1 U15924 ( .A1(n15372), .A2(n13853), .A3(n13841), .ZN(n13842) );
  NAND3_X1 U15925 ( .A1(n13844), .A2(n13843), .A3(n13842), .ZN(P2_U3221) );
  NOR2_X1 U15926 ( .A1(n15379), .A2(n13850), .ZN(n13845) );
  AOI211_X1 U15927 ( .C1(n15371), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n13846), .B(
        n13845), .ZN(n13858) );
  OAI211_X1 U15928 ( .C1(n13849), .C2(n13848), .A(n15364), .B(n13847), .ZN(
        n13857) );
  MUX2_X1 U15929 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10814), .S(n13850), .Z(
        n13851) );
  NAND3_X1 U15930 ( .A1(n13853), .A2(n13852), .A3(n13851), .ZN(n13854) );
  NAND3_X1 U15931 ( .A1(n15372), .A2(n13855), .A3(n13854), .ZN(n13856) );
  NAND3_X1 U15932 ( .A1(n13858), .A2(n13857), .A3(n13856), .ZN(P2_U3222) );
  NOR2_X1 U15933 ( .A1(n13860), .A2(n13859), .ZN(n13861) );
  XOR2_X1 U15934 ( .A(n13861), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13870) );
  NOR2_X1 U15935 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  XNOR2_X1 U15936 ( .A(n13864), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13869) );
  INV_X1 U15937 ( .A(n13869), .ZN(n13865) );
  NAND2_X1 U15938 ( .A1(n13865), .A2(n15364), .ZN(n13866) );
  OAI211_X1 U15939 ( .C1(n13870), .C2(n13867), .A(n13866), .B(n15379), .ZN(
        n13868) );
  INV_X1 U15940 ( .A(n13868), .ZN(n13873) );
  AOI22_X1 U15941 ( .A1(n13870), .A2(n15372), .B1(n15364), .B2(n13869), .ZN(
        n13872) );
  MUX2_X1 U15942 ( .A(n13873), .B(n13872), .S(n13871), .Z(n13875) );
  OAI211_X1 U15943 ( .C1(n7801), .C2(n15363), .A(n13875), .B(n13874), .ZN(
        P2_U3233) );
  INV_X1 U15944 ( .A(n14145), .ZN(n13937) );
  NAND2_X1 U15945 ( .A1(n14112), .A2(n14120), .ZN(n14113) );
  NOR2_X1 U15946 ( .A1(n14113), .A2(n14195), .ZN(n14099) );
  INV_X1 U15947 ( .A(n14191), .ZN(n14084) );
  NAND2_X1 U15948 ( .A1(n14099), .A2(n14084), .ZN(n14078) );
  INV_X1 U15949 ( .A(n14159), .ZN(n13991) );
  AND2_X2 U15950 ( .A1(n14007), .A2(n13991), .ZN(n13992) );
  INV_X1 U15951 ( .A(n14154), .ZN(n13974) );
  NAND2_X1 U15952 ( .A1(n14138), .A2(n13904), .ZN(n13882) );
  XNOR2_X1 U15953 ( .A(n14135), .B(n13882), .ZN(n13877) );
  NAND2_X1 U15954 ( .A1(n13877), .A2(n8580), .ZN(n14134) );
  AOI21_X1 U15955 ( .B1(n13878), .B2(P2_B_REG_SCAN_IN), .A(n15388), .ZN(n13929) );
  NAND2_X1 U15956 ( .A1(n13929), .A2(n13879), .ZN(n14136) );
  NOR2_X1 U15957 ( .A1(n15394), .A2(n14136), .ZN(n13884) );
  NOR2_X1 U15958 ( .A1(n14135), .A2(n14102), .ZN(n13880) );
  AOI211_X1 U15959 ( .C1(n15394), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13884), 
        .B(n13880), .ZN(n13881) );
  OAI21_X1 U15960 ( .B1(n13886), .B2(n14134), .A(n13881), .ZN(P2_U3234) );
  OAI211_X1 U15961 ( .C1(n14138), .C2(n13904), .A(n13882), .B(n8580), .ZN(
        n14137) );
  NOR2_X1 U15962 ( .A1(n14138), .A2(n14102), .ZN(n13883) );
  AOI211_X1 U15963 ( .C1(n15394), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13884), 
        .B(n13883), .ZN(n13885) );
  OAI21_X1 U15964 ( .B1(n13886), .B2(n14137), .A(n13885), .ZN(P2_U3235) );
  INV_X1 U15965 ( .A(n14175), .ZN(n13916) );
  INV_X1 U15966 ( .A(n14207), .ZN(n13909) );
  NAND2_X1 U15967 ( .A1(n14089), .A2(n14093), .ZN(n14088) );
  INV_X1 U15968 ( .A(n14185), .ZN(n14066) );
  INV_X1 U15969 ( .A(n13895), .ZN(n13897) );
  INV_X1 U15970 ( .A(n13998), .ZN(n14004) );
  NAND2_X1 U15971 ( .A1(n13986), .A2(n13985), .ZN(n13984) );
  NOR2_X1 U15972 ( .A1(n14154), .A2(n13960), .ZN(n13901) );
  AOI211_X1 U15973 ( .C1(n14140), .C2(n13933), .A(n6678), .B(n13904), .ZN(
        n14139) );
  INV_X1 U15974 ( .A(n13905), .ZN(n13906) );
  AOI22_X1 U15975 ( .A1(n15394), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13906), 
        .B2(n14117), .ZN(n13907) );
  OAI21_X1 U15976 ( .B1(n7340), .B2(n14102), .A(n13907), .ZN(n13931) );
  INV_X1 U15977 ( .A(n14195), .ZN(n14103) );
  INV_X1 U15978 ( .A(n13908), .ZN(n13910) );
  INV_X1 U15979 ( .A(n14110), .ZN(n14123) );
  NAND2_X1 U15980 ( .A1(n14122), .A2(n14123), .ZN(n14121) );
  NAND2_X1 U15981 ( .A1(n14121), .A2(n13912), .ZN(n14094) );
  INV_X1 U15982 ( .A(n14074), .ZN(n14072) );
  INV_X1 U15983 ( .A(n14170), .ZN(n14020) );
  NAND2_X1 U15984 ( .A1(n14020), .A2(n14030), .ZN(n13919) );
  INV_X1 U15985 ( .A(n13985), .ZN(n13980) );
  AOI22_X1 U15986 ( .A1(n13981), .A2(n13980), .B1(n13922), .B2(n14159), .ZN(
        n13965) );
  INV_X1 U15987 ( .A(n13923), .ZN(n13925) );
  NAND2_X1 U15988 ( .A1(n14149), .A2(n13926), .ZN(n13941) );
  INV_X1 U15989 ( .A(n13952), .ZN(n13935) );
  INV_X1 U15990 ( .A(n13933), .ZN(n13934) );
  AOI211_X1 U15991 ( .C1(n14145), .C2(n13935), .A(n6678), .B(n13934), .ZN(
        n14144) );
  INV_X1 U15992 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13936) );
  OAI22_X1 U15993 ( .A1(n13937), .A2(n14102), .B1(n15392), .B2(n13936), .ZN(
        n13938) );
  AOI21_X1 U15994 ( .B1(n14144), .B2(n14108), .A(n13938), .ZN(n13950) );
  NAND2_X1 U15995 ( .A1(n13939), .A2(n14129), .ZN(n13946) );
  AOI21_X1 U15996 ( .B1(n13956), .B2(n13941), .A(n13940), .ZN(n13945) );
  AOI22_X1 U15997 ( .A1(n14126), .A2(n13943), .B1(n14124), .B2(n13942), .ZN(
        n13944) );
  NOR2_X1 U15998 ( .A1(n15384), .A2(n13947), .ZN(n13948) );
  OAI211_X1 U15999 ( .C1(n14147), .C2(n14133), .A(n13950), .B(n13949), .ZN(
        P2_U3237) );
  XNOR2_X1 U16000 ( .A(n13951), .B(n7024), .ZN(n14152) );
  AOI211_X1 U16001 ( .C1(n14149), .C2(n13968), .A(n6678), .B(n13952), .ZN(
        n14148) );
  INV_X1 U16002 ( .A(n13953), .ZN(n13954) );
  AOI22_X1 U16003 ( .A1(n15394), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13954), 
        .B2(n14117), .ZN(n13955) );
  OAI21_X1 U16004 ( .B1(n7344), .B2(n14102), .A(n13955), .ZN(n13963) );
  OAI21_X1 U16005 ( .B1(n13958), .B2(n13957), .A(n13956), .ZN(n13961) );
  AOI211_X1 U16006 ( .C1(n14148), .C2(n14108), .A(n13963), .B(n13962), .ZN(
        n13964) );
  OAI21_X1 U16007 ( .B1(n14152), .B2(n14133), .A(n13964), .ZN(P2_U3238) );
  XNOR2_X1 U16008 ( .A(n13965), .B(n13976), .ZN(n13967) );
  AOI21_X1 U16009 ( .B1(n13967), .B2(n14129), .A(n13966), .ZN(n14156) );
  INV_X1 U16010 ( .A(n13992), .ZN(n13970) );
  INV_X1 U16011 ( .A(n13968), .ZN(n13969) );
  AOI211_X1 U16012 ( .C1(n14154), .C2(n13970), .A(n6678), .B(n13969), .ZN(
        n14153) );
  INV_X1 U16013 ( .A(n13971), .ZN(n13972) );
  AOI22_X1 U16014 ( .A1(n15394), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13972), 
        .B2(n14117), .ZN(n13973) );
  OAI21_X1 U16015 ( .B1(n13974), .B2(n14102), .A(n13973), .ZN(n13978) );
  XOR2_X1 U16016 ( .A(n13976), .B(n13975), .Z(n14157) );
  NOR2_X1 U16017 ( .A1(n14157), .A2(n14133), .ZN(n13977) );
  AOI211_X1 U16018 ( .C1(n14153), .C2(n14108), .A(n13978), .B(n13977), .ZN(
        n13979) );
  OAI21_X1 U16019 ( .B1(n15394), .B2(n14156), .A(n13979), .ZN(P2_U3239) );
  XNOR2_X1 U16020 ( .A(n13981), .B(n13980), .ZN(n13983) );
  AOI21_X1 U16021 ( .B1(n13983), .B2(n14129), .A(n13982), .ZN(n14161) );
  OAI21_X1 U16022 ( .B1(n13986), .B2(n13985), .A(n13984), .ZN(n13987) );
  INV_X1 U16023 ( .A(n13987), .ZN(n14162) );
  OAI22_X1 U16024 ( .A1(n15392), .A2(n13989), .B1(n13988), .B2(n15384), .ZN(
        n13990) );
  AOI21_X1 U16025 ( .B1(n14159), .B2(n14038), .A(n13990), .ZN(n13995) );
  OAI21_X1 U16026 ( .B1(n14007), .B2(n13991), .A(n8580), .ZN(n13993) );
  NOR2_X1 U16027 ( .A1(n13993), .A2(n13992), .ZN(n14158) );
  NAND2_X1 U16028 ( .A1(n14158), .A2(n14108), .ZN(n13994) );
  OAI211_X1 U16029 ( .C1(n14162), .C2(n14133), .A(n13995), .B(n13994), .ZN(
        n13996) );
  INV_X1 U16030 ( .A(n13996), .ZN(n13997) );
  OAI21_X1 U16031 ( .B1(n15394), .B2(n14161), .A(n13997), .ZN(P2_U3240) );
  XNOR2_X1 U16032 ( .A(n13999), .B(n13998), .ZN(n14002) );
  INV_X1 U16033 ( .A(n14000), .ZN(n14001) );
  AOI21_X1 U16034 ( .B1(n14002), .B2(n14129), .A(n14001), .ZN(n14167) );
  AOI21_X1 U16035 ( .B1(n14004), .B2(n14003), .A(n6748), .ZN(n14163) );
  NAND2_X1 U16036 ( .A1(n14016), .A2(n14165), .ZN(n14005) );
  NAND2_X1 U16037 ( .A1(n14005), .A2(n8580), .ZN(n14006) );
  NOR2_X1 U16038 ( .A1(n14007), .A2(n14006), .ZN(n14164) );
  NAND2_X1 U16039 ( .A1(n14164), .A2(n14108), .ZN(n14012) );
  OAI22_X1 U16040 ( .A1(n15392), .A2(n14009), .B1(n14008), .B2(n15384), .ZN(
        n14010) );
  AOI21_X1 U16041 ( .B1(n14165), .B2(n14038), .A(n14010), .ZN(n14011) );
  NAND2_X1 U16042 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  AOI21_X1 U16043 ( .B1(n14163), .B2(n12324), .A(n14013), .ZN(n14014) );
  OAI21_X1 U16044 ( .B1(n15394), .B2(n14167), .A(n14014), .ZN(P2_U3241) );
  XOR2_X1 U16045 ( .A(n14015), .B(n14022), .Z(n14173) );
  INV_X1 U16046 ( .A(n14016), .ZN(n14017) );
  AOI211_X1 U16047 ( .C1(n14170), .C2(n14039), .A(n14018), .B(n14017), .ZN(
        n14169) );
  INV_X1 U16048 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14019) );
  OAI22_X1 U16049 ( .A1(n14020), .A2(n14102), .B1(n15392), .B2(n14019), .ZN(
        n14021) );
  AOI21_X1 U16050 ( .B1(n14169), .B2(n14108), .A(n14021), .ZN(n14028) );
  XNOR2_X1 U16051 ( .A(n6795), .B(n14022), .ZN(n14024) );
  AOI21_X1 U16052 ( .B1(n14024), .B2(n14129), .A(n14023), .ZN(n14172) );
  OAI21_X1 U16053 ( .B1(n14025), .B2(n15384), .A(n14172), .ZN(n14026) );
  NAND2_X1 U16054 ( .A1(n14026), .A2(n15392), .ZN(n14027) );
  OAI211_X1 U16055 ( .C1(n14173), .C2(n14133), .A(n14028), .B(n14027), .ZN(
        P2_U3242) );
  XNOR2_X1 U16056 ( .A(n14029), .B(n7493), .ZN(n14032) );
  AOI222_X1 U16057 ( .A1(n14129), .A2(n14032), .B1(n14031), .B2(n14124), .C1(
        n14030), .C2(n14126), .ZN(n14177) );
  OAI21_X1 U16058 ( .B1(n14034), .B2(n7493), .A(n6995), .ZN(n14178) );
  OAI22_X1 U16059 ( .A1(n15392), .A2(n14036), .B1(n14035), .B2(n15384), .ZN(
        n14037) );
  AOI21_X1 U16060 ( .B1(n14175), .B2(n14038), .A(n14037), .ZN(n14042) );
  AOI21_X1 U16061 ( .B1(n14049), .B2(n14175), .A(n6678), .ZN(n14040) );
  AND2_X1 U16062 ( .A1(n14040), .A2(n14039), .ZN(n14174) );
  NAND2_X1 U16063 ( .A1(n14174), .A2(n14108), .ZN(n14041) );
  OAI211_X1 U16064 ( .C1(n14178), .C2(n14133), .A(n14042), .B(n14041), .ZN(
        n14043) );
  INV_X1 U16065 ( .A(n14043), .ZN(n14044) );
  OAI21_X1 U16066 ( .B1(n15394), .B2(n14177), .A(n14044), .ZN(P2_U3243) );
  XNOR2_X1 U16067 ( .A(n14045), .B(n14054), .ZN(n14048) );
  INV_X1 U16068 ( .A(n14046), .ZN(n14047) );
  AOI21_X1 U16069 ( .B1(n14048), .B2(n14129), .A(n14047), .ZN(n14182) );
  INV_X1 U16070 ( .A(n14049), .ZN(n14050) );
  AOI211_X1 U16071 ( .C1(n14180), .C2(n14062), .A(n6678), .B(n14050), .ZN(
        n14179) );
  AOI22_X1 U16072 ( .A1(n15394), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14051), 
        .B2(n14117), .ZN(n14052) );
  OAI21_X1 U16073 ( .B1(n14053), .B2(n14102), .A(n14052), .ZN(n14057) );
  XNOR2_X1 U16074 ( .A(n14055), .B(n14054), .ZN(n14183) );
  NOR2_X1 U16075 ( .A1(n14183), .A2(n14133), .ZN(n14056) );
  AOI211_X1 U16076 ( .C1(n14179), .C2(n14108), .A(n14057), .B(n14056), .ZN(
        n14058) );
  OAI21_X1 U16077 ( .B1(n15394), .B2(n14182), .A(n14058), .ZN(P2_U3244) );
  XNOR2_X1 U16078 ( .A(n14059), .B(n14068), .ZN(n14061) );
  AOI21_X1 U16079 ( .B1(n14061), .B2(n14129), .A(n14060), .ZN(n14187) );
  AOI211_X1 U16080 ( .C1(n14185), .C2(n14078), .A(n6678), .B(n7350), .ZN(
        n14184) );
  INV_X1 U16081 ( .A(n14063), .ZN(n14064) );
  AOI22_X1 U16082 ( .A1(n15394), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14064), 
        .B2(n14117), .ZN(n14065) );
  OAI21_X1 U16083 ( .B1(n14066), .B2(n14102), .A(n14065), .ZN(n14070) );
  XOR2_X1 U16084 ( .A(n14068), .B(n14067), .Z(n14188) );
  NOR2_X1 U16085 ( .A1(n14188), .A2(n14133), .ZN(n14069) );
  AOI211_X1 U16086 ( .C1(n14184), .C2(n14108), .A(n14070), .B(n14069), .ZN(
        n14071) );
  OAI21_X1 U16087 ( .B1(n15394), .B2(n14187), .A(n14071), .ZN(P2_U3245) );
  XNOR2_X1 U16088 ( .A(n14073), .B(n14072), .ZN(n14193) );
  XNOR2_X1 U16089 ( .A(n14075), .B(n14074), .ZN(n14077) );
  OAI21_X1 U16090 ( .B1(n14077), .B2(n14095), .A(n14076), .ZN(n14189) );
  NAND2_X1 U16091 ( .A1(n14189), .A2(n15392), .ZN(n14087) );
  INV_X1 U16092 ( .A(n14099), .ZN(n14080) );
  INV_X1 U16093 ( .A(n14078), .ZN(n14079) );
  AOI211_X1 U16094 ( .C1(n14191), .C2(n14080), .A(n6678), .B(n14079), .ZN(
        n14190) );
  INV_X1 U16095 ( .A(n14081), .ZN(n14082) );
  AOI22_X1 U16096 ( .A1(n15394), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14082), 
        .B2(n14117), .ZN(n14083) );
  OAI21_X1 U16097 ( .B1(n14084), .B2(n14102), .A(n14083), .ZN(n14085) );
  AOI21_X1 U16098 ( .B1(n14190), .B2(n14108), .A(n14085), .ZN(n14086) );
  OAI211_X1 U16099 ( .C1(n14133), .C2(n14193), .A(n14087), .B(n14086), .ZN(
        P2_U3246) );
  INV_X1 U16100 ( .A(n15471), .ZN(n15460) );
  OAI21_X1 U16101 ( .B1(n14089), .B2(n14093), .A(n14088), .ZN(n14104) );
  OAI22_X1 U16102 ( .A1(n14092), .A2(n15388), .B1(n14091), .B2(n14090), .ZN(
        n14098) );
  XNOR2_X1 U16103 ( .A(n14094), .B(n14093), .ZN(n14096) );
  NOR2_X1 U16104 ( .A1(n14096), .A2(n14095), .ZN(n14097) );
  AOI211_X1 U16105 ( .C1(n15460), .C2(n14104), .A(n14098), .B(n14097), .ZN(
        n14197) );
  AOI211_X1 U16106 ( .C1(n14195), .C2(n14113), .A(n6678), .B(n14099), .ZN(
        n14194) );
  AOI22_X1 U16107 ( .A1(n15394), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14100), 
        .B2(n14117), .ZN(n14101) );
  OAI21_X1 U16108 ( .B1(n14103), .B2(n14102), .A(n14101), .ZN(n14107) );
  INV_X1 U16109 ( .A(n14104), .ZN(n14198) );
  NOR2_X1 U16110 ( .A1(n14198), .A2(n14105), .ZN(n14106) );
  AOI211_X1 U16111 ( .C1(n14194), .C2(n14108), .A(n14107), .B(n14106), .ZN(
        n14109) );
  OAI21_X1 U16112 ( .B1(n15394), .B2(n14197), .A(n14109), .ZN(P2_U3247) );
  XNOR2_X1 U16113 ( .A(n14111), .B(n14110), .ZN(n14203) );
  INV_X1 U16114 ( .A(n14112), .ZN(n14115) );
  INV_X1 U16115 ( .A(n14113), .ZN(n14114) );
  AOI211_X1 U16116 ( .C1(n14200), .C2(n14115), .A(n6678), .B(n14114), .ZN(
        n14199) );
  INV_X1 U16117 ( .A(n14116), .ZN(n14118) );
  AOI22_X1 U16118 ( .A1(n15394), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14118), 
        .B2(n14117), .ZN(n14119) );
  OAI21_X1 U16119 ( .B1(n14120), .B2(n14102), .A(n14119), .ZN(n14131) );
  OAI21_X1 U16120 ( .B1(n14123), .B2(n14122), .A(n14121), .ZN(n14128) );
  AOI222_X1 U16121 ( .A1(n14129), .A2(n14128), .B1(n14127), .B2(n14126), .C1(
        n14125), .C2(n14124), .ZN(n14202) );
  NOR2_X1 U16122 ( .A1(n14202), .A2(n15394), .ZN(n14130) );
  AOI211_X1 U16123 ( .C1(n14199), .C2(n14108), .A(n14131), .B(n14130), .ZN(
        n14132) );
  OAI21_X1 U16124 ( .B1(n14133), .B2(n14203), .A(n14132), .ZN(P2_U3248) );
  OAI211_X1 U16125 ( .C1(n14135), .C2(n15467), .A(n14134), .B(n14136), .ZN(
        n14217) );
  MUX2_X1 U16126 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14217), .S(n15489), .Z(
        P2_U3530) );
  OAI211_X1 U16127 ( .C1(n14138), .C2(n15467), .A(n14137), .B(n14136), .ZN(
        n14218) );
  MUX2_X1 U16128 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14218), .S(n15489), .Z(
        P2_U3529) );
  AOI21_X1 U16129 ( .B1(n15450), .B2(n14140), .A(n14139), .ZN(n14141) );
  MUX2_X1 U16130 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14219), .S(n15489), .Z(
        P2_U3528) );
  OAI21_X1 U16131 ( .B1(n14147), .B2(n15454), .A(n14146), .ZN(n14220) );
  MUX2_X1 U16132 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14220), .S(n15489), .Z(
        P2_U3527) );
  AOI21_X1 U16133 ( .B1(n15450), .B2(n14149), .A(n14148), .ZN(n14150) );
  OAI211_X1 U16134 ( .C1(n14152), .C2(n15454), .A(n14151), .B(n14150), .ZN(
        n14221) );
  MUX2_X1 U16135 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14221), .S(n15489), .Z(
        P2_U3526) );
  AOI21_X1 U16136 ( .B1(n15450), .B2(n14154), .A(n14153), .ZN(n14155) );
  OAI211_X1 U16137 ( .C1(n14157), .C2(n15454), .A(n14156), .B(n14155), .ZN(
        n14222) );
  MUX2_X1 U16138 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14222), .S(n15489), .Z(
        P2_U3525) );
  AOI21_X1 U16139 ( .B1(n15450), .B2(n14159), .A(n14158), .ZN(n14160) );
  OAI211_X1 U16140 ( .C1(n14162), .C2(n15454), .A(n14161), .B(n14160), .ZN(
        n14223) );
  MUX2_X1 U16141 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14223), .S(n15489), .Z(
        P2_U3524) );
  INV_X1 U16142 ( .A(n14163), .ZN(n14168) );
  AOI21_X1 U16143 ( .B1(n15450), .B2(n14165), .A(n14164), .ZN(n14166) );
  OAI211_X1 U16144 ( .C1(n14168), .C2(n15454), .A(n14167), .B(n14166), .ZN(
        n14224) );
  MUX2_X1 U16145 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14224), .S(n15489), .Z(
        P2_U3523) );
  AOI21_X1 U16146 ( .B1(n15450), .B2(n14170), .A(n14169), .ZN(n14171) );
  OAI211_X1 U16147 ( .C1(n14173), .C2(n15454), .A(n14172), .B(n14171), .ZN(
        n14225) );
  MUX2_X1 U16148 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14225), .S(n15489), .Z(
        P2_U3522) );
  AOI21_X1 U16149 ( .B1(n15450), .B2(n14175), .A(n14174), .ZN(n14176) );
  OAI211_X1 U16150 ( .C1(n14178), .C2(n15454), .A(n14177), .B(n14176), .ZN(
        n14226) );
  MUX2_X1 U16151 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14226), .S(n15489), .Z(
        P2_U3521) );
  AOI21_X1 U16152 ( .B1(n15450), .B2(n14180), .A(n14179), .ZN(n14181) );
  OAI211_X1 U16153 ( .C1(n14183), .C2(n15454), .A(n14182), .B(n14181), .ZN(
        n14227) );
  MUX2_X1 U16154 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14227), .S(n15489), .Z(
        P2_U3520) );
  AOI21_X1 U16155 ( .B1(n15450), .B2(n14185), .A(n14184), .ZN(n14186) );
  OAI211_X1 U16156 ( .C1(n14188), .C2(n15454), .A(n14187), .B(n14186), .ZN(
        n14228) );
  MUX2_X1 U16157 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14228), .S(n15489), .Z(
        P2_U3519) );
  AOI211_X1 U16158 ( .C1(n15450), .C2(n14191), .A(n14190), .B(n14189), .ZN(
        n14192) );
  OAI21_X1 U16159 ( .B1(n15454), .B2(n14193), .A(n14192), .ZN(n14229) );
  MUX2_X1 U16160 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14229), .S(n15489), .Z(
        P2_U3518) );
  AOI21_X1 U16161 ( .B1(n15450), .B2(n14195), .A(n14194), .ZN(n14196) );
  OAI211_X1 U16162 ( .C1(n14198), .C2(n15470), .A(n14197), .B(n14196), .ZN(
        n14230) );
  MUX2_X1 U16163 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14230), .S(n15489), .Z(
        P2_U3517) );
  AOI21_X1 U16164 ( .B1(n15450), .B2(n14200), .A(n14199), .ZN(n14201) );
  OAI211_X1 U16165 ( .C1(n15454), .C2(n14203), .A(n14202), .B(n14201), .ZN(
        n14231) );
  MUX2_X1 U16166 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14231), .S(n15489), .Z(
        P2_U3516) );
  INV_X1 U16167 ( .A(n14204), .ZN(n14206) );
  AOI211_X1 U16168 ( .C1(n15450), .C2(n14207), .A(n14206), .B(n14205), .ZN(
        n14209) );
  OAI211_X1 U16169 ( .C1(n14210), .C2(n15454), .A(n14209), .B(n14208), .ZN(
        n14232) );
  MUX2_X1 U16170 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14232), .S(n15489), .Z(
        P2_U3515) );
  AND2_X1 U16171 ( .A1(n14211), .A2(n15077), .ZN(n14216) );
  OAI21_X1 U16172 ( .B1(n7001), .B2(n15467), .A(n14212), .ZN(n14214) );
  OR3_X1 U16173 ( .A1(n14216), .A2(n14215), .A3(n14214), .ZN(n15406) );
  MUX2_X1 U16174 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n15406), .S(n15489), .Z(
        P2_U3500) );
  MUX2_X1 U16175 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14217), .S(n15475), .Z(
        P2_U3498) );
  MUX2_X1 U16176 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14218), .S(n15475), .Z(
        P2_U3497) );
  MUX2_X1 U16177 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14219), .S(n15475), .Z(
        P2_U3496) );
  MUX2_X1 U16178 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14220), .S(n15475), .Z(
        P2_U3495) );
  MUX2_X1 U16179 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14221), .S(n15475), .Z(
        P2_U3494) );
  MUX2_X1 U16180 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14222), .S(n15475), .Z(
        P2_U3493) );
  MUX2_X1 U16181 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14223), .S(n15475), .Z(
        P2_U3492) );
  MUX2_X1 U16182 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14224), .S(n15475), .Z(
        P2_U3491) );
  MUX2_X1 U16183 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14225), .S(n15475), .Z(
        P2_U3490) );
  MUX2_X1 U16184 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14226), .S(n15475), .Z(
        P2_U3489) );
  MUX2_X1 U16185 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14227), .S(n15475), .Z(
        P2_U3488) );
  MUX2_X1 U16186 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14228), .S(n15475), .Z(
        P2_U3487) );
  MUX2_X1 U16187 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14229), .S(n15475), .Z(
        P2_U3486) );
  MUX2_X1 U16188 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14230), .S(n15475), .Z(
        P2_U3484) );
  MUX2_X1 U16189 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14231), .S(n15475), .Z(
        P2_U3481) );
  MUX2_X1 U16190 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14232), .S(n15475), .Z(
        P2_U3478) );
  NAND3_X1 U16191 ( .A1(n14233), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14234) );
  OAI22_X1 U16192 ( .A1(n14235), .A2(n14234), .B1(n10585), .B2(n14249), .ZN(
        n14236) );
  AOI21_X1 U16193 ( .B1(n14237), .B2(n14246), .A(n14236), .ZN(n14238) );
  INV_X1 U16194 ( .A(n14238), .ZN(P2_U3296) );
  INV_X1 U16195 ( .A(n14239), .ZN(n14943) );
  OAI222_X1 U16196 ( .A1(n14254), .A2(n14943), .B1(P2_U3088), .B2(n14241), 
        .C1(n14240), .C2(n14252), .ZN(P2_U3298) );
  NAND2_X1 U16197 ( .A1(n14242), .A2(n14246), .ZN(n14244) );
  OAI211_X1 U16198 ( .C1(n14252), .C2(n14245), .A(n14244), .B(n14243), .ZN(
        P2_U3299) );
  NAND2_X1 U16199 ( .A1(n14945), .A2(n14246), .ZN(n14248) );
  OAI211_X1 U16200 ( .C1(n14250), .C2(n14249), .A(n14248), .B(n14247), .ZN(
        P2_U3300) );
  INV_X1 U16201 ( .A(n14251), .ZN(n14951) );
  OAI222_X1 U16202 ( .A1(n14255), .A2(P2_U3088), .B1(n14254), .B2(n14951), 
        .C1(n14253), .C2(n14252), .ZN(P2_U3301) );
  INV_X1 U16203 ( .A(n14256), .ZN(n14257) );
  MUX2_X1 U16204 ( .A(n14257), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16205 ( .A(n14837), .ZN(n14625) );
  OAI21_X1 U16206 ( .B1(n14260), .B2(n14259), .A(n14258), .ZN(n14261) );
  NAND2_X1 U16207 ( .A1(n14261), .A2(n15081), .ZN(n14265) );
  OAI22_X1 U16208 ( .A1(n14551), .A2(n15097), .B1(n14309), .B2(n15095), .ZN(
        n14836) );
  INV_X1 U16209 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14262) );
  OAI22_X1 U16210 ( .A1(n15090), .A2(n14620), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14262), .ZN(n14263) );
  AOI21_X1 U16211 ( .B1(n14836), .B2(n15105), .A(n14263), .ZN(n14264) );
  OAI211_X1 U16212 ( .C1(n14625), .C2(n14388), .A(n14265), .B(n14264), .ZN(
        P1_U3214) );
  INV_X1 U16213 ( .A(n14266), .ZN(n14267) );
  AOI21_X1 U16214 ( .B1(n14269), .B2(n14268), .A(n14267), .ZN(n14274) );
  NAND2_X1 U16215 ( .A1(n14920), .A2(n15105), .ZN(n14270) );
  NAND2_X1 U16216 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14472)
         );
  OAI211_X1 U16217 ( .C1(n15090), .C2(n14271), .A(n14270), .B(n14472), .ZN(
        n14272) );
  AOI21_X1 U16218 ( .B1(n14921), .B2(n15088), .A(n14272), .ZN(n14273) );
  OAI21_X1 U16219 ( .B1(n14274), .B2(n15101), .A(n14273), .ZN(P1_U3215) );
  INV_X1 U16220 ( .A(n14334), .ZN(n14278) );
  NOR3_X1 U16221 ( .A1(n14354), .A2(n14276), .A3(n14275), .ZN(n14277) );
  OAI21_X1 U16222 ( .B1(n14278), .B2(n14277), .A(n15081), .ZN(n14285) );
  NAND2_X1 U16223 ( .A1(n14548), .A2(n14986), .ZN(n14280) );
  NAND2_X1 U16224 ( .A1(n14577), .A2(n14987), .ZN(n14279) );
  NAND2_X1 U16225 ( .A1(n14280), .A2(n14279), .ZN(n14865) );
  INV_X1 U16226 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14281) );
  OAI22_X1 U16227 ( .A1(n14282), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14281), .ZN(n14283) );
  AOI21_X1 U16228 ( .B1(n14865), .B2(n15105), .A(n14283), .ZN(n14284) );
  OAI211_X1 U16229 ( .C1(n14679), .C2(n14388), .A(n14285), .B(n14284), .ZN(
        P1_U3216) );
  AND2_X1 U16230 ( .A1(n14359), .A2(n14286), .ZN(n14289) );
  OAI211_X1 U16231 ( .C1(n14289), .C2(n14288), .A(n15081), .B(n14287), .ZN(
        n14292) );
  OAI22_X1 U16232 ( .A1(n14571), .A2(n15097), .B1(n14542), .B2(n15095), .ZN(
        n14735) );
  NAND2_X1 U16233 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14519)
         );
  OAI21_X1 U16234 ( .B1(n15090), .B2(n14738), .A(n14519), .ZN(n14290) );
  AOI21_X1 U16235 ( .B1(n14735), .B2(n15105), .A(n14290), .ZN(n14291) );
  OAI211_X1 U16236 ( .C1(n14742), .C2(n14388), .A(n14292), .B(n14291), .ZN(
        P1_U3219) );
  OAI21_X1 U16237 ( .B1(n14294), .B2(n14293), .A(n14352), .ZN(n14295) );
  NAND2_X1 U16238 ( .A1(n14295), .A2(n15081), .ZN(n14302) );
  NAND2_X1 U16239 ( .A1(n14548), .A2(n14987), .ZN(n14297) );
  NAND2_X1 U16240 ( .A1(n14396), .A2(n14986), .ZN(n14296) );
  NAND2_X1 U16241 ( .A1(n14297), .A2(n14296), .ZN(n14704) );
  INV_X1 U16242 ( .A(n14298), .ZN(n14709) );
  OAI22_X1 U16243 ( .A1(n14709), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14299), .ZN(n14300) );
  AOI21_X1 U16244 ( .B1(n14704), .B2(n15105), .A(n14300), .ZN(n14301) );
  OAI211_X1 U16245 ( .C1(n14303), .C2(n14388), .A(n14302), .B(n14301), .ZN(
        P1_U3223) );
  NAND2_X1 U16246 ( .A1(n14647), .A2(n15283), .ZN(n14850) );
  INV_X1 U16247 ( .A(n14304), .ZN(n14308) );
  NOR3_X1 U16248 ( .A1(n14336), .A2(n14306), .A3(n14305), .ZN(n14307) );
  OAI21_X1 U16249 ( .B1(n14308), .B2(n14307), .A(n15081), .ZN(n14316) );
  OR2_X1 U16250 ( .A1(n14309), .A2(n15097), .ZN(n14311) );
  NAND2_X1 U16251 ( .A1(n14577), .A2(n14986), .ZN(n14310) );
  AND2_X1 U16252 ( .A1(n14311), .A2(n14310), .ZN(n14851) );
  INV_X1 U16253 ( .A(n14851), .ZN(n14314) );
  INV_X1 U16254 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14312) );
  OAI22_X1 U16255 ( .A1(n15090), .A2(n14644), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14312), .ZN(n14313) );
  AOI21_X1 U16256 ( .B1(n14314), .B2(n15105), .A(n14313), .ZN(n14315) );
  OAI211_X1 U16257 ( .C1(n14850), .C2(n15093), .A(n14316), .B(n14315), .ZN(
        P1_U3225) );
  AOI21_X1 U16258 ( .B1(n14318), .B2(n6996), .A(n14317), .ZN(n14323) );
  OAI22_X1 U16259 ( .A1(n14566), .A2(n15097), .B1(n14562), .B2(n15095), .ZN(
        n14774) );
  NAND2_X1 U16260 ( .A1(n14774), .A2(n15105), .ZN(n14320) );
  OAI211_X1 U16261 ( .C1(n15090), .C2(n14777), .A(n14320), .B(n14319), .ZN(
        n14321) );
  AOI21_X1 U16262 ( .B1(n14905), .B2(n15088), .A(n14321), .ZN(n14322) );
  OAI21_X1 U16263 ( .B1(n14323), .B2(n15101), .A(n14322), .ZN(P1_U3226) );
  XNOR2_X1 U16264 ( .A(n14325), .B(n14324), .ZN(n14326) );
  XNOR2_X1 U16265 ( .A(n6731), .B(n14326), .ZN(n14327) );
  NAND2_X1 U16266 ( .A1(n14327), .A2(n15081), .ZN(n14331) );
  OAI22_X1 U16267 ( .A1(n14542), .A2(n15097), .B1(n14541), .B2(n15095), .ZN(
        n14898) );
  OAI21_X1 U16268 ( .B1(n15090), .B2(n14763), .A(n14328), .ZN(n14329) );
  AOI21_X1 U16269 ( .B1(n14898), .B2(n15105), .A(n14329), .ZN(n14330) );
  OAI211_X1 U16270 ( .C1(n8244), .C2(n14388), .A(n14331), .B(n14330), .ZN(
        P1_U3228) );
  AND3_X1 U16271 ( .A1(n14334), .A2(n14333), .A3(n14332), .ZN(n14335) );
  OAI21_X1 U16272 ( .B1(n14336), .B2(n14335), .A(n15081), .ZN(n14340) );
  OAI22_X1 U16273 ( .A1(n14576), .A2(n15095), .B1(n14579), .B2(n15097), .ZN(
        n14657) );
  INV_X1 U16274 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14337) );
  OAI22_X1 U16275 ( .A1(n15090), .A2(n14663), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14337), .ZN(n14338) );
  AOI21_X1 U16276 ( .B1(n14657), .B2(n15105), .A(n14338), .ZN(n14339) );
  OAI211_X1 U16277 ( .C1(n7267), .C2(n14388), .A(n14340), .B(n14339), .ZN(
        P1_U3229) );
  XOR2_X1 U16278 ( .A(n14342), .B(n14341), .Z(n14343) );
  NAND2_X1 U16279 ( .A1(n14343), .A2(n15081), .ZN(n14349) );
  NAND2_X1 U16280 ( .A1(n14573), .A2(n14987), .ZN(n14345) );
  INV_X1 U16281 ( .A(n14570), .ZN(n14397) );
  NAND2_X1 U16282 ( .A1(n14397), .A2(n14986), .ZN(n14344) );
  NAND2_X1 U16283 ( .A1(n14345), .A2(n14344), .ZN(n14717) );
  OAI22_X1 U16284 ( .A1(n14722), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14346), .ZN(n14347) );
  AOI21_X1 U16285 ( .B1(n14717), .B2(n15105), .A(n14347), .ZN(n14348) );
  OAI211_X1 U16286 ( .C1(n10382), .C2(n14388), .A(n14349), .B(n14348), .ZN(
        P1_U3233) );
  AND3_X1 U16287 ( .A1(n14352), .A2(n14351), .A3(n14350), .ZN(n14353) );
  OAI21_X1 U16288 ( .B1(n14354), .B2(n14353), .A(n15081), .ZN(n14358) );
  OAI22_X1 U16289 ( .A1(n14576), .A2(n15097), .B1(n14546), .B2(n15095), .ZN(
        n14871) );
  INV_X1 U16290 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14355) );
  OAI22_X1 U16291 ( .A1(n14690), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14355), .ZN(n14356) );
  AOI21_X1 U16292 ( .B1(n14871), .B2(n15105), .A(n14356), .ZN(n14357) );
  OAI211_X1 U16293 ( .C1(n14388), .C2(n14692), .A(n14358), .B(n14357), .ZN(
        P1_U3235) );
  OAI21_X1 U16294 ( .B1(n14361), .B2(n14360), .A(n14359), .ZN(n14362) );
  NAND2_X1 U16295 ( .A1(n14362), .A2(n15081), .ZN(n14367) );
  NAND2_X1 U16296 ( .A1(n14565), .A2(n14986), .ZN(n14363) );
  OAI21_X1 U16297 ( .B1(n14570), .B2(n15097), .A(n14363), .ZN(n14755) );
  INV_X1 U16298 ( .A(n14749), .ZN(n14364) );
  NAND2_X1 U16299 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14486)
         );
  OAI21_X1 U16300 ( .B1(n14364), .B2(n15090), .A(n14486), .ZN(n14365) );
  AOI21_X1 U16301 ( .B1(n14755), .B2(n15105), .A(n14365), .ZN(n14366) );
  OAI211_X1 U16302 ( .C1(n14751), .C2(n14388), .A(n14367), .B(n14366), .ZN(
        P1_U3238) );
  OAI21_X1 U16303 ( .B1(n14370), .B2(n14369), .A(n14368), .ZN(n14371) );
  NAND2_X1 U16304 ( .A1(n14371), .A2(n15081), .ZN(n14377) );
  OR2_X1 U16305 ( .A1(n14550), .A2(n15097), .ZN(n14373) );
  OR2_X1 U16306 ( .A1(n14579), .A2(n15095), .ZN(n14372) );
  NAND2_X1 U16307 ( .A1(n14373), .A2(n14372), .ZN(n14842) );
  INV_X1 U16308 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14374) );
  OAI22_X1 U16309 ( .A1(n15090), .A2(n14633), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14374), .ZN(n14375) );
  AOI21_X1 U16310 ( .B1(n14842), .B2(n15105), .A(n14375), .ZN(n14376) );
  OAI211_X1 U16311 ( .C1(n7265), .C2(n14388), .A(n14377), .B(n14376), .ZN(
        P1_U3240) );
  INV_X1 U16312 ( .A(n6996), .ZN(n14385) );
  INV_X1 U16313 ( .A(n14379), .ZN(n14381) );
  NAND2_X1 U16314 ( .A1(n14381), .A2(n14380), .ZN(n14383) );
  AOI22_X1 U16315 ( .A1(n14385), .A2(n14384), .B1(n14383), .B2(n14382), .ZN(
        n14392) );
  OR2_X1 U16316 ( .A1(n14560), .A2(n15095), .ZN(n14387) );
  NAND2_X1 U16317 ( .A1(n14564), .A2(n14987), .ZN(n14386) );
  NAND2_X1 U16318 ( .A1(n14387), .A2(n14386), .ZN(n14910) );
  NAND2_X1 U16319 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15195)
         );
  OAI21_X1 U16320 ( .B1(n15090), .B2(n14792), .A(n15195), .ZN(n14390) );
  NOR2_X1 U16321 ( .A1(n14563), .A2(n14388), .ZN(n14389) );
  AOI211_X1 U16322 ( .C1(n15105), .C2(n14910), .A(n14390), .B(n14389), .ZN(
        n14391) );
  OAI21_X1 U16323 ( .B1(n14392), .B2(n15101), .A(n14391), .ZN(P1_U3241) );
  MUX2_X1 U16324 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14820), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16325 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14393), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16326 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14557), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16327 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14582), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16328 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14580), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16329 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14394), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16330 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14577), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16331 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14395), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16332 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14548), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16333 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14573), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16334 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14396), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16335 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14397), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16336 ( .A(n14398), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14409), .Z(
        P1_U3578) );
  MUX2_X1 U16337 ( .A(n14565), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14409), .Z(
        P1_U3577) );
  MUX2_X1 U16338 ( .A(n14564), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14409), .Z(
        P1_U3576) );
  MUX2_X1 U16339 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14988), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16340 ( .A(n14399), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14409), .Z(
        P1_U3572) );
  MUX2_X1 U16341 ( .A(n14985), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14409), .Z(
        P1_U3571) );
  MUX2_X1 U16342 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14400), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16343 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14401), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16344 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14402), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16345 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14403), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16346 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14404), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16347 ( .A(n14405), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14409), .Z(
        P1_U3565) );
  MUX2_X1 U16348 ( .A(n14406), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14409), .Z(
        P1_U3564) );
  MUX2_X1 U16349 ( .A(n14407), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14409), .Z(
        P1_U3563) );
  MUX2_X1 U16350 ( .A(n14408), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14409), .Z(
        P1_U3562) );
  MUX2_X1 U16351 ( .A(n14410), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14409), .Z(
        P1_U3561) );
  MUX2_X1 U16352 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14411), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16353 ( .C1(n14414), .C2(n14413), .A(n15188), .B(n14412), .ZN(
        n14421) );
  NAND2_X1 U16354 ( .A1(n14955), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14423) );
  OAI211_X1 U16355 ( .C1(n10600), .C2(n14416), .A(n14515), .B(n14415), .ZN(
        n14420) );
  AOI22_X1 U16356 ( .A1(n15177), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14419) );
  NAND2_X1 U16357 ( .A1(n14489), .A2(n14417), .ZN(n14418) );
  NAND4_X1 U16358 ( .A1(n14421), .A2(n14420), .A3(n14419), .A4(n14418), .ZN(
        P1_U3244) );
  MUX2_X1 U16359 ( .A(n14423), .B(n14422), .S(n6988), .Z(n14425) );
  NOR2_X1 U16360 ( .A1(n6988), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14424) );
  OR2_X1 U16361 ( .A1(n8555), .A2(n14424), .ZN(n15170) );
  INV_X1 U16362 ( .A(n14955), .ZN(n15172) );
  NAND2_X1 U16363 ( .A1(n15170), .A2(n15172), .ZN(n15175) );
  OAI211_X1 U16364 ( .C1(n14425), .C2(n8555), .A(P1_U4016), .B(n15175), .ZN(
        n14471) );
  NOR2_X1 U16365 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7913), .ZN(n14427) );
  AOI21_X1 U16366 ( .B1(n15177), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n14427), .ZN(
        n14428) );
  OAI21_X1 U16367 ( .B1(n15193), .B2(n14429), .A(n14428), .ZN(n14430) );
  INV_X1 U16368 ( .A(n14430), .ZN(n14439) );
  INV_X1 U16369 ( .A(n14431), .ZN(n14449) );
  OAI211_X1 U16370 ( .C1(n14433), .C2(n14432), .A(n14515), .B(n14449), .ZN(
        n14438) );
  OAI211_X1 U16371 ( .C1(n14436), .C2(n14435), .A(n15188), .B(n14434), .ZN(
        n14437) );
  NAND4_X1 U16372 ( .A1(n14471), .A2(n14439), .A3(n14438), .A4(n14437), .ZN(
        P1_U3245) );
  AND2_X1 U16373 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14441) );
  NOR2_X1 U16374 ( .A1(n15193), .A2(n14446), .ZN(n14440) );
  AOI211_X1 U16375 ( .C1(n15177), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n14441), .B(
        n14440), .ZN(n14453) );
  OAI211_X1 U16376 ( .C1(n14444), .C2(n14443), .A(n15188), .B(n14442), .ZN(
        n14452) );
  INV_X1 U16377 ( .A(n14445), .ZN(n14448) );
  MUX2_X1 U16378 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11179), .S(n14446), .Z(
        n14447) );
  NAND3_X1 U16379 ( .A1(n14449), .A2(n14448), .A3(n14447), .ZN(n14450) );
  NAND3_X1 U16380 ( .A1(n14515), .A2(n14465), .A3(n14450), .ZN(n14451) );
  NAND3_X1 U16381 ( .A1(n14453), .A2(n14452), .A3(n14451), .ZN(P1_U3246) );
  NAND2_X1 U16382 ( .A1(n15177), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14454) );
  OAI211_X1 U16383 ( .C1(n15193), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        n14457) );
  INV_X1 U16384 ( .A(n14457), .ZN(n14470) );
  INV_X1 U16385 ( .A(n14458), .ZN(n14459) );
  OAI211_X1 U16386 ( .C1(n14461), .C2(n14460), .A(n15188), .B(n14459), .ZN(
        n14469) );
  INV_X1 U16387 ( .A(n14462), .ZN(n14467) );
  NAND3_X1 U16388 ( .A1(n14465), .A2(n14464), .A3(n14463), .ZN(n14466) );
  NAND3_X1 U16389 ( .A1(n14515), .A2(n14467), .A3(n14466), .ZN(n14468) );
  NAND4_X1 U16390 ( .A1(n14471), .A2(n14470), .A3(n14469), .A4(n14468), .ZN(
        P1_U3247) );
  INV_X1 U16391 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14473) );
  OAI21_X1 U16392 ( .B1(n15197), .B2(n14473), .A(n14472), .ZN(n14474) );
  AOI21_X1 U16393 ( .B1(n14475), .B2(n14489), .A(n14474), .ZN(n14485) );
  OAI211_X1 U16394 ( .C1(n14478), .C2(n14477), .A(n14515), .B(n14476), .ZN(
        n14484) );
  OAI21_X1 U16395 ( .B1(n14481), .B2(n14480), .A(n14479), .ZN(n14482) );
  NAND2_X1 U16396 ( .A1(n15188), .A2(n14482), .ZN(n14483) );
  NAND3_X1 U16397 ( .A1(n14485), .A2(n14484), .A3(n14483), .ZN(P1_U3257) );
  INV_X1 U16398 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14487) );
  OAI21_X1 U16399 ( .B1(n15197), .B2(n14487), .A(n14486), .ZN(n14488) );
  AOI21_X1 U16400 ( .B1(n14508), .B2(n14489), .A(n14488), .ZN(n14501) );
  OAI21_X1 U16401 ( .B1(n14767), .B2(n14491), .A(n14490), .ZN(n14507) );
  XNOR2_X1 U16402 ( .A(n14502), .B(n14507), .ZN(n14492) );
  NAND2_X1 U16403 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14492), .ZN(n14510) );
  OAI211_X1 U16404 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14492), .A(n14515), 
        .B(n14510), .ZN(n14500) );
  XNOR2_X1 U16405 ( .A(n14502), .B(n14503), .ZN(n14495) );
  INV_X1 U16406 ( .A(n14495), .ZN(n14498) );
  NOR2_X1 U16407 ( .A1(n14496), .A2(n14495), .ZN(n14504) );
  INV_X1 U16408 ( .A(n14504), .ZN(n14497) );
  OAI211_X1 U16409 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14498), .A(n15188), 
        .B(n14497), .ZN(n14499) );
  NAND3_X1 U16410 ( .A1(n14501), .A2(n14500), .A3(n14499), .ZN(P1_U3261) );
  INV_X1 U16411 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14521) );
  NOR2_X1 U16412 ( .A1(n14503), .A2(n14502), .ZN(n14505) );
  XNOR2_X1 U16413 ( .A(n14506), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14516) );
  INV_X1 U16414 ( .A(n14516), .ZN(n14513) );
  NAND2_X1 U16415 ( .A1(n14508), .A2(n14507), .ZN(n14509) );
  NAND2_X1 U16416 ( .A1(n14510), .A2(n14509), .ZN(n14511) );
  XOR2_X1 U16417 ( .A(n14511), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14514) );
  OAI21_X1 U16418 ( .B1(n14514), .B2(n15183), .A(n15193), .ZN(n14512) );
  AOI21_X1 U16419 ( .B1(n14513), .B2(n15188), .A(n14512), .ZN(n14518) );
  AOI22_X1 U16420 ( .A1(n14516), .A2(n15188), .B1(n14515), .B2(n14514), .ZN(
        n14517) );
  MUX2_X1 U16421 ( .A(n14518), .B(n14517), .S(n6966), .Z(n14520) );
  OAI211_X1 U16422 ( .C1(n14521), .C2(n15197), .A(n14520), .B(n14519), .ZN(
        P1_U3262) );
  NAND2_X1 U16423 ( .A1(n15220), .A2(n15209), .ZN(n14805) );
  NAND2_X1 U16424 ( .A1(n15169), .A2(P1_B_REG_SCAN_IN), .ZN(n14523) );
  AND2_X1 U16425 ( .A1(n14987), .A2(n14523), .ZN(n14821) );
  INV_X1 U16426 ( .A(n14821), .ZN(n14524) );
  NOR2_X1 U16427 ( .A1(n14525), .A2(n14524), .ZN(n14815) );
  NAND2_X1 U16428 ( .A1(n14815), .A2(n15120), .ZN(n14531) );
  OAI21_X1 U16429 ( .B1(n15120), .B2(n14526), .A(n14531), .ZN(n14527) );
  AOI21_X1 U16430 ( .B1(n7262), .B2(n15215), .A(n14527), .ZN(n14528) );
  OAI21_X1 U16431 ( .B1(n14814), .B2(n14805), .A(n14528), .ZN(P1_U3263) );
  INV_X1 U16432 ( .A(n14587), .ZN(n14529) );
  OAI211_X1 U16433 ( .C1(n14818), .C2(n14529), .A(n7263), .B(n15209), .ZN(
        n14817) );
  NAND2_X1 U16434 ( .A1(n6676), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U16435 ( .A1(n14531), .A2(n14530), .ZN(n14532) );
  AOI21_X1 U16436 ( .B1(n14533), .B2(n15215), .A(n14532), .ZN(n14534) );
  OAI21_X1 U16437 ( .B1(n14817), .B2(n15124), .A(n14534), .ZN(P1_U3264) );
  INV_X1 U16438 ( .A(n14535), .ZN(n14537) );
  INV_X1 U16439 ( .A(n14787), .ZN(n14797) );
  INV_X1 U16440 ( .A(n14539), .ZN(n14540) );
  AOI22_X1 U16441 ( .A1(n14773), .A2(n14781), .B1(n14541), .B2(n14905), .ZN(
        n14769) );
  NOR2_X1 U16442 ( .A1(n14893), .A2(n14542), .ZN(n14733) );
  NAND2_X1 U16443 ( .A1(n14716), .A2(n14544), .ZN(n14718) );
  NAND2_X1 U16444 ( .A1(n14718), .A2(n14545), .ZN(n14701) );
  NAND2_X1 U16445 ( .A1(n14701), .A2(n14702), .ZN(n14705) );
  INV_X1 U16446 ( .A(n14661), .ZN(n14655) );
  AOI22_X2 U16447 ( .A1(n14617), .A2(n14616), .B1(n14550), .B2(n14837), .ZN(
        n14599) );
  NAND2_X1 U16448 ( .A1(n14830), .A2(n14551), .ZN(n14552) );
  NAND2_X1 U16449 ( .A1(n14599), .A2(n14552), .ZN(n14554) );
  NAND2_X1 U16450 ( .A1(n14554), .A2(n14553), .ZN(n14556) );
  INV_X1 U16451 ( .A(n14585), .ZN(n14555) );
  XNOR2_X1 U16452 ( .A(n14556), .B(n14555), .ZN(n14558) );
  INV_X1 U16453 ( .A(n14921), .ZN(n14561) );
  NOR2_X2 U16454 ( .A1(n14786), .A2(n14787), .ZN(n14785) );
  NOR2_X1 U16455 ( .A1(n14899), .A2(n14565), .ZN(n14567) );
  AOI22_X1 U16456 ( .A1(n14731), .A2(n14732), .B1(n14570), .B2(n14742), .ZN(
        n14727) );
  INV_X1 U16457 ( .A(n14577), .ZN(n14578) );
  NAND2_X1 U16458 ( .A1(n14843), .A2(n14580), .ZN(n14581) );
  XNOR2_X1 U16459 ( .A(n14586), .B(n14585), .ZN(n14819) );
  NAND2_X1 U16460 ( .A1(n14819), .A2(n15126), .ZN(n14598) );
  OAI211_X1 U16461 ( .C1(n14594), .C2(n14603), .A(n15209), .B(n14587), .ZN(
        n14824) );
  INV_X1 U16462 ( .A(n14824), .ZN(n14596) );
  INV_X1 U16463 ( .A(n14588), .ZN(n14589) );
  AOI22_X1 U16464 ( .A1(n6676), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n14589), 
        .B2(n15217), .ZN(n14593) );
  INV_X1 U16465 ( .A(n14590), .ZN(n14591) );
  NAND3_X1 U16466 ( .A1(n14820), .A2(n14821), .A3(n14591), .ZN(n14592) );
  OAI211_X1 U16467 ( .C1(n14594), .C2(n14780), .A(n14593), .B(n14592), .ZN(
        n14595) );
  AOI21_X1 U16468 ( .B1(n14596), .B2(n15220), .A(n14595), .ZN(n14597) );
  OAI211_X1 U16469 ( .C1(n14826), .C2(n6676), .A(n14598), .B(n14597), .ZN(
        P1_U3356) );
  XNOR2_X1 U16470 ( .A(n14599), .B(n14601), .ZN(n14831) );
  INV_X1 U16471 ( .A(n14831), .ZN(n14614) );
  OAI21_X1 U16472 ( .B1(n14602), .B2(n14601), .A(n14600), .ZN(n14834) );
  INV_X1 U16473 ( .A(n14834), .ZN(n14612) );
  OAI21_X1 U16474 ( .B1(n14610), .B2(n14618), .A(n15209), .ZN(n14604) );
  NOR2_X1 U16475 ( .A1(n14604), .A2(n14603), .ZN(n14828) );
  NAND2_X1 U16476 ( .A1(n14828), .A2(n15220), .ZN(n14609) );
  NAND2_X1 U16477 ( .A1(n6676), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14605) );
  OAI21_X1 U16478 ( .B1(n15117), .B2(n14606), .A(n14605), .ZN(n14607) );
  AOI21_X1 U16479 ( .B1(n14829), .B2(n15120), .A(n14607), .ZN(n14608) );
  OAI211_X1 U16480 ( .C1(n14610), .C2(n14780), .A(n14609), .B(n14608), .ZN(
        n14611) );
  AOI21_X1 U16481 ( .B1(n14612), .B2(n15126), .A(n14611), .ZN(n14613) );
  OAI21_X1 U16482 ( .B1(n14614), .B2(n14697), .A(n14613), .ZN(P1_U3265) );
  XNOR2_X1 U16483 ( .A(n14615), .B(n14616), .ZN(n14841) );
  XNOR2_X1 U16484 ( .A(n14617), .B(n14616), .ZN(n14838) );
  INV_X1 U16485 ( .A(n14634), .ZN(n14619) );
  AOI211_X1 U16486 ( .C1(n14837), .C2(n14619), .A(n14862), .B(n14618), .ZN(
        n14835) );
  NAND2_X1 U16487 ( .A1(n14835), .A2(n15220), .ZN(n14624) );
  OAI22_X1 U16488 ( .A1(n15120), .A2(n14621), .B1(n14620), .B2(n15117), .ZN(
        n14622) );
  AOI21_X1 U16489 ( .B1(n14836), .B2(n15120), .A(n14622), .ZN(n14623) );
  OAI211_X1 U16490 ( .C1(n14625), .C2(n14780), .A(n14624), .B(n14623), .ZN(
        n14626) );
  AOI21_X1 U16491 ( .B1(n14838), .B2(n14804), .A(n14626), .ZN(n14627) );
  OAI21_X1 U16492 ( .B1(n14841), .B2(n14802), .A(n14627), .ZN(P1_U3266) );
  XOR2_X1 U16493 ( .A(n14630), .B(n14628), .Z(n14849) );
  OAI21_X1 U16494 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14632) );
  INV_X1 U16495 ( .A(n14632), .ZN(n14847) );
  INV_X1 U16496 ( .A(n14633), .ZN(n14637) );
  AND2_X1 U16497 ( .A1(n14648), .A2(n14843), .ZN(n14635) );
  OR2_X1 U16498 ( .A1(n14635), .A2(n14634), .ZN(n14845) );
  NOR2_X1 U16499 ( .A1(n14845), .A2(n14710), .ZN(n14636) );
  AOI211_X1 U16500 ( .C1(n15217), .C2(n14637), .A(n14842), .B(n14636), .ZN(
        n14639) );
  AOI22_X1 U16501 ( .A1(n14843), .A2(n15215), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n6676), .ZN(n14638) );
  OAI21_X1 U16502 ( .B1(n14639), .B2(n6676), .A(n14638), .ZN(n14640) );
  AOI21_X1 U16503 ( .B1(n14847), .B2(n15126), .A(n14640), .ZN(n14641) );
  OAI21_X1 U16504 ( .B1(n14849), .B2(n14697), .A(n14641), .ZN(P1_U3267) );
  OAI21_X1 U16505 ( .B1(n6747), .B2(n14643), .A(n14642), .ZN(n14855) );
  OAI22_X1 U16506 ( .A1(n15120), .A2(n14645), .B1(n14644), .B2(n15117), .ZN(
        n14646) );
  AOI21_X1 U16507 ( .B1(n14647), .B2(n15215), .A(n14646), .ZN(n14654) );
  AOI21_X1 U16508 ( .B1(n14665), .B2(n14647), .A(n14862), .ZN(n14649) );
  NAND2_X1 U16509 ( .A1(n14649), .A2(n14648), .ZN(n14852) );
  XNOR2_X1 U16510 ( .A(n14650), .B(n7380), .ZN(n14651) );
  NAND2_X1 U16511 ( .A1(n14651), .A2(n15253), .ZN(n14853) );
  OAI211_X1 U16512 ( .C1(n6681), .C2(n14852), .A(n14853), .B(n14851), .ZN(
        n14652) );
  NAND2_X1 U16513 ( .A1(n14652), .A2(n15120), .ZN(n14653) );
  OAI211_X1 U16514 ( .C1(n14855), .C2(n14802), .A(n14654), .B(n14653), .ZN(
        P1_U3268) );
  XNOR2_X1 U16515 ( .A(n14656), .B(n14655), .ZN(n14658) );
  AOI21_X1 U16516 ( .B1(n14658), .B2(n15253), .A(n14657), .ZN(n14859) );
  AOI21_X1 U16517 ( .B1(n14661), .B2(n14660), .A(n14659), .ZN(n14860) );
  NAND2_X1 U16518 ( .A1(n6676), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n14662) );
  OAI21_X1 U16519 ( .B1(n15117), .B2(n14663), .A(n14662), .ZN(n14664) );
  AOI21_X1 U16520 ( .B1(n14857), .B2(n15215), .A(n14664), .ZN(n14668) );
  AOI21_X1 U16521 ( .B1(n14678), .B2(n14857), .A(n14862), .ZN(n14666) );
  AND2_X1 U16522 ( .A1(n14666), .A2(n14665), .ZN(n14856) );
  NAND2_X1 U16523 ( .A1(n14856), .A2(n15220), .ZN(n14667) );
  OAI211_X1 U16524 ( .C1(n14860), .C2(n14802), .A(n14668), .B(n14667), .ZN(
        n14669) );
  INV_X1 U16525 ( .A(n14669), .ZN(n14670) );
  OAI21_X1 U16526 ( .B1(n6676), .B2(n14859), .A(n14670), .ZN(P1_U3269) );
  XNOR2_X1 U16527 ( .A(n14671), .B(n14672), .ZN(n14869) );
  OR2_X1 U16528 ( .A1(n14673), .A2(n14672), .ZN(n14861) );
  NAND3_X1 U16529 ( .A1(n14861), .A2(n14674), .A3(n15126), .ZN(n14683) );
  INV_X1 U16530 ( .A(n14865), .ZN(n14677) );
  AOI22_X1 U16531 ( .A1(n14675), .A2(n15217), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n6676), .ZN(n14676) );
  OAI21_X1 U16532 ( .B1(n14677), .B2(n6676), .A(n14676), .ZN(n14681) );
  OAI21_X1 U16533 ( .B1(n14687), .B2(n14679), .A(n14678), .ZN(n14863) );
  NOR2_X1 U16534 ( .A1(n14863), .A2(n14805), .ZN(n14680) );
  AOI211_X1 U16535 ( .C1(n15215), .C2(n14866), .A(n14681), .B(n14680), .ZN(
        n14682) );
  OAI211_X1 U16536 ( .C1(n14869), .C2(n14697), .A(n14683), .B(n14682), .ZN(
        P1_U3270) );
  XOR2_X1 U16537 ( .A(n14684), .B(n14685), .Z(n14876) );
  XNOR2_X1 U16538 ( .A(n14686), .B(n14685), .ZN(n14873) );
  NAND2_X1 U16539 ( .A1(n14873), .A2(n15126), .ZN(n14696) );
  AOI211_X1 U16540 ( .C1(n14872), .C2(n14707), .A(n14862), .B(n14687), .ZN(
        n14870) );
  NAND2_X1 U16541 ( .A1(n14870), .A2(n6966), .ZN(n14689) );
  INV_X1 U16542 ( .A(n14871), .ZN(n14688) );
  OAI211_X1 U16543 ( .C1(n15117), .C2(n14690), .A(n14689), .B(n14688), .ZN(
        n14694) );
  INV_X1 U16544 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14691) );
  OAI22_X1 U16545 ( .A1(n14692), .A2(n14780), .B1(n14691), .B2(n15120), .ZN(
        n14693) );
  AOI21_X1 U16546 ( .B1(n14694), .B2(n15120), .A(n14693), .ZN(n14695) );
  OAI211_X1 U16547 ( .C1(n14876), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        P1_U3271) );
  INV_X1 U16548 ( .A(n14698), .ZN(n14699) );
  AOI21_X1 U16549 ( .B1(n14702), .B2(n14700), .A(n14699), .ZN(n14881) );
  AOI22_X1 U16550 ( .A1(n14877), .A2(n15215), .B1(n6676), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14715) );
  INV_X1 U16551 ( .A(n14701), .ZN(n14703) );
  AOI21_X1 U16552 ( .B1(n14703), .B2(n14572), .A(n15260), .ZN(n14706) );
  AOI21_X1 U16553 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14880) );
  INV_X1 U16554 ( .A(n14880), .ZN(n14713) );
  INV_X1 U16555 ( .A(n14707), .ZN(n14708) );
  AOI21_X1 U16556 ( .B1(n14877), .B2(n14720), .A(n14708), .ZN(n14878) );
  INV_X1 U16557 ( .A(n14878), .ZN(n14711) );
  OAI22_X1 U16558 ( .A1(n14711), .A2(n14710), .B1(n14709), .B2(n15117), .ZN(
        n14712) );
  OAI21_X1 U16559 ( .B1(n14713), .B2(n14712), .A(n15120), .ZN(n14714) );
  OAI211_X1 U16560 ( .C1(n14881), .C2(n14802), .A(n14715), .B(n14714), .ZN(
        P1_U3272) );
  AOI21_X1 U16561 ( .B1(n7714), .B2(n14726), .A(n15260), .ZN(n14719) );
  AOI21_X1 U16562 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14885) );
  AOI21_X1 U16563 ( .B1(n14883), .B2(n6715), .A(n14862), .ZN(n14721) );
  AND2_X1 U16564 ( .A1(n14721), .A2(n14720), .ZN(n14882) );
  INV_X1 U16565 ( .A(n14722), .ZN(n14723) );
  AOI22_X1 U16566 ( .A1(n14723), .A2(n15217), .B1(n6676), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14724) );
  OAI21_X1 U16567 ( .B1(n10382), .B2(n14780), .A(n14724), .ZN(n14729) );
  OAI21_X1 U16568 ( .B1(n14727), .B2(n14726), .A(n14725), .ZN(n14886) );
  NOR2_X1 U16569 ( .A1(n14886), .A2(n14802), .ZN(n14728) );
  AOI211_X1 U16570 ( .C1(n14882), .C2(n15220), .A(n14729), .B(n14728), .ZN(
        n14730) );
  OAI21_X1 U16571 ( .B1(n6676), .B2(n14885), .A(n14730), .ZN(P1_U3273) );
  XNOR2_X1 U16572 ( .A(n14731), .B(n7726), .ZN(n14891) );
  OAI21_X1 U16573 ( .B1(n14752), .B2(n14733), .A(n14732), .ZN(n14734) );
  AOI21_X1 U16574 ( .B1(n6761), .B2(n14734), .A(n15260), .ZN(n14736) );
  NOR2_X1 U16575 ( .A1(n14736), .A2(n14735), .ZN(n14890) );
  INV_X1 U16576 ( .A(n14890), .ZN(n14744) );
  OR2_X1 U16577 ( .A1(n14747), .A2(n14742), .ZN(n14737) );
  AND3_X1 U16578 ( .A1(n6715), .A2(n14737), .A3(n15209), .ZN(n14887) );
  NAND2_X1 U16579 ( .A1(n14887), .A2(n15220), .ZN(n14741) );
  INV_X1 U16580 ( .A(n14738), .ZN(n14739) );
  AOI22_X1 U16581 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n6676), .B1(n14739), 
        .B2(n15217), .ZN(n14740) );
  OAI211_X1 U16582 ( .C1(n14742), .C2(n14780), .A(n14741), .B(n14740), .ZN(
        n14743) );
  AOI21_X1 U16583 ( .B1(n14744), .B2(n15120), .A(n14743), .ZN(n14745) );
  OAI21_X1 U16584 ( .B1(n14891), .B2(n14802), .A(n14745), .ZN(P1_U3274) );
  XNOR2_X1 U16585 ( .A(n14746), .B(n14754), .ZN(n14896) );
  OAI21_X1 U16586 ( .B1(n14751), .B2(n14761), .A(n15209), .ZN(n14748) );
  NOR2_X1 U16587 ( .A1(n14748), .A2(n14747), .ZN(n14892) );
  AOI22_X1 U16588 ( .A1(n6676), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14749), 
        .B2(n15217), .ZN(n14750) );
  OAI21_X1 U16589 ( .B1(n14751), .B2(n14780), .A(n14750), .ZN(n14758) );
  AOI211_X1 U16590 ( .C1(n14754), .C2(n14753), .A(n15260), .B(n14752), .ZN(
        n14756) );
  NOR2_X1 U16591 ( .A1(n14756), .A2(n14755), .ZN(n14895) );
  NOR2_X1 U16592 ( .A1(n14895), .A2(n6676), .ZN(n14757) );
  AOI211_X1 U16593 ( .C1(n14892), .C2(n15220), .A(n14758), .B(n14757), .ZN(
        n14759) );
  OAI21_X1 U16594 ( .B1(n14802), .B2(n14896), .A(n14759), .ZN(P1_U3275) );
  XNOR2_X1 U16595 ( .A(n14760), .B(n14770), .ZN(n14903) );
  OAI21_X1 U16596 ( .B1(n14776), .B2(n8244), .A(n15209), .ZN(n14762) );
  NOR2_X1 U16597 ( .A1(n14762), .A2(n14761), .ZN(n14897) );
  NAND2_X1 U16598 ( .A1(n14899), .A2(n15215), .ZN(n14766) );
  NOR2_X1 U16599 ( .A1(n14763), .A2(n15117), .ZN(n14764) );
  OAI21_X1 U16600 ( .B1(n14898), .B2(n14764), .A(n15120), .ZN(n14765) );
  OAI211_X1 U16601 ( .C1(n15120), .C2(n14767), .A(n14766), .B(n14765), .ZN(
        n14768) );
  AOI21_X1 U16602 ( .B1(n14897), .B2(n15220), .A(n14768), .ZN(n14772) );
  XOR2_X1 U16603 ( .A(n14770), .B(n14769), .Z(n14900) );
  NAND2_X1 U16604 ( .A1(n14900), .A2(n14804), .ZN(n14771) );
  OAI211_X1 U16605 ( .C1(n14903), .C2(n14802), .A(n14772), .B(n14771), .ZN(
        P1_U3276) );
  XNOR2_X1 U16606 ( .A(n14773), .B(n14781), .ZN(n14775) );
  AOI21_X1 U16607 ( .B1(n14775), .B2(n15253), .A(n14774), .ZN(n14907) );
  AOI211_X1 U16608 ( .C1(n14905), .C2(n14789), .A(n14862), .B(n14776), .ZN(
        n14904) );
  INV_X1 U16609 ( .A(n14777), .ZN(n14778) );
  AOI22_X1 U16610 ( .A1(n6676), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n14778), 
        .B2(n15217), .ZN(n14779) );
  OAI21_X1 U16611 ( .B1(n7272), .B2(n14780), .A(n14779), .ZN(n14783) );
  XOR2_X1 U16612 ( .A(n14781), .B(n6821), .Z(n14908) );
  NOR2_X1 U16613 ( .A1(n14908), .A2(n14802), .ZN(n14782) );
  AOI211_X1 U16614 ( .C1(n14904), .C2(n15220), .A(n14783), .B(n14782), .ZN(
        n14784) );
  OAI21_X1 U16615 ( .B1(n6676), .B2(n14907), .A(n14784), .ZN(P1_U3277) );
  AOI21_X1 U16616 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14918) );
  AOI21_X1 U16617 ( .B1(n14911), .B2(n14788), .A(n14862), .ZN(n14790) );
  NAND2_X1 U16618 ( .A1(n14790), .A2(n14789), .ZN(n14912) );
  NAND2_X1 U16619 ( .A1(n6676), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n14791) );
  OAI21_X1 U16620 ( .B1(n15117), .B2(n14792), .A(n14791), .ZN(n14793) );
  AOI21_X1 U16621 ( .B1(n14910), .B2(n15120), .A(n14793), .ZN(n14795) );
  NAND2_X1 U16622 ( .A1(n14911), .A2(n15215), .ZN(n14794) );
  OAI211_X1 U16623 ( .C1(n14912), .C2(n15124), .A(n14795), .B(n14794), .ZN(
        n14796) );
  INV_X1 U16624 ( .A(n14796), .ZN(n14801) );
  INV_X1 U16625 ( .A(n14915), .ZN(n14799) );
  NAND2_X1 U16626 ( .A1(n14798), .A2(n14797), .ZN(n14909) );
  NAND3_X1 U16627 ( .A1(n14799), .A2(n14804), .A3(n14909), .ZN(n14800) );
  OAI211_X1 U16628 ( .C1(n14918), .C2(n14802), .A(n14801), .B(n14800), .ZN(
        P1_U3278) );
  OAI21_X1 U16629 ( .B1(n14804), .B2(n15126), .A(n14803), .ZN(n14812) );
  INV_X1 U16630 ( .A(n14805), .ZN(n14807) );
  OAI21_X1 U16631 ( .B1(n15215), .B2(n14807), .A(n14806), .ZN(n14811) );
  AOI22_X1 U16632 ( .A1(n6676), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15217), .ZN(n14810) );
  NAND2_X1 U16633 ( .A1(n14808), .A2(n15120), .ZN(n14809) );
  NAND4_X1 U16634 ( .A1(n14812), .A2(n14811), .A3(n14810), .A4(n14809), .ZN(
        P1_U3293) );
  AOI21_X1 U16635 ( .B1(n7262), .B2(n15283), .A(n14815), .ZN(n14813) );
  OAI21_X1 U16636 ( .B1(n14814), .B2(n14862), .A(n14813), .ZN(n14925) );
  MUX2_X1 U16637 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14925), .S(n15140), .Z(
        P1_U3559) );
  INV_X1 U16638 ( .A(n14815), .ZN(n14816) );
  OAI211_X1 U16639 ( .C1(n14818), .C2(n15246), .A(n14817), .B(n14816), .ZN(
        n14926) );
  MUX2_X1 U16640 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14926), .S(n15296), .Z(
        P1_U3558) );
  NAND2_X1 U16641 ( .A1(n14819), .A2(n15289), .ZN(n14827) );
  AOI22_X1 U16642 ( .A1(n14822), .A2(n15283), .B1(n14821), .B2(n14820), .ZN(
        n14823) );
  MUX2_X1 U16643 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14927), .S(n15296), .Z(
        P1_U3557) );
  AOI211_X1 U16644 ( .C1(n14830), .C2(n15283), .A(n14829), .B(n14828), .ZN(
        n14833) );
  NAND2_X1 U16645 ( .A1(n14831), .A2(n15253), .ZN(n14832) );
  OAI211_X1 U16646 ( .C1(n14834), .C2(n15248), .A(n14833), .B(n14832), .ZN(
        n14928) );
  MUX2_X1 U16647 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14928), .S(n15296), .Z(
        P1_U3556) );
  AOI211_X1 U16648 ( .C1(n14837), .C2(n15283), .A(n14836), .B(n14835), .ZN(
        n14840) );
  NAND2_X1 U16649 ( .A1(n14838), .A2(n15253), .ZN(n14839) );
  OAI211_X1 U16650 ( .C1(n14841), .C2(n15248), .A(n14840), .B(n14839), .ZN(
        n14929) );
  MUX2_X1 U16651 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14929), .S(n15296), .Z(
        P1_U3555) );
  AOI21_X1 U16652 ( .B1(n14843), .B2(n15283), .A(n14842), .ZN(n14844) );
  OAI21_X1 U16653 ( .B1(n14845), .B2(n14862), .A(n14844), .ZN(n14846) );
  AOI21_X1 U16654 ( .B1(n14847), .B2(n15289), .A(n14846), .ZN(n14848) );
  OAI21_X1 U16655 ( .B1(n15260), .B2(n14849), .A(n14848), .ZN(n14930) );
  MUX2_X1 U16656 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14930), .S(n15296), .Z(
        P1_U3554) );
  OAI211_X1 U16657 ( .C1(n14855), .C2(n15248), .A(n14854), .B(n14853), .ZN(
        n14931) );
  MUX2_X1 U16658 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14931), .S(n15296), .Z(
        P1_U3553) );
  AOI21_X1 U16659 ( .B1(n14857), .B2(n15283), .A(n14856), .ZN(n14858) );
  OAI211_X1 U16660 ( .C1(n14860), .C2(n15248), .A(n14859), .B(n14858), .ZN(
        n14932) );
  MUX2_X1 U16661 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14932), .S(n15296), .Z(
        P1_U3552) );
  NAND3_X1 U16662 ( .A1(n14861), .A2(n14674), .A3(n15289), .ZN(n14868) );
  NOR2_X1 U16663 ( .A1(n14863), .A2(n14862), .ZN(n14864) );
  AOI211_X1 U16664 ( .C1(n14866), .C2(n15283), .A(n14865), .B(n14864), .ZN(
        n14867) );
  OAI211_X1 U16665 ( .C1(n15260), .C2(n14869), .A(n14868), .B(n14867), .ZN(
        n14933) );
  MUX2_X1 U16666 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14933), .S(n15296), .Z(
        P1_U3551) );
  AOI211_X1 U16667 ( .C1(n14872), .C2(n15283), .A(n14871), .B(n14870), .ZN(
        n14875) );
  NAND2_X1 U16668 ( .A1(n14873), .A2(n15289), .ZN(n14874) );
  OAI211_X1 U16669 ( .C1(n14876), .C2(n15260), .A(n14875), .B(n14874), .ZN(
        n14934) );
  MUX2_X1 U16670 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14934), .S(n15296), .Z(
        P1_U3550) );
  AOI22_X1 U16671 ( .A1(n14878), .A2(n15209), .B1(n14877), .B2(n15283), .ZN(
        n14879) );
  OAI211_X1 U16672 ( .C1(n14881), .C2(n15248), .A(n14880), .B(n14879), .ZN(
        n14935) );
  MUX2_X1 U16673 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14935), .S(n15296), .Z(
        P1_U3549) );
  AOI21_X1 U16674 ( .B1(n14883), .B2(n15283), .A(n14882), .ZN(n14884) );
  OAI211_X1 U16675 ( .C1(n14886), .C2(n15248), .A(n14885), .B(n14884), .ZN(
        n14936) );
  MUX2_X1 U16676 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14936), .S(n15140), .Z(
        P1_U3548) );
  AOI21_X1 U16677 ( .B1(n14888), .B2(n15283), .A(n14887), .ZN(n14889) );
  OAI211_X1 U16678 ( .C1(n14891), .C2(n15248), .A(n14890), .B(n14889), .ZN(
        n14937) );
  MUX2_X1 U16679 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14937), .S(n15140), .Z(
        P1_U3547) );
  AOI21_X1 U16680 ( .B1(n14893), .B2(n15283), .A(n14892), .ZN(n14894) );
  OAI211_X1 U16681 ( .C1(n15248), .C2(n14896), .A(n14895), .B(n14894), .ZN(
        n14938) );
  MUX2_X1 U16682 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14938), .S(n15140), .Z(
        P1_U3546) );
  AOI211_X1 U16683 ( .C1(n14899), .C2(n15283), .A(n14898), .B(n14897), .ZN(
        n14902) );
  NAND2_X1 U16684 ( .A1(n14900), .A2(n15253), .ZN(n14901) );
  OAI211_X1 U16685 ( .C1(n14903), .C2(n15248), .A(n14902), .B(n14901), .ZN(
        n14939) );
  MUX2_X1 U16686 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14939), .S(n15140), .Z(
        P1_U3545) );
  AOI21_X1 U16687 ( .B1(n14905), .B2(n15283), .A(n14904), .ZN(n14906) );
  OAI211_X1 U16688 ( .C1(n14908), .C2(n15248), .A(n14907), .B(n14906), .ZN(
        n14940) );
  MUX2_X1 U16689 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14940), .S(n15140), .Z(
        P1_U3544) );
  NAND2_X1 U16690 ( .A1(n14909), .A2(n15253), .ZN(n14914) );
  AOI21_X1 U16691 ( .B1(n14911), .B2(n15283), .A(n14910), .ZN(n14913) );
  OAI211_X1 U16692 ( .C1(n14915), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        n14916) );
  INV_X1 U16693 ( .A(n14916), .ZN(n14917) );
  OAI21_X1 U16694 ( .B1(n14918), .B2(n15248), .A(n14917), .ZN(n14941) );
  MUX2_X1 U16695 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14941), .S(n15140), .Z(
        P1_U3543) );
  AOI211_X1 U16696 ( .C1(n14921), .C2(n15283), .A(n14920), .B(n14919), .ZN(
        n14923) );
  OAI211_X1 U16697 ( .C1(n14924), .C2(n15248), .A(n14923), .B(n14922), .ZN(
        n14942) );
  MUX2_X1 U16698 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14942), .S(n15140), .Z(
        P1_U3542) );
  MUX2_X1 U16699 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14925), .S(n15291), .Z(
        P1_U3527) );
  INV_X2 U16700 ( .A(n15290), .ZN(n15291) );
  MUX2_X1 U16701 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14926), .S(n15291), .Z(
        P1_U3526) );
  MUX2_X1 U16702 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14927), .S(n15291), .Z(
        P1_U3525) );
  MUX2_X1 U16703 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14928), .S(n15291), .Z(
        P1_U3524) );
  MUX2_X1 U16704 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14929), .S(n15291), .Z(
        P1_U3523) );
  MUX2_X1 U16705 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14930), .S(n15291), .Z(
        P1_U3522) );
  MUX2_X1 U16706 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14931), .S(n15291), .Z(
        P1_U3521) );
  MUX2_X1 U16707 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14932), .S(n15291), .Z(
        P1_U3520) );
  MUX2_X1 U16708 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14933), .S(n15291), .Z(
        P1_U3519) );
  MUX2_X1 U16709 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14934), .S(n15291), .Z(
        P1_U3518) );
  MUX2_X1 U16710 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14935), .S(n15291), .Z(
        P1_U3517) );
  MUX2_X1 U16711 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14936), .S(n15291), .Z(
        P1_U3516) );
  MUX2_X1 U16712 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14937), .S(n15291), .Z(
        P1_U3515) );
  MUX2_X1 U16713 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14938), .S(n15291), .Z(
        P1_U3513) );
  MUX2_X1 U16714 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14939), .S(n15291), .Z(
        P1_U3510) );
  MUX2_X1 U16715 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14940), .S(n15291), .Z(
        P1_U3507) );
  MUX2_X1 U16716 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14941), .S(n15291), .Z(
        P1_U3504) );
  MUX2_X1 U16717 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n14942), .S(n15291), .Z(
        P1_U3501) );
  OAI222_X1 U16718 ( .A1(n14949), .A2(n14944), .B1(P1_U3086), .B2(n7788), .C1(
        n12208), .C2(n14943), .ZN(P1_U3326) );
  INV_X1 U16719 ( .A(n14945), .ZN(n14948) );
  OAI222_X1 U16720 ( .A1(n14949), .A2(n7617), .B1(n12208), .B2(n14948), .C1(
        n6988), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16721 ( .A1(n14952), .A2(P1_U3086), .B1(n12208), .B2(n14951), 
        .C1(n14950), .C2(n14949), .ZN(P1_U3329) );
  MUX2_X1 U16722 ( .A(n14954), .B(n14953), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16723 ( .A(n14956), .B(n14955), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  AOI21_X1 U16724 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14959) );
  OAI21_X1 U16725 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14959), 
        .ZN(U28) );
  INV_X1 U16726 ( .A(P2_RD_REG_SCAN_IN), .ZN(n14962) );
  INV_X1 U16727 ( .A(P1_RD_REG_SCAN_IN), .ZN(n14961) );
  OAI221_X1 U16728 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n14962), .C2(n14961), .A(n14960), .ZN(U29) );
  AOI21_X1 U16729 ( .B1(n14965), .B2(n14964), .A(n14963), .ZN(n14966) );
  XOR2_X1 U16730 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n14966), .Z(SUB_1596_U61) );
  AOI21_X1 U16731 ( .B1(n14969), .B2(n14968), .A(n14967), .ZN(SUB_1596_U57) );
  AOI21_X1 U16732 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(SUB_1596_U55) );
  AOI21_X1 U16733 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n14976) );
  XOR2_X1 U16734 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14976), .Z(SUB_1596_U54) );
  OAI21_X1 U16735 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14980) );
  XNOR2_X1 U16736 ( .A(n14980), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI22_X1 U16737 ( .A1(n15120), .A2(n14981), .B1(n15091), .B2(n15117), .ZN(
        n14992) );
  XNOR2_X1 U16738 ( .A(n14982), .B(n14983), .ZN(n15001) );
  XNOR2_X1 U16739 ( .A(n14984), .B(n14983), .ZN(n14989) );
  AOI22_X1 U16740 ( .A1(n14988), .A2(n14987), .B1(n14986), .B2(n14985), .ZN(
        n15080) );
  OAI21_X1 U16741 ( .B1(n14989), .B2(n15260), .A(n15080), .ZN(n14999) );
  AOI21_X1 U16742 ( .B1(n15001), .B2(n15271), .A(n14999), .ZN(n14990) );
  NOR2_X1 U16743 ( .A1(n14990), .A2(n6676), .ZN(n14991) );
  AOI211_X1 U16744 ( .C1(n15215), .C2(n15087), .A(n14992), .B(n14991), .ZN(
        n14996) );
  OAI211_X1 U16745 ( .C1(n15113), .C2(n14998), .A(n15209), .B(n14993), .ZN(
        n14997) );
  INV_X1 U16746 ( .A(n14997), .ZN(n14994) );
  AOI22_X1 U16747 ( .A1(n15001), .A2(n15221), .B1(n15220), .B2(n14994), .ZN(
        n14995) );
  NAND2_X1 U16748 ( .A1(n14996), .A2(n14995), .ZN(P1_U3281) );
  OAI21_X1 U16749 ( .B1(n14998), .B2(n15246), .A(n14997), .ZN(n15000) );
  AOI211_X1 U16750 ( .C1(n15001), .C2(n15289), .A(n15000), .B(n14999), .ZN(
        n15003) );
  INV_X1 U16751 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U16752 ( .A1(n15291), .A2(n15003), .B1(n15002), .B2(n15290), .ZN(
        P1_U3495) );
  AOI22_X1 U16753 ( .A1(n15140), .A2(n15003), .B1(n10947), .B2(n15300), .ZN(
        P1_U3540) );
  AOI21_X1 U16754 ( .B1(n15006), .B2(n15005), .A(n15004), .ZN(n15007) );
  XOR2_X1 U16755 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n15007), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16756 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15026) );
  OAI22_X1 U16757 ( .A1(n15535), .A2(n15012), .B1(n15011), .B2(n15532), .ZN(
        n15023) );
  AOI21_X1 U16758 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15021) );
  NOR2_X1 U16759 ( .A1(n15017), .A2(n15016), .ZN(n15018) );
  OAI21_X1 U16760 ( .B1(n15019), .B2(n15018), .A(n15550), .ZN(n15020) );
  OAI21_X1 U16761 ( .B1(n15021), .B2(n15547), .A(n15020), .ZN(n15022) );
  NOR3_X1 U16762 ( .A1(n15024), .A2(n15023), .A3(n15022), .ZN(n15025) );
  OAI21_X1 U16763 ( .B1(n15026), .B2(n15515), .A(n15025), .ZN(P3_U3197) );
  INV_X1 U16764 ( .A(n15027), .ZN(n15028) );
  AOI22_X1 U16765 ( .A1(n15030), .A2(n15622), .B1(n15039), .B2(n15625), .ZN(
        n15035) );
  AOI22_X1 U16766 ( .A1(n15031), .A2(n15033), .B1(P3_REG2_REG_31__SCAN_IN), 
        .B2(n15627), .ZN(n15032) );
  NAND2_X1 U16767 ( .A1(n15035), .A2(n15032), .ZN(P3_U3202) );
  AOI22_X1 U16768 ( .A1(n15040), .A2(n15033), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15627), .ZN(n15034) );
  NAND2_X1 U16769 ( .A1(n15035), .A2(n15034), .ZN(P3_U3203) );
  OR2_X1 U16770 ( .A1(n15036), .A2(n15607), .ZN(n15038) );
  INV_X1 U16771 ( .A(n15039), .ZN(n15037) );
  AOI22_X1 U16772 ( .A1(n15693), .A2(n15060), .B1(n9626), .B2(n15691), .ZN(
        P3_U3490) );
  AOI21_X1 U16773 ( .B1(n15040), .B2(n15650), .A(n15039), .ZN(n15062) );
  AOI22_X1 U16774 ( .A1(n15693), .A2(n15062), .B1(n9615), .B2(n15691), .ZN(
        P3_U3489) );
  AOI21_X1 U16775 ( .B1(n15042), .B2(n15051), .A(n15041), .ZN(n15043) );
  AND2_X1 U16776 ( .A1(n15044), .A2(n15043), .ZN(n15064) );
  INV_X1 U16777 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n15045) );
  AOI22_X1 U16778 ( .A1(n15693), .A2(n15064), .B1(n15045), .B2(n15691), .ZN(
        P3_U3473) );
  OAI22_X1 U16779 ( .A1(n15047), .A2(n15675), .B1(n15607), .B2(n15046), .ZN(
        n15048) );
  NOR2_X1 U16780 ( .A1(n15049), .A2(n15048), .ZN(n15066) );
  AOI22_X1 U16781 ( .A1(n15693), .A2(n15066), .B1(n9815), .B2(n15691), .ZN(
        P3_U3472) );
  AOI21_X1 U16782 ( .B1(n15052), .B2(n15051), .A(n15050), .ZN(n15053) );
  AND2_X1 U16783 ( .A1(n15054), .A2(n15053), .ZN(n15068) );
  INV_X1 U16784 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U16785 ( .A1(n15693), .A2(n15068), .B1(n15055), .B2(n15691), .ZN(
        P3_U3471) );
  OAI22_X1 U16786 ( .A1(n15057), .A2(n15675), .B1(n15607), .B2(n15056), .ZN(
        n15058) );
  NOR2_X1 U16787 ( .A1(n15059), .A2(n15058), .ZN(n15070) );
  AOI22_X1 U16788 ( .A1(n15693), .A2(n15070), .B1(n12259), .B2(n15691), .ZN(
        P3_U3470) );
  INV_X1 U16789 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n15061) );
  AOI22_X1 U16790 ( .A1(n15681), .A2(n15061), .B1(n15060), .B2(n15679), .ZN(
        P3_U3458) );
  INV_X1 U16791 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n15063) );
  AOI22_X1 U16792 ( .A1(n15681), .A2(n15063), .B1(n15062), .B2(n15679), .ZN(
        P3_U3457) );
  INV_X1 U16793 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U16794 ( .A1(n15681), .A2(n15065), .B1(n15064), .B2(n15679), .ZN(
        P3_U3432) );
  INV_X1 U16795 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15067) );
  AOI22_X1 U16796 ( .A1(n15681), .A2(n15067), .B1(n15066), .B2(n15679), .ZN(
        P3_U3429) );
  INV_X1 U16797 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U16798 ( .A1(n15681), .A2(n15069), .B1(n15068), .B2(n15679), .ZN(
        P3_U3426) );
  INV_X1 U16799 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15071) );
  AOI22_X1 U16800 ( .A1(n15681), .A2(n15071), .B1(n15070), .B2(n15679), .ZN(
        P3_U3423) );
  OAI211_X1 U16801 ( .C1(n15074), .C2(n15467), .A(n15073), .B(n15072), .ZN(
        n15075) );
  AOI21_X1 U16802 ( .B1(n15077), .B2(n15076), .A(n15075), .ZN(n15078) );
  AOI22_X1 U16803 ( .A1(n15489), .A2(n15078), .B1(n10912), .B2(n15487), .ZN(
        P2_U3511) );
  AOI22_X1 U16804 ( .A1(n15475), .A2(n15078), .B1(n8838), .B2(n15474), .ZN(
        P2_U3466) );
  OAI22_X1 U16805 ( .A1(n15080), .A2(n15079), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10953), .ZN(n15086) );
  OAI211_X1 U16806 ( .C1(n6830), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15084) );
  INV_X1 U16807 ( .A(n15084), .ZN(n15085) );
  AOI211_X1 U16808 ( .C1(n15088), .C2(n15087), .A(n15086), .B(n15085), .ZN(
        n15089) );
  OAI21_X1 U16809 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(P1_U3224) );
  NAND2_X1 U16810 ( .A1(n15122), .A2(n15283), .ZN(n15135) );
  OAI22_X1 U16811 ( .A1(n15135), .A2(n15093), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15092), .ZN(n15094) );
  INV_X1 U16812 ( .A(n15094), .ZN(n15107) );
  OAI22_X1 U16813 ( .A1(n15098), .A2(n15097), .B1(n15096), .B2(n15095), .ZN(
        n15109) );
  NAND2_X1 U16814 ( .A1(n15100), .A2(n15099), .ZN(n15102) );
  AOI21_X1 U16815 ( .B1(n15103), .B2(n15102), .A(n15101), .ZN(n15104) );
  AOI21_X1 U16816 ( .B1(n15105), .B2(n15109), .A(n15104), .ZN(n15106) );
  OAI211_X1 U16817 ( .C1(n15118), .C2(n15090), .A(n15107), .B(n15106), .ZN(
        P1_U3236) );
  XOR2_X1 U16818 ( .A(n15112), .B(n15108), .Z(n15110) );
  AOI21_X1 U16819 ( .B1(n15110), .B2(n15253), .A(n15109), .ZN(n15137) );
  XOR2_X1 U16820 ( .A(n15112), .B(n15111), .Z(n15139) );
  INV_X1 U16821 ( .A(n15113), .ZN(n15114) );
  OAI211_X1 U16822 ( .C1(n15116), .C2(n15115), .A(n15114), .B(n15209), .ZN(
        n15136) );
  OAI22_X1 U16823 ( .A1(n15120), .A2(n15119), .B1(n15118), .B2(n15117), .ZN(
        n15121) );
  AOI21_X1 U16824 ( .B1(n15122), .B2(n15215), .A(n15121), .ZN(n15123) );
  OAI21_X1 U16825 ( .B1(n15136), .B2(n15124), .A(n15123), .ZN(n15125) );
  AOI21_X1 U16826 ( .B1(n15139), .B2(n15126), .A(n15125), .ZN(n15127) );
  OAI21_X1 U16827 ( .B1(n6676), .B2(n15137), .A(n15127), .ZN(P1_U3282) );
  AOI211_X1 U16828 ( .C1(n15130), .C2(n15283), .A(n15129), .B(n15128), .ZN(
        n15131) );
  OAI21_X1 U16829 ( .B1(n15132), .B2(n15260), .A(n15131), .ZN(n15133) );
  AOI21_X1 U16830 ( .B1(n15134), .B2(n15289), .A(n15133), .ZN(n15141) );
  AOI22_X1 U16831 ( .A1(n15296), .A2(n15141), .B1(n11090), .B2(n15300), .ZN(
        P1_U3541) );
  NAND3_X1 U16832 ( .A1(n15137), .A2(n15136), .A3(n15135), .ZN(n15138) );
  AOI21_X1 U16833 ( .B1(n15139), .B2(n15289), .A(n15138), .ZN(n15143) );
  AOI22_X1 U16834 ( .A1(n15140), .A2(n15143), .B1(n10834), .B2(n15300), .ZN(
        P1_U3539) );
  AOI22_X1 U16835 ( .A1(n15291), .A2(n15141), .B1(n8122), .B2(n15290), .ZN(
        P1_U3498) );
  INV_X1 U16836 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U16837 ( .A1(n15291), .A2(n15143), .B1(n15142), .B2(n15290), .ZN(
        P1_U3492) );
  AOI21_X1 U16838 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n15147) );
  XOR2_X1 U16839 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15147), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16840 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(n15151) );
  XNOR2_X1 U16841 ( .A(n15151), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI222_X1 U16842 ( .A1(n15156), .A2(n15155), .B1(n15156), .B2(n15154), .C1(
        n15153), .C2(n15152), .ZN(SUB_1596_U67) );
  OAI21_X1 U16843 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15160) );
  XNOR2_X1 U16844 ( .A(n15160), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16845 ( .B1(n15163), .B2(n15162), .A(n15161), .ZN(n15164) );
  XOR2_X1 U16846 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15164), .Z(SUB_1596_U65)
         );
  OAI21_X1 U16847 ( .B1(n15167), .B2(n15166), .A(n15165), .ZN(n15168) );
  XNOR2_X1 U16848 ( .A(n15168), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U16849 ( .A1(n15169), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15171) );
  OR2_X1 U16850 ( .A1(n15170), .A2(n15171), .ZN(n15174) );
  INV_X1 U16851 ( .A(n15171), .ZN(n15173) );
  MUX2_X1 U16852 ( .A(n15174), .B(n15173), .S(n15172), .Z(n15176) );
  NAND2_X1 U16853 ( .A1(n15176), .A2(n15175), .ZN(n15179) );
  AOI22_X1 U16854 ( .A1(n15177), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15178) );
  OAI21_X1 U16855 ( .B1(n15180), .B2(n15179), .A(n15178), .ZN(P1_U3243) );
  INV_X1 U16856 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15198) );
  AOI21_X1 U16857 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15182), .A(n15181), 
        .ZN(n15184) );
  OR2_X1 U16858 ( .A1(n15184), .A2(n15183), .ZN(n15191) );
  OAI21_X1 U16859 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n15189) );
  NAND2_X1 U16860 ( .A1(n15189), .A2(n15188), .ZN(n15190) );
  OAI211_X1 U16861 ( .C1(n15193), .C2(n15192), .A(n15191), .B(n15190), .ZN(
        n15194) );
  INV_X1 U16862 ( .A(n15194), .ZN(n15196) );
  OAI211_X1 U16863 ( .C1(n15198), .C2(n15197), .A(n15196), .B(n15195), .ZN(
        P1_U3258) );
  XNOR2_X1 U16864 ( .A(n15199), .B(n15200), .ZN(n15236) );
  XNOR2_X1 U16865 ( .A(n15202), .B(n15201), .ZN(n15203) );
  NOR2_X1 U16866 ( .A1(n15203), .A2(n15260), .ZN(n15204) );
  AOI211_X1 U16867 ( .C1(n15271), .C2(n15236), .A(n15205), .B(n15204), .ZN(
        n15233) );
  AOI222_X1 U16868 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n6676), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15217), .C1(n15206), .C2(n15215), .ZN(
        n15214) );
  INV_X1 U16869 ( .A(n15207), .ZN(n15211) );
  INV_X1 U16870 ( .A(n15208), .ZN(n15210) );
  OAI211_X1 U16871 ( .C1(n15232), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15231) );
  INV_X1 U16872 ( .A(n15231), .ZN(n15212) );
  AOI22_X1 U16873 ( .A1(n15236), .A2(n15221), .B1(n15220), .B2(n15212), .ZN(
        n15213) );
  OAI211_X1 U16874 ( .C1(n6676), .C2(n15233), .A(n15214), .B(n15213), .ZN(
        P1_U3291) );
  AOI222_X1 U16875 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n6676), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n15217), .C1(n15216), .C2(n15215), .ZN(
        n15224) );
  INV_X1 U16876 ( .A(n15218), .ZN(n15219) );
  AOI22_X1 U16877 ( .A1(n15222), .A2(n15221), .B1(n15220), .B2(n15219), .ZN(
        n15223) );
  OAI211_X1 U16878 ( .C1(n6676), .C2(n15225), .A(n15224), .B(n15223), .ZN(
        P1_U3292) );
  AND2_X1 U16879 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15226), .ZN(P1_U3294) );
  AND2_X1 U16880 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15226), .ZN(P1_U3295) );
  AND2_X1 U16881 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15226), .ZN(P1_U3296) );
  AND2_X1 U16882 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15226), .ZN(P1_U3297) );
  AND2_X1 U16883 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15226), .ZN(P1_U3298) );
  AND2_X1 U16884 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15226), .ZN(P1_U3299) );
  AND2_X1 U16885 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15226), .ZN(P1_U3300) );
  AND2_X1 U16886 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15226), .ZN(P1_U3301) );
  AND2_X1 U16887 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15226), .ZN(P1_U3302) );
  AND2_X1 U16888 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15226), .ZN(P1_U3303) );
  AND2_X1 U16889 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15226), .ZN(P1_U3304) );
  AND2_X1 U16890 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15226), .ZN(P1_U3305) );
  AND2_X1 U16891 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15226), .ZN(P1_U3306) );
  AND2_X1 U16892 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15226), .ZN(P1_U3307) );
  AND2_X1 U16893 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15226), .ZN(P1_U3308) );
  AND2_X1 U16894 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15226), .ZN(P1_U3309) );
  AND2_X1 U16895 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15226), .ZN(P1_U3310) );
  AND2_X1 U16896 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15226), .ZN(P1_U3311) );
  AND2_X1 U16897 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15226), .ZN(P1_U3312) );
  AND2_X1 U16898 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15226), .ZN(P1_U3313) );
  AND2_X1 U16899 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15226), .ZN(P1_U3314) );
  AND2_X1 U16900 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15226), .ZN(P1_U3315) );
  AND2_X1 U16901 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15226), .ZN(P1_U3316) );
  AND2_X1 U16902 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15226), .ZN(P1_U3317) );
  AND2_X1 U16903 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15226), .ZN(P1_U3318) );
  AND2_X1 U16904 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15226), .ZN(P1_U3319) );
  AND2_X1 U16905 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15226), .ZN(P1_U3320) );
  AND2_X1 U16906 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15226), .ZN(P1_U3321) );
  AND2_X1 U16907 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15226), .ZN(P1_U3322) );
  AND2_X1 U16908 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15226), .ZN(P1_U3323) );
  INV_X1 U16909 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U16910 ( .A1(n15291), .A2(n15228), .B1(n15227), .B2(n15290), .ZN(
        P1_U3459) );
  INV_X1 U16911 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U16912 ( .A1(n15291), .A2(n15230), .B1(n15229), .B2(n15290), .ZN(
        P1_U3462) );
  OAI21_X1 U16913 ( .B1(n15232), .B2(n15246), .A(n15231), .ZN(n15235) );
  INV_X1 U16914 ( .A(n15233), .ZN(n15234) );
  AOI211_X1 U16915 ( .C1(n15279), .C2(n15236), .A(n15235), .B(n15234), .ZN(
        n15292) );
  AOI22_X1 U16916 ( .A1(n15291), .A2(n15292), .B1(n7914), .B2(n15290), .ZN(
        P1_U3465) );
  OAI211_X1 U16917 ( .C1(n15239), .C2(n15246), .A(n15238), .B(n15237), .ZN(
        n15242) );
  AOI21_X1 U16918 ( .B1(n15274), .B2(n15266), .A(n15240), .ZN(n15241) );
  NOR2_X1 U16919 ( .A1(n15242), .A2(n15241), .ZN(n15293) );
  AOI22_X1 U16920 ( .A1(n15291), .A2(n15293), .B1(n7930), .B2(n15290), .ZN(
        P1_U3468) );
  INV_X1 U16921 ( .A(n15243), .ZN(n15244) );
  OAI211_X1 U16922 ( .C1(n15247), .C2(n15246), .A(n15245), .B(n15244), .ZN(
        n15251) );
  NOR2_X1 U16923 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  AOI211_X1 U16924 ( .C1(n15253), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15295) );
  AOI22_X1 U16925 ( .A1(n15291), .A2(n15295), .B1(n7954), .B2(n15290), .ZN(
        P1_U3471) );
  AOI211_X1 U16926 ( .C1(n15256), .C2(n15279), .A(n15255), .B(n15254), .ZN(
        n15258) );
  AND2_X1 U16927 ( .A1(n15258), .A2(n15257), .ZN(n15297) );
  INV_X1 U16928 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15259) );
  AOI22_X1 U16929 ( .A1(n15291), .A2(n15297), .B1(n15259), .B2(n15290), .ZN(
        P1_U3474) );
  NOR2_X1 U16930 ( .A1(n15261), .A2(n15260), .ZN(n15269) );
  INV_X1 U16931 ( .A(n15270), .ZN(n15267) );
  AOI21_X1 U16932 ( .B1(n15263), .B2(n15283), .A(n15262), .ZN(n15265) );
  OAI211_X1 U16933 ( .C1(n15267), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        n15268) );
  AOI211_X1 U16934 ( .C1(n15271), .C2(n15270), .A(n15269), .B(n15268), .ZN(
        n15298) );
  AOI22_X1 U16935 ( .A1(n15291), .A2(n15298), .B1(n8019), .B2(n15290), .ZN(
        P1_U3480) );
  OAI211_X1 U16936 ( .C1(n15275), .C2(n15274), .A(n15273), .B(n15272), .ZN(
        n15276) );
  AOI211_X1 U16937 ( .C1(n15279), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15299) );
  INV_X1 U16938 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U16939 ( .A1(n15291), .A2(n15299), .B1(n15280), .B2(n15290), .ZN(
        P1_U3486) );
  AOI211_X1 U16940 ( .C1(n15284), .C2(n15283), .A(n15282), .B(n15281), .ZN(
        n15285) );
  NAND2_X1 U16941 ( .A1(n15286), .A2(n15285), .ZN(n15287) );
  AOI21_X1 U16942 ( .B1(n15289), .B2(n15288), .A(n15287), .ZN(n15301) );
  AOI22_X1 U16943 ( .A1(n15291), .A2(n15301), .B1(n8080), .B2(n15290), .ZN(
        P1_U3489) );
  AOI22_X1 U16944 ( .A1(n15296), .A2(n15292), .B1(n10590), .B2(n15300), .ZN(
        P1_U3530) );
  AOI22_X1 U16945 ( .A1(n15296), .A2(n15293), .B1(n10591), .B2(n15300), .ZN(
        P1_U3531) );
  AOI22_X1 U16946 ( .A1(n15296), .A2(n15295), .B1(n15294), .B2(n15300), .ZN(
        P1_U3532) );
  AOI22_X1 U16947 ( .A1(n15296), .A2(n15297), .B1(n10593), .B2(n15300), .ZN(
        P1_U3533) );
  AOI22_X1 U16948 ( .A1(n15296), .A2(n15298), .B1(n10616), .B2(n15300), .ZN(
        P1_U3535) );
  AOI22_X1 U16949 ( .A1(n15296), .A2(n15299), .B1(n10669), .B2(n15300), .ZN(
        P1_U3537) );
  AOI22_X1 U16950 ( .A1(n15296), .A2(n15301), .B1(n10727), .B2(n15300), .ZN(
        P1_U3538) );
  NOR2_X1 U16951 ( .A1(n15371), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16952 ( .A(n15302), .ZN(n15304) );
  OAI21_X1 U16953 ( .B1(n15304), .B2(n15303), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15305) );
  OAI21_X1 U16954 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15305), .ZN(n15316) );
  OAI211_X1 U16955 ( .C1(n15308), .C2(n15307), .A(n15364), .B(n15306), .ZN(
        n15309) );
  INV_X1 U16956 ( .A(n15309), .ZN(n15310) );
  AOI21_X1 U16957 ( .B1(n15371), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n15310), .ZN(
        n15315) );
  OAI211_X1 U16958 ( .C1(n15313), .C2(n15312), .A(n15372), .B(n15311), .ZN(
        n15314) );
  NAND3_X1 U16959 ( .A1(n15316), .A2(n15315), .A3(n15314), .ZN(P2_U3216) );
  OAI211_X1 U16960 ( .C1(n15319), .C2(n15318), .A(n15364), .B(n15317), .ZN(
        n15322) );
  INV_X1 U16961 ( .A(n15320), .ZN(n15321) );
  OAI211_X1 U16962 ( .C1(n15379), .C2(n15323), .A(n15322), .B(n15321), .ZN(
        n15324) );
  INV_X1 U16963 ( .A(n15324), .ZN(n15329) );
  OAI211_X1 U16964 ( .C1(n15327), .C2(n15326), .A(n15372), .B(n15325), .ZN(
        n15328) );
  OAI211_X1 U16965 ( .C1(n15363), .C2(n15698), .A(n15329), .B(n15328), .ZN(
        P2_U3219) );
  NAND2_X1 U16966 ( .A1(n15331), .A2(n15330), .ZN(n15332) );
  NAND2_X1 U16967 ( .A1(n15333), .A2(n15332), .ZN(n15334) );
  NAND2_X1 U16968 ( .A1(n15372), .A2(n15334), .ZN(n15341) );
  NAND2_X1 U16969 ( .A1(n15336), .A2(n15335), .ZN(n15337) );
  NAND2_X1 U16970 ( .A1(n15338), .A2(n15337), .ZN(n15339) );
  NAND2_X1 U16971 ( .A1(n15339), .A2(n15364), .ZN(n15340) );
  OAI211_X1 U16972 ( .C1(n15379), .C2(n15342), .A(n15341), .B(n15340), .ZN(
        n15343) );
  INV_X1 U16973 ( .A(n15343), .ZN(n15345) );
  OAI211_X1 U16974 ( .C1(n6938), .C2(n15363), .A(n15345), .B(n15344), .ZN(
        P2_U3223) );
  INV_X1 U16975 ( .A(n15346), .ZN(n15351) );
  NAND3_X1 U16976 ( .A1(n15349), .A2(n15348), .A3(n15347), .ZN(n15350) );
  NAND2_X1 U16977 ( .A1(n15351), .A2(n15350), .ZN(n15360) );
  NAND2_X1 U16978 ( .A1(n15353), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n15352) );
  OAI21_X1 U16979 ( .B1(n15353), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15352), 
        .ZN(n15355) );
  OAI21_X1 U16980 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15357) );
  AOI222_X1 U16981 ( .A1(n15360), .A2(n15372), .B1(n15359), .B2(n15358), .C1(
        n15357), .C2(n15364), .ZN(n15362) );
  OAI211_X1 U16982 ( .C1(n6927), .C2(n15363), .A(n15362), .B(n15361), .ZN(
        P2_U3226) );
  OAI21_X1 U16983 ( .B1(n15366), .B2(n15365), .A(n15364), .ZN(n15368) );
  NOR2_X1 U16984 ( .A1(n15368), .A2(n15367), .ZN(n15369) );
  AOI211_X1 U16985 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n15371), .A(n15370), 
        .B(n15369), .ZN(n15377) );
  OAI211_X1 U16986 ( .C1(n15375), .C2(n15374), .A(n15373), .B(n15372), .ZN(
        n15376) );
  OAI211_X1 U16987 ( .C1(n15379), .C2(n15378), .A(n15377), .B(n15376), .ZN(
        P2_U3231) );
  INV_X1 U16988 ( .A(n15380), .ZN(n15382) );
  NOR2_X1 U16989 ( .A1(n15382), .A2(n15381), .ZN(n15404) );
  INV_X1 U16990 ( .A(n15404), .ZN(n15386) );
  OAI22_X1 U16991 ( .A1(n15386), .A2(n15385), .B1(n15384), .B2(n15383), .ZN(
        n15390) );
  OAI21_X1 U16992 ( .B1(n15460), .B2(n14129), .A(n15405), .ZN(n15387) );
  OAI21_X1 U16993 ( .B1(n15389), .B2(n15388), .A(n15387), .ZN(n15403) );
  AOI211_X1 U16994 ( .C1(n15391), .C2(n15405), .A(n15390), .B(n15403), .ZN(
        n15393) );
  AOI22_X1 U16995 ( .A1(n15394), .A2(n8640), .B1(n15393), .B2(n15392), .ZN(
        P2_U3265) );
  AND2_X1 U16996 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15397), .ZN(P2_U3266) );
  AND2_X1 U16997 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15397), .ZN(P2_U3267) );
  AND2_X1 U16998 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15397), .ZN(P2_U3268) );
  AND2_X1 U16999 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15397), .ZN(P2_U3269) );
  AND2_X1 U17000 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15397), .ZN(P2_U3270) );
  AND2_X1 U17001 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15397), .ZN(P2_U3271) );
  AND2_X1 U17002 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15397), .ZN(P2_U3272) );
  AND2_X1 U17003 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15397), .ZN(P2_U3273) );
  AND2_X1 U17004 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15397), .ZN(P2_U3274) );
  AND2_X1 U17005 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15397), .ZN(P2_U3275) );
  AND2_X1 U17006 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15397), .ZN(P2_U3276) );
  AND2_X1 U17007 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15397), .ZN(P2_U3277) );
  AND2_X1 U17008 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15397), .ZN(P2_U3278) );
  AND2_X1 U17009 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15397), .ZN(P2_U3279) );
  AND2_X1 U17010 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15397), .ZN(P2_U3280) );
  AND2_X1 U17011 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15397), .ZN(P2_U3281) );
  AND2_X1 U17012 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15397), .ZN(P2_U3282) );
  AND2_X1 U17013 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15397), .ZN(P2_U3283) );
  AND2_X1 U17014 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15397), .ZN(P2_U3284) );
  AND2_X1 U17015 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15397), .ZN(P2_U3285) );
  AND2_X1 U17016 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15397), .ZN(P2_U3286) );
  AND2_X1 U17017 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15397), .ZN(P2_U3287) );
  AND2_X1 U17018 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15397), .ZN(P2_U3288) );
  AND2_X1 U17019 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15397), .ZN(P2_U3289) );
  AND2_X1 U17020 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15397), .ZN(P2_U3290) );
  AND2_X1 U17021 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15397), .ZN(P2_U3291) );
  AND2_X1 U17022 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15397), .ZN(P2_U3292) );
  AND2_X1 U17023 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15397), .ZN(P2_U3293) );
  AND2_X1 U17024 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15397), .ZN(P2_U3294) );
  AND2_X1 U17025 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15397), .ZN(P2_U3295) );
  INV_X1 U17026 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15399) );
  OAI21_X1 U17027 ( .B1(n15401), .B2(n15399), .A(n15398), .ZN(P2_U3416) );
  INV_X1 U17028 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15402) );
  OAI21_X1 U17029 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(P2_U3417) );
  INV_X1 U17030 ( .A(n15470), .ZN(n15459) );
  AOI211_X1 U17031 ( .C1(n15459), .C2(n15405), .A(n15404), .B(n15403), .ZN(
        n15476) );
  AOI22_X1 U17032 ( .A1(n15475), .A2(n15476), .B1(n7157), .B2(n15474), .ZN(
        P2_U3430) );
  INV_X1 U17033 ( .A(n15406), .ZN(n15407) );
  AOI22_X1 U17034 ( .A1(n15475), .A2(n15407), .B1(n8634), .B2(n15474), .ZN(
        P2_U3433) );
  AOI22_X1 U17035 ( .A1(n15475), .A2(n15408), .B1(n8654), .B2(n15474), .ZN(
        P2_U3436) );
  AOI21_X1 U17036 ( .B1(n15450), .B2(n15410), .A(n15409), .ZN(n15411) );
  OAI211_X1 U17037 ( .C1(n15454), .C2(n15413), .A(n15412), .B(n15411), .ZN(
        n15414) );
  INV_X1 U17038 ( .A(n15414), .ZN(n15477) );
  INV_X1 U17039 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U17040 ( .A1(n15475), .A2(n15477), .B1(n15415), .B2(n15474), .ZN(
        P2_U3439) );
  AOI21_X1 U17041 ( .B1(n15450), .B2(n15417), .A(n15416), .ZN(n15418) );
  OAI211_X1 U17042 ( .C1(n15454), .C2(n15420), .A(n15419), .B(n15418), .ZN(
        n15421) );
  INV_X1 U17043 ( .A(n15421), .ZN(n15479) );
  AOI22_X1 U17044 ( .A1(n15475), .A2(n15479), .B1(n8686), .B2(n15474), .ZN(
        P2_U3442) );
  AOI21_X1 U17045 ( .B1(n15450), .B2(n15423), .A(n15422), .ZN(n15424) );
  OAI211_X1 U17046 ( .C1(n15426), .C2(n15470), .A(n15425), .B(n15424), .ZN(
        n15427) );
  INV_X1 U17047 ( .A(n15427), .ZN(n15481) );
  AOI22_X1 U17048 ( .A1(n15475), .A2(n15481), .B1(n8705), .B2(n15474), .ZN(
        P2_U3445) );
  AOI21_X1 U17049 ( .B1(n15450), .B2(n15429), .A(n15428), .ZN(n15430) );
  OAI211_X1 U17050 ( .C1(n15432), .C2(n15470), .A(n15431), .B(n15430), .ZN(
        n15433) );
  INV_X1 U17051 ( .A(n15433), .ZN(n15482) );
  AOI22_X1 U17052 ( .A1(n15475), .A2(n15482), .B1(n8726), .B2(n15474), .ZN(
        P2_U3448) );
  NAND2_X1 U17053 ( .A1(n15434), .A2(n15450), .ZN(n15437) );
  INV_X1 U17054 ( .A(n15435), .ZN(n15436) );
  OAI211_X1 U17055 ( .C1(n15438), .C2(n15454), .A(n15437), .B(n15436), .ZN(
        n15439) );
  INV_X1 U17056 ( .A(n15439), .ZN(n15441) );
  AND2_X1 U17057 ( .A1(n15441), .A2(n15440), .ZN(n15483) );
  AOI22_X1 U17058 ( .A1(n15475), .A2(n15483), .B1(n8745), .B2(n15474), .ZN(
        P2_U3451) );
  INV_X1 U17059 ( .A(n15442), .ZN(n15447) );
  INV_X1 U17060 ( .A(n15443), .ZN(n15444) );
  OAI21_X1 U17061 ( .B1(n7347), .B2(n15467), .A(n15444), .ZN(n15446) );
  AOI211_X1 U17062 ( .C1(n15459), .C2(n15447), .A(n15446), .B(n15445), .ZN(
        n15484) );
  AOI22_X1 U17063 ( .A1(n15475), .A2(n15484), .B1(n8764), .B2(n15474), .ZN(
        P2_U3454) );
  AOI21_X1 U17064 ( .B1(n15450), .B2(n15449), .A(n15448), .ZN(n15452) );
  OAI211_X1 U17065 ( .C1(n15454), .C2(n15453), .A(n15452), .B(n15451), .ZN(
        n15455) );
  INV_X1 U17066 ( .A(n15455), .ZN(n15485) );
  AOI22_X1 U17067 ( .A1(n15475), .A2(n15485), .B1(n8783), .B2(n15474), .ZN(
        P2_U3457) );
  OAI21_X1 U17068 ( .B1(n15457), .B2(n15467), .A(n15456), .ZN(n15458) );
  AOI21_X1 U17069 ( .B1(n15461), .B2(n15459), .A(n15458), .ZN(n15464) );
  NAND2_X1 U17070 ( .A1(n15461), .A2(n15460), .ZN(n15462) );
  AOI22_X1 U17071 ( .A1(n15475), .A2(n15486), .B1(n8804), .B2(n15474), .ZN(
        P2_U3460) );
  OAI211_X1 U17072 ( .C1(n15468), .C2(n15467), .A(n15466), .B(n15465), .ZN(
        n15473) );
  AOI21_X1 U17073 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(n15472) );
  NOR2_X1 U17074 ( .A1(n15473), .A2(n15472), .ZN(n15488) );
  AOI22_X1 U17075 ( .A1(n15475), .A2(n15488), .B1(n8820), .B2(n15474), .ZN(
        P2_U3463) );
  AOI22_X1 U17076 ( .A1(n15489), .A2(n15476), .B1(n10797), .B2(n15487), .ZN(
        P2_U3499) );
  AOI22_X1 U17077 ( .A1(n15489), .A2(n15477), .B1(n10777), .B2(n15487), .ZN(
        P2_U3502) );
  INV_X1 U17078 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U17079 ( .A1(n15489), .A2(n15479), .B1(n15478), .B2(n15487), .ZN(
        P2_U3503) );
  AOI22_X1 U17080 ( .A1(n15489), .A2(n15481), .B1(n15480), .B2(n15487), .ZN(
        P2_U3504) );
  AOI22_X1 U17081 ( .A1(n15489), .A2(n15482), .B1(n8720), .B2(n15487), .ZN(
        P2_U3505) );
  AOI22_X1 U17082 ( .A1(n15489), .A2(n15483), .B1(n8741), .B2(n15487), .ZN(
        P2_U3506) );
  AOI22_X1 U17083 ( .A1(n15489), .A2(n15484), .B1(n8760), .B2(n15487), .ZN(
        P2_U3507) );
  AOI22_X1 U17084 ( .A1(n15489), .A2(n15485), .B1(n8778), .B2(n15487), .ZN(
        P2_U3508) );
  AOI22_X1 U17085 ( .A1(n15489), .A2(n15486), .B1(n10804), .B2(n15487), .ZN(
        P2_U3509) );
  AOI22_X1 U17086 ( .A1(n15489), .A2(n15488), .B1(n10855), .B2(n15487), .ZN(
        P2_U3510) );
  NOR2_X1 U17087 ( .A1(P3_U3897), .A2(n15538), .ZN(P3_U3150) );
  AOI22_X1 U17088 ( .A1(n15492), .A2(n15491), .B1(n11366), .B2(n15490), .ZN(
        n15496) );
  NAND2_X1 U17089 ( .A1(n15494), .A2(n15493), .ZN(n15495) );
  AND2_X1 U17090 ( .A1(n15496), .A2(n15495), .ZN(n15497) );
  OAI21_X1 U17091 ( .B1(n15498), .B2(n15505), .A(n15497), .ZN(P3_U3172) );
  NOR3_X1 U17092 ( .A1(n15539), .A2(n15500), .A3(n15550), .ZN(n15512) );
  AOI22_X1 U17093 ( .A1(n15539), .A2(n15501), .B1(n15500), .B2(n15499), .ZN(
        n15510) );
  NOR2_X1 U17094 ( .A1(n15520), .A2(n15502), .ZN(n15504) );
  MUX2_X1 U17095 ( .A(n15504), .B(n15503), .S(P3_IR_REG_0__SCAN_IN), .Z(n15508) );
  OAI22_X1 U17096 ( .A1(n15532), .A2(n15506), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15505), .ZN(n15507) );
  NOR2_X1 U17097 ( .A1(n15508), .A2(n15507), .ZN(n15509) );
  OAI211_X1 U17098 ( .C1(n15512), .C2(n15511), .A(n15510), .B(n15509), .ZN(
        P3_U3182) );
  NAND2_X1 U17099 ( .A1(n15514), .A2(n15513), .ZN(n15516) );
  AOI21_X1 U17100 ( .B1(n15517), .B2(n15516), .A(n15515), .ZN(n15529) );
  XOR2_X1 U17101 ( .A(n15519), .B(n15518), .Z(n15521) );
  OAI22_X1 U17102 ( .A1(n15535), .A2(n15522), .B1(n15521), .B2(n15520), .ZN(
        n15528) );
  NAND2_X1 U17103 ( .A1(n15524), .A2(n15523), .ZN(n15525) );
  AOI21_X1 U17104 ( .B1(n15526), .B2(n15525), .A(n15547), .ZN(n15527) );
  NOR3_X1 U17105 ( .A1(n15529), .A2(n15528), .A3(n15527), .ZN(n15531) );
  OAI211_X1 U17106 ( .C1(n15533), .C2(n15532), .A(n15531), .B(n15530), .ZN(
        P3_U3190) );
  NOR2_X1 U17107 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  AOI211_X1 U17108 ( .C1(n15538), .C2(P3_ADDR_REG_12__SCAN_IN), .A(n15537), 
        .B(n15536), .ZN(n15556) );
  OAI221_X1 U17109 ( .B1(n15542), .B2(n15541), .C1(n15542), .C2(n15540), .A(
        n15539), .ZN(n15555) );
  INV_X1 U17110 ( .A(n15543), .ZN(n15544) );
  AOI21_X1 U17111 ( .B1(n15546), .B2(n15545), .A(n15544), .ZN(n15548) );
  OR2_X1 U17112 ( .A1(n15548), .A2(n15547), .ZN(n15554) );
  OAI211_X1 U17113 ( .C1(n15552), .C2(n15551), .A(n15550), .B(n15549), .ZN(
        n15553) );
  NAND4_X1 U17114 ( .A1(n15556), .A2(n15555), .A3(n15554), .A4(n15553), .ZN(
        P3_U3194) );
  XNOR2_X1 U17115 ( .A(n15557), .B(n15561), .ZN(n15647) );
  INV_X1 U17116 ( .A(n15558), .ZN(n15559) );
  AOI21_X1 U17117 ( .B1(n15561), .B2(n15560), .A(n15559), .ZN(n15566) );
  AOI22_X1 U17118 ( .A1(n15615), .A2(n15563), .B1(n15562), .B2(n15613), .ZN(
        n15565) );
  NAND2_X1 U17119 ( .A1(n15647), .A2(n15656), .ZN(n15564) );
  OAI211_X1 U17120 ( .C1(n15566), .C2(n15619), .A(n15565), .B(n15564), .ZN(
        n15645) );
  AOI21_X1 U17121 ( .B1(n15605), .B2(n15647), .A(n15645), .ZN(n15571) );
  AND2_X1 U17122 ( .A1(n15650), .A2(n15567), .ZN(n15646) );
  AOI22_X1 U17123 ( .A1(n15583), .A2(n15646), .B1(n15622), .B2(n15568), .ZN(
        n15569) );
  OAI221_X1 U17124 ( .B1(n15627), .B2(n15571), .C1(n15625), .C2(n15570), .A(
        n15569), .ZN(P3_U3228) );
  XNOR2_X1 U17125 ( .A(n15576), .B(n15572), .ZN(n15580) );
  INV_X1 U17126 ( .A(n15580), .ZN(n15643) );
  AOI22_X1 U17127 ( .A1(n15613), .A2(n15574), .B1(n15573), .B2(n15615), .ZN(
        n15579) );
  OAI211_X1 U17128 ( .C1(n15577), .C2(n15576), .A(n15575), .B(n15599), .ZN(
        n15578) );
  OAI211_X1 U17129 ( .C1(n15580), .C2(n15602), .A(n15579), .B(n15578), .ZN(
        n15641) );
  AOI21_X1 U17130 ( .B1(n15605), .B2(n15643), .A(n15641), .ZN(n15586) );
  AND2_X1 U17131 ( .A1(n15650), .A2(n15581), .ZN(n15642) );
  AOI22_X1 U17132 ( .A1(n15583), .A2(n15642), .B1(n15622), .B2(n15582), .ZN(
        n15584) );
  OAI221_X1 U17133 ( .B1(n15627), .B2(n15586), .C1(n15625), .C2(n15585), .A(
        n15584), .ZN(P3_U3229) );
  XNOR2_X1 U17134 ( .A(n15587), .B(n15593), .ZN(n15603) );
  INV_X1 U17135 ( .A(n15603), .ZN(n15634) );
  INV_X1 U17136 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15590) );
  NOR2_X1 U17137 ( .A1(n15607), .A2(n15588), .ZN(n15633) );
  INV_X1 U17138 ( .A(n15633), .ZN(n15589) );
  OAI22_X1 U17139 ( .A1(n15591), .A2(n15590), .B1(n15589), .B2(n15609), .ZN(
        n15604) );
  XNOR2_X1 U17140 ( .A(n15592), .B(n15593), .ZN(n15600) );
  OAI22_X1 U17141 ( .A1(n15597), .A2(n15596), .B1(n15595), .B2(n15594), .ZN(
        n15598) );
  AOI21_X1 U17142 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n15601) );
  OAI21_X1 U17143 ( .B1(n15603), .B2(n15602), .A(n15601), .ZN(n15632) );
  AOI211_X1 U17144 ( .C1(n15605), .C2(n15634), .A(n15604), .B(n15632), .ZN(
        n15606) );
  AOI22_X1 U17145 ( .A1(n15627), .A2(n11562), .B1(n15606), .B2(n15625), .ZN(
        P3_U3231) );
  NOR2_X1 U17146 ( .A1(n15608), .A2(n15607), .ZN(n15629) );
  INV_X1 U17147 ( .A(n15609), .ZN(n15621) );
  XNOR2_X1 U17148 ( .A(n15611), .B(n15610), .ZN(n15620) );
  AOI22_X1 U17149 ( .A1(n15615), .A2(n15614), .B1(n15613), .B2(n15612), .ZN(
        n15618) );
  XNOR2_X1 U17150 ( .A(n15616), .B(n11492), .ZN(n15630) );
  NAND2_X1 U17151 ( .A1(n15630), .A2(n15656), .ZN(n15617) );
  OAI211_X1 U17152 ( .C1(n15620), .C2(n15619), .A(n15618), .B(n15617), .ZN(
        n15628) );
  AOI21_X1 U17153 ( .B1(n15629), .B2(n15621), .A(n15628), .ZN(n15626) );
  AOI22_X1 U17154 ( .A1(n15623), .A2(n15630), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15622), .ZN(n15624) );
  OAI221_X1 U17155 ( .B1(n15627), .B2(n15626), .C1(n15625), .C2(n11535), .A(
        n15624), .ZN(P3_U3232) );
  INV_X1 U17156 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15631) );
  AOI211_X1 U17157 ( .C1(n15672), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        n15682) );
  AOI22_X1 U17158 ( .A1(n15681), .A2(n15631), .B1(n15682), .B2(n15679), .ZN(
        P3_U3393) );
  INV_X1 U17159 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15635) );
  AOI211_X1 U17160 ( .C1(n15634), .C2(n15672), .A(n15633), .B(n15632), .ZN(
        n15683) );
  AOI22_X1 U17161 ( .A1(n15681), .A2(n15635), .B1(n15683), .B2(n15679), .ZN(
        P3_U3396) );
  INV_X1 U17162 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15640) );
  INV_X1 U17163 ( .A(n15636), .ZN(n15637) );
  AOI211_X1 U17164 ( .C1(n15639), .C2(n15672), .A(n15638), .B(n15637), .ZN(
        n15684) );
  AOI22_X1 U17165 ( .A1(n15681), .A2(n15640), .B1(n15684), .B2(n15679), .ZN(
        P3_U3399) );
  INV_X1 U17166 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15644) );
  AOI211_X1 U17167 ( .C1(n15643), .C2(n15672), .A(n15642), .B(n15641), .ZN(
        n15685) );
  AOI22_X1 U17168 ( .A1(n15681), .A2(n15644), .B1(n15685), .B2(n15679), .ZN(
        P3_U3402) );
  INV_X1 U17169 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15648) );
  AOI211_X1 U17170 ( .C1(n15647), .C2(n15672), .A(n15646), .B(n15645), .ZN(
        n15686) );
  AOI22_X1 U17171 ( .A1(n15681), .A2(n15648), .B1(n15686), .B2(n15679), .ZN(
        P3_U3405) );
  INV_X1 U17172 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15658) );
  INV_X1 U17173 ( .A(n15653), .ZN(n15657) );
  NAND2_X1 U17174 ( .A1(n15650), .A2(n15649), .ZN(n15651) );
  OAI211_X1 U17175 ( .C1(n15654), .C2(n15653), .A(n15652), .B(n15651), .ZN(
        n15655) );
  AOI21_X1 U17176 ( .B1(n15657), .B2(n15656), .A(n15655), .ZN(n15687) );
  AOI22_X1 U17177 ( .A1(n15681), .A2(n15658), .B1(n15687), .B2(n15679), .ZN(
        P3_U3408) );
  INV_X1 U17178 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15662) );
  AOI211_X1 U17179 ( .C1(n15661), .C2(n15672), .A(n15660), .B(n15659), .ZN(
        n15688) );
  AOI22_X1 U17180 ( .A1(n15681), .A2(n15662), .B1(n15688), .B2(n15679), .ZN(
        P3_U3411) );
  INV_X1 U17181 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15667) );
  INV_X1 U17182 ( .A(n15663), .ZN(n15666) );
  AOI211_X1 U17183 ( .C1(n15666), .C2(n15672), .A(n15665), .B(n15664), .ZN(
        n15689) );
  AOI22_X1 U17184 ( .A1(n15681), .A2(n15667), .B1(n15689), .B2(n15679), .ZN(
        P3_U3414) );
  INV_X1 U17185 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15673) );
  INV_X1 U17186 ( .A(n15668), .ZN(n15671) );
  AOI211_X1 U17187 ( .C1(n15672), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15690) );
  AOI22_X1 U17188 ( .A1(n15681), .A2(n15673), .B1(n15690), .B2(n15679), .ZN(
        P3_U3417) );
  INV_X1 U17189 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15680) );
  OAI21_X1 U17190 ( .B1(n15676), .B2(n15675), .A(n15674), .ZN(n15677) );
  NOR2_X1 U17191 ( .A1(n15678), .A2(n15677), .ZN(n15692) );
  AOI22_X1 U17192 ( .A1(n15681), .A2(n15680), .B1(n15692), .B2(n15679), .ZN(
        P3_U3420) );
  AOI22_X1 U17193 ( .A1(n15693), .A2(n15682), .B1(n11534), .B2(n15691), .ZN(
        P3_U3460) );
  AOI22_X1 U17194 ( .A1(n15693), .A2(n15683), .B1(n11574), .B2(n15691), .ZN(
        P3_U3461) );
  AOI22_X1 U17195 ( .A1(n15693), .A2(n15684), .B1(n11545), .B2(n15691), .ZN(
        P3_U3462) );
  AOI22_X1 U17196 ( .A1(n15693), .A2(n15685), .B1(n9671), .B2(n15691), .ZN(
        P3_U3463) );
  AOI22_X1 U17197 ( .A1(n15693), .A2(n15686), .B1(n9691), .B2(n15691), .ZN(
        P3_U3464) );
  AOI22_X1 U17198 ( .A1(n15693), .A2(n15687), .B1(n9706), .B2(n15691), .ZN(
        P3_U3465) );
  AOI22_X1 U17199 ( .A1(n15693), .A2(n15688), .B1(n11860), .B2(n15691), .ZN(
        P3_U3466) );
  AOI22_X1 U17200 ( .A1(n15693), .A2(n15689), .B1(n9734), .B2(n15691), .ZN(
        P3_U3467) );
  AOI22_X1 U17201 ( .A1(n15693), .A2(n15690), .B1(n9752), .B2(n15691), .ZN(
        P3_U3468) );
  AOI22_X1 U17202 ( .A1(n15693), .A2(n15692), .B1(n12000), .B2(n15691), .ZN(
        P3_U3469) );
  AOI21_X1 U17203 ( .B1(n15696), .B2(n15695), .A(n15694), .ZN(SUB_1596_U59) );
  OAI21_X1 U17204 ( .B1(n15699), .B2(n15698), .A(n15697), .ZN(SUB_1596_U58) );
  XOR2_X1 U17205 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15700), .Z(SUB_1596_U53) );
  AOI21_X1 U17206 ( .B1(n15703), .B2(n15702), .A(n15701), .ZN(SUB_1596_U56) );
  OAI21_X1 U17207 ( .B1(n15706), .B2(n15705), .A(n15704), .ZN(n15707) );
  XNOR2_X1 U17208 ( .A(n15707), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17209 ( .B1(n15710), .B2(n15709), .A(n15708), .ZN(SUB_1596_U5) );
  NAND2_X1 U9375 ( .A1(n8590), .A2(n8597), .ZN(n8721) );
  CLKBUF_X1 U7462 ( .A(n10417), .Z(n6967) );
  NAND2_X1 U7481 ( .A1(n11104), .A2(n8774), .ZN(n11165) );
  CLKBUF_X1 U7482 ( .A(n13729), .Z(n6990) );
  NAND2_X1 U7537 ( .A1(n8597), .A2(n14241), .ZN(n8656) );
  CLKBUF_X1 U7560 ( .A(n14033), .Z(n6995) );
  CLKBUF_X1 U7616 ( .A(n8263), .Z(n6681) );
  NAND2_X1 U7644 ( .A1(n7482), .A2(n7481), .ZN(n13774) );
  CLKBUF_X1 U8133 ( .A(n14213), .Z(n7001) );
  OR2_X2 U8646 ( .A1(n13162), .A2(n11535), .ZN(n13164) );
  XNOR2_X1 U9507 ( .A(n13190), .B(n13173), .ZN(n12270) );
endmodule

